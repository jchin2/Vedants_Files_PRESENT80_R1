magic
tech sky130A
timestamp 1670909827
<< nmoslvt >>
rect -935 10 -885 485
rect -825 10 -775 485
rect -715 10 -665 485
rect -605 10 -555 485
<< ndiff >>
rect -995 470 -935 485
rect -995 25 -975 470
rect -955 25 -935 470
rect -995 10 -935 25
rect -885 470 -825 485
rect -885 25 -865 470
rect -845 25 -825 470
rect -885 10 -825 25
rect -775 470 -715 485
rect -775 25 -755 470
rect -735 25 -715 470
rect -775 10 -715 25
rect -665 470 -605 485
rect -665 25 -645 470
rect -625 25 -605 470
rect -665 10 -605 25
rect -555 470 -495 485
rect -555 25 -535 470
rect -515 25 -495 470
rect -555 10 -495 25
<< ndiffc >>
rect -975 25 -955 470
rect -865 25 -845 470
rect -755 25 -735 470
rect -645 25 -625 470
rect -535 25 -515 470
<< psubdiff >>
rect -1055 465 -995 485
rect -1055 30 -1035 465
rect -1015 30 -995 465
rect -1055 10 -995 30
<< psubdiffcont >>
rect -1035 30 -1015 465
<< poly >>
rect -935 510 -555 525
rect -935 485 -885 510
rect -825 485 -775 510
rect -715 485 -665 510
rect -605 485 -555 510
rect -935 -5 -885 10
rect -825 -5 -775 10
rect -715 -5 -665 10
rect -605 -5 -555 10
<< locali >>
rect -865 495 -625 515
rect -865 475 -845 495
rect -645 475 -625 495
rect -1045 465 -1005 475
rect -1045 30 -1035 465
rect -1015 30 -1005 465
rect -1045 20 -1005 30
rect -985 470 -945 475
rect -985 25 -975 470
rect -955 25 -945 470
rect -985 20 -945 25
rect -875 470 -835 475
rect -875 25 -865 470
rect -845 25 -835 470
rect -875 20 -835 25
rect -765 470 -725 475
rect -765 25 -755 470
rect -735 25 -725 470
rect -765 20 -725 25
rect -655 470 -615 475
rect -655 25 -645 470
rect -625 25 -615 470
rect -655 20 -615 25
rect -545 470 -505 475
rect -545 25 -535 470
rect -515 25 -505 470
rect -545 20 -505 25
rect -975 0 -955 20
rect -755 0 -735 20
rect -535 0 -515 20
rect -975 -20 -515 0
<< end >>
