magic
tech sky130A
magscale 1 2
timestamp 1670968230
<< poly >>
rect -2850 7904 -2784 7970
rect 1250 7917 1316 7983
rect -2838 7885 -2784 7904
rect 1268 7855 1298 7917
rect 2756 7904 2822 7970
rect 2768 7885 2822 7904
rect -1338 6753 -1308 6824
rect -1356 6687 -1290 6753
<< locali >>
rect -37898 17197 -3290 17220
rect -37898 17163 -37852 17197
rect -37818 17163 -37772 17197
rect -37738 17163 -37692 17197
rect -37658 17163 -37612 17197
rect -37578 17163 -37532 17197
rect -37498 17163 -37452 17197
rect -37418 17163 -37372 17197
rect -37338 17163 -37292 17197
rect -37258 17163 -37212 17197
rect -37178 17163 -37132 17197
rect -37098 17163 -37052 17197
rect -37018 17163 -36972 17197
rect -36938 17163 -36892 17197
rect -36858 17163 -36812 17197
rect -36778 17163 -36732 17197
rect -36698 17163 -36652 17197
rect -36618 17163 -36572 17197
rect -36538 17163 -36492 17197
rect -36458 17163 -36412 17197
rect -36378 17163 -36332 17197
rect -36298 17163 -36252 17197
rect -36218 17163 -36172 17197
rect -36138 17163 -36092 17197
rect -36058 17163 -36012 17197
rect -35978 17163 -35932 17197
rect -35898 17163 -35852 17197
rect -35818 17163 -35772 17197
rect -35738 17163 -35692 17197
rect -35658 17163 -35612 17197
rect -35578 17163 -35532 17197
rect -35498 17163 -35452 17197
rect -35418 17163 -35372 17197
rect -35338 17163 -35292 17197
rect -35258 17163 -35212 17197
rect -35178 17163 -35132 17197
rect -35098 17163 -35052 17197
rect -35018 17163 -34972 17197
rect -34938 17163 -34892 17197
rect -34858 17163 -34812 17197
rect -34778 17163 -34732 17197
rect -34698 17163 -34652 17197
rect -34618 17163 -34572 17197
rect -34538 17163 -34492 17197
rect -34458 17163 -34412 17197
rect -34378 17163 -34332 17197
rect -34298 17163 -34252 17197
rect -34218 17163 -34172 17197
rect -34138 17163 -34092 17197
rect -34058 17163 -34012 17197
rect -33978 17163 -33932 17197
rect -33898 17163 -33852 17197
rect -33818 17163 -33772 17197
rect -33738 17163 -33692 17197
rect -33658 17163 -33612 17197
rect -33578 17163 -33532 17197
rect -33498 17163 -33452 17197
rect -33418 17163 -33372 17197
rect -33338 17163 -33292 17197
rect -33258 17163 -33212 17197
rect -33178 17163 -33132 17197
rect -33098 17163 -33052 17197
rect -33018 17163 -32972 17197
rect -32938 17163 -32892 17197
rect -32858 17163 -32812 17197
rect -32778 17163 -32732 17197
rect -32698 17163 -32652 17197
rect -32618 17163 -32572 17197
rect -32538 17163 -32492 17197
rect -32458 17163 -32412 17197
rect -32378 17163 -32332 17197
rect -32298 17163 -32252 17197
rect -32218 17163 -32172 17197
rect -32138 17163 -32092 17197
rect -32058 17163 -32012 17197
rect -31978 17163 -31932 17197
rect -31898 17163 -31852 17197
rect -31818 17163 -31772 17197
rect -31738 17163 -31692 17197
rect -31658 17163 -31612 17197
rect -31578 17163 -31532 17197
rect -31498 17163 -31452 17197
rect -31418 17163 -31372 17197
rect -31338 17163 -31292 17197
rect -31258 17163 -31212 17197
rect -31178 17163 -31132 17197
rect -31098 17163 -31052 17197
rect -31018 17163 -30972 17197
rect -30938 17163 -30892 17197
rect -30858 17163 -30812 17197
rect -30778 17163 -30732 17197
rect -30698 17163 -30652 17197
rect -30618 17163 -30572 17197
rect -30538 17163 -30492 17197
rect -30458 17163 -30412 17197
rect -30378 17163 -30332 17197
rect -30298 17163 -30252 17197
rect -30218 17163 -30172 17197
rect -30138 17163 -30092 17197
rect -30058 17163 -30012 17197
rect -29978 17163 -29932 17197
rect -29898 17163 -29852 17197
rect -29818 17163 -29772 17197
rect -29738 17163 -29692 17197
rect -29658 17163 -29612 17197
rect -29578 17163 -29532 17197
rect -29498 17163 -29452 17197
rect -29418 17163 -29372 17197
rect -29338 17163 -29292 17197
rect -29258 17163 -29212 17197
rect -29178 17163 -29132 17197
rect -29098 17163 -29052 17197
rect -29018 17163 -28972 17197
rect -28938 17163 -28892 17197
rect -28858 17163 -28812 17197
rect -28778 17163 -28732 17197
rect -28698 17163 -28652 17197
rect -28618 17163 -28572 17197
rect -28538 17163 -28492 17197
rect -28458 17163 -28412 17197
rect -28378 17163 -28332 17197
rect -28298 17163 -28252 17197
rect -28218 17163 -28172 17197
rect -28138 17163 -28092 17197
rect -28058 17163 -28012 17197
rect -27978 17163 -27932 17197
rect -27898 17163 -27852 17197
rect -27818 17163 -27772 17197
rect -27738 17163 -27692 17197
rect -27658 17163 -27612 17197
rect -27578 17163 -27532 17197
rect -27498 17163 -27452 17197
rect -27418 17163 -27372 17197
rect -27338 17163 -27292 17197
rect -27258 17163 -27212 17197
rect -27178 17163 -27132 17197
rect -27098 17163 -27052 17197
rect -27018 17163 -26972 17197
rect -26938 17163 -26892 17197
rect -26858 17163 -26812 17197
rect -26778 17163 -26732 17197
rect -26698 17163 -26652 17197
rect -26618 17163 -26572 17197
rect -26538 17163 -26492 17197
rect -26458 17163 -26412 17197
rect -26378 17163 -26332 17197
rect -26298 17163 -26252 17197
rect -26218 17163 -26172 17197
rect -26138 17163 -26092 17197
rect -26058 17163 -26012 17197
rect -25978 17163 -25932 17197
rect -25898 17163 -25852 17197
rect -25818 17163 -25772 17197
rect -25738 17163 -25692 17197
rect -25658 17163 -25612 17197
rect -25578 17163 -25532 17197
rect -25498 17163 -25452 17197
rect -25418 17163 -25372 17197
rect -25338 17163 -25292 17197
rect -25258 17163 -25212 17197
rect -25178 17163 -25132 17197
rect -25098 17163 -25052 17197
rect -25018 17163 -24972 17197
rect -24938 17163 -24891 17197
rect -24857 17163 -24811 17197
rect -24777 17163 -24731 17197
rect -24697 17163 -24651 17197
rect -24617 17163 -24571 17197
rect -24537 17163 -24491 17197
rect -24457 17163 -24411 17197
rect -24377 17163 -24331 17197
rect -24297 17163 -24251 17197
rect -24217 17163 -24171 17197
rect -24137 17163 -24091 17197
rect -24057 17163 -24011 17197
rect -23977 17163 -23931 17197
rect -23897 17163 -23851 17197
rect -23817 17163 -23771 17197
rect -23737 17163 -23691 17197
rect -23657 17163 -23611 17197
rect -23577 17163 -23531 17197
rect -23497 17163 -23451 17197
rect -23417 17163 -23371 17197
rect -23337 17163 -23291 17197
rect -23257 17163 -23211 17197
rect -23177 17163 -23131 17197
rect -23097 17163 -23051 17197
rect -23017 17163 -22971 17197
rect -22937 17163 -22891 17197
rect -22857 17163 -22811 17197
rect -22777 17163 -22731 17197
rect -22697 17163 -22651 17197
rect -22617 17163 -22571 17197
rect -22537 17163 -22491 17197
rect -22457 17163 -22411 17197
rect -22377 17163 -22331 17197
rect -22297 17163 -22251 17197
rect -22217 17163 -22171 17197
rect -22137 17163 -22091 17197
rect -22057 17163 -22011 17197
rect -21977 17163 -21931 17197
rect -21897 17163 -21851 17197
rect -21817 17163 -21771 17197
rect -21737 17163 -21691 17197
rect -21657 17163 -21611 17197
rect -21577 17163 -21531 17197
rect -21497 17163 -21451 17197
rect -21417 17163 -21371 17197
rect -21337 17163 -21291 17197
rect -21257 17163 -21211 17197
rect -21177 17163 -21131 17197
rect -21097 17163 -21051 17197
rect -21017 17163 -20971 17197
rect -20937 17163 -20891 17197
rect -20857 17163 -20811 17197
rect -20777 17163 -20731 17197
rect -20697 17163 -20651 17197
rect -20617 17163 -20571 17197
rect -20537 17163 -20491 17197
rect -20457 17163 -20411 17197
rect -20377 17163 -20331 17197
rect -20297 17163 -20251 17197
rect -20217 17163 -20171 17197
rect -20137 17163 -20091 17197
rect -20057 17163 -20011 17197
rect -19977 17163 -19931 17197
rect -19897 17163 -19851 17197
rect -19817 17163 -19771 17197
rect -19737 17163 -19691 17197
rect -19657 17163 -19611 17197
rect -19577 17163 -19531 17197
rect -19497 17163 -19451 17197
rect -19417 17163 -19371 17197
rect -19337 17163 -19291 17197
rect -19257 17163 -19211 17197
rect -19177 17163 -19131 17197
rect -19097 17163 -19051 17197
rect -19017 17163 -18971 17197
rect -18937 17163 -18891 17197
rect -18857 17163 -18811 17197
rect -18777 17163 -18731 17197
rect -18697 17163 -18651 17197
rect -18617 17163 -18571 17197
rect -18537 17163 -18491 17197
rect -18457 17163 -18411 17197
rect -18377 17163 -18331 17197
rect -18297 17163 -18251 17197
rect -18217 17163 -18171 17197
rect -18137 17163 -18091 17197
rect -18057 17163 -18011 17197
rect -17977 17163 -17931 17197
rect -17897 17163 -17851 17197
rect -17817 17163 -17771 17197
rect -17737 17163 -17691 17197
rect -17657 17163 -17611 17197
rect -17577 17163 -17531 17197
rect -17497 17163 -17451 17197
rect -17417 17163 -17371 17197
rect -17337 17163 -17291 17197
rect -17257 17163 -17211 17197
rect -17177 17163 -17131 17197
rect -17097 17163 -17051 17197
rect -17017 17163 -16971 17197
rect -16937 17163 -16891 17197
rect -16857 17163 -16811 17197
rect -16777 17163 -16731 17197
rect -16697 17163 -16651 17197
rect -16617 17163 -16571 17197
rect -16537 17163 -16491 17197
rect -16457 17163 -16411 17197
rect -16377 17163 -16331 17197
rect -16297 17163 -16251 17197
rect -16217 17163 -16171 17197
rect -16137 17163 -16091 17197
rect -16057 17163 -16011 17197
rect -15977 17163 -15931 17197
rect -15897 17163 -15851 17197
rect -15817 17163 -15771 17197
rect -15737 17163 -15691 17197
rect -15657 17163 -15611 17197
rect -15577 17163 -15531 17197
rect -15497 17163 -15451 17197
rect -15417 17163 -15371 17197
rect -15337 17163 -15291 17197
rect -15257 17163 -15211 17197
rect -15177 17163 -15131 17197
rect -15097 17163 -15051 17197
rect -15017 17163 -14971 17197
rect -14937 17163 -14891 17197
rect -14857 17163 -14811 17197
rect -14777 17163 -14731 17197
rect -14697 17163 -14651 17197
rect -14617 17163 -14571 17197
rect -14537 17163 -14491 17197
rect -14457 17163 -14411 17197
rect -14377 17163 -14331 17197
rect -14297 17163 -14251 17197
rect -14217 17163 -14171 17197
rect -14137 17163 -14091 17197
rect -14057 17163 -14011 17197
rect -13977 17163 -13931 17197
rect -13897 17163 -13851 17197
rect -13817 17163 -13771 17197
rect -13737 17163 -13691 17197
rect -13657 17163 -13611 17197
rect -13577 17163 -13531 17197
rect -13497 17163 -13451 17197
rect -13417 17163 -13371 17197
rect -13337 17163 -13291 17197
rect -13257 17163 -13211 17197
rect -13177 17163 -13131 17197
rect -13097 17163 -13051 17197
rect -13017 17163 -12971 17197
rect -12937 17163 -12891 17197
rect -12857 17163 -12811 17197
rect -12777 17163 -12731 17197
rect -12697 17163 -12651 17197
rect -12617 17163 -12571 17197
rect -12537 17163 -12491 17197
rect -12457 17163 -12411 17197
rect -12377 17163 -12331 17197
rect -12297 17163 -12251 17197
rect -12217 17163 -12171 17197
rect -12137 17163 -12091 17197
rect -12057 17163 -12011 17197
rect -11977 17163 -11930 17197
rect -11896 17163 -11850 17197
rect -11816 17163 -11770 17197
rect -11736 17163 -11690 17197
rect -11656 17163 -11610 17197
rect -11576 17163 -11530 17197
rect -11496 17163 -11450 17197
rect -11416 17163 -11370 17197
rect -11336 17163 -11290 17197
rect -11256 17163 -11210 17197
rect -11176 17163 -11130 17197
rect -11096 17163 -11050 17197
rect -11016 17163 -10970 17197
rect -10936 17163 -10890 17197
rect -10856 17163 -10810 17197
rect -10776 17163 -10730 17197
rect -10696 17163 -10650 17197
rect -10616 17163 -10570 17197
rect -10536 17163 -10490 17197
rect -10456 17163 -10410 17197
rect -10376 17163 -10330 17197
rect -10296 17163 -10250 17197
rect -10216 17163 -10170 17197
rect -10136 17163 -10090 17197
rect -10056 17163 -10010 17197
rect -9976 17163 -9930 17197
rect -9896 17163 -9850 17197
rect -9816 17163 -9770 17197
rect -9736 17163 -9690 17197
rect -9656 17163 -9610 17197
rect -9576 17163 -9530 17197
rect -9496 17163 -9450 17197
rect -9416 17163 -9370 17197
rect -9336 17163 -9290 17197
rect -9256 17163 -9210 17197
rect -9176 17163 -9130 17197
rect -9096 17163 -9050 17197
rect -9016 17163 -8970 17197
rect -8936 17163 -8890 17197
rect -8856 17163 -8810 17197
rect -8776 17163 -8730 17197
rect -8696 17163 -8650 17197
rect -8616 17163 -8570 17197
rect -8536 17163 -8490 17197
rect -8456 17163 -8410 17197
rect -8376 17163 -8330 17197
rect -8296 17163 -8250 17197
rect -8216 17163 -8170 17197
rect -8136 17163 -8090 17197
rect -8056 17163 -8010 17197
rect -7976 17163 -7930 17197
rect -7896 17163 -7850 17197
rect -7816 17163 -7770 17197
rect -7736 17163 -7690 17197
rect -7656 17163 -7610 17197
rect -7576 17163 -7530 17197
rect -7496 17163 -7450 17197
rect -7416 17163 -7370 17197
rect -7336 17163 -7290 17197
rect -7256 17163 -7210 17197
rect -7176 17163 -7130 17197
rect -7096 17163 -7050 17197
rect -7016 17163 -6970 17197
rect -6936 17163 -6890 17197
rect -6856 17163 -6810 17197
rect -6776 17163 -6730 17197
rect -6696 17163 -6650 17197
rect -6616 17163 -6570 17197
rect -6536 17163 -6490 17197
rect -6456 17163 -6410 17197
rect -6376 17163 -6330 17197
rect -6296 17163 -6250 17197
rect -6216 17163 -6170 17197
rect -6136 17163 -6090 17197
rect -6056 17163 -6010 17197
rect -5976 17163 -5930 17197
rect -5896 17163 -5850 17197
rect -5816 17163 -5770 17197
rect -5736 17163 -5690 17197
rect -5656 17163 -5610 17197
rect -5576 17163 -5530 17197
rect -5496 17163 -5450 17197
rect -5416 17163 -5370 17197
rect -5336 17163 -5290 17197
rect -5256 17163 -5210 17197
rect -5176 17163 -5130 17197
rect -5096 17163 -5050 17197
rect -5016 17163 -4970 17197
rect -4936 17163 -4890 17197
rect -4856 17163 -4810 17197
rect -4776 17163 -4730 17197
rect -4696 17163 -4650 17197
rect -4616 17163 -4570 17197
rect -4536 17163 -4490 17197
rect -4456 17163 -4410 17197
rect -4376 17163 -4330 17197
rect -4296 17163 -4250 17197
rect -4216 17163 -4170 17197
rect -4136 17163 -4090 17197
rect -4056 17163 -4010 17197
rect -3976 17163 -3930 17197
rect -3896 17163 -3850 17197
rect -3816 17163 -3770 17197
rect -3736 17163 -3690 17197
rect -3656 17163 -3610 17197
rect -3576 17163 -3530 17197
rect -3496 17163 -3450 17197
rect -3416 17163 -3370 17197
rect -3336 17163 -3290 17197
rect -37898 17140 -3290 17163
rect -1942 17197 2397 17220
rect -1942 17163 -1929 17197
rect -1895 17163 -1849 17197
rect -1815 17163 -1769 17197
rect -1735 17163 -1689 17197
rect -1655 17163 -1609 17197
rect -1575 17163 -1529 17197
rect -1495 17163 -1449 17197
rect -1415 17163 -1369 17197
rect -1335 17163 -1289 17197
rect -1255 17163 -1209 17197
rect -1175 17163 -1129 17197
rect -1095 17163 -1049 17197
rect -1015 17163 -969 17197
rect -935 17163 -889 17197
rect -855 17163 -809 17197
rect -775 17163 -729 17197
rect -695 17163 -649 17197
rect -615 17163 -569 17197
rect -535 17163 -489 17197
rect -455 17163 -409 17197
rect -375 17163 -329 17197
rect -295 17163 -249 17197
rect -215 17163 -169 17197
rect -135 17163 -89 17197
rect -55 17163 -9 17197
rect 25 17163 71 17197
rect 105 17163 151 17197
rect 185 17163 231 17197
rect 265 17163 311 17197
rect 345 17163 391 17197
rect 425 17163 471 17197
rect 505 17163 551 17197
rect 585 17163 631 17197
rect 665 17163 711 17197
rect 745 17163 791 17197
rect 825 17163 871 17197
rect 905 17163 951 17197
rect 985 17163 1031 17197
rect 1065 17163 1111 17197
rect 1145 17163 1191 17197
rect 1225 17163 1271 17197
rect 1305 17163 1351 17197
rect 1385 17163 1431 17197
rect 1465 17163 1511 17197
rect 1545 17163 1591 17197
rect 1625 17163 1671 17197
rect 1705 17163 1751 17197
rect 1785 17163 1831 17197
rect 1865 17163 1911 17197
rect 1945 17163 1991 17197
rect 2025 17163 2071 17197
rect 2105 17163 2151 17197
rect 2185 17163 2231 17197
rect 2265 17163 2311 17197
rect 2345 17163 2397 17197
rect -1942 17140 2397 17163
rect 3744 17197 38351 17220
rect 3744 17163 3790 17197
rect 3824 17163 3870 17197
rect 3904 17163 3950 17197
rect 3984 17163 4030 17197
rect 4064 17163 4110 17197
rect 4144 17163 4190 17197
rect 4224 17163 4270 17197
rect 4304 17163 4350 17197
rect 4384 17163 4430 17197
rect 4464 17163 4510 17197
rect 4544 17163 4590 17197
rect 4624 17163 4670 17197
rect 4704 17163 4750 17197
rect 4784 17163 4830 17197
rect 4864 17163 4910 17197
rect 4944 17163 4990 17197
rect 5024 17163 5070 17197
rect 5104 17163 5150 17197
rect 5184 17163 5230 17197
rect 5264 17163 5310 17197
rect 5344 17163 5390 17197
rect 5424 17163 5470 17197
rect 5504 17163 5550 17197
rect 5584 17163 5630 17197
rect 5664 17163 5710 17197
rect 5744 17163 5790 17197
rect 5824 17163 5870 17197
rect 5904 17163 5950 17197
rect 5984 17163 6030 17197
rect 6064 17163 6110 17197
rect 6144 17163 6190 17197
rect 6224 17163 6270 17197
rect 6304 17163 6350 17197
rect 6384 17163 6430 17197
rect 6464 17163 6510 17197
rect 6544 17163 6590 17197
rect 6624 17163 6670 17197
rect 6704 17163 6750 17197
rect 6784 17163 6830 17197
rect 6864 17163 6910 17197
rect 6944 17163 6990 17197
rect 7024 17163 7070 17197
rect 7104 17163 7150 17197
rect 7184 17163 7230 17197
rect 7264 17163 7310 17197
rect 7344 17163 7390 17197
rect 7424 17163 7470 17197
rect 7504 17163 7550 17197
rect 7584 17163 7630 17197
rect 7664 17163 7710 17197
rect 7744 17163 7790 17197
rect 7824 17163 7870 17197
rect 7904 17163 7950 17197
rect 7984 17163 8030 17197
rect 8064 17163 8110 17197
rect 8144 17163 8190 17197
rect 8224 17163 8270 17197
rect 8304 17163 8350 17197
rect 8384 17163 8430 17197
rect 8464 17163 8510 17197
rect 8544 17163 8590 17197
rect 8624 17163 8670 17197
rect 8704 17163 8750 17197
rect 8784 17163 8830 17197
rect 8864 17163 8910 17197
rect 8944 17163 8990 17197
rect 9024 17163 9070 17197
rect 9104 17163 9150 17197
rect 9184 17163 9230 17197
rect 9264 17163 9310 17197
rect 9344 17163 9390 17197
rect 9424 17163 9470 17197
rect 9504 17163 9550 17197
rect 9584 17163 9630 17197
rect 9664 17163 9710 17197
rect 9744 17163 9790 17197
rect 9824 17163 9870 17197
rect 9904 17163 9950 17197
rect 9984 17163 10030 17197
rect 10064 17163 10110 17197
rect 10144 17163 10190 17197
rect 10224 17163 10270 17197
rect 10304 17163 10350 17197
rect 10384 17163 10430 17197
rect 10464 17163 10510 17197
rect 10544 17163 10590 17197
rect 10624 17163 10670 17197
rect 10704 17163 10750 17197
rect 10784 17163 10830 17197
rect 10864 17163 10910 17197
rect 10944 17163 10990 17197
rect 11024 17163 11070 17197
rect 11104 17163 11150 17197
rect 11184 17163 11230 17197
rect 11264 17163 11310 17197
rect 11344 17163 11390 17197
rect 11424 17163 11470 17197
rect 11504 17163 11550 17197
rect 11584 17163 11630 17197
rect 11664 17163 11710 17197
rect 11744 17163 11790 17197
rect 11824 17163 11870 17197
rect 11904 17163 11950 17197
rect 11984 17163 12030 17197
rect 12064 17163 12110 17197
rect 12144 17163 12190 17197
rect 12224 17163 12270 17197
rect 12304 17163 12350 17197
rect 12384 17163 12430 17197
rect 12464 17163 12510 17197
rect 12544 17163 12590 17197
rect 12624 17163 12670 17197
rect 12704 17163 12750 17197
rect 12784 17163 12830 17197
rect 12864 17163 12910 17197
rect 12944 17163 12990 17197
rect 13024 17163 13070 17197
rect 13104 17163 13150 17197
rect 13184 17163 13230 17197
rect 13264 17163 13310 17197
rect 13344 17163 13390 17197
rect 13424 17163 13470 17197
rect 13504 17163 13550 17197
rect 13584 17163 13630 17197
rect 13664 17163 13710 17197
rect 13744 17163 13790 17197
rect 13824 17163 13870 17197
rect 13904 17163 13950 17197
rect 13984 17163 14030 17197
rect 14064 17163 14110 17197
rect 14144 17163 14190 17197
rect 14224 17163 14270 17197
rect 14304 17163 14350 17197
rect 14384 17163 14430 17197
rect 14464 17163 14510 17197
rect 14544 17163 14590 17197
rect 14624 17163 14670 17197
rect 14704 17163 14750 17197
rect 14784 17163 14830 17197
rect 14864 17163 14910 17197
rect 14944 17163 14990 17197
rect 15024 17163 15070 17197
rect 15104 17163 15150 17197
rect 15184 17163 15230 17197
rect 15264 17163 15310 17197
rect 15344 17163 15390 17197
rect 15424 17163 15470 17197
rect 15504 17163 15550 17197
rect 15584 17163 15630 17197
rect 15664 17163 15710 17197
rect 15744 17163 15790 17197
rect 15824 17163 15870 17197
rect 15904 17163 15950 17197
rect 15984 17163 16030 17197
rect 16064 17163 16110 17197
rect 16144 17163 16190 17197
rect 16224 17163 16270 17197
rect 16304 17163 16350 17197
rect 16384 17163 16430 17197
rect 16464 17163 16510 17197
rect 16544 17163 16590 17197
rect 16624 17163 16670 17197
rect 16704 17163 16751 17197
rect 16785 17163 16831 17197
rect 16865 17163 16911 17197
rect 16945 17163 16991 17197
rect 17025 17163 17071 17197
rect 17105 17163 17151 17197
rect 17185 17163 17231 17197
rect 17265 17163 17311 17197
rect 17345 17163 17391 17197
rect 17425 17163 17471 17197
rect 17505 17163 17551 17197
rect 17585 17163 17631 17197
rect 17665 17163 17711 17197
rect 17745 17163 17791 17197
rect 17825 17163 17871 17197
rect 17905 17163 17951 17197
rect 17985 17163 18031 17197
rect 18065 17163 18111 17197
rect 18145 17163 18191 17197
rect 18225 17163 18271 17197
rect 18305 17163 18351 17197
rect 18385 17163 18431 17197
rect 18465 17163 18511 17197
rect 18545 17163 18591 17197
rect 18625 17163 18671 17197
rect 18705 17163 18751 17197
rect 18785 17163 18831 17197
rect 18865 17163 18911 17197
rect 18945 17163 18991 17197
rect 19025 17163 19071 17197
rect 19105 17163 19151 17197
rect 19185 17163 19231 17197
rect 19265 17163 19311 17197
rect 19345 17163 19391 17197
rect 19425 17163 19471 17197
rect 19505 17163 19551 17197
rect 19585 17163 19631 17197
rect 19665 17163 19711 17197
rect 19745 17163 19791 17197
rect 19825 17163 19871 17197
rect 19905 17163 19951 17197
rect 19985 17163 20031 17197
rect 20065 17163 20111 17197
rect 20145 17163 20191 17197
rect 20225 17163 20271 17197
rect 20305 17163 20351 17197
rect 20385 17163 20431 17197
rect 20465 17163 20511 17197
rect 20545 17163 20591 17197
rect 20625 17163 20671 17197
rect 20705 17163 20751 17197
rect 20785 17163 20831 17197
rect 20865 17163 20911 17197
rect 20945 17163 20991 17197
rect 21025 17163 21071 17197
rect 21105 17163 21151 17197
rect 21185 17163 21231 17197
rect 21265 17163 21311 17197
rect 21345 17163 21391 17197
rect 21425 17163 21471 17197
rect 21505 17163 21551 17197
rect 21585 17163 21631 17197
rect 21665 17163 21711 17197
rect 21745 17163 21791 17197
rect 21825 17163 21871 17197
rect 21905 17163 21951 17197
rect 21985 17163 22031 17197
rect 22065 17163 22111 17197
rect 22145 17163 22191 17197
rect 22225 17163 22271 17197
rect 22305 17163 22351 17197
rect 22385 17163 22431 17197
rect 22465 17163 22511 17197
rect 22545 17163 22591 17197
rect 22625 17163 22671 17197
rect 22705 17163 22751 17197
rect 22785 17163 22831 17197
rect 22865 17163 22911 17197
rect 22945 17163 22991 17197
rect 23025 17163 23071 17197
rect 23105 17163 23151 17197
rect 23185 17163 23231 17197
rect 23265 17163 23311 17197
rect 23345 17163 23391 17197
rect 23425 17163 23471 17197
rect 23505 17163 23551 17197
rect 23585 17163 23631 17197
rect 23665 17163 23711 17197
rect 23745 17163 23791 17197
rect 23825 17163 23871 17197
rect 23905 17163 23951 17197
rect 23985 17163 24031 17197
rect 24065 17163 24111 17197
rect 24145 17163 24191 17197
rect 24225 17163 24271 17197
rect 24305 17163 24351 17197
rect 24385 17163 24431 17197
rect 24465 17163 24511 17197
rect 24545 17163 24591 17197
rect 24625 17163 24671 17197
rect 24705 17163 24751 17197
rect 24785 17163 24831 17197
rect 24865 17163 24911 17197
rect 24945 17163 24991 17197
rect 25025 17163 25071 17197
rect 25105 17163 25151 17197
rect 25185 17163 25231 17197
rect 25265 17163 25311 17197
rect 25345 17163 25391 17197
rect 25425 17163 25471 17197
rect 25505 17163 25551 17197
rect 25585 17163 25631 17197
rect 25665 17163 25711 17197
rect 25745 17163 25791 17197
rect 25825 17163 25871 17197
rect 25905 17163 25951 17197
rect 25985 17163 26031 17197
rect 26065 17163 26111 17197
rect 26145 17163 26191 17197
rect 26225 17163 26271 17197
rect 26305 17163 26351 17197
rect 26385 17163 26431 17197
rect 26465 17163 26511 17197
rect 26545 17163 26591 17197
rect 26625 17163 26671 17197
rect 26705 17163 26751 17197
rect 26785 17163 26831 17197
rect 26865 17163 26911 17197
rect 26945 17163 26991 17197
rect 27025 17163 27071 17197
rect 27105 17163 27151 17197
rect 27185 17163 27231 17197
rect 27265 17163 27311 17197
rect 27345 17163 27391 17197
rect 27425 17163 27471 17197
rect 27505 17163 27551 17197
rect 27585 17163 27631 17197
rect 27665 17163 27711 17197
rect 27745 17163 27791 17197
rect 27825 17163 27871 17197
rect 27905 17163 27951 17197
rect 27985 17163 28031 17197
rect 28065 17163 28111 17197
rect 28145 17163 28191 17197
rect 28225 17163 28271 17197
rect 28305 17163 28351 17197
rect 28385 17163 28431 17197
rect 28465 17163 28511 17197
rect 28545 17163 28591 17197
rect 28625 17163 28671 17197
rect 28705 17163 28751 17197
rect 28785 17163 28831 17197
rect 28865 17163 28911 17197
rect 28945 17163 28991 17197
rect 29025 17163 29071 17197
rect 29105 17163 29151 17197
rect 29185 17163 29231 17197
rect 29265 17163 29311 17197
rect 29345 17163 29391 17197
rect 29425 17163 29471 17197
rect 29505 17163 29551 17197
rect 29585 17163 29631 17197
rect 29665 17163 29711 17197
rect 29745 17163 29791 17197
rect 29825 17163 29871 17197
rect 29905 17163 29951 17197
rect 29985 17163 30031 17197
rect 30065 17163 30111 17197
rect 30145 17163 30191 17197
rect 30225 17163 30271 17197
rect 30305 17163 30351 17197
rect 30385 17163 30431 17197
rect 30465 17163 30511 17197
rect 30545 17163 30591 17197
rect 30625 17163 30671 17197
rect 30705 17163 30751 17197
rect 30785 17163 30831 17197
rect 30865 17163 30911 17197
rect 30945 17163 30991 17197
rect 31025 17163 31071 17197
rect 31105 17163 31151 17197
rect 31185 17163 31231 17197
rect 31265 17163 31311 17197
rect 31345 17163 31391 17197
rect 31425 17163 31471 17197
rect 31505 17163 31551 17197
rect 31585 17163 31631 17197
rect 31665 17163 31711 17197
rect 31745 17163 31791 17197
rect 31825 17163 31871 17197
rect 31905 17163 31951 17197
rect 31985 17163 32031 17197
rect 32065 17163 32111 17197
rect 32145 17163 32191 17197
rect 32225 17163 32271 17197
rect 32305 17163 32351 17197
rect 32385 17163 32431 17197
rect 32465 17163 32511 17197
rect 32545 17163 32591 17197
rect 32625 17163 32671 17197
rect 32705 17163 32751 17197
rect 32785 17163 32831 17197
rect 32865 17163 32911 17197
rect 32945 17163 32991 17197
rect 33025 17163 33071 17197
rect 33105 17163 33151 17197
rect 33185 17163 33231 17197
rect 33265 17163 33311 17197
rect 33345 17163 33391 17197
rect 33425 17163 33471 17197
rect 33505 17163 33551 17197
rect 33585 17163 33631 17197
rect 33665 17163 33711 17197
rect 33745 17163 33791 17197
rect 33825 17163 33871 17197
rect 33905 17163 33951 17197
rect 33985 17163 34031 17197
rect 34065 17163 34111 17197
rect 34145 17163 34191 17197
rect 34225 17163 34271 17197
rect 34305 17163 34351 17197
rect 34385 17163 34431 17197
rect 34465 17163 34511 17197
rect 34545 17163 34591 17197
rect 34625 17163 34671 17197
rect 34705 17163 34751 17197
rect 34785 17163 34831 17197
rect 34865 17163 34911 17197
rect 34945 17163 34991 17197
rect 35025 17163 35071 17197
rect 35105 17163 35151 17197
rect 35185 17163 35231 17197
rect 35265 17163 35311 17197
rect 35345 17163 35391 17197
rect 35425 17163 35471 17197
rect 35505 17163 35551 17197
rect 35585 17163 35631 17197
rect 35665 17163 35711 17197
rect 35745 17163 35791 17197
rect 35825 17163 35871 17197
rect 35905 17163 35951 17197
rect 35985 17163 36031 17197
rect 36065 17163 36111 17197
rect 36145 17163 36191 17197
rect 36225 17163 36271 17197
rect 36305 17163 36351 17197
rect 36385 17163 36431 17197
rect 36465 17163 36511 17197
rect 36545 17163 36591 17197
rect 36625 17163 36671 17197
rect 36705 17163 36751 17197
rect 36785 17163 36831 17197
rect 36865 17163 36911 17197
rect 36945 17163 36991 17197
rect 37025 17163 37071 17197
rect 37105 17163 37151 17197
rect 37185 17163 37231 17197
rect 37265 17163 37311 17197
rect 37345 17163 37391 17197
rect 37425 17163 37471 17197
rect 37505 17163 37551 17197
rect 37585 17163 37631 17197
rect 37665 17163 37711 17197
rect 37745 17163 37791 17197
rect 37825 17163 37871 17197
rect 37905 17163 37951 17197
rect 37985 17163 38031 17197
rect 38065 17163 38111 17197
rect 38145 17163 38191 17197
rect 38225 17163 38271 17197
rect 38305 17163 38351 17197
rect 3744 17140 38351 17163
rect -37898 9338 -3290 9361
rect -37898 9304 -37852 9338
rect -37818 9304 -37772 9338
rect -37738 9304 -37692 9338
rect -37658 9304 -37612 9338
rect -37578 9304 -37532 9338
rect -37498 9304 -37452 9338
rect -37418 9304 -37372 9338
rect -37338 9304 -37292 9338
rect -37258 9304 -37212 9338
rect -37178 9304 -37132 9338
rect -37098 9304 -37052 9338
rect -37018 9304 -36972 9338
rect -36938 9304 -36892 9338
rect -36858 9304 -36812 9338
rect -36778 9304 -36732 9338
rect -36698 9304 -36652 9338
rect -36618 9304 -36572 9338
rect -36538 9304 -36492 9338
rect -36458 9304 -36412 9338
rect -36378 9304 -36332 9338
rect -36298 9304 -36252 9338
rect -36218 9304 -36172 9338
rect -36138 9304 -36092 9338
rect -36058 9304 -36012 9338
rect -35978 9304 -35932 9338
rect -35898 9304 -35852 9338
rect -35818 9304 -35772 9338
rect -35738 9304 -35692 9338
rect -35658 9304 -35612 9338
rect -35578 9304 -35532 9338
rect -35498 9304 -35452 9338
rect -35418 9304 -35372 9338
rect -35338 9304 -35292 9338
rect -35258 9304 -35212 9338
rect -35178 9304 -35132 9338
rect -35098 9304 -35052 9338
rect -35018 9304 -34972 9338
rect -34938 9304 -34892 9338
rect -34858 9304 -34812 9338
rect -34778 9304 -34732 9338
rect -34698 9304 -34652 9338
rect -34618 9304 -34572 9338
rect -34538 9304 -34492 9338
rect -34458 9304 -34412 9338
rect -34378 9304 -34332 9338
rect -34298 9304 -34252 9338
rect -34218 9304 -34172 9338
rect -34138 9304 -34092 9338
rect -34058 9304 -34012 9338
rect -33978 9304 -33932 9338
rect -33898 9304 -33852 9338
rect -33818 9304 -33772 9338
rect -33738 9304 -33692 9338
rect -33658 9304 -33612 9338
rect -33578 9304 -33532 9338
rect -33498 9304 -33452 9338
rect -33418 9304 -33372 9338
rect -33338 9304 -33292 9338
rect -33258 9304 -33212 9338
rect -33178 9304 -33132 9338
rect -33098 9304 -33052 9338
rect -33018 9304 -32972 9338
rect -32938 9304 -32892 9338
rect -32858 9304 -32812 9338
rect -32778 9304 -32732 9338
rect -32698 9304 -32652 9338
rect -32618 9304 -32572 9338
rect -32538 9304 -32492 9338
rect -32458 9304 -32412 9338
rect -32378 9304 -32332 9338
rect -32298 9304 -32252 9338
rect -32218 9304 -32172 9338
rect -32138 9304 -32092 9338
rect -32058 9304 -32012 9338
rect -31978 9304 -31932 9338
rect -31898 9304 -31852 9338
rect -31818 9304 -31772 9338
rect -31738 9304 -31692 9338
rect -31658 9304 -31612 9338
rect -31578 9304 -31532 9338
rect -31498 9304 -31452 9338
rect -31418 9304 -31372 9338
rect -31338 9304 -31292 9338
rect -31258 9304 -31212 9338
rect -31178 9304 -31132 9338
rect -31098 9304 -31052 9338
rect -31018 9304 -30972 9338
rect -30938 9304 -30892 9338
rect -30858 9304 -30812 9338
rect -30778 9304 -30732 9338
rect -30698 9304 -30652 9338
rect -30618 9304 -30572 9338
rect -30538 9304 -30492 9338
rect -30458 9304 -30412 9338
rect -30378 9304 -30332 9338
rect -30298 9304 -30252 9338
rect -30218 9304 -30172 9338
rect -30138 9304 -30092 9338
rect -30058 9304 -30012 9338
rect -29978 9304 -29932 9338
rect -29898 9304 -29852 9338
rect -29818 9304 -29772 9338
rect -29738 9304 -29692 9338
rect -29658 9304 -29612 9338
rect -29578 9304 -29532 9338
rect -29498 9304 -29452 9338
rect -29418 9304 -29372 9338
rect -29338 9304 -29292 9338
rect -29258 9304 -29212 9338
rect -29178 9304 -29132 9338
rect -29098 9304 -29052 9338
rect -29018 9304 -28972 9338
rect -28938 9304 -28892 9338
rect -28858 9304 -28812 9338
rect -28778 9304 -28732 9338
rect -28698 9304 -28652 9338
rect -28618 9304 -28572 9338
rect -28538 9304 -28492 9338
rect -28458 9304 -28412 9338
rect -28378 9304 -28332 9338
rect -28298 9304 -28252 9338
rect -28218 9304 -28172 9338
rect -28138 9304 -28092 9338
rect -28058 9304 -28012 9338
rect -27978 9304 -27932 9338
rect -27898 9304 -27852 9338
rect -27818 9304 -27772 9338
rect -27738 9304 -27692 9338
rect -27658 9304 -27612 9338
rect -27578 9304 -27532 9338
rect -27498 9304 -27452 9338
rect -27418 9304 -27372 9338
rect -27338 9304 -27292 9338
rect -27258 9304 -27212 9338
rect -27178 9304 -27132 9338
rect -27098 9304 -27052 9338
rect -27018 9304 -26972 9338
rect -26938 9304 -26892 9338
rect -26858 9304 -26812 9338
rect -26778 9304 -26732 9338
rect -26698 9304 -26652 9338
rect -26618 9304 -26572 9338
rect -26538 9304 -26492 9338
rect -26458 9304 -26412 9338
rect -26378 9304 -26332 9338
rect -26298 9304 -26252 9338
rect -26218 9304 -26172 9338
rect -26138 9304 -26092 9338
rect -26058 9304 -26012 9338
rect -25978 9304 -25932 9338
rect -25898 9304 -25852 9338
rect -25818 9304 -25772 9338
rect -25738 9304 -25692 9338
rect -25658 9304 -25612 9338
rect -25578 9304 -25532 9338
rect -25498 9304 -25452 9338
rect -25418 9304 -25372 9338
rect -25338 9304 -25292 9338
rect -25258 9304 -25212 9338
rect -25178 9304 -25132 9338
rect -25098 9304 -25052 9338
rect -25018 9304 -24972 9338
rect -24938 9304 -24891 9338
rect -24857 9304 -24811 9338
rect -24777 9304 -24731 9338
rect -24697 9304 -24651 9338
rect -24617 9304 -24571 9338
rect -24537 9304 -24491 9338
rect -24457 9304 -24411 9338
rect -24377 9304 -24331 9338
rect -24297 9304 -24251 9338
rect -24217 9304 -24171 9338
rect -24137 9304 -24091 9338
rect -24057 9304 -24011 9338
rect -23977 9304 -23931 9338
rect -23897 9304 -23851 9338
rect -23817 9304 -23771 9338
rect -23737 9304 -23691 9338
rect -23657 9304 -23611 9338
rect -23577 9304 -23531 9338
rect -23497 9304 -23451 9338
rect -23417 9304 -23371 9338
rect -23337 9304 -23291 9338
rect -23257 9304 -23211 9338
rect -23177 9304 -23131 9338
rect -23097 9304 -23051 9338
rect -23017 9304 -22971 9338
rect -22937 9304 -22891 9338
rect -22857 9304 -22811 9338
rect -22777 9304 -22731 9338
rect -22697 9304 -22651 9338
rect -22617 9304 -22571 9338
rect -22537 9304 -22491 9338
rect -22457 9304 -22411 9338
rect -22377 9304 -22331 9338
rect -22297 9304 -22251 9338
rect -22217 9304 -22171 9338
rect -22137 9304 -22091 9338
rect -22057 9304 -22011 9338
rect -21977 9304 -21931 9338
rect -21897 9304 -21851 9338
rect -21817 9304 -21771 9338
rect -21737 9304 -21691 9338
rect -21657 9304 -21611 9338
rect -21577 9304 -21531 9338
rect -21497 9304 -21451 9338
rect -21417 9304 -21371 9338
rect -21337 9304 -21291 9338
rect -21257 9304 -21211 9338
rect -21177 9304 -21131 9338
rect -21097 9304 -21051 9338
rect -21017 9304 -20971 9338
rect -20937 9304 -20891 9338
rect -20857 9304 -20811 9338
rect -20777 9304 -20731 9338
rect -20697 9304 -20651 9338
rect -20617 9304 -20571 9338
rect -20537 9304 -20491 9338
rect -20457 9304 -20411 9338
rect -20377 9304 -20331 9338
rect -20297 9304 -20251 9338
rect -20217 9304 -20171 9338
rect -20137 9304 -20091 9338
rect -20057 9304 -20011 9338
rect -19977 9304 -19931 9338
rect -19897 9304 -19851 9338
rect -19817 9304 -19771 9338
rect -19737 9304 -19691 9338
rect -19657 9304 -19611 9338
rect -19577 9304 -19531 9338
rect -19497 9304 -19451 9338
rect -19417 9304 -19371 9338
rect -19337 9304 -19291 9338
rect -19257 9304 -19211 9338
rect -19177 9304 -19131 9338
rect -19097 9304 -19051 9338
rect -19017 9304 -18971 9338
rect -18937 9304 -18891 9338
rect -18857 9304 -18811 9338
rect -18777 9304 -18731 9338
rect -18697 9304 -18651 9338
rect -18617 9304 -18571 9338
rect -18537 9304 -18491 9338
rect -18457 9304 -18411 9338
rect -18377 9304 -18331 9338
rect -18297 9304 -18251 9338
rect -18217 9304 -18171 9338
rect -18137 9304 -18091 9338
rect -18057 9304 -18011 9338
rect -17977 9304 -17931 9338
rect -17897 9304 -17851 9338
rect -17817 9304 -17771 9338
rect -17737 9304 -17691 9338
rect -17657 9304 -17611 9338
rect -17577 9304 -17531 9338
rect -17497 9304 -17451 9338
rect -17417 9304 -17371 9338
rect -17337 9304 -17291 9338
rect -17257 9304 -17211 9338
rect -17177 9304 -17131 9338
rect -17097 9304 -17051 9338
rect -17017 9304 -16971 9338
rect -16937 9304 -16891 9338
rect -16857 9304 -16811 9338
rect -16777 9304 -16731 9338
rect -16697 9304 -16651 9338
rect -16617 9304 -16571 9338
rect -16537 9304 -16491 9338
rect -16457 9304 -16411 9338
rect -16377 9304 -16331 9338
rect -16297 9304 -16251 9338
rect -16217 9304 -16171 9338
rect -16137 9304 -16091 9338
rect -16057 9304 -16011 9338
rect -15977 9304 -15931 9338
rect -15897 9304 -15851 9338
rect -15817 9304 -15771 9338
rect -15737 9304 -15691 9338
rect -15657 9304 -15611 9338
rect -15577 9304 -15531 9338
rect -15497 9304 -15451 9338
rect -15417 9304 -15371 9338
rect -15337 9304 -15291 9338
rect -15257 9304 -15211 9338
rect -15177 9304 -15131 9338
rect -15097 9304 -15051 9338
rect -15017 9304 -14971 9338
rect -14937 9304 -14891 9338
rect -14857 9304 -14811 9338
rect -14777 9304 -14731 9338
rect -14697 9304 -14651 9338
rect -14617 9304 -14571 9338
rect -14537 9304 -14491 9338
rect -14457 9304 -14411 9338
rect -14377 9304 -14331 9338
rect -14297 9304 -14251 9338
rect -14217 9304 -14171 9338
rect -14137 9304 -14091 9338
rect -14057 9304 -14011 9338
rect -13977 9304 -13931 9338
rect -13897 9304 -13851 9338
rect -13817 9304 -13771 9338
rect -13737 9304 -13691 9338
rect -13657 9304 -13611 9338
rect -13577 9304 -13531 9338
rect -13497 9304 -13451 9338
rect -13417 9304 -13371 9338
rect -13337 9304 -13291 9338
rect -13257 9304 -13211 9338
rect -13177 9304 -13131 9338
rect -13097 9304 -13051 9338
rect -13017 9304 -12971 9338
rect -12937 9304 -12891 9338
rect -12857 9304 -12811 9338
rect -12777 9304 -12731 9338
rect -12697 9304 -12651 9338
rect -12617 9304 -12571 9338
rect -12537 9304 -12491 9338
rect -12457 9304 -12411 9338
rect -12377 9304 -12331 9338
rect -12297 9304 -12251 9338
rect -12217 9304 -12171 9338
rect -12137 9304 -12091 9338
rect -12057 9304 -12011 9338
rect -11977 9304 -11930 9338
rect -11896 9304 -11850 9338
rect -11816 9304 -11770 9338
rect -11736 9304 -11690 9338
rect -11656 9304 -11610 9338
rect -11576 9304 -11530 9338
rect -11496 9304 -11450 9338
rect -11416 9304 -11370 9338
rect -11336 9304 -11290 9338
rect -11256 9304 -11210 9338
rect -11176 9304 -11130 9338
rect -11096 9304 -11050 9338
rect -11016 9304 -10970 9338
rect -10936 9304 -10890 9338
rect -10856 9304 -10810 9338
rect -10776 9304 -10730 9338
rect -10696 9304 -10650 9338
rect -10616 9304 -10570 9338
rect -10536 9304 -10490 9338
rect -10456 9304 -10410 9338
rect -10376 9304 -10330 9338
rect -10296 9304 -10250 9338
rect -10216 9304 -10170 9338
rect -10136 9304 -10090 9338
rect -10056 9304 -10010 9338
rect -9976 9304 -9930 9338
rect -9896 9304 -9850 9338
rect -9816 9304 -9770 9338
rect -9736 9304 -9690 9338
rect -9656 9304 -9610 9338
rect -9576 9304 -9530 9338
rect -9496 9304 -9450 9338
rect -9416 9304 -9370 9338
rect -9336 9304 -9290 9338
rect -9256 9304 -9210 9338
rect -9176 9304 -9130 9338
rect -9096 9304 -9050 9338
rect -9016 9304 -8970 9338
rect -8936 9304 -8890 9338
rect -8856 9304 -8810 9338
rect -8776 9304 -8730 9338
rect -8696 9304 -8650 9338
rect -8616 9304 -8570 9338
rect -8536 9304 -8490 9338
rect -8456 9304 -8410 9338
rect -8376 9304 -8330 9338
rect -8296 9304 -8250 9338
rect -8216 9304 -8170 9338
rect -8136 9304 -8090 9338
rect -8056 9304 -8010 9338
rect -7976 9304 -7930 9338
rect -7896 9304 -7850 9338
rect -7816 9304 -7770 9338
rect -7736 9304 -7690 9338
rect -7656 9304 -7610 9338
rect -7576 9304 -7530 9338
rect -7496 9304 -7450 9338
rect -7416 9304 -7370 9338
rect -7336 9304 -7290 9338
rect -7256 9304 -7210 9338
rect -7176 9304 -7130 9338
rect -7096 9304 -7050 9338
rect -7016 9304 -6970 9338
rect -6936 9304 -6890 9338
rect -6856 9304 -6810 9338
rect -6776 9304 -6730 9338
rect -6696 9304 -6650 9338
rect -6616 9304 -6570 9338
rect -6536 9304 -6490 9338
rect -6456 9304 -6410 9338
rect -6376 9304 -6330 9338
rect -6296 9304 -6250 9338
rect -6216 9304 -6170 9338
rect -6136 9304 -6090 9338
rect -6056 9304 -6010 9338
rect -5976 9304 -5930 9338
rect -5896 9304 -5850 9338
rect -5816 9304 -5770 9338
rect -5736 9304 -5690 9338
rect -5656 9304 -5610 9338
rect -5576 9304 -5530 9338
rect -5496 9304 -5450 9338
rect -5416 9304 -5370 9338
rect -5336 9304 -5290 9338
rect -5256 9304 -5210 9338
rect -5176 9304 -5130 9338
rect -5096 9304 -5050 9338
rect -5016 9304 -4970 9338
rect -4936 9304 -4890 9338
rect -4856 9304 -4810 9338
rect -4776 9304 -4730 9338
rect -4696 9304 -4650 9338
rect -4616 9304 -4570 9338
rect -4536 9304 -4490 9338
rect -4456 9304 -4410 9338
rect -4376 9304 -4330 9338
rect -4296 9304 -4250 9338
rect -4216 9304 -4170 9338
rect -4136 9304 -4090 9338
rect -4056 9304 -4010 9338
rect -3976 9304 -3930 9338
rect -3896 9304 -3850 9338
rect -3816 9304 -3770 9338
rect -3736 9304 -3690 9338
rect -3656 9304 -3610 9338
rect -3576 9304 -3530 9338
rect -3496 9304 -3450 9338
rect -3416 9304 -3370 9338
rect -3336 9304 -3290 9338
rect -37898 9281 -3290 9304
rect -1942 9338 2397 9361
rect -1942 9304 -1929 9338
rect -1895 9304 -1849 9338
rect -1815 9304 -1769 9338
rect -1735 9304 -1689 9338
rect -1655 9304 -1609 9338
rect -1575 9304 -1529 9338
rect -1495 9304 -1449 9338
rect -1415 9304 -1369 9338
rect -1335 9304 -1289 9338
rect -1255 9304 -1209 9338
rect -1175 9304 -1129 9338
rect -1095 9304 -1049 9338
rect -1015 9304 -969 9338
rect -935 9304 -889 9338
rect -855 9304 -809 9338
rect -775 9304 -729 9338
rect -695 9304 -649 9338
rect -615 9304 -569 9338
rect -535 9304 -489 9338
rect -455 9304 -409 9338
rect -375 9304 -329 9338
rect -295 9304 -249 9338
rect -215 9304 -169 9338
rect -135 9304 -89 9338
rect -55 9304 -9 9338
rect 25 9304 71 9338
rect 105 9304 151 9338
rect 185 9304 231 9338
rect 265 9304 311 9338
rect 345 9304 391 9338
rect 425 9304 471 9338
rect 505 9304 551 9338
rect 585 9304 631 9338
rect 665 9304 711 9338
rect 745 9304 791 9338
rect 825 9304 871 9338
rect 905 9304 951 9338
rect 985 9304 1031 9338
rect 1065 9304 1111 9338
rect 1145 9304 1191 9338
rect 1225 9304 1271 9338
rect 1305 9304 1351 9338
rect 1385 9304 1431 9338
rect 1465 9304 1511 9338
rect 1545 9304 1591 9338
rect 1625 9304 1671 9338
rect 1705 9304 1751 9338
rect 1785 9304 1831 9338
rect 1865 9304 1911 9338
rect 1945 9304 1991 9338
rect 2025 9304 2071 9338
rect 2105 9304 2151 9338
rect 2185 9304 2231 9338
rect 2265 9304 2311 9338
rect 2345 9304 2397 9338
rect -1942 9281 2397 9304
rect 3744 9338 38351 9361
rect 3744 9304 3790 9338
rect 3824 9304 3870 9338
rect 3904 9304 3950 9338
rect 3984 9304 4030 9338
rect 4064 9304 4110 9338
rect 4144 9304 4190 9338
rect 4224 9304 4270 9338
rect 4304 9304 4350 9338
rect 4384 9304 4430 9338
rect 4464 9304 4510 9338
rect 4544 9304 4590 9338
rect 4624 9304 4670 9338
rect 4704 9304 4750 9338
rect 4784 9304 4830 9338
rect 4864 9304 4910 9338
rect 4944 9304 4990 9338
rect 5024 9304 5070 9338
rect 5104 9304 5150 9338
rect 5184 9304 5230 9338
rect 5264 9304 5310 9338
rect 5344 9304 5390 9338
rect 5424 9304 5470 9338
rect 5504 9304 5550 9338
rect 5584 9304 5630 9338
rect 5664 9304 5710 9338
rect 5744 9304 5790 9338
rect 5824 9304 5870 9338
rect 5904 9304 5950 9338
rect 5984 9304 6030 9338
rect 6064 9304 6110 9338
rect 6144 9304 6190 9338
rect 6224 9304 6270 9338
rect 6304 9304 6350 9338
rect 6384 9304 6430 9338
rect 6464 9304 6510 9338
rect 6544 9304 6590 9338
rect 6624 9304 6670 9338
rect 6704 9304 6750 9338
rect 6784 9304 6830 9338
rect 6864 9304 6910 9338
rect 6944 9304 6990 9338
rect 7024 9304 7070 9338
rect 7104 9304 7150 9338
rect 7184 9304 7230 9338
rect 7264 9304 7310 9338
rect 7344 9304 7390 9338
rect 7424 9304 7470 9338
rect 7504 9304 7550 9338
rect 7584 9304 7630 9338
rect 7664 9304 7710 9338
rect 7744 9304 7790 9338
rect 7824 9304 7870 9338
rect 7904 9304 7950 9338
rect 7984 9304 8030 9338
rect 8064 9304 8110 9338
rect 8144 9304 8190 9338
rect 8224 9304 8270 9338
rect 8304 9304 8350 9338
rect 8384 9304 8430 9338
rect 8464 9304 8510 9338
rect 8544 9304 8590 9338
rect 8624 9304 8670 9338
rect 8704 9304 8750 9338
rect 8784 9304 8830 9338
rect 8864 9304 8910 9338
rect 8944 9304 8990 9338
rect 9024 9304 9070 9338
rect 9104 9304 9150 9338
rect 9184 9304 9230 9338
rect 9264 9304 9310 9338
rect 9344 9304 9390 9338
rect 9424 9304 9470 9338
rect 9504 9304 9550 9338
rect 9584 9304 9630 9338
rect 9664 9304 9710 9338
rect 9744 9304 9790 9338
rect 9824 9304 9870 9338
rect 9904 9304 9950 9338
rect 9984 9304 10030 9338
rect 10064 9304 10110 9338
rect 10144 9304 10190 9338
rect 10224 9304 10270 9338
rect 10304 9304 10350 9338
rect 10384 9304 10430 9338
rect 10464 9304 10510 9338
rect 10544 9304 10590 9338
rect 10624 9304 10670 9338
rect 10704 9304 10750 9338
rect 10784 9304 10830 9338
rect 10864 9304 10910 9338
rect 10944 9304 10990 9338
rect 11024 9304 11070 9338
rect 11104 9304 11150 9338
rect 11184 9304 11230 9338
rect 11264 9304 11310 9338
rect 11344 9304 11390 9338
rect 11424 9304 11470 9338
rect 11504 9304 11550 9338
rect 11584 9304 11630 9338
rect 11664 9304 11710 9338
rect 11744 9304 11790 9338
rect 11824 9304 11870 9338
rect 11904 9304 11950 9338
rect 11984 9304 12030 9338
rect 12064 9304 12110 9338
rect 12144 9304 12190 9338
rect 12224 9304 12270 9338
rect 12304 9304 12350 9338
rect 12384 9304 12430 9338
rect 12464 9304 12510 9338
rect 12544 9304 12590 9338
rect 12624 9304 12670 9338
rect 12704 9304 12750 9338
rect 12784 9304 12830 9338
rect 12864 9304 12910 9338
rect 12944 9304 12990 9338
rect 13024 9304 13070 9338
rect 13104 9304 13150 9338
rect 13184 9304 13230 9338
rect 13264 9304 13310 9338
rect 13344 9304 13390 9338
rect 13424 9304 13470 9338
rect 13504 9304 13550 9338
rect 13584 9304 13630 9338
rect 13664 9304 13710 9338
rect 13744 9304 13790 9338
rect 13824 9304 13870 9338
rect 13904 9304 13950 9338
rect 13984 9304 14030 9338
rect 14064 9304 14110 9338
rect 14144 9304 14190 9338
rect 14224 9304 14270 9338
rect 14304 9304 14350 9338
rect 14384 9304 14430 9338
rect 14464 9304 14510 9338
rect 14544 9304 14590 9338
rect 14624 9304 14670 9338
rect 14704 9304 14750 9338
rect 14784 9304 14830 9338
rect 14864 9304 14910 9338
rect 14944 9304 14990 9338
rect 15024 9304 15070 9338
rect 15104 9304 15150 9338
rect 15184 9304 15230 9338
rect 15264 9304 15310 9338
rect 15344 9304 15390 9338
rect 15424 9304 15470 9338
rect 15504 9304 15550 9338
rect 15584 9304 15630 9338
rect 15664 9304 15710 9338
rect 15744 9304 15790 9338
rect 15824 9304 15870 9338
rect 15904 9304 15950 9338
rect 15984 9304 16030 9338
rect 16064 9304 16110 9338
rect 16144 9304 16190 9338
rect 16224 9304 16270 9338
rect 16304 9304 16350 9338
rect 16384 9304 16430 9338
rect 16464 9304 16510 9338
rect 16544 9304 16590 9338
rect 16624 9304 16670 9338
rect 16704 9304 16751 9338
rect 16785 9304 16831 9338
rect 16865 9304 16911 9338
rect 16945 9304 16991 9338
rect 17025 9304 17071 9338
rect 17105 9304 17151 9338
rect 17185 9304 17231 9338
rect 17265 9304 17311 9338
rect 17345 9304 17391 9338
rect 17425 9304 17471 9338
rect 17505 9304 17551 9338
rect 17585 9304 17631 9338
rect 17665 9304 17711 9338
rect 17745 9304 17791 9338
rect 17825 9304 17871 9338
rect 17905 9304 17951 9338
rect 17985 9304 18031 9338
rect 18065 9304 18111 9338
rect 18145 9304 18191 9338
rect 18225 9304 18271 9338
rect 18305 9304 18351 9338
rect 18385 9304 18431 9338
rect 18465 9304 18511 9338
rect 18545 9304 18591 9338
rect 18625 9304 18671 9338
rect 18705 9304 18751 9338
rect 18785 9304 18831 9338
rect 18865 9304 18911 9338
rect 18945 9304 18991 9338
rect 19025 9304 19071 9338
rect 19105 9304 19151 9338
rect 19185 9304 19231 9338
rect 19265 9304 19311 9338
rect 19345 9304 19391 9338
rect 19425 9304 19471 9338
rect 19505 9304 19551 9338
rect 19585 9304 19631 9338
rect 19665 9304 19711 9338
rect 19745 9304 19791 9338
rect 19825 9304 19871 9338
rect 19905 9304 19951 9338
rect 19985 9304 20031 9338
rect 20065 9304 20111 9338
rect 20145 9304 20191 9338
rect 20225 9304 20271 9338
rect 20305 9304 20351 9338
rect 20385 9304 20431 9338
rect 20465 9304 20511 9338
rect 20545 9304 20591 9338
rect 20625 9304 20671 9338
rect 20705 9304 20751 9338
rect 20785 9304 20831 9338
rect 20865 9304 20911 9338
rect 20945 9304 20991 9338
rect 21025 9304 21071 9338
rect 21105 9304 21151 9338
rect 21185 9304 21231 9338
rect 21265 9304 21311 9338
rect 21345 9304 21391 9338
rect 21425 9304 21471 9338
rect 21505 9304 21551 9338
rect 21585 9304 21631 9338
rect 21665 9304 21711 9338
rect 21745 9304 21791 9338
rect 21825 9304 21871 9338
rect 21905 9304 21951 9338
rect 21985 9304 22031 9338
rect 22065 9304 22111 9338
rect 22145 9304 22191 9338
rect 22225 9304 22271 9338
rect 22305 9304 22351 9338
rect 22385 9304 22431 9338
rect 22465 9304 22511 9338
rect 22545 9304 22591 9338
rect 22625 9304 22671 9338
rect 22705 9304 22751 9338
rect 22785 9304 22831 9338
rect 22865 9304 22911 9338
rect 22945 9304 22991 9338
rect 23025 9304 23071 9338
rect 23105 9304 23151 9338
rect 23185 9304 23231 9338
rect 23265 9304 23311 9338
rect 23345 9304 23391 9338
rect 23425 9304 23471 9338
rect 23505 9304 23551 9338
rect 23585 9304 23631 9338
rect 23665 9304 23711 9338
rect 23745 9304 23791 9338
rect 23825 9304 23871 9338
rect 23905 9304 23951 9338
rect 23985 9304 24031 9338
rect 24065 9304 24111 9338
rect 24145 9304 24191 9338
rect 24225 9304 24271 9338
rect 24305 9304 24351 9338
rect 24385 9304 24431 9338
rect 24465 9304 24511 9338
rect 24545 9304 24591 9338
rect 24625 9304 24671 9338
rect 24705 9304 24751 9338
rect 24785 9304 24831 9338
rect 24865 9304 24911 9338
rect 24945 9304 24991 9338
rect 25025 9304 25071 9338
rect 25105 9304 25151 9338
rect 25185 9304 25231 9338
rect 25265 9304 25311 9338
rect 25345 9304 25391 9338
rect 25425 9304 25471 9338
rect 25505 9304 25551 9338
rect 25585 9304 25631 9338
rect 25665 9304 25711 9338
rect 25745 9304 25791 9338
rect 25825 9304 25871 9338
rect 25905 9304 25951 9338
rect 25985 9304 26031 9338
rect 26065 9304 26111 9338
rect 26145 9304 26191 9338
rect 26225 9304 26271 9338
rect 26305 9304 26351 9338
rect 26385 9304 26431 9338
rect 26465 9304 26511 9338
rect 26545 9304 26591 9338
rect 26625 9304 26671 9338
rect 26705 9304 26751 9338
rect 26785 9304 26831 9338
rect 26865 9304 26911 9338
rect 26945 9304 26991 9338
rect 27025 9304 27071 9338
rect 27105 9304 27151 9338
rect 27185 9304 27231 9338
rect 27265 9304 27311 9338
rect 27345 9304 27391 9338
rect 27425 9304 27471 9338
rect 27505 9304 27551 9338
rect 27585 9304 27631 9338
rect 27665 9304 27711 9338
rect 27745 9304 27791 9338
rect 27825 9304 27871 9338
rect 27905 9304 27951 9338
rect 27985 9304 28031 9338
rect 28065 9304 28111 9338
rect 28145 9304 28191 9338
rect 28225 9304 28271 9338
rect 28305 9304 28351 9338
rect 28385 9304 28431 9338
rect 28465 9304 28511 9338
rect 28545 9304 28591 9338
rect 28625 9304 28671 9338
rect 28705 9304 28751 9338
rect 28785 9304 28831 9338
rect 28865 9304 28911 9338
rect 28945 9304 28991 9338
rect 29025 9304 29071 9338
rect 29105 9304 29151 9338
rect 29185 9304 29231 9338
rect 29265 9304 29311 9338
rect 29345 9304 29391 9338
rect 29425 9304 29471 9338
rect 29505 9304 29551 9338
rect 29585 9304 29631 9338
rect 29665 9304 29711 9338
rect 29745 9304 29791 9338
rect 29825 9304 29871 9338
rect 29905 9304 29951 9338
rect 29985 9304 30031 9338
rect 30065 9304 30111 9338
rect 30145 9304 30191 9338
rect 30225 9304 30271 9338
rect 30305 9304 30351 9338
rect 30385 9304 30431 9338
rect 30465 9304 30511 9338
rect 30545 9304 30591 9338
rect 30625 9304 30671 9338
rect 30705 9304 30751 9338
rect 30785 9304 30831 9338
rect 30865 9304 30911 9338
rect 30945 9304 30991 9338
rect 31025 9304 31071 9338
rect 31105 9304 31151 9338
rect 31185 9304 31231 9338
rect 31265 9304 31311 9338
rect 31345 9304 31391 9338
rect 31425 9304 31471 9338
rect 31505 9304 31551 9338
rect 31585 9304 31631 9338
rect 31665 9304 31711 9338
rect 31745 9304 31791 9338
rect 31825 9304 31871 9338
rect 31905 9304 31951 9338
rect 31985 9304 32031 9338
rect 32065 9304 32111 9338
rect 32145 9304 32191 9338
rect 32225 9304 32271 9338
rect 32305 9304 32351 9338
rect 32385 9304 32431 9338
rect 32465 9304 32511 9338
rect 32545 9304 32591 9338
rect 32625 9304 32671 9338
rect 32705 9304 32751 9338
rect 32785 9304 32831 9338
rect 32865 9304 32911 9338
rect 32945 9304 32991 9338
rect 33025 9304 33071 9338
rect 33105 9304 33151 9338
rect 33185 9304 33231 9338
rect 33265 9304 33311 9338
rect 33345 9304 33391 9338
rect 33425 9304 33471 9338
rect 33505 9304 33551 9338
rect 33585 9304 33631 9338
rect 33665 9304 33711 9338
rect 33745 9304 33791 9338
rect 33825 9304 33871 9338
rect 33905 9304 33951 9338
rect 33985 9304 34031 9338
rect 34065 9304 34111 9338
rect 34145 9304 34191 9338
rect 34225 9304 34271 9338
rect 34305 9304 34351 9338
rect 34385 9304 34431 9338
rect 34465 9304 34511 9338
rect 34545 9304 34591 9338
rect 34625 9304 34671 9338
rect 34705 9304 34751 9338
rect 34785 9304 34831 9338
rect 34865 9304 34911 9338
rect 34945 9304 34991 9338
rect 35025 9304 35071 9338
rect 35105 9304 35151 9338
rect 35185 9304 35231 9338
rect 35265 9304 35311 9338
rect 35345 9304 35391 9338
rect 35425 9304 35471 9338
rect 35505 9304 35551 9338
rect 35585 9304 35631 9338
rect 35665 9304 35711 9338
rect 35745 9304 35791 9338
rect 35825 9304 35871 9338
rect 35905 9304 35951 9338
rect 35985 9304 36031 9338
rect 36065 9304 36111 9338
rect 36145 9304 36191 9338
rect 36225 9304 36271 9338
rect 36305 9304 36351 9338
rect 36385 9304 36431 9338
rect 36465 9304 36511 9338
rect 36545 9304 36591 9338
rect 36625 9304 36671 9338
rect 36705 9304 36751 9338
rect 36785 9304 36831 9338
rect 36865 9304 36911 9338
rect 36945 9304 36991 9338
rect 37025 9304 37071 9338
rect 37105 9304 37151 9338
rect 37185 9304 37231 9338
rect 37265 9304 37311 9338
rect 37345 9304 37391 9338
rect 37425 9304 37471 9338
rect 37505 9304 37551 9338
rect 37585 9304 37631 9338
rect 37665 9304 37711 9338
rect 37745 9304 37791 9338
rect 37825 9304 37871 9338
rect 37905 9304 37951 9338
rect 37985 9304 38031 9338
rect 38065 9304 38111 9338
rect 38145 9304 38191 9338
rect 38225 9304 38271 9338
rect 38305 9304 38351 9338
rect 3744 9281 38351 9304
rect -3860 7826 -3600 8086
rect -2850 7970 -2784 9281
rect -317 9106 -283 9281
rect -1562 8709 -1289 8743
rect -2188 8132 -1988 8332
rect -2172 7865 -2012 8132
rect -1562 7865 -1528 8709
rect 2756 7970 2822 9281
rect 5230 9105 5264 9281
rect 4044 8727 4256 8761
rect 3393 8132 3593 8332
rect 3413 7865 3573 8132
rect 4044 7865 4078 8727
rect -3860 6588 -3600 6848
rect -3058 6383 -2978 6925
rect -288 6493 -28 6845
rect 1338 6493 1598 6845
rect 4288 6383 4368 6925
rect -37897 6360 35594 6383
rect -37897 6326 -37851 6360
rect -37817 6326 -37771 6360
rect -37737 6326 -37691 6360
rect -37657 6326 -37611 6360
rect -37577 6326 -37531 6360
rect -37497 6326 -37451 6360
rect -37417 6326 -37371 6360
rect -37337 6326 -37291 6360
rect -37257 6326 -37211 6360
rect -37177 6326 -37131 6360
rect -37097 6326 -37051 6360
rect -37017 6326 -36971 6360
rect -36937 6326 -36891 6360
rect -36857 6326 -36811 6360
rect -36777 6326 -36731 6360
rect -36697 6326 -36651 6360
rect -36617 6326 -36571 6360
rect -36537 6326 -36491 6360
rect -36457 6326 -36411 6360
rect -36377 6326 -36331 6360
rect -36297 6326 -36251 6360
rect -36217 6326 -36171 6360
rect -36137 6326 -36091 6360
rect -36057 6326 -36011 6360
rect -35977 6326 -35931 6360
rect -35897 6326 -35851 6360
rect -35817 6326 -35771 6360
rect -35737 6326 -35691 6360
rect -35657 6326 -35611 6360
rect -35577 6326 -35531 6360
rect -35497 6326 -35451 6360
rect -35417 6326 -35371 6360
rect -35337 6326 -35291 6360
rect -35257 6326 -35211 6360
rect -35177 6326 -35131 6360
rect -35097 6326 -35051 6360
rect -35017 6326 -34971 6360
rect -34937 6326 -34891 6360
rect -34857 6326 -34811 6360
rect -34777 6326 -34731 6360
rect -34697 6326 -34651 6360
rect -34617 6326 -34571 6360
rect -34537 6326 -34491 6360
rect -34457 6326 -34411 6360
rect -34377 6326 -34331 6360
rect -34297 6326 -34251 6360
rect -34217 6326 -34171 6360
rect -34137 6326 -34091 6360
rect -34057 6326 -34011 6360
rect -33977 6326 -33931 6360
rect -33897 6326 -33851 6360
rect -33817 6326 -33771 6360
rect -33737 6326 -33691 6360
rect -33657 6326 -33611 6360
rect -33577 6326 -33531 6360
rect -33497 6326 -33451 6360
rect -33417 6326 -33371 6360
rect -33337 6326 -33291 6360
rect -33257 6326 -33211 6360
rect -33177 6326 -33131 6360
rect -33097 6326 -33051 6360
rect -33017 6326 -32971 6360
rect -32937 6326 -32891 6360
rect -32857 6326 -32811 6360
rect -32777 6326 -32731 6360
rect -32697 6326 -32651 6360
rect -32617 6326 -32571 6360
rect -32537 6326 -32491 6360
rect -32457 6326 -32411 6360
rect -32377 6326 -32331 6360
rect -32297 6326 -32251 6360
rect -32217 6326 -32171 6360
rect -32137 6326 -32091 6360
rect -32057 6326 -32011 6360
rect -31977 6326 -31931 6360
rect -31897 6326 -31851 6360
rect -31817 6326 -31771 6360
rect -31737 6326 -31691 6360
rect -31657 6326 -31611 6360
rect -31577 6326 -31531 6360
rect -31497 6326 -31451 6360
rect -31417 6326 -31371 6360
rect -31337 6326 -31291 6360
rect -31257 6326 -31211 6360
rect -31177 6326 -31131 6360
rect -31097 6326 -31051 6360
rect -31017 6326 -30971 6360
rect -30937 6326 -30891 6360
rect -30857 6326 -30811 6360
rect -30777 6326 -30731 6360
rect -30697 6326 -30651 6360
rect -30617 6326 -30571 6360
rect -30537 6326 -30491 6360
rect -30457 6326 -30411 6360
rect -30377 6326 -30331 6360
rect -30297 6326 -30251 6360
rect -30217 6326 -30171 6360
rect -30137 6326 -30091 6360
rect -30057 6326 -30011 6360
rect -29977 6326 -29931 6360
rect -29897 6326 -29851 6360
rect -29817 6326 -29771 6360
rect -29737 6326 -29691 6360
rect -29657 6326 -29611 6360
rect -29577 6326 -29531 6360
rect -29497 6326 -29451 6360
rect -29417 6326 -29371 6360
rect -29337 6326 -29291 6360
rect -29257 6326 -29211 6360
rect -29177 6326 -29131 6360
rect -29097 6326 -29051 6360
rect -29017 6326 -28971 6360
rect -28937 6326 -28891 6360
rect -28857 6326 -28811 6360
rect -28777 6326 -28731 6360
rect -28697 6326 -28651 6360
rect -28617 6326 -28571 6360
rect -28537 6326 -28491 6360
rect -28457 6326 -28411 6360
rect -28377 6326 -28331 6360
rect -28297 6326 -28251 6360
rect -28217 6326 -28171 6360
rect -28137 6326 -28091 6360
rect -28057 6326 -28011 6360
rect -27977 6326 -27931 6360
rect -27897 6326 -27851 6360
rect -27817 6326 -27771 6360
rect -27737 6326 -27691 6360
rect -27657 6326 -27611 6360
rect -27577 6326 -27531 6360
rect -27497 6326 -27451 6360
rect -27417 6326 -27371 6360
rect -27337 6326 -27291 6360
rect -27257 6326 -27211 6360
rect -27177 6326 -27131 6360
rect -27097 6326 -27051 6360
rect -27017 6326 -26971 6360
rect -26937 6326 -26891 6360
rect -26857 6326 -26811 6360
rect -26777 6326 -26731 6360
rect -26697 6326 -26651 6360
rect -26617 6326 -26571 6360
rect -26537 6326 -26491 6360
rect -26457 6326 -26411 6360
rect -26377 6326 -26331 6360
rect -26297 6326 -26251 6360
rect -26217 6326 -26171 6360
rect -26137 6326 -26091 6360
rect -26057 6326 -26011 6360
rect -25977 6326 -25931 6360
rect -25897 6326 -25851 6360
rect -25817 6326 -25771 6360
rect -25737 6326 -25691 6360
rect -25657 6326 -25611 6360
rect -25577 6326 -25531 6360
rect -25497 6326 -25451 6360
rect -25417 6326 -25371 6360
rect -25337 6326 -25291 6360
rect -25257 6326 -25211 6360
rect -25177 6326 -25131 6360
rect -25097 6326 -25051 6360
rect -25017 6326 -24971 6360
rect -24937 6326 -24890 6360
rect -24856 6326 -24810 6360
rect -24776 6326 -24730 6360
rect -24696 6326 -24650 6360
rect -24616 6326 -24570 6360
rect -24536 6326 -24490 6360
rect -24456 6326 -24410 6360
rect -24376 6326 -24330 6360
rect -24296 6326 -24250 6360
rect -24216 6326 -24170 6360
rect -24136 6326 -24090 6360
rect -24056 6326 -24010 6360
rect -23976 6326 -23930 6360
rect -23896 6326 -23850 6360
rect -23816 6326 -23770 6360
rect -23736 6326 -23690 6360
rect -23656 6326 -23610 6360
rect -23576 6326 -23530 6360
rect -23496 6326 -23450 6360
rect -23416 6326 -23370 6360
rect -23336 6326 -23290 6360
rect -23256 6326 -23210 6360
rect -23176 6326 -23130 6360
rect -23096 6326 -23050 6360
rect -23016 6326 -22970 6360
rect -22936 6326 -22890 6360
rect -22856 6326 -22810 6360
rect -22776 6326 -22730 6360
rect -22696 6326 -22650 6360
rect -22616 6326 -22570 6360
rect -22536 6326 -22490 6360
rect -22456 6326 -22410 6360
rect -22376 6326 -22330 6360
rect -22296 6326 -22250 6360
rect -22216 6326 -22170 6360
rect -22136 6326 -22090 6360
rect -22056 6326 -22010 6360
rect -21976 6326 -21930 6360
rect -21896 6326 -21850 6360
rect -21816 6326 -21770 6360
rect -21736 6326 -21690 6360
rect -21656 6326 -21610 6360
rect -21576 6326 -21530 6360
rect -21496 6326 -21450 6360
rect -21416 6326 -21370 6360
rect -21336 6326 -21290 6360
rect -21256 6326 -21210 6360
rect -21176 6326 -21130 6360
rect -21096 6326 -21050 6360
rect -21016 6326 -20970 6360
rect -20936 6326 -20890 6360
rect -20856 6326 -20810 6360
rect -20776 6326 -20730 6360
rect -20696 6326 -20650 6360
rect -20616 6326 -20570 6360
rect -20536 6326 -20490 6360
rect -20456 6326 -20410 6360
rect -20376 6326 -20330 6360
rect -20296 6326 -20250 6360
rect -20216 6326 -20170 6360
rect -20136 6326 -20090 6360
rect -20056 6326 -20010 6360
rect -19976 6326 -19930 6360
rect -19896 6326 -19850 6360
rect -19816 6326 -19770 6360
rect -19736 6326 -19690 6360
rect -19656 6326 -19610 6360
rect -19576 6326 -19530 6360
rect -19496 6326 -19450 6360
rect -19416 6326 -19370 6360
rect -19336 6326 -19290 6360
rect -19256 6326 -19210 6360
rect -19176 6326 -19130 6360
rect -19096 6326 -19050 6360
rect -19016 6326 -18970 6360
rect -18936 6326 -18890 6360
rect -18856 6326 -18810 6360
rect -18776 6326 -18730 6360
rect -18696 6326 -18650 6360
rect -18616 6326 -18570 6360
rect -18536 6326 -18490 6360
rect -18456 6326 -18410 6360
rect -18376 6326 -18330 6360
rect -18296 6326 -18250 6360
rect -18216 6326 -18170 6360
rect -18136 6326 -18090 6360
rect -18056 6326 -18010 6360
rect -17976 6326 -17930 6360
rect -17896 6326 -17850 6360
rect -17816 6326 -17770 6360
rect -17736 6326 -17690 6360
rect -17656 6326 -17610 6360
rect -17576 6326 -17530 6360
rect -17496 6326 -17450 6360
rect -17416 6326 -17370 6360
rect -17336 6326 -17290 6360
rect -17256 6326 -17210 6360
rect -17176 6326 -17130 6360
rect -17096 6326 -17050 6360
rect -17016 6326 -16970 6360
rect -16936 6326 -16890 6360
rect -16856 6326 -16810 6360
rect -16776 6326 -16730 6360
rect -16696 6326 -16650 6360
rect -16616 6326 -16570 6360
rect -16536 6326 -16490 6360
rect -16456 6326 -16410 6360
rect -16376 6326 -16330 6360
rect -16296 6326 -16250 6360
rect -16216 6326 -16170 6360
rect -16136 6326 -16090 6360
rect -16056 6326 -16010 6360
rect -15976 6326 -15930 6360
rect -15896 6326 -15850 6360
rect -15816 6326 -15770 6360
rect -15736 6326 -15690 6360
rect -15656 6326 -15610 6360
rect -15576 6326 -15530 6360
rect -15496 6326 -15450 6360
rect -15416 6326 -15370 6360
rect -15336 6326 -15290 6360
rect -15256 6326 -15210 6360
rect -15176 6326 -15130 6360
rect -15096 6326 -15050 6360
rect -15016 6326 -14970 6360
rect -14936 6326 -14890 6360
rect -14856 6326 -14810 6360
rect -14776 6326 -14730 6360
rect -14696 6326 -14650 6360
rect -14616 6326 -14570 6360
rect -14536 6326 -14490 6360
rect -14456 6326 -14410 6360
rect -14376 6326 -14330 6360
rect -14296 6326 -14250 6360
rect -14216 6326 -14170 6360
rect -14136 6326 -14090 6360
rect -14056 6326 -14010 6360
rect -13976 6326 -13930 6360
rect -13896 6326 -13850 6360
rect -13816 6326 -13770 6360
rect -13736 6326 -13690 6360
rect -13656 6326 -13610 6360
rect -13576 6326 -13530 6360
rect -13496 6326 -13450 6360
rect -13416 6326 -13370 6360
rect -13336 6326 -13290 6360
rect -13256 6326 -13210 6360
rect -13176 6326 -13130 6360
rect -13096 6326 -13050 6360
rect -13016 6326 -12970 6360
rect -12936 6326 -12890 6360
rect -12856 6326 -12810 6360
rect -12776 6326 -12730 6360
rect -12696 6326 -12650 6360
rect -12616 6326 -12570 6360
rect -12536 6326 -12490 6360
rect -12456 6326 -12410 6360
rect -12376 6326 -12330 6360
rect -12296 6326 -12250 6360
rect -12216 6326 -12170 6360
rect -12136 6326 -12090 6360
rect -12056 6326 -12010 6360
rect -11976 6326 -11929 6360
rect -11895 6326 -11849 6360
rect -11815 6326 -11769 6360
rect -11735 6326 -11689 6360
rect -11655 6326 -11609 6360
rect -11575 6326 -11529 6360
rect -11495 6326 -11449 6360
rect -11415 6326 -11369 6360
rect -11335 6326 -11289 6360
rect -11255 6326 -11209 6360
rect -11175 6326 -11129 6360
rect -11095 6326 -11049 6360
rect -11015 6326 -10969 6360
rect -10935 6326 -10889 6360
rect -10855 6326 -10809 6360
rect -10775 6326 -10729 6360
rect -10695 6326 -10649 6360
rect -10615 6326 -10569 6360
rect -10535 6326 -10489 6360
rect -10455 6326 -10409 6360
rect -10375 6326 -10329 6360
rect -10295 6326 -10249 6360
rect -10215 6326 -10169 6360
rect -10135 6326 -10089 6360
rect -10055 6326 -10009 6360
rect -9975 6326 -9929 6360
rect -9895 6326 -9849 6360
rect -9815 6326 -9769 6360
rect -9735 6326 -9689 6360
rect -9655 6326 -9609 6360
rect -9575 6326 -9529 6360
rect -9495 6326 -9449 6360
rect -9415 6326 -9369 6360
rect -9335 6326 -9289 6360
rect -9255 6326 -9209 6360
rect -9175 6326 -9129 6360
rect -9095 6326 -9049 6360
rect -9015 6326 -8969 6360
rect -8935 6326 -8889 6360
rect -8855 6326 -8809 6360
rect -8775 6326 -8729 6360
rect -8695 6326 -8649 6360
rect -8615 6326 -8569 6360
rect -8535 6326 -8489 6360
rect -8455 6326 -8409 6360
rect -8375 6326 -8329 6360
rect -8295 6326 -8249 6360
rect -8215 6326 -8169 6360
rect -8135 6326 -8089 6360
rect -8055 6326 -8009 6360
rect -7975 6326 -7929 6360
rect -7895 6326 -7849 6360
rect -7815 6326 -7769 6360
rect -7735 6326 -7689 6360
rect -7655 6326 -7609 6360
rect -7575 6326 -7529 6360
rect -7495 6326 -7449 6360
rect -7415 6326 -7369 6360
rect -7335 6326 -7289 6360
rect -7255 6326 -7209 6360
rect -7175 6326 -7129 6360
rect -7095 6326 -7049 6360
rect -7015 6326 -6969 6360
rect -6935 6326 -6889 6360
rect -6855 6326 -6809 6360
rect -6775 6326 -6729 6360
rect -6695 6326 -6649 6360
rect -6615 6326 -6569 6360
rect -6535 6326 -6489 6360
rect -6455 6326 -6409 6360
rect -6375 6326 -6329 6360
rect -6295 6326 -6249 6360
rect -6215 6326 -6169 6360
rect -6135 6326 -6089 6360
rect -6055 6326 -6009 6360
rect -5975 6326 -5929 6360
rect -5895 6326 -5849 6360
rect -5815 6326 -5769 6360
rect -5735 6326 -5689 6360
rect -5655 6326 -5609 6360
rect -5575 6326 -5529 6360
rect -5495 6326 -5449 6360
rect -5415 6326 -5369 6360
rect -5335 6326 -5289 6360
rect -5255 6326 -5209 6360
rect -5175 6326 -5129 6360
rect -5095 6326 -5049 6360
rect -5015 6326 -4969 6360
rect -4935 6326 -4889 6360
rect -4855 6326 -4809 6360
rect -4775 6326 -4729 6360
rect -4695 6326 -4649 6360
rect -4615 6326 -4569 6360
rect -4535 6326 -4489 6360
rect -4455 6326 -4409 6360
rect -4375 6326 -4329 6360
rect -4295 6326 -4249 6360
rect -4215 6326 -4169 6360
rect -4135 6326 -4089 6360
rect -4055 6326 -4009 6360
rect -3975 6326 -3929 6360
rect -3895 6326 -3849 6360
rect -3815 6326 -3769 6360
rect -3735 6326 -3689 6360
rect -3655 6326 -3609 6360
rect -3575 6326 -3529 6360
rect -3495 6326 -3449 6360
rect -3415 6326 -3369 6360
rect -3335 6326 -3289 6360
rect -3255 6326 -3209 6360
rect -3175 6326 -3129 6360
rect -3095 6326 -3049 6360
rect -3015 6326 -2969 6360
rect -2935 6326 -2889 6360
rect -2855 6326 -2809 6360
rect -2775 6326 -2729 6360
rect -2695 6326 -2649 6360
rect -2615 6326 -2569 6360
rect -2535 6326 -2489 6360
rect -2455 6326 -2409 6360
rect -2375 6326 -2329 6360
rect -2295 6326 -2249 6360
rect -2215 6326 -2169 6360
rect -2135 6326 -2089 6360
rect -2055 6326 -2009 6360
rect -1975 6326 -1929 6360
rect -1895 6326 -1849 6360
rect -1815 6326 -1769 6360
rect -1735 6326 -1689 6360
rect -1655 6326 -1609 6360
rect -1575 6326 -1529 6360
rect -1495 6326 -1449 6360
rect -1415 6326 -1369 6360
rect -1335 6326 -1289 6360
rect -1255 6326 -1209 6360
rect -1175 6326 -1129 6360
rect -1095 6326 -1049 6360
rect -1015 6326 -969 6360
rect -935 6326 -889 6360
rect -855 6326 -809 6360
rect -775 6326 -729 6360
rect -695 6326 -649 6360
rect -615 6326 -569 6360
rect -535 6326 -489 6360
rect -455 6326 -409 6360
rect -375 6326 -329 6360
rect -295 6326 -249 6360
rect -215 6326 -169 6360
rect -135 6326 -89 6360
rect -55 6326 -9 6360
rect 25 6326 71 6360
rect 105 6326 151 6360
rect 185 6326 231 6360
rect 265 6326 311 6360
rect 345 6326 391 6360
rect 425 6326 471 6360
rect 505 6326 551 6360
rect 585 6326 631 6360
rect 665 6326 711 6360
rect 745 6326 791 6360
rect 825 6326 871 6360
rect 905 6326 951 6360
rect 985 6326 1031 6360
rect 1065 6326 1111 6360
rect 1145 6326 1191 6360
rect 1225 6326 1271 6360
rect 1305 6326 1351 6360
rect 1385 6326 1431 6360
rect 1465 6326 1511 6360
rect 1545 6326 1591 6360
rect 1625 6326 1671 6360
rect 1705 6326 1751 6360
rect 1785 6326 1831 6360
rect 1865 6326 1911 6360
rect 1945 6326 1991 6360
rect 2025 6326 2071 6360
rect 2105 6326 2151 6360
rect 2185 6326 2231 6360
rect 2265 6326 2311 6360
rect 2345 6326 2391 6360
rect 2425 6326 2471 6360
rect 2505 6326 2551 6360
rect 2585 6326 2631 6360
rect 2665 6326 2711 6360
rect 2745 6326 2791 6360
rect 2825 6326 2871 6360
rect 2905 6326 2951 6360
rect 2985 6326 3031 6360
rect 3065 6326 3111 6360
rect 3145 6326 3191 6360
rect 3225 6326 3271 6360
rect 3305 6326 3351 6360
rect 3385 6326 3431 6360
rect 3465 6326 3511 6360
rect 3545 6326 3591 6360
rect 3625 6326 3671 6360
rect 3705 6326 3751 6360
rect 3785 6326 3831 6360
rect 3865 6326 3911 6360
rect 3945 6326 3991 6360
rect 4025 6326 4071 6360
rect 4105 6326 4151 6360
rect 4185 6326 4231 6360
rect 4265 6326 4311 6360
rect 4345 6326 4391 6360
rect 4425 6326 4471 6360
rect 4505 6326 4551 6360
rect 4585 6326 4631 6360
rect 4665 6326 4711 6360
rect 4745 6326 4791 6360
rect 4825 6326 4871 6360
rect 4905 6326 4951 6360
rect 4985 6326 5031 6360
rect 5065 6326 5111 6360
rect 5145 6326 5191 6360
rect 5225 6326 5271 6360
rect 5305 6326 5351 6360
rect 5385 6326 5431 6360
rect 5465 6326 5511 6360
rect 5545 6326 5591 6360
rect 5625 6326 5671 6360
rect 5705 6326 5751 6360
rect 5785 6326 5831 6360
rect 5865 6326 5911 6360
rect 5945 6326 5991 6360
rect 6025 6326 6071 6360
rect 6105 6326 6151 6360
rect 6185 6326 6231 6360
rect 6265 6326 6311 6360
rect 6345 6326 6391 6360
rect 6425 6326 6471 6360
rect 6505 6326 6551 6360
rect 6585 6326 6631 6360
rect 6665 6326 6711 6360
rect 6745 6326 6791 6360
rect 6825 6326 6871 6360
rect 6905 6326 6951 6360
rect 6985 6326 7031 6360
rect 7065 6326 7111 6360
rect 7145 6326 7191 6360
rect 7225 6326 7271 6360
rect 7305 6326 7351 6360
rect 7385 6326 7431 6360
rect 7465 6326 7511 6360
rect 7545 6326 7591 6360
rect 7625 6326 7671 6360
rect 7705 6326 7751 6360
rect 7785 6326 7831 6360
rect 7865 6326 7911 6360
rect 7945 6326 7991 6360
rect 8025 6326 8071 6360
rect 8105 6326 8151 6360
rect 8185 6326 8231 6360
rect 8265 6326 8311 6360
rect 8345 6326 8391 6360
rect 8425 6326 8471 6360
rect 8505 6326 8551 6360
rect 8585 6326 8631 6360
rect 8665 6326 8711 6360
rect 8745 6326 8791 6360
rect 8825 6326 8871 6360
rect 8905 6326 8951 6360
rect 8985 6326 9031 6360
rect 9065 6326 9111 6360
rect 9145 6326 9191 6360
rect 9225 6326 9271 6360
rect 9305 6326 9351 6360
rect 9385 6326 9431 6360
rect 9465 6326 9511 6360
rect 9545 6326 9591 6360
rect 9625 6326 9672 6360
rect 9706 6326 9752 6360
rect 9786 6326 9832 6360
rect 9866 6326 9912 6360
rect 9946 6326 9992 6360
rect 10026 6326 10072 6360
rect 10106 6326 10152 6360
rect 10186 6326 10232 6360
rect 10266 6326 10312 6360
rect 10346 6326 10392 6360
rect 10426 6326 10472 6360
rect 10506 6326 10552 6360
rect 10586 6326 10632 6360
rect 10666 6326 10712 6360
rect 10746 6326 10792 6360
rect 10826 6326 10872 6360
rect 10906 6326 10952 6360
rect 10986 6326 11032 6360
rect 11066 6326 11112 6360
rect 11146 6326 11192 6360
rect 11226 6326 11272 6360
rect 11306 6326 11352 6360
rect 11386 6326 11432 6360
rect 11466 6326 11512 6360
rect 11546 6326 11592 6360
rect 11626 6326 11672 6360
rect 11706 6326 11752 6360
rect 11786 6326 11832 6360
rect 11866 6326 11912 6360
rect 11946 6326 11992 6360
rect 12026 6326 12072 6360
rect 12106 6326 12152 6360
rect 12186 6326 12232 6360
rect 12266 6326 12312 6360
rect 12346 6326 12392 6360
rect 12426 6326 12472 6360
rect 12506 6326 12552 6360
rect 12586 6326 12632 6360
rect 12666 6326 12712 6360
rect 12746 6326 12792 6360
rect 12826 6326 12872 6360
rect 12906 6326 12952 6360
rect 12986 6326 13032 6360
rect 13066 6326 13112 6360
rect 13146 6326 13192 6360
rect 13226 6326 13272 6360
rect 13306 6326 13352 6360
rect 13386 6326 13432 6360
rect 13466 6326 13512 6360
rect 13546 6326 13592 6360
rect 13626 6326 13672 6360
rect 13706 6326 13752 6360
rect 13786 6326 13832 6360
rect 13866 6326 13912 6360
rect 13946 6326 13992 6360
rect 14026 6326 14072 6360
rect 14106 6326 14152 6360
rect 14186 6326 14232 6360
rect 14266 6326 14312 6360
rect 14346 6326 14392 6360
rect 14426 6326 14472 6360
rect 14506 6326 14552 6360
rect 14586 6326 14632 6360
rect 14666 6326 14712 6360
rect 14746 6326 14792 6360
rect 14826 6326 14872 6360
rect 14906 6326 14952 6360
rect 14986 6326 15032 6360
rect 15066 6326 15112 6360
rect 15146 6326 15192 6360
rect 15226 6326 15272 6360
rect 15306 6326 15352 6360
rect 15386 6326 15432 6360
rect 15466 6326 15512 6360
rect 15546 6326 15592 6360
rect 15626 6326 15672 6360
rect 15706 6326 15752 6360
rect 15786 6326 15832 6360
rect 15866 6326 15912 6360
rect 15946 6326 15992 6360
rect 16026 6326 16072 6360
rect 16106 6326 16152 6360
rect 16186 6326 16232 6360
rect 16266 6326 16312 6360
rect 16346 6326 16392 6360
rect 16426 6326 16472 6360
rect 16506 6326 16552 6360
rect 16586 6326 16632 6360
rect 16666 6326 16712 6360
rect 16746 6326 16792 6360
rect 16826 6326 16872 6360
rect 16906 6326 16952 6360
rect 16986 6326 17032 6360
rect 17066 6326 17112 6360
rect 17146 6326 17192 6360
rect 17226 6326 17272 6360
rect 17306 6326 17352 6360
rect 17386 6326 17432 6360
rect 17466 6326 17512 6360
rect 17546 6326 17592 6360
rect 17626 6326 17672 6360
rect 17706 6326 17752 6360
rect 17786 6326 17832 6360
rect 17866 6326 17912 6360
rect 17946 6326 17992 6360
rect 18026 6326 18072 6360
rect 18106 6326 18152 6360
rect 18186 6326 18232 6360
rect 18266 6326 18312 6360
rect 18346 6326 18392 6360
rect 18426 6326 18472 6360
rect 18506 6326 18552 6360
rect 18586 6326 18632 6360
rect 18666 6326 18712 6360
rect 18746 6326 18792 6360
rect 18826 6326 18872 6360
rect 18906 6326 18952 6360
rect 18986 6326 19032 6360
rect 19066 6326 19112 6360
rect 19146 6326 19192 6360
rect 19226 6326 19272 6360
rect 19306 6326 19352 6360
rect 19386 6326 19432 6360
rect 19466 6326 19512 6360
rect 19546 6326 19592 6360
rect 19626 6326 19672 6360
rect 19706 6326 19752 6360
rect 19786 6326 19832 6360
rect 19866 6326 19912 6360
rect 19946 6326 19992 6360
rect 20026 6326 20072 6360
rect 20106 6326 20152 6360
rect 20186 6326 20232 6360
rect 20266 6326 20312 6360
rect 20346 6326 20392 6360
rect 20426 6326 20472 6360
rect 20506 6326 20552 6360
rect 20586 6326 20632 6360
rect 20666 6326 20712 6360
rect 20746 6326 20792 6360
rect 20826 6326 20872 6360
rect 20906 6326 20952 6360
rect 20986 6326 21032 6360
rect 21066 6326 21112 6360
rect 21146 6326 21192 6360
rect 21226 6326 21272 6360
rect 21306 6326 21352 6360
rect 21386 6326 21432 6360
rect 21466 6326 21512 6360
rect 21546 6326 21592 6360
rect 21626 6326 21672 6360
rect 21706 6326 21752 6360
rect 21786 6326 21832 6360
rect 21866 6326 21912 6360
rect 21946 6326 21992 6360
rect 22026 6326 22072 6360
rect 22106 6326 22152 6360
rect 22186 6326 22232 6360
rect 22266 6326 22312 6360
rect 22346 6326 22392 6360
rect 22426 6326 22472 6360
rect 22506 6326 22552 6360
rect 22586 6326 22633 6360
rect 22667 6326 22713 6360
rect 22747 6326 22793 6360
rect 22827 6326 22873 6360
rect 22907 6326 22953 6360
rect 22987 6326 23033 6360
rect 23067 6326 23113 6360
rect 23147 6326 23193 6360
rect 23227 6326 23273 6360
rect 23307 6326 23353 6360
rect 23387 6326 23433 6360
rect 23467 6326 23513 6360
rect 23547 6326 23593 6360
rect 23627 6326 23673 6360
rect 23707 6326 23753 6360
rect 23787 6326 23833 6360
rect 23867 6326 23913 6360
rect 23947 6326 23993 6360
rect 24027 6326 24073 6360
rect 24107 6326 24153 6360
rect 24187 6326 24233 6360
rect 24267 6326 24313 6360
rect 24347 6326 24393 6360
rect 24427 6326 24473 6360
rect 24507 6326 24553 6360
rect 24587 6326 24633 6360
rect 24667 6326 24713 6360
rect 24747 6326 24793 6360
rect 24827 6326 24873 6360
rect 24907 6326 24953 6360
rect 24987 6326 25033 6360
rect 25067 6326 25113 6360
rect 25147 6326 25193 6360
rect 25227 6326 25273 6360
rect 25307 6326 25353 6360
rect 25387 6326 25433 6360
rect 25467 6326 25513 6360
rect 25547 6326 25593 6360
rect 25627 6326 25673 6360
rect 25707 6326 25753 6360
rect 25787 6326 25833 6360
rect 25867 6326 25913 6360
rect 25947 6326 25993 6360
rect 26027 6326 26073 6360
rect 26107 6326 26153 6360
rect 26187 6326 26233 6360
rect 26267 6326 26313 6360
rect 26347 6326 26393 6360
rect 26427 6326 26473 6360
rect 26507 6326 26553 6360
rect 26587 6326 26633 6360
rect 26667 6326 26713 6360
rect 26747 6326 26793 6360
rect 26827 6326 26873 6360
rect 26907 6326 26953 6360
rect 26987 6326 27033 6360
rect 27067 6326 27113 6360
rect 27147 6326 27193 6360
rect 27227 6326 27273 6360
rect 27307 6326 27353 6360
rect 27387 6326 27433 6360
rect 27467 6326 27513 6360
rect 27547 6326 27593 6360
rect 27627 6326 27673 6360
rect 27707 6326 27753 6360
rect 27787 6326 27833 6360
rect 27867 6326 27913 6360
rect 27947 6326 27993 6360
rect 28027 6326 28073 6360
rect 28107 6326 28153 6360
rect 28187 6326 28233 6360
rect 28267 6326 28313 6360
rect 28347 6326 28393 6360
rect 28427 6326 28473 6360
rect 28507 6326 28553 6360
rect 28587 6326 28633 6360
rect 28667 6326 28713 6360
rect 28747 6326 28793 6360
rect 28827 6326 28873 6360
rect 28907 6326 28953 6360
rect 28987 6326 29033 6360
rect 29067 6326 29113 6360
rect 29147 6326 29193 6360
rect 29227 6326 29273 6360
rect 29307 6326 29353 6360
rect 29387 6326 29433 6360
rect 29467 6326 29513 6360
rect 29547 6326 29593 6360
rect 29627 6326 29673 6360
rect 29707 6326 29753 6360
rect 29787 6326 29833 6360
rect 29867 6326 29913 6360
rect 29947 6326 29993 6360
rect 30027 6326 30073 6360
rect 30107 6326 30153 6360
rect 30187 6326 30233 6360
rect 30267 6326 30313 6360
rect 30347 6326 30393 6360
rect 30427 6326 30473 6360
rect 30507 6326 30553 6360
rect 30587 6326 30633 6360
rect 30667 6326 30713 6360
rect 30747 6326 30793 6360
rect 30827 6326 30873 6360
rect 30907 6326 30953 6360
rect 30987 6326 31033 6360
rect 31067 6326 31113 6360
rect 31147 6326 31193 6360
rect 31227 6326 31274 6360
rect 31308 6326 31354 6360
rect 31388 6326 31434 6360
rect 31468 6326 31514 6360
rect 31548 6326 31594 6360
rect 31628 6326 31674 6360
rect 31708 6326 31754 6360
rect 31788 6326 31834 6360
rect 31868 6326 31914 6360
rect 31948 6326 31994 6360
rect 32028 6326 32074 6360
rect 32108 6326 32154 6360
rect 32188 6326 32234 6360
rect 32268 6326 32314 6360
rect 32348 6326 32394 6360
rect 32428 6326 32474 6360
rect 32508 6326 32554 6360
rect 32588 6326 32634 6360
rect 32668 6326 32714 6360
rect 32748 6326 32794 6360
rect 32828 6326 32874 6360
rect 32908 6326 32954 6360
rect 32988 6326 33034 6360
rect 33068 6326 33114 6360
rect 33148 6326 33194 6360
rect 33228 6326 33274 6360
rect 33308 6326 33354 6360
rect 33388 6326 33434 6360
rect 33468 6326 33514 6360
rect 33548 6326 33594 6360
rect 33628 6326 33674 6360
rect 33708 6326 33754 6360
rect 33788 6326 33834 6360
rect 33868 6326 33914 6360
rect 33948 6326 33994 6360
rect 34028 6326 34074 6360
rect 34108 6326 34154 6360
rect 34188 6326 34234 6360
rect 34268 6326 34314 6360
rect 34348 6326 34394 6360
rect 34428 6326 34474 6360
rect 34508 6326 34554 6360
rect 34588 6326 34634 6360
rect 34668 6326 34714 6360
rect 34748 6326 34794 6360
rect 34828 6326 34874 6360
rect 34908 6326 34954 6360
rect 34988 6326 35034 6360
rect 35068 6326 35114 6360
rect 35148 6326 35194 6360
rect 35228 6326 35274 6360
rect 35308 6326 35354 6360
rect 35388 6326 35434 6360
rect 35468 6326 35514 6360
rect 35548 6326 35594 6360
rect -37897 6303 35594 6326
rect -285 5631 -25 5891
rect 1341 5631 1601 5891
rect -34951 4821 -343 4844
rect -34951 4787 -34905 4821
rect -34871 4787 -34825 4821
rect -34791 4787 -34745 4821
rect -34711 4787 -34665 4821
rect -34631 4787 -34585 4821
rect -34551 4787 -34505 4821
rect -34471 4787 -34425 4821
rect -34391 4787 -34345 4821
rect -34311 4787 -34265 4821
rect -34231 4787 -34185 4821
rect -34151 4787 -34105 4821
rect -34071 4787 -34025 4821
rect -33991 4787 -33945 4821
rect -33911 4787 -33865 4821
rect -33831 4787 -33785 4821
rect -33751 4787 -33705 4821
rect -33671 4787 -33625 4821
rect -33591 4787 -33545 4821
rect -33511 4787 -33465 4821
rect -33431 4787 -33385 4821
rect -33351 4787 -33305 4821
rect -33271 4787 -33225 4821
rect -33191 4787 -33145 4821
rect -33111 4787 -33065 4821
rect -33031 4787 -32985 4821
rect -32951 4787 -32905 4821
rect -32871 4787 -32825 4821
rect -32791 4787 -32745 4821
rect -32711 4787 -32665 4821
rect -32631 4787 -32585 4821
rect -32551 4787 -32505 4821
rect -32471 4787 -32425 4821
rect -32391 4787 -32345 4821
rect -32311 4787 -32265 4821
rect -32231 4787 -32185 4821
rect -32151 4787 -32105 4821
rect -32071 4787 -32025 4821
rect -31991 4787 -31945 4821
rect -31911 4787 -31865 4821
rect -31831 4787 -31785 4821
rect -31751 4787 -31705 4821
rect -31671 4787 -31625 4821
rect -31591 4787 -31545 4821
rect -31511 4787 -31465 4821
rect -31431 4787 -31385 4821
rect -31351 4787 -31305 4821
rect -31271 4787 -31225 4821
rect -31191 4787 -31145 4821
rect -31111 4787 -31065 4821
rect -31031 4787 -30985 4821
rect -30951 4787 -30905 4821
rect -30871 4787 -30825 4821
rect -30791 4787 -30745 4821
rect -30711 4787 -30665 4821
rect -30631 4787 -30585 4821
rect -30551 4787 -30505 4821
rect -30471 4787 -30425 4821
rect -30391 4787 -30345 4821
rect -30311 4787 -30265 4821
rect -30231 4787 -30185 4821
rect -30151 4787 -30105 4821
rect -30071 4787 -30025 4821
rect -29991 4787 -29945 4821
rect -29911 4787 -29865 4821
rect -29831 4787 -29785 4821
rect -29751 4787 -29705 4821
rect -29671 4787 -29625 4821
rect -29591 4787 -29545 4821
rect -29511 4787 -29465 4821
rect -29431 4787 -29385 4821
rect -29351 4787 -29305 4821
rect -29271 4787 -29225 4821
rect -29191 4787 -29145 4821
rect -29111 4787 -29065 4821
rect -29031 4787 -28985 4821
rect -28951 4787 -28905 4821
rect -28871 4787 -28825 4821
rect -28791 4787 -28745 4821
rect -28711 4787 -28665 4821
rect -28631 4787 -28585 4821
rect -28551 4787 -28505 4821
rect -28471 4787 -28425 4821
rect -28391 4787 -28345 4821
rect -28311 4787 -28265 4821
rect -28231 4787 -28185 4821
rect -28151 4787 -28105 4821
rect -28071 4787 -28025 4821
rect -27991 4787 -27945 4821
rect -27911 4787 -27865 4821
rect -27831 4787 -27785 4821
rect -27751 4787 -27705 4821
rect -27671 4787 -27625 4821
rect -27591 4787 -27545 4821
rect -27511 4787 -27465 4821
rect -27431 4787 -27385 4821
rect -27351 4787 -27305 4821
rect -27271 4787 -27225 4821
rect -27191 4787 -27145 4821
rect -27111 4787 -27065 4821
rect -27031 4787 -26985 4821
rect -26951 4787 -26905 4821
rect -26871 4787 -26825 4821
rect -26791 4787 -26745 4821
rect -26711 4787 -26665 4821
rect -26631 4787 -26585 4821
rect -26551 4787 -26505 4821
rect -26471 4787 -26425 4821
rect -26391 4787 -26345 4821
rect -26311 4787 -26265 4821
rect -26231 4787 -26185 4821
rect -26151 4787 -26105 4821
rect -26071 4787 -26025 4821
rect -25991 4787 -25945 4821
rect -25911 4787 -25865 4821
rect -25831 4787 -25785 4821
rect -25751 4787 -25705 4821
rect -25671 4787 -25625 4821
rect -25591 4787 -25545 4821
rect -25511 4787 -25465 4821
rect -25431 4787 -25385 4821
rect -25351 4787 -25305 4821
rect -25271 4787 -25225 4821
rect -25191 4787 -25145 4821
rect -25111 4787 -25065 4821
rect -25031 4787 -24985 4821
rect -24951 4787 -24905 4821
rect -24871 4787 -24825 4821
rect -24791 4787 -24745 4821
rect -24711 4787 -24665 4821
rect -24631 4787 -24585 4821
rect -24551 4787 -24505 4821
rect -24471 4787 -24425 4821
rect -24391 4787 -24345 4821
rect -24311 4787 -24265 4821
rect -24231 4787 -24185 4821
rect -24151 4787 -24105 4821
rect -24071 4787 -24025 4821
rect -23991 4787 -23945 4821
rect -23911 4787 -23865 4821
rect -23831 4787 -23785 4821
rect -23751 4787 -23705 4821
rect -23671 4787 -23625 4821
rect -23591 4787 -23545 4821
rect -23511 4787 -23465 4821
rect -23431 4787 -23385 4821
rect -23351 4787 -23305 4821
rect -23271 4787 -23225 4821
rect -23191 4787 -23145 4821
rect -23111 4787 -23065 4821
rect -23031 4787 -22985 4821
rect -22951 4787 -22905 4821
rect -22871 4787 -22825 4821
rect -22791 4787 -22745 4821
rect -22711 4787 -22665 4821
rect -22631 4787 -22585 4821
rect -22551 4787 -22505 4821
rect -22471 4787 -22425 4821
rect -22391 4787 -22345 4821
rect -22311 4787 -22265 4821
rect -22231 4787 -22185 4821
rect -22151 4787 -22105 4821
rect -22071 4787 -22025 4821
rect -21991 4787 -21944 4821
rect -21910 4787 -21864 4821
rect -21830 4787 -21784 4821
rect -21750 4787 -21704 4821
rect -21670 4787 -21624 4821
rect -21590 4787 -21544 4821
rect -21510 4787 -21464 4821
rect -21430 4787 -21384 4821
rect -21350 4787 -21304 4821
rect -21270 4787 -21224 4821
rect -21190 4787 -21144 4821
rect -21110 4787 -21064 4821
rect -21030 4787 -20984 4821
rect -20950 4787 -20904 4821
rect -20870 4787 -20824 4821
rect -20790 4787 -20744 4821
rect -20710 4787 -20664 4821
rect -20630 4787 -20584 4821
rect -20550 4787 -20504 4821
rect -20470 4787 -20424 4821
rect -20390 4787 -20344 4821
rect -20310 4787 -20264 4821
rect -20230 4787 -20184 4821
rect -20150 4787 -20104 4821
rect -20070 4787 -20024 4821
rect -19990 4787 -19944 4821
rect -19910 4787 -19864 4821
rect -19830 4787 -19784 4821
rect -19750 4787 -19704 4821
rect -19670 4787 -19624 4821
rect -19590 4787 -19544 4821
rect -19510 4787 -19464 4821
rect -19430 4787 -19384 4821
rect -19350 4787 -19304 4821
rect -19270 4787 -19224 4821
rect -19190 4787 -19144 4821
rect -19110 4787 -19064 4821
rect -19030 4787 -18984 4821
rect -18950 4787 -18904 4821
rect -18870 4787 -18824 4821
rect -18790 4787 -18744 4821
rect -18710 4787 -18664 4821
rect -18630 4787 -18584 4821
rect -18550 4787 -18504 4821
rect -18470 4787 -18424 4821
rect -18390 4787 -18344 4821
rect -18310 4787 -18264 4821
rect -18230 4787 -18184 4821
rect -18150 4787 -18104 4821
rect -18070 4787 -18024 4821
rect -17990 4787 -17944 4821
rect -17910 4787 -17864 4821
rect -17830 4787 -17784 4821
rect -17750 4787 -17704 4821
rect -17670 4787 -17624 4821
rect -17590 4787 -17544 4821
rect -17510 4787 -17464 4821
rect -17430 4787 -17384 4821
rect -17350 4787 -17304 4821
rect -17270 4787 -17224 4821
rect -17190 4787 -17144 4821
rect -17110 4787 -17064 4821
rect -17030 4787 -16984 4821
rect -16950 4787 -16904 4821
rect -16870 4787 -16824 4821
rect -16790 4787 -16744 4821
rect -16710 4787 -16664 4821
rect -16630 4787 -16584 4821
rect -16550 4787 -16504 4821
rect -16470 4787 -16424 4821
rect -16390 4787 -16344 4821
rect -16310 4787 -16264 4821
rect -16230 4787 -16184 4821
rect -16150 4787 -16104 4821
rect -16070 4787 -16024 4821
rect -15990 4787 -15944 4821
rect -15910 4787 -15864 4821
rect -15830 4787 -15784 4821
rect -15750 4787 -15704 4821
rect -15670 4787 -15624 4821
rect -15590 4787 -15544 4821
rect -15510 4787 -15464 4821
rect -15430 4787 -15384 4821
rect -15350 4787 -15304 4821
rect -15270 4787 -15224 4821
rect -15190 4787 -15144 4821
rect -15110 4787 -15064 4821
rect -15030 4787 -14984 4821
rect -14950 4787 -14904 4821
rect -14870 4787 -14824 4821
rect -14790 4787 -14744 4821
rect -14710 4787 -14664 4821
rect -14630 4787 -14584 4821
rect -14550 4787 -14504 4821
rect -14470 4787 -14424 4821
rect -14390 4787 -14344 4821
rect -14310 4787 -14264 4821
rect -14230 4787 -14184 4821
rect -14150 4787 -14104 4821
rect -14070 4787 -14024 4821
rect -13990 4787 -13944 4821
rect -13910 4787 -13864 4821
rect -13830 4787 -13784 4821
rect -13750 4787 -13704 4821
rect -13670 4787 -13624 4821
rect -13590 4787 -13544 4821
rect -13510 4787 -13464 4821
rect -13430 4787 -13384 4821
rect -13350 4787 -13304 4821
rect -13270 4787 -13224 4821
rect -13190 4787 -13144 4821
rect -13110 4787 -13064 4821
rect -13030 4787 -12984 4821
rect -12950 4787 -12904 4821
rect -12870 4787 -12824 4821
rect -12790 4787 -12744 4821
rect -12710 4787 -12664 4821
rect -12630 4787 -12584 4821
rect -12550 4787 -12504 4821
rect -12470 4787 -12424 4821
rect -12390 4787 -12344 4821
rect -12310 4787 -12264 4821
rect -12230 4787 -12184 4821
rect -12150 4787 -12104 4821
rect -12070 4787 -12024 4821
rect -11990 4787 -11944 4821
rect -11910 4787 -11864 4821
rect -11830 4787 -11784 4821
rect -11750 4787 -11704 4821
rect -11670 4787 -11624 4821
rect -11590 4787 -11544 4821
rect -11510 4787 -11464 4821
rect -11430 4787 -11384 4821
rect -11350 4787 -11304 4821
rect -11270 4787 -11224 4821
rect -11190 4787 -11144 4821
rect -11110 4787 -11064 4821
rect -11030 4787 -10984 4821
rect -10950 4787 -10904 4821
rect -10870 4787 -10824 4821
rect -10790 4787 -10744 4821
rect -10710 4787 -10664 4821
rect -10630 4787 -10584 4821
rect -10550 4787 -10504 4821
rect -10470 4787 -10424 4821
rect -10390 4787 -10344 4821
rect -10310 4787 -10264 4821
rect -10230 4787 -10184 4821
rect -10150 4787 -10104 4821
rect -10070 4787 -10024 4821
rect -9990 4787 -9944 4821
rect -9910 4787 -9864 4821
rect -9830 4787 -9784 4821
rect -9750 4787 -9704 4821
rect -9670 4787 -9624 4821
rect -9590 4787 -9544 4821
rect -9510 4787 -9464 4821
rect -9430 4787 -9384 4821
rect -9350 4787 -9304 4821
rect -9270 4787 -9224 4821
rect -9190 4787 -9144 4821
rect -9110 4787 -9064 4821
rect -9030 4787 -8983 4821
rect -8949 4787 -8903 4821
rect -8869 4787 -8823 4821
rect -8789 4787 -8743 4821
rect -8709 4787 -8663 4821
rect -8629 4787 -8583 4821
rect -8549 4787 -8503 4821
rect -8469 4787 -8423 4821
rect -8389 4787 -8343 4821
rect -8309 4787 -8263 4821
rect -8229 4787 -8183 4821
rect -8149 4787 -8103 4821
rect -8069 4787 -8023 4821
rect -7989 4787 -7943 4821
rect -7909 4787 -7863 4821
rect -7829 4787 -7783 4821
rect -7749 4787 -7703 4821
rect -7669 4787 -7623 4821
rect -7589 4787 -7543 4821
rect -7509 4787 -7463 4821
rect -7429 4787 -7383 4821
rect -7349 4787 -7303 4821
rect -7269 4787 -7223 4821
rect -7189 4787 -7143 4821
rect -7109 4787 -7063 4821
rect -7029 4787 -6983 4821
rect -6949 4787 -6903 4821
rect -6869 4787 -6823 4821
rect -6789 4787 -6743 4821
rect -6709 4787 -6663 4821
rect -6629 4787 -6583 4821
rect -6549 4787 -6503 4821
rect -6469 4787 -6423 4821
rect -6389 4787 -6343 4821
rect -6309 4787 -6263 4821
rect -6229 4787 -6183 4821
rect -6149 4787 -6103 4821
rect -6069 4787 -6023 4821
rect -5989 4787 -5943 4821
rect -5909 4787 -5863 4821
rect -5829 4787 -5783 4821
rect -5749 4787 -5703 4821
rect -5669 4787 -5623 4821
rect -5589 4787 -5543 4821
rect -5509 4787 -5463 4821
rect -5429 4787 -5383 4821
rect -5349 4787 -5303 4821
rect -5269 4787 -5223 4821
rect -5189 4787 -5143 4821
rect -5109 4787 -5063 4821
rect -5029 4787 -4983 4821
rect -4949 4787 -4903 4821
rect -4869 4787 -4823 4821
rect -4789 4787 -4743 4821
rect -4709 4787 -4663 4821
rect -4629 4787 -4583 4821
rect -4549 4787 -4503 4821
rect -4469 4787 -4423 4821
rect -4389 4787 -4343 4821
rect -4309 4787 -4263 4821
rect -4229 4787 -4183 4821
rect -4149 4787 -4103 4821
rect -4069 4787 -4023 4821
rect -3989 4787 -3943 4821
rect -3909 4787 -3863 4821
rect -3829 4787 -3783 4821
rect -3749 4787 -3703 4821
rect -3669 4787 -3623 4821
rect -3589 4787 -3543 4821
rect -3509 4787 -3463 4821
rect -3429 4787 -3383 4821
rect -3349 4787 -3303 4821
rect -3269 4787 -3223 4821
rect -3189 4787 -3143 4821
rect -3109 4787 -3063 4821
rect -3029 4787 -2983 4821
rect -2949 4787 -2903 4821
rect -2869 4787 -2823 4821
rect -2789 4787 -2743 4821
rect -2709 4787 -2663 4821
rect -2629 4787 -2583 4821
rect -2549 4787 -2503 4821
rect -2469 4787 -2423 4821
rect -2389 4787 -2343 4821
rect -2309 4787 -2263 4821
rect -2229 4787 -2183 4821
rect -2149 4787 -2103 4821
rect -2069 4787 -2023 4821
rect -1989 4787 -1943 4821
rect -1909 4787 -1863 4821
rect -1829 4787 -1783 4821
rect -1749 4787 -1703 4821
rect -1669 4787 -1623 4821
rect -1589 4787 -1543 4821
rect -1509 4787 -1463 4821
rect -1429 4787 -1383 4821
rect -1349 4787 -1303 4821
rect -1269 4787 -1223 4821
rect -1189 4787 -1143 4821
rect -1109 4787 -1063 4821
rect -1029 4787 -983 4821
rect -949 4787 -903 4821
rect -869 4787 -823 4821
rect -789 4787 -743 4821
rect -709 4787 -663 4821
rect -629 4787 -583 4821
rect -549 4787 -503 4821
rect -469 4787 -423 4821
rect -389 4787 -343 4821
rect -34951 4764 -343 4787
rect 1635 4821 36243 4844
rect 1635 4787 1681 4821
rect 1715 4787 1761 4821
rect 1795 4787 1841 4821
rect 1875 4787 1921 4821
rect 1955 4787 2001 4821
rect 2035 4787 2081 4821
rect 2115 4787 2161 4821
rect 2195 4787 2241 4821
rect 2275 4787 2321 4821
rect 2355 4787 2401 4821
rect 2435 4787 2481 4821
rect 2515 4787 2561 4821
rect 2595 4787 2641 4821
rect 2675 4787 2721 4821
rect 2755 4787 2801 4821
rect 2835 4787 2881 4821
rect 2915 4787 2961 4821
rect 2995 4787 3041 4821
rect 3075 4787 3121 4821
rect 3155 4787 3201 4821
rect 3235 4787 3281 4821
rect 3315 4787 3361 4821
rect 3395 4787 3441 4821
rect 3475 4787 3521 4821
rect 3555 4787 3601 4821
rect 3635 4787 3681 4821
rect 3715 4787 3761 4821
rect 3795 4787 3841 4821
rect 3875 4787 3921 4821
rect 3955 4787 4001 4821
rect 4035 4787 4081 4821
rect 4115 4787 4161 4821
rect 4195 4787 4241 4821
rect 4275 4787 4321 4821
rect 4355 4787 4401 4821
rect 4435 4787 4481 4821
rect 4515 4787 4561 4821
rect 4595 4787 4641 4821
rect 4675 4787 4721 4821
rect 4755 4787 4801 4821
rect 4835 4787 4881 4821
rect 4915 4787 4961 4821
rect 4995 4787 5041 4821
rect 5075 4787 5121 4821
rect 5155 4787 5201 4821
rect 5235 4787 5281 4821
rect 5315 4787 5361 4821
rect 5395 4787 5441 4821
rect 5475 4787 5521 4821
rect 5555 4787 5601 4821
rect 5635 4787 5681 4821
rect 5715 4787 5761 4821
rect 5795 4787 5841 4821
rect 5875 4787 5921 4821
rect 5955 4787 6001 4821
rect 6035 4787 6081 4821
rect 6115 4787 6161 4821
rect 6195 4787 6241 4821
rect 6275 4787 6321 4821
rect 6355 4787 6401 4821
rect 6435 4787 6481 4821
rect 6515 4787 6561 4821
rect 6595 4787 6641 4821
rect 6675 4787 6721 4821
rect 6755 4787 6801 4821
rect 6835 4787 6881 4821
rect 6915 4787 6961 4821
rect 6995 4787 7041 4821
rect 7075 4787 7121 4821
rect 7155 4787 7201 4821
rect 7235 4787 7281 4821
rect 7315 4787 7361 4821
rect 7395 4787 7441 4821
rect 7475 4787 7521 4821
rect 7555 4787 7601 4821
rect 7635 4787 7681 4821
rect 7715 4787 7761 4821
rect 7795 4787 7841 4821
rect 7875 4787 7921 4821
rect 7955 4787 8001 4821
rect 8035 4787 8081 4821
rect 8115 4787 8161 4821
rect 8195 4787 8241 4821
rect 8275 4787 8321 4821
rect 8355 4787 8401 4821
rect 8435 4787 8481 4821
rect 8515 4787 8561 4821
rect 8595 4787 8641 4821
rect 8675 4787 8721 4821
rect 8755 4787 8801 4821
rect 8835 4787 8881 4821
rect 8915 4787 8961 4821
rect 8995 4787 9041 4821
rect 9075 4787 9121 4821
rect 9155 4787 9201 4821
rect 9235 4787 9281 4821
rect 9315 4787 9361 4821
rect 9395 4787 9441 4821
rect 9475 4787 9521 4821
rect 9555 4787 9601 4821
rect 9635 4787 9681 4821
rect 9715 4787 9761 4821
rect 9795 4787 9841 4821
rect 9875 4787 9921 4821
rect 9955 4787 10001 4821
rect 10035 4787 10081 4821
rect 10115 4787 10161 4821
rect 10195 4787 10241 4821
rect 10275 4787 10321 4821
rect 10355 4787 10401 4821
rect 10435 4787 10481 4821
rect 10515 4787 10561 4821
rect 10595 4787 10641 4821
rect 10675 4787 10721 4821
rect 10755 4787 10801 4821
rect 10835 4787 10881 4821
rect 10915 4787 10961 4821
rect 10995 4787 11041 4821
rect 11075 4787 11121 4821
rect 11155 4787 11201 4821
rect 11235 4787 11281 4821
rect 11315 4787 11361 4821
rect 11395 4787 11441 4821
rect 11475 4787 11521 4821
rect 11555 4787 11601 4821
rect 11635 4787 11681 4821
rect 11715 4787 11761 4821
rect 11795 4787 11841 4821
rect 11875 4787 11921 4821
rect 11955 4787 12001 4821
rect 12035 4787 12081 4821
rect 12115 4787 12161 4821
rect 12195 4787 12241 4821
rect 12275 4787 12321 4821
rect 12355 4787 12401 4821
rect 12435 4787 12481 4821
rect 12515 4787 12561 4821
rect 12595 4787 12641 4821
rect 12675 4787 12721 4821
rect 12755 4787 12801 4821
rect 12835 4787 12881 4821
rect 12915 4787 12961 4821
rect 12995 4787 13041 4821
rect 13075 4787 13121 4821
rect 13155 4787 13201 4821
rect 13235 4787 13281 4821
rect 13315 4787 13361 4821
rect 13395 4787 13441 4821
rect 13475 4787 13521 4821
rect 13555 4787 13601 4821
rect 13635 4787 13681 4821
rect 13715 4787 13761 4821
rect 13795 4787 13841 4821
rect 13875 4787 13921 4821
rect 13955 4787 14001 4821
rect 14035 4787 14081 4821
rect 14115 4787 14161 4821
rect 14195 4787 14241 4821
rect 14275 4787 14321 4821
rect 14355 4787 14401 4821
rect 14435 4787 14481 4821
rect 14515 4787 14561 4821
rect 14595 4787 14642 4821
rect 14676 4787 14722 4821
rect 14756 4787 14802 4821
rect 14836 4787 14882 4821
rect 14916 4787 14962 4821
rect 14996 4787 15042 4821
rect 15076 4787 15122 4821
rect 15156 4787 15202 4821
rect 15236 4787 15282 4821
rect 15316 4787 15362 4821
rect 15396 4787 15442 4821
rect 15476 4787 15522 4821
rect 15556 4787 15602 4821
rect 15636 4787 15682 4821
rect 15716 4787 15762 4821
rect 15796 4787 15842 4821
rect 15876 4787 15922 4821
rect 15956 4787 16002 4821
rect 16036 4787 16082 4821
rect 16116 4787 16162 4821
rect 16196 4787 16242 4821
rect 16276 4787 16322 4821
rect 16356 4787 16402 4821
rect 16436 4787 16482 4821
rect 16516 4787 16562 4821
rect 16596 4787 16642 4821
rect 16676 4787 16722 4821
rect 16756 4787 16802 4821
rect 16836 4787 16882 4821
rect 16916 4787 16962 4821
rect 16996 4787 17042 4821
rect 17076 4787 17122 4821
rect 17156 4787 17202 4821
rect 17236 4787 17282 4821
rect 17316 4787 17362 4821
rect 17396 4787 17442 4821
rect 17476 4787 17522 4821
rect 17556 4787 17602 4821
rect 17636 4787 17682 4821
rect 17716 4787 17762 4821
rect 17796 4787 17842 4821
rect 17876 4787 17922 4821
rect 17956 4787 18002 4821
rect 18036 4787 18082 4821
rect 18116 4787 18162 4821
rect 18196 4787 18242 4821
rect 18276 4787 18322 4821
rect 18356 4787 18402 4821
rect 18436 4787 18482 4821
rect 18516 4787 18562 4821
rect 18596 4787 18642 4821
rect 18676 4787 18722 4821
rect 18756 4787 18802 4821
rect 18836 4787 18882 4821
rect 18916 4787 18962 4821
rect 18996 4787 19042 4821
rect 19076 4787 19122 4821
rect 19156 4787 19202 4821
rect 19236 4787 19282 4821
rect 19316 4787 19362 4821
rect 19396 4787 19442 4821
rect 19476 4787 19522 4821
rect 19556 4787 19602 4821
rect 19636 4787 19682 4821
rect 19716 4787 19762 4821
rect 19796 4787 19842 4821
rect 19876 4787 19922 4821
rect 19956 4787 20002 4821
rect 20036 4787 20082 4821
rect 20116 4787 20162 4821
rect 20196 4787 20242 4821
rect 20276 4787 20322 4821
rect 20356 4787 20402 4821
rect 20436 4787 20482 4821
rect 20516 4787 20562 4821
rect 20596 4787 20642 4821
rect 20676 4787 20722 4821
rect 20756 4787 20802 4821
rect 20836 4787 20882 4821
rect 20916 4787 20962 4821
rect 20996 4787 21042 4821
rect 21076 4787 21122 4821
rect 21156 4787 21202 4821
rect 21236 4787 21282 4821
rect 21316 4787 21362 4821
rect 21396 4787 21442 4821
rect 21476 4787 21522 4821
rect 21556 4787 21602 4821
rect 21636 4787 21682 4821
rect 21716 4787 21762 4821
rect 21796 4787 21842 4821
rect 21876 4787 21922 4821
rect 21956 4787 22002 4821
rect 22036 4787 22082 4821
rect 22116 4787 22162 4821
rect 22196 4787 22242 4821
rect 22276 4787 22322 4821
rect 22356 4787 22402 4821
rect 22436 4787 22482 4821
rect 22516 4787 22562 4821
rect 22596 4787 22642 4821
rect 22676 4787 22722 4821
rect 22756 4787 22802 4821
rect 22836 4787 22882 4821
rect 22916 4787 22962 4821
rect 22996 4787 23042 4821
rect 23076 4787 23122 4821
rect 23156 4787 23202 4821
rect 23236 4787 23282 4821
rect 23316 4787 23362 4821
rect 23396 4787 23442 4821
rect 23476 4787 23522 4821
rect 23556 4787 23602 4821
rect 23636 4787 23682 4821
rect 23716 4787 23762 4821
rect 23796 4787 23842 4821
rect 23876 4787 23922 4821
rect 23956 4787 24002 4821
rect 24036 4787 24082 4821
rect 24116 4787 24162 4821
rect 24196 4787 24242 4821
rect 24276 4787 24322 4821
rect 24356 4787 24402 4821
rect 24436 4787 24482 4821
rect 24516 4787 24562 4821
rect 24596 4787 24642 4821
rect 24676 4787 24722 4821
rect 24756 4787 24802 4821
rect 24836 4787 24882 4821
rect 24916 4787 24962 4821
rect 24996 4787 25042 4821
rect 25076 4787 25122 4821
rect 25156 4787 25202 4821
rect 25236 4787 25282 4821
rect 25316 4787 25362 4821
rect 25396 4787 25442 4821
rect 25476 4787 25522 4821
rect 25556 4787 25602 4821
rect 25636 4787 25682 4821
rect 25716 4787 25762 4821
rect 25796 4787 25842 4821
rect 25876 4787 25922 4821
rect 25956 4787 26002 4821
rect 26036 4787 26082 4821
rect 26116 4787 26162 4821
rect 26196 4787 26242 4821
rect 26276 4787 26322 4821
rect 26356 4787 26402 4821
rect 26436 4787 26482 4821
rect 26516 4787 26562 4821
rect 26596 4787 26642 4821
rect 26676 4787 26722 4821
rect 26756 4787 26802 4821
rect 26836 4787 26882 4821
rect 26916 4787 26962 4821
rect 26996 4787 27042 4821
rect 27076 4787 27122 4821
rect 27156 4787 27202 4821
rect 27236 4787 27282 4821
rect 27316 4787 27362 4821
rect 27396 4787 27442 4821
rect 27476 4787 27522 4821
rect 27556 4787 27603 4821
rect 27637 4787 27683 4821
rect 27717 4787 27763 4821
rect 27797 4787 27843 4821
rect 27877 4787 27923 4821
rect 27957 4787 28003 4821
rect 28037 4787 28083 4821
rect 28117 4787 28163 4821
rect 28197 4787 28243 4821
rect 28277 4787 28323 4821
rect 28357 4787 28403 4821
rect 28437 4787 28483 4821
rect 28517 4787 28563 4821
rect 28597 4787 28643 4821
rect 28677 4787 28723 4821
rect 28757 4787 28803 4821
rect 28837 4787 28883 4821
rect 28917 4787 28963 4821
rect 28997 4787 29043 4821
rect 29077 4787 29123 4821
rect 29157 4787 29203 4821
rect 29237 4787 29283 4821
rect 29317 4787 29363 4821
rect 29397 4787 29443 4821
rect 29477 4787 29523 4821
rect 29557 4787 29603 4821
rect 29637 4787 29683 4821
rect 29717 4787 29763 4821
rect 29797 4787 29843 4821
rect 29877 4787 29923 4821
rect 29957 4787 30003 4821
rect 30037 4787 30083 4821
rect 30117 4787 30163 4821
rect 30197 4787 30243 4821
rect 30277 4787 30323 4821
rect 30357 4787 30403 4821
rect 30437 4787 30483 4821
rect 30517 4787 30563 4821
rect 30597 4787 30643 4821
rect 30677 4787 30723 4821
rect 30757 4787 30803 4821
rect 30837 4787 30883 4821
rect 30917 4787 30963 4821
rect 30997 4787 31043 4821
rect 31077 4787 31123 4821
rect 31157 4787 31203 4821
rect 31237 4787 31283 4821
rect 31317 4787 31363 4821
rect 31397 4787 31443 4821
rect 31477 4787 31523 4821
rect 31557 4787 31603 4821
rect 31637 4787 31683 4821
rect 31717 4787 31763 4821
rect 31797 4787 31843 4821
rect 31877 4787 31923 4821
rect 31957 4787 32003 4821
rect 32037 4787 32083 4821
rect 32117 4787 32163 4821
rect 32197 4787 32243 4821
rect 32277 4787 32323 4821
rect 32357 4787 32403 4821
rect 32437 4787 32483 4821
rect 32517 4787 32563 4821
rect 32597 4787 32643 4821
rect 32677 4787 32723 4821
rect 32757 4787 32803 4821
rect 32837 4787 32883 4821
rect 32917 4787 32963 4821
rect 32997 4787 33043 4821
rect 33077 4787 33123 4821
rect 33157 4787 33203 4821
rect 33237 4787 33283 4821
rect 33317 4787 33363 4821
rect 33397 4787 33443 4821
rect 33477 4787 33523 4821
rect 33557 4787 33603 4821
rect 33637 4787 33683 4821
rect 33717 4787 33763 4821
rect 33797 4787 33843 4821
rect 33877 4787 33923 4821
rect 33957 4787 34003 4821
rect 34037 4787 34083 4821
rect 34117 4787 34163 4821
rect 34197 4787 34243 4821
rect 34277 4787 34323 4821
rect 34357 4787 34403 4821
rect 34437 4787 34483 4821
rect 34517 4787 34563 4821
rect 34597 4787 34643 4821
rect 34677 4787 34723 4821
rect 34757 4787 34803 4821
rect 34837 4787 34883 4821
rect 34917 4787 34963 4821
rect 34997 4787 35043 4821
rect 35077 4787 35123 4821
rect 35157 4787 35203 4821
rect 35237 4787 35283 4821
rect 35317 4787 35363 4821
rect 35397 4787 35443 4821
rect 35477 4787 35523 4821
rect 35557 4787 35603 4821
rect 35637 4787 35683 4821
rect 35717 4787 35763 4821
rect 35797 4787 35843 4821
rect 35877 4787 35923 4821
rect 35957 4787 36003 4821
rect 36037 4787 36083 4821
rect 36117 4787 36163 4821
rect 36197 4787 36243 4821
rect 1635 4764 36243 4787
<< viali >>
rect -37852 17163 -37818 17197
rect -37772 17163 -37738 17197
rect -37692 17163 -37658 17197
rect -37612 17163 -37578 17197
rect -37532 17163 -37498 17197
rect -37452 17163 -37418 17197
rect -37372 17163 -37338 17197
rect -37292 17163 -37258 17197
rect -37212 17163 -37178 17197
rect -37132 17163 -37098 17197
rect -37052 17163 -37018 17197
rect -36972 17163 -36938 17197
rect -36892 17163 -36858 17197
rect -36812 17163 -36778 17197
rect -36732 17163 -36698 17197
rect -36652 17163 -36618 17197
rect -36572 17163 -36538 17197
rect -36492 17163 -36458 17197
rect -36412 17163 -36378 17197
rect -36332 17163 -36298 17197
rect -36252 17163 -36218 17197
rect -36172 17163 -36138 17197
rect -36092 17163 -36058 17197
rect -36012 17163 -35978 17197
rect -35932 17163 -35898 17197
rect -35852 17163 -35818 17197
rect -35772 17163 -35738 17197
rect -35692 17163 -35658 17197
rect -35612 17163 -35578 17197
rect -35532 17163 -35498 17197
rect -35452 17163 -35418 17197
rect -35372 17163 -35338 17197
rect -35292 17163 -35258 17197
rect -35212 17163 -35178 17197
rect -35132 17163 -35098 17197
rect -35052 17163 -35018 17197
rect -34972 17163 -34938 17197
rect -34892 17163 -34858 17197
rect -34812 17163 -34778 17197
rect -34732 17163 -34698 17197
rect -34652 17163 -34618 17197
rect -34572 17163 -34538 17197
rect -34492 17163 -34458 17197
rect -34412 17163 -34378 17197
rect -34332 17163 -34298 17197
rect -34252 17163 -34218 17197
rect -34172 17163 -34138 17197
rect -34092 17163 -34058 17197
rect -34012 17163 -33978 17197
rect -33932 17163 -33898 17197
rect -33852 17163 -33818 17197
rect -33772 17163 -33738 17197
rect -33692 17163 -33658 17197
rect -33612 17163 -33578 17197
rect -33532 17163 -33498 17197
rect -33452 17163 -33418 17197
rect -33372 17163 -33338 17197
rect -33292 17163 -33258 17197
rect -33212 17163 -33178 17197
rect -33132 17163 -33098 17197
rect -33052 17163 -33018 17197
rect -32972 17163 -32938 17197
rect -32892 17163 -32858 17197
rect -32812 17163 -32778 17197
rect -32732 17163 -32698 17197
rect -32652 17163 -32618 17197
rect -32572 17163 -32538 17197
rect -32492 17163 -32458 17197
rect -32412 17163 -32378 17197
rect -32332 17163 -32298 17197
rect -32252 17163 -32218 17197
rect -32172 17163 -32138 17197
rect -32092 17163 -32058 17197
rect -32012 17163 -31978 17197
rect -31932 17163 -31898 17197
rect -31852 17163 -31818 17197
rect -31772 17163 -31738 17197
rect -31692 17163 -31658 17197
rect -31612 17163 -31578 17197
rect -31532 17163 -31498 17197
rect -31452 17163 -31418 17197
rect -31372 17163 -31338 17197
rect -31292 17163 -31258 17197
rect -31212 17163 -31178 17197
rect -31132 17163 -31098 17197
rect -31052 17163 -31018 17197
rect -30972 17163 -30938 17197
rect -30892 17163 -30858 17197
rect -30812 17163 -30778 17197
rect -30732 17163 -30698 17197
rect -30652 17163 -30618 17197
rect -30572 17163 -30538 17197
rect -30492 17163 -30458 17197
rect -30412 17163 -30378 17197
rect -30332 17163 -30298 17197
rect -30252 17163 -30218 17197
rect -30172 17163 -30138 17197
rect -30092 17163 -30058 17197
rect -30012 17163 -29978 17197
rect -29932 17163 -29898 17197
rect -29852 17163 -29818 17197
rect -29772 17163 -29738 17197
rect -29692 17163 -29658 17197
rect -29612 17163 -29578 17197
rect -29532 17163 -29498 17197
rect -29452 17163 -29418 17197
rect -29372 17163 -29338 17197
rect -29292 17163 -29258 17197
rect -29212 17163 -29178 17197
rect -29132 17163 -29098 17197
rect -29052 17163 -29018 17197
rect -28972 17163 -28938 17197
rect -28892 17163 -28858 17197
rect -28812 17163 -28778 17197
rect -28732 17163 -28698 17197
rect -28652 17163 -28618 17197
rect -28572 17163 -28538 17197
rect -28492 17163 -28458 17197
rect -28412 17163 -28378 17197
rect -28332 17163 -28298 17197
rect -28252 17163 -28218 17197
rect -28172 17163 -28138 17197
rect -28092 17163 -28058 17197
rect -28012 17163 -27978 17197
rect -27932 17163 -27898 17197
rect -27852 17163 -27818 17197
rect -27772 17163 -27738 17197
rect -27692 17163 -27658 17197
rect -27612 17163 -27578 17197
rect -27532 17163 -27498 17197
rect -27452 17163 -27418 17197
rect -27372 17163 -27338 17197
rect -27292 17163 -27258 17197
rect -27212 17163 -27178 17197
rect -27132 17163 -27098 17197
rect -27052 17163 -27018 17197
rect -26972 17163 -26938 17197
rect -26892 17163 -26858 17197
rect -26812 17163 -26778 17197
rect -26732 17163 -26698 17197
rect -26652 17163 -26618 17197
rect -26572 17163 -26538 17197
rect -26492 17163 -26458 17197
rect -26412 17163 -26378 17197
rect -26332 17163 -26298 17197
rect -26252 17163 -26218 17197
rect -26172 17163 -26138 17197
rect -26092 17163 -26058 17197
rect -26012 17163 -25978 17197
rect -25932 17163 -25898 17197
rect -25852 17163 -25818 17197
rect -25772 17163 -25738 17197
rect -25692 17163 -25658 17197
rect -25612 17163 -25578 17197
rect -25532 17163 -25498 17197
rect -25452 17163 -25418 17197
rect -25372 17163 -25338 17197
rect -25292 17163 -25258 17197
rect -25212 17163 -25178 17197
rect -25132 17163 -25098 17197
rect -25052 17163 -25018 17197
rect -24972 17163 -24938 17197
rect -24891 17163 -24857 17197
rect -24811 17163 -24777 17197
rect -24731 17163 -24697 17197
rect -24651 17163 -24617 17197
rect -24571 17163 -24537 17197
rect -24491 17163 -24457 17197
rect -24411 17163 -24377 17197
rect -24331 17163 -24297 17197
rect -24251 17163 -24217 17197
rect -24171 17163 -24137 17197
rect -24091 17163 -24057 17197
rect -24011 17163 -23977 17197
rect -23931 17163 -23897 17197
rect -23851 17163 -23817 17197
rect -23771 17163 -23737 17197
rect -23691 17163 -23657 17197
rect -23611 17163 -23577 17197
rect -23531 17163 -23497 17197
rect -23451 17163 -23417 17197
rect -23371 17163 -23337 17197
rect -23291 17163 -23257 17197
rect -23211 17163 -23177 17197
rect -23131 17163 -23097 17197
rect -23051 17163 -23017 17197
rect -22971 17163 -22937 17197
rect -22891 17163 -22857 17197
rect -22811 17163 -22777 17197
rect -22731 17163 -22697 17197
rect -22651 17163 -22617 17197
rect -22571 17163 -22537 17197
rect -22491 17163 -22457 17197
rect -22411 17163 -22377 17197
rect -22331 17163 -22297 17197
rect -22251 17163 -22217 17197
rect -22171 17163 -22137 17197
rect -22091 17163 -22057 17197
rect -22011 17163 -21977 17197
rect -21931 17163 -21897 17197
rect -21851 17163 -21817 17197
rect -21771 17163 -21737 17197
rect -21691 17163 -21657 17197
rect -21611 17163 -21577 17197
rect -21531 17163 -21497 17197
rect -21451 17163 -21417 17197
rect -21371 17163 -21337 17197
rect -21291 17163 -21257 17197
rect -21211 17163 -21177 17197
rect -21131 17163 -21097 17197
rect -21051 17163 -21017 17197
rect -20971 17163 -20937 17197
rect -20891 17163 -20857 17197
rect -20811 17163 -20777 17197
rect -20731 17163 -20697 17197
rect -20651 17163 -20617 17197
rect -20571 17163 -20537 17197
rect -20491 17163 -20457 17197
rect -20411 17163 -20377 17197
rect -20331 17163 -20297 17197
rect -20251 17163 -20217 17197
rect -20171 17163 -20137 17197
rect -20091 17163 -20057 17197
rect -20011 17163 -19977 17197
rect -19931 17163 -19897 17197
rect -19851 17163 -19817 17197
rect -19771 17163 -19737 17197
rect -19691 17163 -19657 17197
rect -19611 17163 -19577 17197
rect -19531 17163 -19497 17197
rect -19451 17163 -19417 17197
rect -19371 17163 -19337 17197
rect -19291 17163 -19257 17197
rect -19211 17163 -19177 17197
rect -19131 17163 -19097 17197
rect -19051 17163 -19017 17197
rect -18971 17163 -18937 17197
rect -18891 17163 -18857 17197
rect -18811 17163 -18777 17197
rect -18731 17163 -18697 17197
rect -18651 17163 -18617 17197
rect -18571 17163 -18537 17197
rect -18491 17163 -18457 17197
rect -18411 17163 -18377 17197
rect -18331 17163 -18297 17197
rect -18251 17163 -18217 17197
rect -18171 17163 -18137 17197
rect -18091 17163 -18057 17197
rect -18011 17163 -17977 17197
rect -17931 17163 -17897 17197
rect -17851 17163 -17817 17197
rect -17771 17163 -17737 17197
rect -17691 17163 -17657 17197
rect -17611 17163 -17577 17197
rect -17531 17163 -17497 17197
rect -17451 17163 -17417 17197
rect -17371 17163 -17337 17197
rect -17291 17163 -17257 17197
rect -17211 17163 -17177 17197
rect -17131 17163 -17097 17197
rect -17051 17163 -17017 17197
rect -16971 17163 -16937 17197
rect -16891 17163 -16857 17197
rect -16811 17163 -16777 17197
rect -16731 17163 -16697 17197
rect -16651 17163 -16617 17197
rect -16571 17163 -16537 17197
rect -16491 17163 -16457 17197
rect -16411 17163 -16377 17197
rect -16331 17163 -16297 17197
rect -16251 17163 -16217 17197
rect -16171 17163 -16137 17197
rect -16091 17163 -16057 17197
rect -16011 17163 -15977 17197
rect -15931 17163 -15897 17197
rect -15851 17163 -15817 17197
rect -15771 17163 -15737 17197
rect -15691 17163 -15657 17197
rect -15611 17163 -15577 17197
rect -15531 17163 -15497 17197
rect -15451 17163 -15417 17197
rect -15371 17163 -15337 17197
rect -15291 17163 -15257 17197
rect -15211 17163 -15177 17197
rect -15131 17163 -15097 17197
rect -15051 17163 -15017 17197
rect -14971 17163 -14937 17197
rect -14891 17163 -14857 17197
rect -14811 17163 -14777 17197
rect -14731 17163 -14697 17197
rect -14651 17163 -14617 17197
rect -14571 17163 -14537 17197
rect -14491 17163 -14457 17197
rect -14411 17163 -14377 17197
rect -14331 17163 -14297 17197
rect -14251 17163 -14217 17197
rect -14171 17163 -14137 17197
rect -14091 17163 -14057 17197
rect -14011 17163 -13977 17197
rect -13931 17163 -13897 17197
rect -13851 17163 -13817 17197
rect -13771 17163 -13737 17197
rect -13691 17163 -13657 17197
rect -13611 17163 -13577 17197
rect -13531 17163 -13497 17197
rect -13451 17163 -13417 17197
rect -13371 17163 -13337 17197
rect -13291 17163 -13257 17197
rect -13211 17163 -13177 17197
rect -13131 17163 -13097 17197
rect -13051 17163 -13017 17197
rect -12971 17163 -12937 17197
rect -12891 17163 -12857 17197
rect -12811 17163 -12777 17197
rect -12731 17163 -12697 17197
rect -12651 17163 -12617 17197
rect -12571 17163 -12537 17197
rect -12491 17163 -12457 17197
rect -12411 17163 -12377 17197
rect -12331 17163 -12297 17197
rect -12251 17163 -12217 17197
rect -12171 17163 -12137 17197
rect -12091 17163 -12057 17197
rect -12011 17163 -11977 17197
rect -11930 17163 -11896 17197
rect -11850 17163 -11816 17197
rect -11770 17163 -11736 17197
rect -11690 17163 -11656 17197
rect -11610 17163 -11576 17197
rect -11530 17163 -11496 17197
rect -11450 17163 -11416 17197
rect -11370 17163 -11336 17197
rect -11290 17163 -11256 17197
rect -11210 17163 -11176 17197
rect -11130 17163 -11096 17197
rect -11050 17163 -11016 17197
rect -10970 17163 -10936 17197
rect -10890 17163 -10856 17197
rect -10810 17163 -10776 17197
rect -10730 17163 -10696 17197
rect -10650 17163 -10616 17197
rect -10570 17163 -10536 17197
rect -10490 17163 -10456 17197
rect -10410 17163 -10376 17197
rect -10330 17163 -10296 17197
rect -10250 17163 -10216 17197
rect -10170 17163 -10136 17197
rect -10090 17163 -10056 17197
rect -10010 17163 -9976 17197
rect -9930 17163 -9896 17197
rect -9850 17163 -9816 17197
rect -9770 17163 -9736 17197
rect -9690 17163 -9656 17197
rect -9610 17163 -9576 17197
rect -9530 17163 -9496 17197
rect -9450 17163 -9416 17197
rect -9370 17163 -9336 17197
rect -9290 17163 -9256 17197
rect -9210 17163 -9176 17197
rect -9130 17163 -9096 17197
rect -9050 17163 -9016 17197
rect -8970 17163 -8936 17197
rect -8890 17163 -8856 17197
rect -8810 17163 -8776 17197
rect -8730 17163 -8696 17197
rect -8650 17163 -8616 17197
rect -8570 17163 -8536 17197
rect -8490 17163 -8456 17197
rect -8410 17163 -8376 17197
rect -8330 17163 -8296 17197
rect -8250 17163 -8216 17197
rect -8170 17163 -8136 17197
rect -8090 17163 -8056 17197
rect -8010 17163 -7976 17197
rect -7930 17163 -7896 17197
rect -7850 17163 -7816 17197
rect -7770 17163 -7736 17197
rect -7690 17163 -7656 17197
rect -7610 17163 -7576 17197
rect -7530 17163 -7496 17197
rect -7450 17163 -7416 17197
rect -7370 17163 -7336 17197
rect -7290 17163 -7256 17197
rect -7210 17163 -7176 17197
rect -7130 17163 -7096 17197
rect -7050 17163 -7016 17197
rect -6970 17163 -6936 17197
rect -6890 17163 -6856 17197
rect -6810 17163 -6776 17197
rect -6730 17163 -6696 17197
rect -6650 17163 -6616 17197
rect -6570 17163 -6536 17197
rect -6490 17163 -6456 17197
rect -6410 17163 -6376 17197
rect -6330 17163 -6296 17197
rect -6250 17163 -6216 17197
rect -6170 17163 -6136 17197
rect -6090 17163 -6056 17197
rect -6010 17163 -5976 17197
rect -5930 17163 -5896 17197
rect -5850 17163 -5816 17197
rect -5770 17163 -5736 17197
rect -5690 17163 -5656 17197
rect -5610 17163 -5576 17197
rect -5530 17163 -5496 17197
rect -5450 17163 -5416 17197
rect -5370 17163 -5336 17197
rect -5290 17163 -5256 17197
rect -5210 17163 -5176 17197
rect -5130 17163 -5096 17197
rect -5050 17163 -5016 17197
rect -4970 17163 -4936 17197
rect -4890 17163 -4856 17197
rect -4810 17163 -4776 17197
rect -4730 17163 -4696 17197
rect -4650 17163 -4616 17197
rect -4570 17163 -4536 17197
rect -4490 17163 -4456 17197
rect -4410 17163 -4376 17197
rect -4330 17163 -4296 17197
rect -4250 17163 -4216 17197
rect -4170 17163 -4136 17197
rect -4090 17163 -4056 17197
rect -4010 17163 -3976 17197
rect -3930 17163 -3896 17197
rect -3850 17163 -3816 17197
rect -3770 17163 -3736 17197
rect -3690 17163 -3656 17197
rect -3610 17163 -3576 17197
rect -3530 17163 -3496 17197
rect -3450 17163 -3416 17197
rect -3370 17163 -3336 17197
rect -1929 17163 -1895 17197
rect -1849 17163 -1815 17197
rect -1769 17163 -1735 17197
rect -1689 17163 -1655 17197
rect -1609 17163 -1575 17197
rect -1529 17163 -1495 17197
rect -1449 17163 -1415 17197
rect -1369 17163 -1335 17197
rect -1289 17163 -1255 17197
rect -1209 17163 -1175 17197
rect -1129 17163 -1095 17197
rect -1049 17163 -1015 17197
rect -969 17163 -935 17197
rect -889 17163 -855 17197
rect -809 17163 -775 17197
rect -729 17163 -695 17197
rect -649 17163 -615 17197
rect -569 17163 -535 17197
rect -489 17163 -455 17197
rect -409 17163 -375 17197
rect -329 17163 -295 17197
rect -249 17163 -215 17197
rect -169 17163 -135 17197
rect -89 17163 -55 17197
rect -9 17163 25 17197
rect 71 17163 105 17197
rect 151 17163 185 17197
rect 231 17163 265 17197
rect 311 17163 345 17197
rect 391 17163 425 17197
rect 471 17163 505 17197
rect 551 17163 585 17197
rect 631 17163 665 17197
rect 711 17163 745 17197
rect 791 17163 825 17197
rect 871 17163 905 17197
rect 951 17163 985 17197
rect 1031 17163 1065 17197
rect 1111 17163 1145 17197
rect 1191 17163 1225 17197
rect 1271 17163 1305 17197
rect 1351 17163 1385 17197
rect 1431 17163 1465 17197
rect 1511 17163 1545 17197
rect 1591 17163 1625 17197
rect 1671 17163 1705 17197
rect 1751 17163 1785 17197
rect 1831 17163 1865 17197
rect 1911 17163 1945 17197
rect 1991 17163 2025 17197
rect 2071 17163 2105 17197
rect 2151 17163 2185 17197
rect 2231 17163 2265 17197
rect 2311 17163 2345 17197
rect 3790 17163 3824 17197
rect 3870 17163 3904 17197
rect 3950 17163 3984 17197
rect 4030 17163 4064 17197
rect 4110 17163 4144 17197
rect 4190 17163 4224 17197
rect 4270 17163 4304 17197
rect 4350 17163 4384 17197
rect 4430 17163 4464 17197
rect 4510 17163 4544 17197
rect 4590 17163 4624 17197
rect 4670 17163 4704 17197
rect 4750 17163 4784 17197
rect 4830 17163 4864 17197
rect 4910 17163 4944 17197
rect 4990 17163 5024 17197
rect 5070 17163 5104 17197
rect 5150 17163 5184 17197
rect 5230 17163 5264 17197
rect 5310 17163 5344 17197
rect 5390 17163 5424 17197
rect 5470 17163 5504 17197
rect 5550 17163 5584 17197
rect 5630 17163 5664 17197
rect 5710 17163 5744 17197
rect 5790 17163 5824 17197
rect 5870 17163 5904 17197
rect 5950 17163 5984 17197
rect 6030 17163 6064 17197
rect 6110 17163 6144 17197
rect 6190 17163 6224 17197
rect 6270 17163 6304 17197
rect 6350 17163 6384 17197
rect 6430 17163 6464 17197
rect 6510 17163 6544 17197
rect 6590 17163 6624 17197
rect 6670 17163 6704 17197
rect 6750 17163 6784 17197
rect 6830 17163 6864 17197
rect 6910 17163 6944 17197
rect 6990 17163 7024 17197
rect 7070 17163 7104 17197
rect 7150 17163 7184 17197
rect 7230 17163 7264 17197
rect 7310 17163 7344 17197
rect 7390 17163 7424 17197
rect 7470 17163 7504 17197
rect 7550 17163 7584 17197
rect 7630 17163 7664 17197
rect 7710 17163 7744 17197
rect 7790 17163 7824 17197
rect 7870 17163 7904 17197
rect 7950 17163 7984 17197
rect 8030 17163 8064 17197
rect 8110 17163 8144 17197
rect 8190 17163 8224 17197
rect 8270 17163 8304 17197
rect 8350 17163 8384 17197
rect 8430 17163 8464 17197
rect 8510 17163 8544 17197
rect 8590 17163 8624 17197
rect 8670 17163 8704 17197
rect 8750 17163 8784 17197
rect 8830 17163 8864 17197
rect 8910 17163 8944 17197
rect 8990 17163 9024 17197
rect 9070 17163 9104 17197
rect 9150 17163 9184 17197
rect 9230 17163 9264 17197
rect 9310 17163 9344 17197
rect 9390 17163 9424 17197
rect 9470 17163 9504 17197
rect 9550 17163 9584 17197
rect 9630 17163 9664 17197
rect 9710 17163 9744 17197
rect 9790 17163 9824 17197
rect 9870 17163 9904 17197
rect 9950 17163 9984 17197
rect 10030 17163 10064 17197
rect 10110 17163 10144 17197
rect 10190 17163 10224 17197
rect 10270 17163 10304 17197
rect 10350 17163 10384 17197
rect 10430 17163 10464 17197
rect 10510 17163 10544 17197
rect 10590 17163 10624 17197
rect 10670 17163 10704 17197
rect 10750 17163 10784 17197
rect 10830 17163 10864 17197
rect 10910 17163 10944 17197
rect 10990 17163 11024 17197
rect 11070 17163 11104 17197
rect 11150 17163 11184 17197
rect 11230 17163 11264 17197
rect 11310 17163 11344 17197
rect 11390 17163 11424 17197
rect 11470 17163 11504 17197
rect 11550 17163 11584 17197
rect 11630 17163 11664 17197
rect 11710 17163 11744 17197
rect 11790 17163 11824 17197
rect 11870 17163 11904 17197
rect 11950 17163 11984 17197
rect 12030 17163 12064 17197
rect 12110 17163 12144 17197
rect 12190 17163 12224 17197
rect 12270 17163 12304 17197
rect 12350 17163 12384 17197
rect 12430 17163 12464 17197
rect 12510 17163 12544 17197
rect 12590 17163 12624 17197
rect 12670 17163 12704 17197
rect 12750 17163 12784 17197
rect 12830 17163 12864 17197
rect 12910 17163 12944 17197
rect 12990 17163 13024 17197
rect 13070 17163 13104 17197
rect 13150 17163 13184 17197
rect 13230 17163 13264 17197
rect 13310 17163 13344 17197
rect 13390 17163 13424 17197
rect 13470 17163 13504 17197
rect 13550 17163 13584 17197
rect 13630 17163 13664 17197
rect 13710 17163 13744 17197
rect 13790 17163 13824 17197
rect 13870 17163 13904 17197
rect 13950 17163 13984 17197
rect 14030 17163 14064 17197
rect 14110 17163 14144 17197
rect 14190 17163 14224 17197
rect 14270 17163 14304 17197
rect 14350 17163 14384 17197
rect 14430 17163 14464 17197
rect 14510 17163 14544 17197
rect 14590 17163 14624 17197
rect 14670 17163 14704 17197
rect 14750 17163 14784 17197
rect 14830 17163 14864 17197
rect 14910 17163 14944 17197
rect 14990 17163 15024 17197
rect 15070 17163 15104 17197
rect 15150 17163 15184 17197
rect 15230 17163 15264 17197
rect 15310 17163 15344 17197
rect 15390 17163 15424 17197
rect 15470 17163 15504 17197
rect 15550 17163 15584 17197
rect 15630 17163 15664 17197
rect 15710 17163 15744 17197
rect 15790 17163 15824 17197
rect 15870 17163 15904 17197
rect 15950 17163 15984 17197
rect 16030 17163 16064 17197
rect 16110 17163 16144 17197
rect 16190 17163 16224 17197
rect 16270 17163 16304 17197
rect 16350 17163 16384 17197
rect 16430 17163 16464 17197
rect 16510 17163 16544 17197
rect 16590 17163 16624 17197
rect 16670 17163 16704 17197
rect 16751 17163 16785 17197
rect 16831 17163 16865 17197
rect 16911 17163 16945 17197
rect 16991 17163 17025 17197
rect 17071 17163 17105 17197
rect 17151 17163 17185 17197
rect 17231 17163 17265 17197
rect 17311 17163 17345 17197
rect 17391 17163 17425 17197
rect 17471 17163 17505 17197
rect 17551 17163 17585 17197
rect 17631 17163 17665 17197
rect 17711 17163 17745 17197
rect 17791 17163 17825 17197
rect 17871 17163 17905 17197
rect 17951 17163 17985 17197
rect 18031 17163 18065 17197
rect 18111 17163 18145 17197
rect 18191 17163 18225 17197
rect 18271 17163 18305 17197
rect 18351 17163 18385 17197
rect 18431 17163 18465 17197
rect 18511 17163 18545 17197
rect 18591 17163 18625 17197
rect 18671 17163 18705 17197
rect 18751 17163 18785 17197
rect 18831 17163 18865 17197
rect 18911 17163 18945 17197
rect 18991 17163 19025 17197
rect 19071 17163 19105 17197
rect 19151 17163 19185 17197
rect 19231 17163 19265 17197
rect 19311 17163 19345 17197
rect 19391 17163 19425 17197
rect 19471 17163 19505 17197
rect 19551 17163 19585 17197
rect 19631 17163 19665 17197
rect 19711 17163 19745 17197
rect 19791 17163 19825 17197
rect 19871 17163 19905 17197
rect 19951 17163 19985 17197
rect 20031 17163 20065 17197
rect 20111 17163 20145 17197
rect 20191 17163 20225 17197
rect 20271 17163 20305 17197
rect 20351 17163 20385 17197
rect 20431 17163 20465 17197
rect 20511 17163 20545 17197
rect 20591 17163 20625 17197
rect 20671 17163 20705 17197
rect 20751 17163 20785 17197
rect 20831 17163 20865 17197
rect 20911 17163 20945 17197
rect 20991 17163 21025 17197
rect 21071 17163 21105 17197
rect 21151 17163 21185 17197
rect 21231 17163 21265 17197
rect 21311 17163 21345 17197
rect 21391 17163 21425 17197
rect 21471 17163 21505 17197
rect 21551 17163 21585 17197
rect 21631 17163 21665 17197
rect 21711 17163 21745 17197
rect 21791 17163 21825 17197
rect 21871 17163 21905 17197
rect 21951 17163 21985 17197
rect 22031 17163 22065 17197
rect 22111 17163 22145 17197
rect 22191 17163 22225 17197
rect 22271 17163 22305 17197
rect 22351 17163 22385 17197
rect 22431 17163 22465 17197
rect 22511 17163 22545 17197
rect 22591 17163 22625 17197
rect 22671 17163 22705 17197
rect 22751 17163 22785 17197
rect 22831 17163 22865 17197
rect 22911 17163 22945 17197
rect 22991 17163 23025 17197
rect 23071 17163 23105 17197
rect 23151 17163 23185 17197
rect 23231 17163 23265 17197
rect 23311 17163 23345 17197
rect 23391 17163 23425 17197
rect 23471 17163 23505 17197
rect 23551 17163 23585 17197
rect 23631 17163 23665 17197
rect 23711 17163 23745 17197
rect 23791 17163 23825 17197
rect 23871 17163 23905 17197
rect 23951 17163 23985 17197
rect 24031 17163 24065 17197
rect 24111 17163 24145 17197
rect 24191 17163 24225 17197
rect 24271 17163 24305 17197
rect 24351 17163 24385 17197
rect 24431 17163 24465 17197
rect 24511 17163 24545 17197
rect 24591 17163 24625 17197
rect 24671 17163 24705 17197
rect 24751 17163 24785 17197
rect 24831 17163 24865 17197
rect 24911 17163 24945 17197
rect 24991 17163 25025 17197
rect 25071 17163 25105 17197
rect 25151 17163 25185 17197
rect 25231 17163 25265 17197
rect 25311 17163 25345 17197
rect 25391 17163 25425 17197
rect 25471 17163 25505 17197
rect 25551 17163 25585 17197
rect 25631 17163 25665 17197
rect 25711 17163 25745 17197
rect 25791 17163 25825 17197
rect 25871 17163 25905 17197
rect 25951 17163 25985 17197
rect 26031 17163 26065 17197
rect 26111 17163 26145 17197
rect 26191 17163 26225 17197
rect 26271 17163 26305 17197
rect 26351 17163 26385 17197
rect 26431 17163 26465 17197
rect 26511 17163 26545 17197
rect 26591 17163 26625 17197
rect 26671 17163 26705 17197
rect 26751 17163 26785 17197
rect 26831 17163 26865 17197
rect 26911 17163 26945 17197
rect 26991 17163 27025 17197
rect 27071 17163 27105 17197
rect 27151 17163 27185 17197
rect 27231 17163 27265 17197
rect 27311 17163 27345 17197
rect 27391 17163 27425 17197
rect 27471 17163 27505 17197
rect 27551 17163 27585 17197
rect 27631 17163 27665 17197
rect 27711 17163 27745 17197
rect 27791 17163 27825 17197
rect 27871 17163 27905 17197
rect 27951 17163 27985 17197
rect 28031 17163 28065 17197
rect 28111 17163 28145 17197
rect 28191 17163 28225 17197
rect 28271 17163 28305 17197
rect 28351 17163 28385 17197
rect 28431 17163 28465 17197
rect 28511 17163 28545 17197
rect 28591 17163 28625 17197
rect 28671 17163 28705 17197
rect 28751 17163 28785 17197
rect 28831 17163 28865 17197
rect 28911 17163 28945 17197
rect 28991 17163 29025 17197
rect 29071 17163 29105 17197
rect 29151 17163 29185 17197
rect 29231 17163 29265 17197
rect 29311 17163 29345 17197
rect 29391 17163 29425 17197
rect 29471 17163 29505 17197
rect 29551 17163 29585 17197
rect 29631 17163 29665 17197
rect 29711 17163 29745 17197
rect 29791 17163 29825 17197
rect 29871 17163 29905 17197
rect 29951 17163 29985 17197
rect 30031 17163 30065 17197
rect 30111 17163 30145 17197
rect 30191 17163 30225 17197
rect 30271 17163 30305 17197
rect 30351 17163 30385 17197
rect 30431 17163 30465 17197
rect 30511 17163 30545 17197
rect 30591 17163 30625 17197
rect 30671 17163 30705 17197
rect 30751 17163 30785 17197
rect 30831 17163 30865 17197
rect 30911 17163 30945 17197
rect 30991 17163 31025 17197
rect 31071 17163 31105 17197
rect 31151 17163 31185 17197
rect 31231 17163 31265 17197
rect 31311 17163 31345 17197
rect 31391 17163 31425 17197
rect 31471 17163 31505 17197
rect 31551 17163 31585 17197
rect 31631 17163 31665 17197
rect 31711 17163 31745 17197
rect 31791 17163 31825 17197
rect 31871 17163 31905 17197
rect 31951 17163 31985 17197
rect 32031 17163 32065 17197
rect 32111 17163 32145 17197
rect 32191 17163 32225 17197
rect 32271 17163 32305 17197
rect 32351 17163 32385 17197
rect 32431 17163 32465 17197
rect 32511 17163 32545 17197
rect 32591 17163 32625 17197
rect 32671 17163 32705 17197
rect 32751 17163 32785 17197
rect 32831 17163 32865 17197
rect 32911 17163 32945 17197
rect 32991 17163 33025 17197
rect 33071 17163 33105 17197
rect 33151 17163 33185 17197
rect 33231 17163 33265 17197
rect 33311 17163 33345 17197
rect 33391 17163 33425 17197
rect 33471 17163 33505 17197
rect 33551 17163 33585 17197
rect 33631 17163 33665 17197
rect 33711 17163 33745 17197
rect 33791 17163 33825 17197
rect 33871 17163 33905 17197
rect 33951 17163 33985 17197
rect 34031 17163 34065 17197
rect 34111 17163 34145 17197
rect 34191 17163 34225 17197
rect 34271 17163 34305 17197
rect 34351 17163 34385 17197
rect 34431 17163 34465 17197
rect 34511 17163 34545 17197
rect 34591 17163 34625 17197
rect 34671 17163 34705 17197
rect 34751 17163 34785 17197
rect 34831 17163 34865 17197
rect 34911 17163 34945 17197
rect 34991 17163 35025 17197
rect 35071 17163 35105 17197
rect 35151 17163 35185 17197
rect 35231 17163 35265 17197
rect 35311 17163 35345 17197
rect 35391 17163 35425 17197
rect 35471 17163 35505 17197
rect 35551 17163 35585 17197
rect 35631 17163 35665 17197
rect 35711 17163 35745 17197
rect 35791 17163 35825 17197
rect 35871 17163 35905 17197
rect 35951 17163 35985 17197
rect 36031 17163 36065 17197
rect 36111 17163 36145 17197
rect 36191 17163 36225 17197
rect 36271 17163 36305 17197
rect 36351 17163 36385 17197
rect 36431 17163 36465 17197
rect 36511 17163 36545 17197
rect 36591 17163 36625 17197
rect 36671 17163 36705 17197
rect 36751 17163 36785 17197
rect 36831 17163 36865 17197
rect 36911 17163 36945 17197
rect 36991 17163 37025 17197
rect 37071 17163 37105 17197
rect 37151 17163 37185 17197
rect 37231 17163 37265 17197
rect 37311 17163 37345 17197
rect 37391 17163 37425 17197
rect 37471 17163 37505 17197
rect 37551 17163 37585 17197
rect 37631 17163 37665 17197
rect 37711 17163 37745 17197
rect 37791 17163 37825 17197
rect 37871 17163 37905 17197
rect 37951 17163 37985 17197
rect 38031 17163 38065 17197
rect 38111 17163 38145 17197
rect 38191 17163 38225 17197
rect 38271 17163 38305 17197
rect -37852 9304 -37818 9338
rect -37772 9304 -37738 9338
rect -37692 9304 -37658 9338
rect -37612 9304 -37578 9338
rect -37532 9304 -37498 9338
rect -37452 9304 -37418 9338
rect -37372 9304 -37338 9338
rect -37292 9304 -37258 9338
rect -37212 9304 -37178 9338
rect -37132 9304 -37098 9338
rect -37052 9304 -37018 9338
rect -36972 9304 -36938 9338
rect -36892 9304 -36858 9338
rect -36812 9304 -36778 9338
rect -36732 9304 -36698 9338
rect -36652 9304 -36618 9338
rect -36572 9304 -36538 9338
rect -36492 9304 -36458 9338
rect -36412 9304 -36378 9338
rect -36332 9304 -36298 9338
rect -36252 9304 -36218 9338
rect -36172 9304 -36138 9338
rect -36092 9304 -36058 9338
rect -36012 9304 -35978 9338
rect -35932 9304 -35898 9338
rect -35852 9304 -35818 9338
rect -35772 9304 -35738 9338
rect -35692 9304 -35658 9338
rect -35612 9304 -35578 9338
rect -35532 9304 -35498 9338
rect -35452 9304 -35418 9338
rect -35372 9304 -35338 9338
rect -35292 9304 -35258 9338
rect -35212 9304 -35178 9338
rect -35132 9304 -35098 9338
rect -35052 9304 -35018 9338
rect -34972 9304 -34938 9338
rect -34892 9304 -34858 9338
rect -34812 9304 -34778 9338
rect -34732 9304 -34698 9338
rect -34652 9304 -34618 9338
rect -34572 9304 -34538 9338
rect -34492 9304 -34458 9338
rect -34412 9304 -34378 9338
rect -34332 9304 -34298 9338
rect -34252 9304 -34218 9338
rect -34172 9304 -34138 9338
rect -34092 9304 -34058 9338
rect -34012 9304 -33978 9338
rect -33932 9304 -33898 9338
rect -33852 9304 -33818 9338
rect -33772 9304 -33738 9338
rect -33692 9304 -33658 9338
rect -33612 9304 -33578 9338
rect -33532 9304 -33498 9338
rect -33452 9304 -33418 9338
rect -33372 9304 -33338 9338
rect -33292 9304 -33258 9338
rect -33212 9304 -33178 9338
rect -33132 9304 -33098 9338
rect -33052 9304 -33018 9338
rect -32972 9304 -32938 9338
rect -32892 9304 -32858 9338
rect -32812 9304 -32778 9338
rect -32732 9304 -32698 9338
rect -32652 9304 -32618 9338
rect -32572 9304 -32538 9338
rect -32492 9304 -32458 9338
rect -32412 9304 -32378 9338
rect -32332 9304 -32298 9338
rect -32252 9304 -32218 9338
rect -32172 9304 -32138 9338
rect -32092 9304 -32058 9338
rect -32012 9304 -31978 9338
rect -31932 9304 -31898 9338
rect -31852 9304 -31818 9338
rect -31772 9304 -31738 9338
rect -31692 9304 -31658 9338
rect -31612 9304 -31578 9338
rect -31532 9304 -31498 9338
rect -31452 9304 -31418 9338
rect -31372 9304 -31338 9338
rect -31292 9304 -31258 9338
rect -31212 9304 -31178 9338
rect -31132 9304 -31098 9338
rect -31052 9304 -31018 9338
rect -30972 9304 -30938 9338
rect -30892 9304 -30858 9338
rect -30812 9304 -30778 9338
rect -30732 9304 -30698 9338
rect -30652 9304 -30618 9338
rect -30572 9304 -30538 9338
rect -30492 9304 -30458 9338
rect -30412 9304 -30378 9338
rect -30332 9304 -30298 9338
rect -30252 9304 -30218 9338
rect -30172 9304 -30138 9338
rect -30092 9304 -30058 9338
rect -30012 9304 -29978 9338
rect -29932 9304 -29898 9338
rect -29852 9304 -29818 9338
rect -29772 9304 -29738 9338
rect -29692 9304 -29658 9338
rect -29612 9304 -29578 9338
rect -29532 9304 -29498 9338
rect -29452 9304 -29418 9338
rect -29372 9304 -29338 9338
rect -29292 9304 -29258 9338
rect -29212 9304 -29178 9338
rect -29132 9304 -29098 9338
rect -29052 9304 -29018 9338
rect -28972 9304 -28938 9338
rect -28892 9304 -28858 9338
rect -28812 9304 -28778 9338
rect -28732 9304 -28698 9338
rect -28652 9304 -28618 9338
rect -28572 9304 -28538 9338
rect -28492 9304 -28458 9338
rect -28412 9304 -28378 9338
rect -28332 9304 -28298 9338
rect -28252 9304 -28218 9338
rect -28172 9304 -28138 9338
rect -28092 9304 -28058 9338
rect -28012 9304 -27978 9338
rect -27932 9304 -27898 9338
rect -27852 9304 -27818 9338
rect -27772 9304 -27738 9338
rect -27692 9304 -27658 9338
rect -27612 9304 -27578 9338
rect -27532 9304 -27498 9338
rect -27452 9304 -27418 9338
rect -27372 9304 -27338 9338
rect -27292 9304 -27258 9338
rect -27212 9304 -27178 9338
rect -27132 9304 -27098 9338
rect -27052 9304 -27018 9338
rect -26972 9304 -26938 9338
rect -26892 9304 -26858 9338
rect -26812 9304 -26778 9338
rect -26732 9304 -26698 9338
rect -26652 9304 -26618 9338
rect -26572 9304 -26538 9338
rect -26492 9304 -26458 9338
rect -26412 9304 -26378 9338
rect -26332 9304 -26298 9338
rect -26252 9304 -26218 9338
rect -26172 9304 -26138 9338
rect -26092 9304 -26058 9338
rect -26012 9304 -25978 9338
rect -25932 9304 -25898 9338
rect -25852 9304 -25818 9338
rect -25772 9304 -25738 9338
rect -25692 9304 -25658 9338
rect -25612 9304 -25578 9338
rect -25532 9304 -25498 9338
rect -25452 9304 -25418 9338
rect -25372 9304 -25338 9338
rect -25292 9304 -25258 9338
rect -25212 9304 -25178 9338
rect -25132 9304 -25098 9338
rect -25052 9304 -25018 9338
rect -24972 9304 -24938 9338
rect -24891 9304 -24857 9338
rect -24811 9304 -24777 9338
rect -24731 9304 -24697 9338
rect -24651 9304 -24617 9338
rect -24571 9304 -24537 9338
rect -24491 9304 -24457 9338
rect -24411 9304 -24377 9338
rect -24331 9304 -24297 9338
rect -24251 9304 -24217 9338
rect -24171 9304 -24137 9338
rect -24091 9304 -24057 9338
rect -24011 9304 -23977 9338
rect -23931 9304 -23897 9338
rect -23851 9304 -23817 9338
rect -23771 9304 -23737 9338
rect -23691 9304 -23657 9338
rect -23611 9304 -23577 9338
rect -23531 9304 -23497 9338
rect -23451 9304 -23417 9338
rect -23371 9304 -23337 9338
rect -23291 9304 -23257 9338
rect -23211 9304 -23177 9338
rect -23131 9304 -23097 9338
rect -23051 9304 -23017 9338
rect -22971 9304 -22937 9338
rect -22891 9304 -22857 9338
rect -22811 9304 -22777 9338
rect -22731 9304 -22697 9338
rect -22651 9304 -22617 9338
rect -22571 9304 -22537 9338
rect -22491 9304 -22457 9338
rect -22411 9304 -22377 9338
rect -22331 9304 -22297 9338
rect -22251 9304 -22217 9338
rect -22171 9304 -22137 9338
rect -22091 9304 -22057 9338
rect -22011 9304 -21977 9338
rect -21931 9304 -21897 9338
rect -21851 9304 -21817 9338
rect -21771 9304 -21737 9338
rect -21691 9304 -21657 9338
rect -21611 9304 -21577 9338
rect -21531 9304 -21497 9338
rect -21451 9304 -21417 9338
rect -21371 9304 -21337 9338
rect -21291 9304 -21257 9338
rect -21211 9304 -21177 9338
rect -21131 9304 -21097 9338
rect -21051 9304 -21017 9338
rect -20971 9304 -20937 9338
rect -20891 9304 -20857 9338
rect -20811 9304 -20777 9338
rect -20731 9304 -20697 9338
rect -20651 9304 -20617 9338
rect -20571 9304 -20537 9338
rect -20491 9304 -20457 9338
rect -20411 9304 -20377 9338
rect -20331 9304 -20297 9338
rect -20251 9304 -20217 9338
rect -20171 9304 -20137 9338
rect -20091 9304 -20057 9338
rect -20011 9304 -19977 9338
rect -19931 9304 -19897 9338
rect -19851 9304 -19817 9338
rect -19771 9304 -19737 9338
rect -19691 9304 -19657 9338
rect -19611 9304 -19577 9338
rect -19531 9304 -19497 9338
rect -19451 9304 -19417 9338
rect -19371 9304 -19337 9338
rect -19291 9304 -19257 9338
rect -19211 9304 -19177 9338
rect -19131 9304 -19097 9338
rect -19051 9304 -19017 9338
rect -18971 9304 -18937 9338
rect -18891 9304 -18857 9338
rect -18811 9304 -18777 9338
rect -18731 9304 -18697 9338
rect -18651 9304 -18617 9338
rect -18571 9304 -18537 9338
rect -18491 9304 -18457 9338
rect -18411 9304 -18377 9338
rect -18331 9304 -18297 9338
rect -18251 9304 -18217 9338
rect -18171 9304 -18137 9338
rect -18091 9304 -18057 9338
rect -18011 9304 -17977 9338
rect -17931 9304 -17897 9338
rect -17851 9304 -17817 9338
rect -17771 9304 -17737 9338
rect -17691 9304 -17657 9338
rect -17611 9304 -17577 9338
rect -17531 9304 -17497 9338
rect -17451 9304 -17417 9338
rect -17371 9304 -17337 9338
rect -17291 9304 -17257 9338
rect -17211 9304 -17177 9338
rect -17131 9304 -17097 9338
rect -17051 9304 -17017 9338
rect -16971 9304 -16937 9338
rect -16891 9304 -16857 9338
rect -16811 9304 -16777 9338
rect -16731 9304 -16697 9338
rect -16651 9304 -16617 9338
rect -16571 9304 -16537 9338
rect -16491 9304 -16457 9338
rect -16411 9304 -16377 9338
rect -16331 9304 -16297 9338
rect -16251 9304 -16217 9338
rect -16171 9304 -16137 9338
rect -16091 9304 -16057 9338
rect -16011 9304 -15977 9338
rect -15931 9304 -15897 9338
rect -15851 9304 -15817 9338
rect -15771 9304 -15737 9338
rect -15691 9304 -15657 9338
rect -15611 9304 -15577 9338
rect -15531 9304 -15497 9338
rect -15451 9304 -15417 9338
rect -15371 9304 -15337 9338
rect -15291 9304 -15257 9338
rect -15211 9304 -15177 9338
rect -15131 9304 -15097 9338
rect -15051 9304 -15017 9338
rect -14971 9304 -14937 9338
rect -14891 9304 -14857 9338
rect -14811 9304 -14777 9338
rect -14731 9304 -14697 9338
rect -14651 9304 -14617 9338
rect -14571 9304 -14537 9338
rect -14491 9304 -14457 9338
rect -14411 9304 -14377 9338
rect -14331 9304 -14297 9338
rect -14251 9304 -14217 9338
rect -14171 9304 -14137 9338
rect -14091 9304 -14057 9338
rect -14011 9304 -13977 9338
rect -13931 9304 -13897 9338
rect -13851 9304 -13817 9338
rect -13771 9304 -13737 9338
rect -13691 9304 -13657 9338
rect -13611 9304 -13577 9338
rect -13531 9304 -13497 9338
rect -13451 9304 -13417 9338
rect -13371 9304 -13337 9338
rect -13291 9304 -13257 9338
rect -13211 9304 -13177 9338
rect -13131 9304 -13097 9338
rect -13051 9304 -13017 9338
rect -12971 9304 -12937 9338
rect -12891 9304 -12857 9338
rect -12811 9304 -12777 9338
rect -12731 9304 -12697 9338
rect -12651 9304 -12617 9338
rect -12571 9304 -12537 9338
rect -12491 9304 -12457 9338
rect -12411 9304 -12377 9338
rect -12331 9304 -12297 9338
rect -12251 9304 -12217 9338
rect -12171 9304 -12137 9338
rect -12091 9304 -12057 9338
rect -12011 9304 -11977 9338
rect -11930 9304 -11896 9338
rect -11850 9304 -11816 9338
rect -11770 9304 -11736 9338
rect -11690 9304 -11656 9338
rect -11610 9304 -11576 9338
rect -11530 9304 -11496 9338
rect -11450 9304 -11416 9338
rect -11370 9304 -11336 9338
rect -11290 9304 -11256 9338
rect -11210 9304 -11176 9338
rect -11130 9304 -11096 9338
rect -11050 9304 -11016 9338
rect -10970 9304 -10936 9338
rect -10890 9304 -10856 9338
rect -10810 9304 -10776 9338
rect -10730 9304 -10696 9338
rect -10650 9304 -10616 9338
rect -10570 9304 -10536 9338
rect -10490 9304 -10456 9338
rect -10410 9304 -10376 9338
rect -10330 9304 -10296 9338
rect -10250 9304 -10216 9338
rect -10170 9304 -10136 9338
rect -10090 9304 -10056 9338
rect -10010 9304 -9976 9338
rect -9930 9304 -9896 9338
rect -9850 9304 -9816 9338
rect -9770 9304 -9736 9338
rect -9690 9304 -9656 9338
rect -9610 9304 -9576 9338
rect -9530 9304 -9496 9338
rect -9450 9304 -9416 9338
rect -9370 9304 -9336 9338
rect -9290 9304 -9256 9338
rect -9210 9304 -9176 9338
rect -9130 9304 -9096 9338
rect -9050 9304 -9016 9338
rect -8970 9304 -8936 9338
rect -8890 9304 -8856 9338
rect -8810 9304 -8776 9338
rect -8730 9304 -8696 9338
rect -8650 9304 -8616 9338
rect -8570 9304 -8536 9338
rect -8490 9304 -8456 9338
rect -8410 9304 -8376 9338
rect -8330 9304 -8296 9338
rect -8250 9304 -8216 9338
rect -8170 9304 -8136 9338
rect -8090 9304 -8056 9338
rect -8010 9304 -7976 9338
rect -7930 9304 -7896 9338
rect -7850 9304 -7816 9338
rect -7770 9304 -7736 9338
rect -7690 9304 -7656 9338
rect -7610 9304 -7576 9338
rect -7530 9304 -7496 9338
rect -7450 9304 -7416 9338
rect -7370 9304 -7336 9338
rect -7290 9304 -7256 9338
rect -7210 9304 -7176 9338
rect -7130 9304 -7096 9338
rect -7050 9304 -7016 9338
rect -6970 9304 -6936 9338
rect -6890 9304 -6856 9338
rect -6810 9304 -6776 9338
rect -6730 9304 -6696 9338
rect -6650 9304 -6616 9338
rect -6570 9304 -6536 9338
rect -6490 9304 -6456 9338
rect -6410 9304 -6376 9338
rect -6330 9304 -6296 9338
rect -6250 9304 -6216 9338
rect -6170 9304 -6136 9338
rect -6090 9304 -6056 9338
rect -6010 9304 -5976 9338
rect -5930 9304 -5896 9338
rect -5850 9304 -5816 9338
rect -5770 9304 -5736 9338
rect -5690 9304 -5656 9338
rect -5610 9304 -5576 9338
rect -5530 9304 -5496 9338
rect -5450 9304 -5416 9338
rect -5370 9304 -5336 9338
rect -5290 9304 -5256 9338
rect -5210 9304 -5176 9338
rect -5130 9304 -5096 9338
rect -5050 9304 -5016 9338
rect -4970 9304 -4936 9338
rect -4890 9304 -4856 9338
rect -4810 9304 -4776 9338
rect -4730 9304 -4696 9338
rect -4650 9304 -4616 9338
rect -4570 9304 -4536 9338
rect -4490 9304 -4456 9338
rect -4410 9304 -4376 9338
rect -4330 9304 -4296 9338
rect -4250 9304 -4216 9338
rect -4170 9304 -4136 9338
rect -4090 9304 -4056 9338
rect -4010 9304 -3976 9338
rect -3930 9304 -3896 9338
rect -3850 9304 -3816 9338
rect -3770 9304 -3736 9338
rect -3690 9304 -3656 9338
rect -3610 9304 -3576 9338
rect -3530 9304 -3496 9338
rect -3450 9304 -3416 9338
rect -3370 9304 -3336 9338
rect -1929 9304 -1895 9338
rect -1849 9304 -1815 9338
rect -1769 9304 -1735 9338
rect -1689 9304 -1655 9338
rect -1609 9304 -1575 9338
rect -1529 9304 -1495 9338
rect -1449 9304 -1415 9338
rect -1369 9304 -1335 9338
rect -1289 9304 -1255 9338
rect -1209 9304 -1175 9338
rect -1129 9304 -1095 9338
rect -1049 9304 -1015 9338
rect -969 9304 -935 9338
rect -889 9304 -855 9338
rect -809 9304 -775 9338
rect -729 9304 -695 9338
rect -649 9304 -615 9338
rect -569 9304 -535 9338
rect -489 9304 -455 9338
rect -409 9304 -375 9338
rect -329 9304 -295 9338
rect -249 9304 -215 9338
rect -169 9304 -135 9338
rect -89 9304 -55 9338
rect -9 9304 25 9338
rect 71 9304 105 9338
rect 151 9304 185 9338
rect 231 9304 265 9338
rect 311 9304 345 9338
rect 391 9304 425 9338
rect 471 9304 505 9338
rect 551 9304 585 9338
rect 631 9304 665 9338
rect 711 9304 745 9338
rect 791 9304 825 9338
rect 871 9304 905 9338
rect 951 9304 985 9338
rect 1031 9304 1065 9338
rect 1111 9304 1145 9338
rect 1191 9304 1225 9338
rect 1271 9304 1305 9338
rect 1351 9304 1385 9338
rect 1431 9304 1465 9338
rect 1511 9304 1545 9338
rect 1591 9304 1625 9338
rect 1671 9304 1705 9338
rect 1751 9304 1785 9338
rect 1831 9304 1865 9338
rect 1911 9304 1945 9338
rect 1991 9304 2025 9338
rect 2071 9304 2105 9338
rect 2151 9304 2185 9338
rect 2231 9304 2265 9338
rect 2311 9304 2345 9338
rect 3790 9304 3824 9338
rect 3870 9304 3904 9338
rect 3950 9304 3984 9338
rect 4030 9304 4064 9338
rect 4110 9304 4144 9338
rect 4190 9304 4224 9338
rect 4270 9304 4304 9338
rect 4350 9304 4384 9338
rect 4430 9304 4464 9338
rect 4510 9304 4544 9338
rect 4590 9304 4624 9338
rect 4670 9304 4704 9338
rect 4750 9304 4784 9338
rect 4830 9304 4864 9338
rect 4910 9304 4944 9338
rect 4990 9304 5024 9338
rect 5070 9304 5104 9338
rect 5150 9304 5184 9338
rect 5230 9304 5264 9338
rect 5310 9304 5344 9338
rect 5390 9304 5424 9338
rect 5470 9304 5504 9338
rect 5550 9304 5584 9338
rect 5630 9304 5664 9338
rect 5710 9304 5744 9338
rect 5790 9304 5824 9338
rect 5870 9304 5904 9338
rect 5950 9304 5984 9338
rect 6030 9304 6064 9338
rect 6110 9304 6144 9338
rect 6190 9304 6224 9338
rect 6270 9304 6304 9338
rect 6350 9304 6384 9338
rect 6430 9304 6464 9338
rect 6510 9304 6544 9338
rect 6590 9304 6624 9338
rect 6670 9304 6704 9338
rect 6750 9304 6784 9338
rect 6830 9304 6864 9338
rect 6910 9304 6944 9338
rect 6990 9304 7024 9338
rect 7070 9304 7104 9338
rect 7150 9304 7184 9338
rect 7230 9304 7264 9338
rect 7310 9304 7344 9338
rect 7390 9304 7424 9338
rect 7470 9304 7504 9338
rect 7550 9304 7584 9338
rect 7630 9304 7664 9338
rect 7710 9304 7744 9338
rect 7790 9304 7824 9338
rect 7870 9304 7904 9338
rect 7950 9304 7984 9338
rect 8030 9304 8064 9338
rect 8110 9304 8144 9338
rect 8190 9304 8224 9338
rect 8270 9304 8304 9338
rect 8350 9304 8384 9338
rect 8430 9304 8464 9338
rect 8510 9304 8544 9338
rect 8590 9304 8624 9338
rect 8670 9304 8704 9338
rect 8750 9304 8784 9338
rect 8830 9304 8864 9338
rect 8910 9304 8944 9338
rect 8990 9304 9024 9338
rect 9070 9304 9104 9338
rect 9150 9304 9184 9338
rect 9230 9304 9264 9338
rect 9310 9304 9344 9338
rect 9390 9304 9424 9338
rect 9470 9304 9504 9338
rect 9550 9304 9584 9338
rect 9630 9304 9664 9338
rect 9710 9304 9744 9338
rect 9790 9304 9824 9338
rect 9870 9304 9904 9338
rect 9950 9304 9984 9338
rect 10030 9304 10064 9338
rect 10110 9304 10144 9338
rect 10190 9304 10224 9338
rect 10270 9304 10304 9338
rect 10350 9304 10384 9338
rect 10430 9304 10464 9338
rect 10510 9304 10544 9338
rect 10590 9304 10624 9338
rect 10670 9304 10704 9338
rect 10750 9304 10784 9338
rect 10830 9304 10864 9338
rect 10910 9304 10944 9338
rect 10990 9304 11024 9338
rect 11070 9304 11104 9338
rect 11150 9304 11184 9338
rect 11230 9304 11264 9338
rect 11310 9304 11344 9338
rect 11390 9304 11424 9338
rect 11470 9304 11504 9338
rect 11550 9304 11584 9338
rect 11630 9304 11664 9338
rect 11710 9304 11744 9338
rect 11790 9304 11824 9338
rect 11870 9304 11904 9338
rect 11950 9304 11984 9338
rect 12030 9304 12064 9338
rect 12110 9304 12144 9338
rect 12190 9304 12224 9338
rect 12270 9304 12304 9338
rect 12350 9304 12384 9338
rect 12430 9304 12464 9338
rect 12510 9304 12544 9338
rect 12590 9304 12624 9338
rect 12670 9304 12704 9338
rect 12750 9304 12784 9338
rect 12830 9304 12864 9338
rect 12910 9304 12944 9338
rect 12990 9304 13024 9338
rect 13070 9304 13104 9338
rect 13150 9304 13184 9338
rect 13230 9304 13264 9338
rect 13310 9304 13344 9338
rect 13390 9304 13424 9338
rect 13470 9304 13504 9338
rect 13550 9304 13584 9338
rect 13630 9304 13664 9338
rect 13710 9304 13744 9338
rect 13790 9304 13824 9338
rect 13870 9304 13904 9338
rect 13950 9304 13984 9338
rect 14030 9304 14064 9338
rect 14110 9304 14144 9338
rect 14190 9304 14224 9338
rect 14270 9304 14304 9338
rect 14350 9304 14384 9338
rect 14430 9304 14464 9338
rect 14510 9304 14544 9338
rect 14590 9304 14624 9338
rect 14670 9304 14704 9338
rect 14750 9304 14784 9338
rect 14830 9304 14864 9338
rect 14910 9304 14944 9338
rect 14990 9304 15024 9338
rect 15070 9304 15104 9338
rect 15150 9304 15184 9338
rect 15230 9304 15264 9338
rect 15310 9304 15344 9338
rect 15390 9304 15424 9338
rect 15470 9304 15504 9338
rect 15550 9304 15584 9338
rect 15630 9304 15664 9338
rect 15710 9304 15744 9338
rect 15790 9304 15824 9338
rect 15870 9304 15904 9338
rect 15950 9304 15984 9338
rect 16030 9304 16064 9338
rect 16110 9304 16144 9338
rect 16190 9304 16224 9338
rect 16270 9304 16304 9338
rect 16350 9304 16384 9338
rect 16430 9304 16464 9338
rect 16510 9304 16544 9338
rect 16590 9304 16624 9338
rect 16670 9304 16704 9338
rect 16751 9304 16785 9338
rect 16831 9304 16865 9338
rect 16911 9304 16945 9338
rect 16991 9304 17025 9338
rect 17071 9304 17105 9338
rect 17151 9304 17185 9338
rect 17231 9304 17265 9338
rect 17311 9304 17345 9338
rect 17391 9304 17425 9338
rect 17471 9304 17505 9338
rect 17551 9304 17585 9338
rect 17631 9304 17665 9338
rect 17711 9304 17745 9338
rect 17791 9304 17825 9338
rect 17871 9304 17905 9338
rect 17951 9304 17985 9338
rect 18031 9304 18065 9338
rect 18111 9304 18145 9338
rect 18191 9304 18225 9338
rect 18271 9304 18305 9338
rect 18351 9304 18385 9338
rect 18431 9304 18465 9338
rect 18511 9304 18545 9338
rect 18591 9304 18625 9338
rect 18671 9304 18705 9338
rect 18751 9304 18785 9338
rect 18831 9304 18865 9338
rect 18911 9304 18945 9338
rect 18991 9304 19025 9338
rect 19071 9304 19105 9338
rect 19151 9304 19185 9338
rect 19231 9304 19265 9338
rect 19311 9304 19345 9338
rect 19391 9304 19425 9338
rect 19471 9304 19505 9338
rect 19551 9304 19585 9338
rect 19631 9304 19665 9338
rect 19711 9304 19745 9338
rect 19791 9304 19825 9338
rect 19871 9304 19905 9338
rect 19951 9304 19985 9338
rect 20031 9304 20065 9338
rect 20111 9304 20145 9338
rect 20191 9304 20225 9338
rect 20271 9304 20305 9338
rect 20351 9304 20385 9338
rect 20431 9304 20465 9338
rect 20511 9304 20545 9338
rect 20591 9304 20625 9338
rect 20671 9304 20705 9338
rect 20751 9304 20785 9338
rect 20831 9304 20865 9338
rect 20911 9304 20945 9338
rect 20991 9304 21025 9338
rect 21071 9304 21105 9338
rect 21151 9304 21185 9338
rect 21231 9304 21265 9338
rect 21311 9304 21345 9338
rect 21391 9304 21425 9338
rect 21471 9304 21505 9338
rect 21551 9304 21585 9338
rect 21631 9304 21665 9338
rect 21711 9304 21745 9338
rect 21791 9304 21825 9338
rect 21871 9304 21905 9338
rect 21951 9304 21985 9338
rect 22031 9304 22065 9338
rect 22111 9304 22145 9338
rect 22191 9304 22225 9338
rect 22271 9304 22305 9338
rect 22351 9304 22385 9338
rect 22431 9304 22465 9338
rect 22511 9304 22545 9338
rect 22591 9304 22625 9338
rect 22671 9304 22705 9338
rect 22751 9304 22785 9338
rect 22831 9304 22865 9338
rect 22911 9304 22945 9338
rect 22991 9304 23025 9338
rect 23071 9304 23105 9338
rect 23151 9304 23185 9338
rect 23231 9304 23265 9338
rect 23311 9304 23345 9338
rect 23391 9304 23425 9338
rect 23471 9304 23505 9338
rect 23551 9304 23585 9338
rect 23631 9304 23665 9338
rect 23711 9304 23745 9338
rect 23791 9304 23825 9338
rect 23871 9304 23905 9338
rect 23951 9304 23985 9338
rect 24031 9304 24065 9338
rect 24111 9304 24145 9338
rect 24191 9304 24225 9338
rect 24271 9304 24305 9338
rect 24351 9304 24385 9338
rect 24431 9304 24465 9338
rect 24511 9304 24545 9338
rect 24591 9304 24625 9338
rect 24671 9304 24705 9338
rect 24751 9304 24785 9338
rect 24831 9304 24865 9338
rect 24911 9304 24945 9338
rect 24991 9304 25025 9338
rect 25071 9304 25105 9338
rect 25151 9304 25185 9338
rect 25231 9304 25265 9338
rect 25311 9304 25345 9338
rect 25391 9304 25425 9338
rect 25471 9304 25505 9338
rect 25551 9304 25585 9338
rect 25631 9304 25665 9338
rect 25711 9304 25745 9338
rect 25791 9304 25825 9338
rect 25871 9304 25905 9338
rect 25951 9304 25985 9338
rect 26031 9304 26065 9338
rect 26111 9304 26145 9338
rect 26191 9304 26225 9338
rect 26271 9304 26305 9338
rect 26351 9304 26385 9338
rect 26431 9304 26465 9338
rect 26511 9304 26545 9338
rect 26591 9304 26625 9338
rect 26671 9304 26705 9338
rect 26751 9304 26785 9338
rect 26831 9304 26865 9338
rect 26911 9304 26945 9338
rect 26991 9304 27025 9338
rect 27071 9304 27105 9338
rect 27151 9304 27185 9338
rect 27231 9304 27265 9338
rect 27311 9304 27345 9338
rect 27391 9304 27425 9338
rect 27471 9304 27505 9338
rect 27551 9304 27585 9338
rect 27631 9304 27665 9338
rect 27711 9304 27745 9338
rect 27791 9304 27825 9338
rect 27871 9304 27905 9338
rect 27951 9304 27985 9338
rect 28031 9304 28065 9338
rect 28111 9304 28145 9338
rect 28191 9304 28225 9338
rect 28271 9304 28305 9338
rect 28351 9304 28385 9338
rect 28431 9304 28465 9338
rect 28511 9304 28545 9338
rect 28591 9304 28625 9338
rect 28671 9304 28705 9338
rect 28751 9304 28785 9338
rect 28831 9304 28865 9338
rect 28911 9304 28945 9338
rect 28991 9304 29025 9338
rect 29071 9304 29105 9338
rect 29151 9304 29185 9338
rect 29231 9304 29265 9338
rect 29311 9304 29345 9338
rect 29391 9304 29425 9338
rect 29471 9304 29505 9338
rect 29551 9304 29585 9338
rect 29631 9304 29665 9338
rect 29711 9304 29745 9338
rect 29791 9304 29825 9338
rect 29871 9304 29905 9338
rect 29951 9304 29985 9338
rect 30031 9304 30065 9338
rect 30111 9304 30145 9338
rect 30191 9304 30225 9338
rect 30271 9304 30305 9338
rect 30351 9304 30385 9338
rect 30431 9304 30465 9338
rect 30511 9304 30545 9338
rect 30591 9304 30625 9338
rect 30671 9304 30705 9338
rect 30751 9304 30785 9338
rect 30831 9304 30865 9338
rect 30911 9304 30945 9338
rect 30991 9304 31025 9338
rect 31071 9304 31105 9338
rect 31151 9304 31185 9338
rect 31231 9304 31265 9338
rect 31311 9304 31345 9338
rect 31391 9304 31425 9338
rect 31471 9304 31505 9338
rect 31551 9304 31585 9338
rect 31631 9304 31665 9338
rect 31711 9304 31745 9338
rect 31791 9304 31825 9338
rect 31871 9304 31905 9338
rect 31951 9304 31985 9338
rect 32031 9304 32065 9338
rect 32111 9304 32145 9338
rect 32191 9304 32225 9338
rect 32271 9304 32305 9338
rect 32351 9304 32385 9338
rect 32431 9304 32465 9338
rect 32511 9304 32545 9338
rect 32591 9304 32625 9338
rect 32671 9304 32705 9338
rect 32751 9304 32785 9338
rect 32831 9304 32865 9338
rect 32911 9304 32945 9338
rect 32991 9304 33025 9338
rect 33071 9304 33105 9338
rect 33151 9304 33185 9338
rect 33231 9304 33265 9338
rect 33311 9304 33345 9338
rect 33391 9304 33425 9338
rect 33471 9304 33505 9338
rect 33551 9304 33585 9338
rect 33631 9304 33665 9338
rect 33711 9304 33745 9338
rect 33791 9304 33825 9338
rect 33871 9304 33905 9338
rect 33951 9304 33985 9338
rect 34031 9304 34065 9338
rect 34111 9304 34145 9338
rect 34191 9304 34225 9338
rect 34271 9304 34305 9338
rect 34351 9304 34385 9338
rect 34431 9304 34465 9338
rect 34511 9304 34545 9338
rect 34591 9304 34625 9338
rect 34671 9304 34705 9338
rect 34751 9304 34785 9338
rect 34831 9304 34865 9338
rect 34911 9304 34945 9338
rect 34991 9304 35025 9338
rect 35071 9304 35105 9338
rect 35151 9304 35185 9338
rect 35231 9304 35265 9338
rect 35311 9304 35345 9338
rect 35391 9304 35425 9338
rect 35471 9304 35505 9338
rect 35551 9304 35585 9338
rect 35631 9304 35665 9338
rect 35711 9304 35745 9338
rect 35791 9304 35825 9338
rect 35871 9304 35905 9338
rect 35951 9304 35985 9338
rect 36031 9304 36065 9338
rect 36111 9304 36145 9338
rect 36191 9304 36225 9338
rect 36271 9304 36305 9338
rect 36351 9304 36385 9338
rect 36431 9304 36465 9338
rect 36511 9304 36545 9338
rect 36591 9304 36625 9338
rect 36671 9304 36705 9338
rect 36751 9304 36785 9338
rect 36831 9304 36865 9338
rect 36911 9304 36945 9338
rect 36991 9304 37025 9338
rect 37071 9304 37105 9338
rect 37151 9304 37185 9338
rect 37231 9304 37265 9338
rect 37311 9304 37345 9338
rect 37391 9304 37425 9338
rect 37471 9304 37505 9338
rect 37551 9304 37585 9338
rect 37631 9304 37665 9338
rect 37711 9304 37745 9338
rect 37791 9304 37825 9338
rect 37871 9304 37905 9338
rect 37951 9304 37985 9338
rect 38031 9304 38065 9338
rect 38111 9304 38145 9338
rect 38191 9304 38225 9338
rect 38271 9304 38305 9338
rect 1266 7933 1300 7967
rect -1340 6703 -1306 6737
rect -37851 6326 -37817 6360
rect -37771 6326 -37737 6360
rect -37691 6326 -37657 6360
rect -37611 6326 -37577 6360
rect -37531 6326 -37497 6360
rect -37451 6326 -37417 6360
rect -37371 6326 -37337 6360
rect -37291 6326 -37257 6360
rect -37211 6326 -37177 6360
rect -37131 6326 -37097 6360
rect -37051 6326 -37017 6360
rect -36971 6326 -36937 6360
rect -36891 6326 -36857 6360
rect -36811 6326 -36777 6360
rect -36731 6326 -36697 6360
rect -36651 6326 -36617 6360
rect -36571 6326 -36537 6360
rect -36491 6326 -36457 6360
rect -36411 6326 -36377 6360
rect -36331 6326 -36297 6360
rect -36251 6326 -36217 6360
rect -36171 6326 -36137 6360
rect -36091 6326 -36057 6360
rect -36011 6326 -35977 6360
rect -35931 6326 -35897 6360
rect -35851 6326 -35817 6360
rect -35771 6326 -35737 6360
rect -35691 6326 -35657 6360
rect -35611 6326 -35577 6360
rect -35531 6326 -35497 6360
rect -35451 6326 -35417 6360
rect -35371 6326 -35337 6360
rect -35291 6326 -35257 6360
rect -35211 6326 -35177 6360
rect -35131 6326 -35097 6360
rect -35051 6326 -35017 6360
rect -34971 6326 -34937 6360
rect -34891 6326 -34857 6360
rect -34811 6326 -34777 6360
rect -34731 6326 -34697 6360
rect -34651 6326 -34617 6360
rect -34571 6326 -34537 6360
rect -34491 6326 -34457 6360
rect -34411 6326 -34377 6360
rect -34331 6326 -34297 6360
rect -34251 6326 -34217 6360
rect -34171 6326 -34137 6360
rect -34091 6326 -34057 6360
rect -34011 6326 -33977 6360
rect -33931 6326 -33897 6360
rect -33851 6326 -33817 6360
rect -33771 6326 -33737 6360
rect -33691 6326 -33657 6360
rect -33611 6326 -33577 6360
rect -33531 6326 -33497 6360
rect -33451 6326 -33417 6360
rect -33371 6326 -33337 6360
rect -33291 6326 -33257 6360
rect -33211 6326 -33177 6360
rect -33131 6326 -33097 6360
rect -33051 6326 -33017 6360
rect -32971 6326 -32937 6360
rect -32891 6326 -32857 6360
rect -32811 6326 -32777 6360
rect -32731 6326 -32697 6360
rect -32651 6326 -32617 6360
rect -32571 6326 -32537 6360
rect -32491 6326 -32457 6360
rect -32411 6326 -32377 6360
rect -32331 6326 -32297 6360
rect -32251 6326 -32217 6360
rect -32171 6326 -32137 6360
rect -32091 6326 -32057 6360
rect -32011 6326 -31977 6360
rect -31931 6326 -31897 6360
rect -31851 6326 -31817 6360
rect -31771 6326 -31737 6360
rect -31691 6326 -31657 6360
rect -31611 6326 -31577 6360
rect -31531 6326 -31497 6360
rect -31451 6326 -31417 6360
rect -31371 6326 -31337 6360
rect -31291 6326 -31257 6360
rect -31211 6326 -31177 6360
rect -31131 6326 -31097 6360
rect -31051 6326 -31017 6360
rect -30971 6326 -30937 6360
rect -30891 6326 -30857 6360
rect -30811 6326 -30777 6360
rect -30731 6326 -30697 6360
rect -30651 6326 -30617 6360
rect -30571 6326 -30537 6360
rect -30491 6326 -30457 6360
rect -30411 6326 -30377 6360
rect -30331 6326 -30297 6360
rect -30251 6326 -30217 6360
rect -30171 6326 -30137 6360
rect -30091 6326 -30057 6360
rect -30011 6326 -29977 6360
rect -29931 6326 -29897 6360
rect -29851 6326 -29817 6360
rect -29771 6326 -29737 6360
rect -29691 6326 -29657 6360
rect -29611 6326 -29577 6360
rect -29531 6326 -29497 6360
rect -29451 6326 -29417 6360
rect -29371 6326 -29337 6360
rect -29291 6326 -29257 6360
rect -29211 6326 -29177 6360
rect -29131 6326 -29097 6360
rect -29051 6326 -29017 6360
rect -28971 6326 -28937 6360
rect -28891 6326 -28857 6360
rect -28811 6326 -28777 6360
rect -28731 6326 -28697 6360
rect -28651 6326 -28617 6360
rect -28571 6326 -28537 6360
rect -28491 6326 -28457 6360
rect -28411 6326 -28377 6360
rect -28331 6326 -28297 6360
rect -28251 6326 -28217 6360
rect -28171 6326 -28137 6360
rect -28091 6326 -28057 6360
rect -28011 6326 -27977 6360
rect -27931 6326 -27897 6360
rect -27851 6326 -27817 6360
rect -27771 6326 -27737 6360
rect -27691 6326 -27657 6360
rect -27611 6326 -27577 6360
rect -27531 6326 -27497 6360
rect -27451 6326 -27417 6360
rect -27371 6326 -27337 6360
rect -27291 6326 -27257 6360
rect -27211 6326 -27177 6360
rect -27131 6326 -27097 6360
rect -27051 6326 -27017 6360
rect -26971 6326 -26937 6360
rect -26891 6326 -26857 6360
rect -26811 6326 -26777 6360
rect -26731 6326 -26697 6360
rect -26651 6326 -26617 6360
rect -26571 6326 -26537 6360
rect -26491 6326 -26457 6360
rect -26411 6326 -26377 6360
rect -26331 6326 -26297 6360
rect -26251 6326 -26217 6360
rect -26171 6326 -26137 6360
rect -26091 6326 -26057 6360
rect -26011 6326 -25977 6360
rect -25931 6326 -25897 6360
rect -25851 6326 -25817 6360
rect -25771 6326 -25737 6360
rect -25691 6326 -25657 6360
rect -25611 6326 -25577 6360
rect -25531 6326 -25497 6360
rect -25451 6326 -25417 6360
rect -25371 6326 -25337 6360
rect -25291 6326 -25257 6360
rect -25211 6326 -25177 6360
rect -25131 6326 -25097 6360
rect -25051 6326 -25017 6360
rect -24971 6326 -24937 6360
rect -24890 6326 -24856 6360
rect -24810 6326 -24776 6360
rect -24730 6326 -24696 6360
rect -24650 6326 -24616 6360
rect -24570 6326 -24536 6360
rect -24490 6326 -24456 6360
rect -24410 6326 -24376 6360
rect -24330 6326 -24296 6360
rect -24250 6326 -24216 6360
rect -24170 6326 -24136 6360
rect -24090 6326 -24056 6360
rect -24010 6326 -23976 6360
rect -23930 6326 -23896 6360
rect -23850 6326 -23816 6360
rect -23770 6326 -23736 6360
rect -23690 6326 -23656 6360
rect -23610 6326 -23576 6360
rect -23530 6326 -23496 6360
rect -23450 6326 -23416 6360
rect -23370 6326 -23336 6360
rect -23290 6326 -23256 6360
rect -23210 6326 -23176 6360
rect -23130 6326 -23096 6360
rect -23050 6326 -23016 6360
rect -22970 6326 -22936 6360
rect -22890 6326 -22856 6360
rect -22810 6326 -22776 6360
rect -22730 6326 -22696 6360
rect -22650 6326 -22616 6360
rect -22570 6326 -22536 6360
rect -22490 6326 -22456 6360
rect -22410 6326 -22376 6360
rect -22330 6326 -22296 6360
rect -22250 6326 -22216 6360
rect -22170 6326 -22136 6360
rect -22090 6326 -22056 6360
rect -22010 6326 -21976 6360
rect -21930 6326 -21896 6360
rect -21850 6326 -21816 6360
rect -21770 6326 -21736 6360
rect -21690 6326 -21656 6360
rect -21610 6326 -21576 6360
rect -21530 6326 -21496 6360
rect -21450 6326 -21416 6360
rect -21370 6326 -21336 6360
rect -21290 6326 -21256 6360
rect -21210 6326 -21176 6360
rect -21130 6326 -21096 6360
rect -21050 6326 -21016 6360
rect -20970 6326 -20936 6360
rect -20890 6326 -20856 6360
rect -20810 6326 -20776 6360
rect -20730 6326 -20696 6360
rect -20650 6326 -20616 6360
rect -20570 6326 -20536 6360
rect -20490 6326 -20456 6360
rect -20410 6326 -20376 6360
rect -20330 6326 -20296 6360
rect -20250 6326 -20216 6360
rect -20170 6326 -20136 6360
rect -20090 6326 -20056 6360
rect -20010 6326 -19976 6360
rect -19930 6326 -19896 6360
rect -19850 6326 -19816 6360
rect -19770 6326 -19736 6360
rect -19690 6326 -19656 6360
rect -19610 6326 -19576 6360
rect -19530 6326 -19496 6360
rect -19450 6326 -19416 6360
rect -19370 6326 -19336 6360
rect -19290 6326 -19256 6360
rect -19210 6326 -19176 6360
rect -19130 6326 -19096 6360
rect -19050 6326 -19016 6360
rect -18970 6326 -18936 6360
rect -18890 6326 -18856 6360
rect -18810 6326 -18776 6360
rect -18730 6326 -18696 6360
rect -18650 6326 -18616 6360
rect -18570 6326 -18536 6360
rect -18490 6326 -18456 6360
rect -18410 6326 -18376 6360
rect -18330 6326 -18296 6360
rect -18250 6326 -18216 6360
rect -18170 6326 -18136 6360
rect -18090 6326 -18056 6360
rect -18010 6326 -17976 6360
rect -17930 6326 -17896 6360
rect -17850 6326 -17816 6360
rect -17770 6326 -17736 6360
rect -17690 6326 -17656 6360
rect -17610 6326 -17576 6360
rect -17530 6326 -17496 6360
rect -17450 6326 -17416 6360
rect -17370 6326 -17336 6360
rect -17290 6326 -17256 6360
rect -17210 6326 -17176 6360
rect -17130 6326 -17096 6360
rect -17050 6326 -17016 6360
rect -16970 6326 -16936 6360
rect -16890 6326 -16856 6360
rect -16810 6326 -16776 6360
rect -16730 6326 -16696 6360
rect -16650 6326 -16616 6360
rect -16570 6326 -16536 6360
rect -16490 6326 -16456 6360
rect -16410 6326 -16376 6360
rect -16330 6326 -16296 6360
rect -16250 6326 -16216 6360
rect -16170 6326 -16136 6360
rect -16090 6326 -16056 6360
rect -16010 6326 -15976 6360
rect -15930 6326 -15896 6360
rect -15850 6326 -15816 6360
rect -15770 6326 -15736 6360
rect -15690 6326 -15656 6360
rect -15610 6326 -15576 6360
rect -15530 6326 -15496 6360
rect -15450 6326 -15416 6360
rect -15370 6326 -15336 6360
rect -15290 6326 -15256 6360
rect -15210 6326 -15176 6360
rect -15130 6326 -15096 6360
rect -15050 6326 -15016 6360
rect -14970 6326 -14936 6360
rect -14890 6326 -14856 6360
rect -14810 6326 -14776 6360
rect -14730 6326 -14696 6360
rect -14650 6326 -14616 6360
rect -14570 6326 -14536 6360
rect -14490 6326 -14456 6360
rect -14410 6326 -14376 6360
rect -14330 6326 -14296 6360
rect -14250 6326 -14216 6360
rect -14170 6326 -14136 6360
rect -14090 6326 -14056 6360
rect -14010 6326 -13976 6360
rect -13930 6326 -13896 6360
rect -13850 6326 -13816 6360
rect -13770 6326 -13736 6360
rect -13690 6326 -13656 6360
rect -13610 6326 -13576 6360
rect -13530 6326 -13496 6360
rect -13450 6326 -13416 6360
rect -13370 6326 -13336 6360
rect -13290 6326 -13256 6360
rect -13210 6326 -13176 6360
rect -13130 6326 -13096 6360
rect -13050 6326 -13016 6360
rect -12970 6326 -12936 6360
rect -12890 6326 -12856 6360
rect -12810 6326 -12776 6360
rect -12730 6326 -12696 6360
rect -12650 6326 -12616 6360
rect -12570 6326 -12536 6360
rect -12490 6326 -12456 6360
rect -12410 6326 -12376 6360
rect -12330 6326 -12296 6360
rect -12250 6326 -12216 6360
rect -12170 6326 -12136 6360
rect -12090 6326 -12056 6360
rect -12010 6326 -11976 6360
rect -11929 6326 -11895 6360
rect -11849 6326 -11815 6360
rect -11769 6326 -11735 6360
rect -11689 6326 -11655 6360
rect -11609 6326 -11575 6360
rect -11529 6326 -11495 6360
rect -11449 6326 -11415 6360
rect -11369 6326 -11335 6360
rect -11289 6326 -11255 6360
rect -11209 6326 -11175 6360
rect -11129 6326 -11095 6360
rect -11049 6326 -11015 6360
rect -10969 6326 -10935 6360
rect -10889 6326 -10855 6360
rect -10809 6326 -10775 6360
rect -10729 6326 -10695 6360
rect -10649 6326 -10615 6360
rect -10569 6326 -10535 6360
rect -10489 6326 -10455 6360
rect -10409 6326 -10375 6360
rect -10329 6326 -10295 6360
rect -10249 6326 -10215 6360
rect -10169 6326 -10135 6360
rect -10089 6326 -10055 6360
rect -10009 6326 -9975 6360
rect -9929 6326 -9895 6360
rect -9849 6326 -9815 6360
rect -9769 6326 -9735 6360
rect -9689 6326 -9655 6360
rect -9609 6326 -9575 6360
rect -9529 6326 -9495 6360
rect -9449 6326 -9415 6360
rect -9369 6326 -9335 6360
rect -9289 6326 -9255 6360
rect -9209 6326 -9175 6360
rect -9129 6326 -9095 6360
rect -9049 6326 -9015 6360
rect -8969 6326 -8935 6360
rect -8889 6326 -8855 6360
rect -8809 6326 -8775 6360
rect -8729 6326 -8695 6360
rect -8649 6326 -8615 6360
rect -8569 6326 -8535 6360
rect -8489 6326 -8455 6360
rect -8409 6326 -8375 6360
rect -8329 6326 -8295 6360
rect -8249 6326 -8215 6360
rect -8169 6326 -8135 6360
rect -8089 6326 -8055 6360
rect -8009 6326 -7975 6360
rect -7929 6326 -7895 6360
rect -7849 6326 -7815 6360
rect -7769 6326 -7735 6360
rect -7689 6326 -7655 6360
rect -7609 6326 -7575 6360
rect -7529 6326 -7495 6360
rect -7449 6326 -7415 6360
rect -7369 6326 -7335 6360
rect -7289 6326 -7255 6360
rect -7209 6326 -7175 6360
rect -7129 6326 -7095 6360
rect -7049 6326 -7015 6360
rect -6969 6326 -6935 6360
rect -6889 6326 -6855 6360
rect -6809 6326 -6775 6360
rect -6729 6326 -6695 6360
rect -6649 6326 -6615 6360
rect -6569 6326 -6535 6360
rect -6489 6326 -6455 6360
rect -6409 6326 -6375 6360
rect -6329 6326 -6295 6360
rect -6249 6326 -6215 6360
rect -6169 6326 -6135 6360
rect -6089 6326 -6055 6360
rect -6009 6326 -5975 6360
rect -5929 6326 -5895 6360
rect -5849 6326 -5815 6360
rect -5769 6326 -5735 6360
rect -5689 6326 -5655 6360
rect -5609 6326 -5575 6360
rect -5529 6326 -5495 6360
rect -5449 6326 -5415 6360
rect -5369 6326 -5335 6360
rect -5289 6326 -5255 6360
rect -5209 6326 -5175 6360
rect -5129 6326 -5095 6360
rect -5049 6326 -5015 6360
rect -4969 6326 -4935 6360
rect -4889 6326 -4855 6360
rect -4809 6326 -4775 6360
rect -4729 6326 -4695 6360
rect -4649 6326 -4615 6360
rect -4569 6326 -4535 6360
rect -4489 6326 -4455 6360
rect -4409 6326 -4375 6360
rect -4329 6326 -4295 6360
rect -4249 6326 -4215 6360
rect -4169 6326 -4135 6360
rect -4089 6326 -4055 6360
rect -4009 6326 -3975 6360
rect -3929 6326 -3895 6360
rect -3849 6326 -3815 6360
rect -3769 6326 -3735 6360
rect -3689 6326 -3655 6360
rect -3609 6326 -3575 6360
rect -3529 6326 -3495 6360
rect -3449 6326 -3415 6360
rect -3369 6326 -3335 6360
rect -3289 6326 -3255 6360
rect -3209 6326 -3175 6360
rect -3129 6326 -3095 6360
rect -3049 6326 -3015 6360
rect -2969 6326 -2935 6360
rect -2889 6326 -2855 6360
rect -2809 6326 -2775 6360
rect -2729 6326 -2695 6360
rect -2649 6326 -2615 6360
rect -2569 6326 -2535 6360
rect -2489 6326 -2455 6360
rect -2409 6326 -2375 6360
rect -2329 6326 -2295 6360
rect -2249 6326 -2215 6360
rect -2169 6326 -2135 6360
rect -2089 6326 -2055 6360
rect -2009 6326 -1975 6360
rect -1929 6326 -1895 6360
rect -1849 6326 -1815 6360
rect -1769 6326 -1735 6360
rect -1689 6326 -1655 6360
rect -1609 6326 -1575 6360
rect -1529 6326 -1495 6360
rect -1449 6326 -1415 6360
rect -1369 6326 -1335 6360
rect -1289 6326 -1255 6360
rect -1209 6326 -1175 6360
rect -1129 6326 -1095 6360
rect -1049 6326 -1015 6360
rect -969 6326 -935 6360
rect -889 6326 -855 6360
rect -809 6326 -775 6360
rect -729 6326 -695 6360
rect -649 6326 -615 6360
rect -569 6326 -535 6360
rect -489 6326 -455 6360
rect -409 6326 -375 6360
rect -329 6326 -295 6360
rect -249 6326 -215 6360
rect -169 6326 -135 6360
rect -89 6326 -55 6360
rect -9 6326 25 6360
rect 71 6326 105 6360
rect 151 6326 185 6360
rect 231 6326 265 6360
rect 311 6326 345 6360
rect 391 6326 425 6360
rect 471 6326 505 6360
rect 551 6326 585 6360
rect 631 6326 665 6360
rect 711 6326 745 6360
rect 791 6326 825 6360
rect 871 6326 905 6360
rect 951 6326 985 6360
rect 1031 6326 1065 6360
rect 1111 6326 1145 6360
rect 1191 6326 1225 6360
rect 1271 6326 1305 6360
rect 1351 6326 1385 6360
rect 1431 6326 1465 6360
rect 1511 6326 1545 6360
rect 1591 6326 1625 6360
rect 1671 6326 1705 6360
rect 1751 6326 1785 6360
rect 1831 6326 1865 6360
rect 1911 6326 1945 6360
rect 1991 6326 2025 6360
rect 2071 6326 2105 6360
rect 2151 6326 2185 6360
rect 2231 6326 2265 6360
rect 2311 6326 2345 6360
rect 2391 6326 2425 6360
rect 2471 6326 2505 6360
rect 2551 6326 2585 6360
rect 2631 6326 2665 6360
rect 2711 6326 2745 6360
rect 2791 6326 2825 6360
rect 2871 6326 2905 6360
rect 2951 6326 2985 6360
rect 3031 6326 3065 6360
rect 3111 6326 3145 6360
rect 3191 6326 3225 6360
rect 3271 6326 3305 6360
rect 3351 6326 3385 6360
rect 3431 6326 3465 6360
rect 3511 6326 3545 6360
rect 3591 6326 3625 6360
rect 3671 6326 3705 6360
rect 3751 6326 3785 6360
rect 3831 6326 3865 6360
rect 3911 6326 3945 6360
rect 3991 6326 4025 6360
rect 4071 6326 4105 6360
rect 4151 6326 4185 6360
rect 4231 6326 4265 6360
rect 4311 6326 4345 6360
rect 4391 6326 4425 6360
rect 4471 6326 4505 6360
rect 4551 6326 4585 6360
rect 4631 6326 4665 6360
rect 4711 6326 4745 6360
rect 4791 6326 4825 6360
rect 4871 6326 4905 6360
rect 4951 6326 4985 6360
rect 5031 6326 5065 6360
rect 5111 6326 5145 6360
rect 5191 6326 5225 6360
rect 5271 6326 5305 6360
rect 5351 6326 5385 6360
rect 5431 6326 5465 6360
rect 5511 6326 5545 6360
rect 5591 6326 5625 6360
rect 5671 6326 5705 6360
rect 5751 6326 5785 6360
rect 5831 6326 5865 6360
rect 5911 6326 5945 6360
rect 5991 6326 6025 6360
rect 6071 6326 6105 6360
rect 6151 6326 6185 6360
rect 6231 6326 6265 6360
rect 6311 6326 6345 6360
rect 6391 6326 6425 6360
rect 6471 6326 6505 6360
rect 6551 6326 6585 6360
rect 6631 6326 6665 6360
rect 6711 6326 6745 6360
rect 6791 6326 6825 6360
rect 6871 6326 6905 6360
rect 6951 6326 6985 6360
rect 7031 6326 7065 6360
rect 7111 6326 7145 6360
rect 7191 6326 7225 6360
rect 7271 6326 7305 6360
rect 7351 6326 7385 6360
rect 7431 6326 7465 6360
rect 7511 6326 7545 6360
rect 7591 6326 7625 6360
rect 7671 6326 7705 6360
rect 7751 6326 7785 6360
rect 7831 6326 7865 6360
rect 7911 6326 7945 6360
rect 7991 6326 8025 6360
rect 8071 6326 8105 6360
rect 8151 6326 8185 6360
rect 8231 6326 8265 6360
rect 8311 6326 8345 6360
rect 8391 6326 8425 6360
rect 8471 6326 8505 6360
rect 8551 6326 8585 6360
rect 8631 6326 8665 6360
rect 8711 6326 8745 6360
rect 8791 6326 8825 6360
rect 8871 6326 8905 6360
rect 8951 6326 8985 6360
rect 9031 6326 9065 6360
rect 9111 6326 9145 6360
rect 9191 6326 9225 6360
rect 9271 6326 9305 6360
rect 9351 6326 9385 6360
rect 9431 6326 9465 6360
rect 9511 6326 9545 6360
rect 9591 6326 9625 6360
rect 9672 6326 9706 6360
rect 9752 6326 9786 6360
rect 9832 6326 9866 6360
rect 9912 6326 9946 6360
rect 9992 6326 10026 6360
rect 10072 6326 10106 6360
rect 10152 6326 10186 6360
rect 10232 6326 10266 6360
rect 10312 6326 10346 6360
rect 10392 6326 10426 6360
rect 10472 6326 10506 6360
rect 10552 6326 10586 6360
rect 10632 6326 10666 6360
rect 10712 6326 10746 6360
rect 10792 6326 10826 6360
rect 10872 6326 10906 6360
rect 10952 6326 10986 6360
rect 11032 6326 11066 6360
rect 11112 6326 11146 6360
rect 11192 6326 11226 6360
rect 11272 6326 11306 6360
rect 11352 6326 11386 6360
rect 11432 6326 11466 6360
rect 11512 6326 11546 6360
rect 11592 6326 11626 6360
rect 11672 6326 11706 6360
rect 11752 6326 11786 6360
rect 11832 6326 11866 6360
rect 11912 6326 11946 6360
rect 11992 6326 12026 6360
rect 12072 6326 12106 6360
rect 12152 6326 12186 6360
rect 12232 6326 12266 6360
rect 12312 6326 12346 6360
rect 12392 6326 12426 6360
rect 12472 6326 12506 6360
rect 12552 6326 12586 6360
rect 12632 6326 12666 6360
rect 12712 6326 12746 6360
rect 12792 6326 12826 6360
rect 12872 6326 12906 6360
rect 12952 6326 12986 6360
rect 13032 6326 13066 6360
rect 13112 6326 13146 6360
rect 13192 6326 13226 6360
rect 13272 6326 13306 6360
rect 13352 6326 13386 6360
rect 13432 6326 13466 6360
rect 13512 6326 13546 6360
rect 13592 6326 13626 6360
rect 13672 6326 13706 6360
rect 13752 6326 13786 6360
rect 13832 6326 13866 6360
rect 13912 6326 13946 6360
rect 13992 6326 14026 6360
rect 14072 6326 14106 6360
rect 14152 6326 14186 6360
rect 14232 6326 14266 6360
rect 14312 6326 14346 6360
rect 14392 6326 14426 6360
rect 14472 6326 14506 6360
rect 14552 6326 14586 6360
rect 14632 6326 14666 6360
rect 14712 6326 14746 6360
rect 14792 6326 14826 6360
rect 14872 6326 14906 6360
rect 14952 6326 14986 6360
rect 15032 6326 15066 6360
rect 15112 6326 15146 6360
rect 15192 6326 15226 6360
rect 15272 6326 15306 6360
rect 15352 6326 15386 6360
rect 15432 6326 15466 6360
rect 15512 6326 15546 6360
rect 15592 6326 15626 6360
rect 15672 6326 15706 6360
rect 15752 6326 15786 6360
rect 15832 6326 15866 6360
rect 15912 6326 15946 6360
rect 15992 6326 16026 6360
rect 16072 6326 16106 6360
rect 16152 6326 16186 6360
rect 16232 6326 16266 6360
rect 16312 6326 16346 6360
rect 16392 6326 16426 6360
rect 16472 6326 16506 6360
rect 16552 6326 16586 6360
rect 16632 6326 16666 6360
rect 16712 6326 16746 6360
rect 16792 6326 16826 6360
rect 16872 6326 16906 6360
rect 16952 6326 16986 6360
rect 17032 6326 17066 6360
rect 17112 6326 17146 6360
rect 17192 6326 17226 6360
rect 17272 6326 17306 6360
rect 17352 6326 17386 6360
rect 17432 6326 17466 6360
rect 17512 6326 17546 6360
rect 17592 6326 17626 6360
rect 17672 6326 17706 6360
rect 17752 6326 17786 6360
rect 17832 6326 17866 6360
rect 17912 6326 17946 6360
rect 17992 6326 18026 6360
rect 18072 6326 18106 6360
rect 18152 6326 18186 6360
rect 18232 6326 18266 6360
rect 18312 6326 18346 6360
rect 18392 6326 18426 6360
rect 18472 6326 18506 6360
rect 18552 6326 18586 6360
rect 18632 6326 18666 6360
rect 18712 6326 18746 6360
rect 18792 6326 18826 6360
rect 18872 6326 18906 6360
rect 18952 6326 18986 6360
rect 19032 6326 19066 6360
rect 19112 6326 19146 6360
rect 19192 6326 19226 6360
rect 19272 6326 19306 6360
rect 19352 6326 19386 6360
rect 19432 6326 19466 6360
rect 19512 6326 19546 6360
rect 19592 6326 19626 6360
rect 19672 6326 19706 6360
rect 19752 6326 19786 6360
rect 19832 6326 19866 6360
rect 19912 6326 19946 6360
rect 19992 6326 20026 6360
rect 20072 6326 20106 6360
rect 20152 6326 20186 6360
rect 20232 6326 20266 6360
rect 20312 6326 20346 6360
rect 20392 6326 20426 6360
rect 20472 6326 20506 6360
rect 20552 6326 20586 6360
rect 20632 6326 20666 6360
rect 20712 6326 20746 6360
rect 20792 6326 20826 6360
rect 20872 6326 20906 6360
rect 20952 6326 20986 6360
rect 21032 6326 21066 6360
rect 21112 6326 21146 6360
rect 21192 6326 21226 6360
rect 21272 6326 21306 6360
rect 21352 6326 21386 6360
rect 21432 6326 21466 6360
rect 21512 6326 21546 6360
rect 21592 6326 21626 6360
rect 21672 6326 21706 6360
rect 21752 6326 21786 6360
rect 21832 6326 21866 6360
rect 21912 6326 21946 6360
rect 21992 6326 22026 6360
rect 22072 6326 22106 6360
rect 22152 6326 22186 6360
rect 22232 6326 22266 6360
rect 22312 6326 22346 6360
rect 22392 6326 22426 6360
rect 22472 6326 22506 6360
rect 22552 6326 22586 6360
rect 22633 6326 22667 6360
rect 22713 6326 22747 6360
rect 22793 6326 22827 6360
rect 22873 6326 22907 6360
rect 22953 6326 22987 6360
rect 23033 6326 23067 6360
rect 23113 6326 23147 6360
rect 23193 6326 23227 6360
rect 23273 6326 23307 6360
rect 23353 6326 23387 6360
rect 23433 6326 23467 6360
rect 23513 6326 23547 6360
rect 23593 6326 23627 6360
rect 23673 6326 23707 6360
rect 23753 6326 23787 6360
rect 23833 6326 23867 6360
rect 23913 6326 23947 6360
rect 23993 6326 24027 6360
rect 24073 6326 24107 6360
rect 24153 6326 24187 6360
rect 24233 6326 24267 6360
rect 24313 6326 24347 6360
rect 24393 6326 24427 6360
rect 24473 6326 24507 6360
rect 24553 6326 24587 6360
rect 24633 6326 24667 6360
rect 24713 6326 24747 6360
rect 24793 6326 24827 6360
rect 24873 6326 24907 6360
rect 24953 6326 24987 6360
rect 25033 6326 25067 6360
rect 25113 6326 25147 6360
rect 25193 6326 25227 6360
rect 25273 6326 25307 6360
rect 25353 6326 25387 6360
rect 25433 6326 25467 6360
rect 25513 6326 25547 6360
rect 25593 6326 25627 6360
rect 25673 6326 25707 6360
rect 25753 6326 25787 6360
rect 25833 6326 25867 6360
rect 25913 6326 25947 6360
rect 25993 6326 26027 6360
rect 26073 6326 26107 6360
rect 26153 6326 26187 6360
rect 26233 6326 26267 6360
rect 26313 6326 26347 6360
rect 26393 6326 26427 6360
rect 26473 6326 26507 6360
rect 26553 6326 26587 6360
rect 26633 6326 26667 6360
rect 26713 6326 26747 6360
rect 26793 6326 26827 6360
rect 26873 6326 26907 6360
rect 26953 6326 26987 6360
rect 27033 6326 27067 6360
rect 27113 6326 27147 6360
rect 27193 6326 27227 6360
rect 27273 6326 27307 6360
rect 27353 6326 27387 6360
rect 27433 6326 27467 6360
rect 27513 6326 27547 6360
rect 27593 6326 27627 6360
rect 27673 6326 27707 6360
rect 27753 6326 27787 6360
rect 27833 6326 27867 6360
rect 27913 6326 27947 6360
rect 27993 6326 28027 6360
rect 28073 6326 28107 6360
rect 28153 6326 28187 6360
rect 28233 6326 28267 6360
rect 28313 6326 28347 6360
rect 28393 6326 28427 6360
rect 28473 6326 28507 6360
rect 28553 6326 28587 6360
rect 28633 6326 28667 6360
rect 28713 6326 28747 6360
rect 28793 6326 28827 6360
rect 28873 6326 28907 6360
rect 28953 6326 28987 6360
rect 29033 6326 29067 6360
rect 29113 6326 29147 6360
rect 29193 6326 29227 6360
rect 29273 6326 29307 6360
rect 29353 6326 29387 6360
rect 29433 6326 29467 6360
rect 29513 6326 29547 6360
rect 29593 6326 29627 6360
rect 29673 6326 29707 6360
rect 29753 6326 29787 6360
rect 29833 6326 29867 6360
rect 29913 6326 29947 6360
rect 29993 6326 30027 6360
rect 30073 6326 30107 6360
rect 30153 6326 30187 6360
rect 30233 6326 30267 6360
rect 30313 6326 30347 6360
rect 30393 6326 30427 6360
rect 30473 6326 30507 6360
rect 30553 6326 30587 6360
rect 30633 6326 30667 6360
rect 30713 6326 30747 6360
rect 30793 6326 30827 6360
rect 30873 6326 30907 6360
rect 30953 6326 30987 6360
rect 31033 6326 31067 6360
rect 31113 6326 31147 6360
rect 31193 6326 31227 6360
rect 31274 6326 31308 6360
rect 31354 6326 31388 6360
rect 31434 6326 31468 6360
rect 31514 6326 31548 6360
rect 31594 6326 31628 6360
rect 31674 6326 31708 6360
rect 31754 6326 31788 6360
rect 31834 6326 31868 6360
rect 31914 6326 31948 6360
rect 31994 6326 32028 6360
rect 32074 6326 32108 6360
rect 32154 6326 32188 6360
rect 32234 6326 32268 6360
rect 32314 6326 32348 6360
rect 32394 6326 32428 6360
rect 32474 6326 32508 6360
rect 32554 6326 32588 6360
rect 32634 6326 32668 6360
rect 32714 6326 32748 6360
rect 32794 6326 32828 6360
rect 32874 6326 32908 6360
rect 32954 6326 32988 6360
rect 33034 6326 33068 6360
rect 33114 6326 33148 6360
rect 33194 6326 33228 6360
rect 33274 6326 33308 6360
rect 33354 6326 33388 6360
rect 33434 6326 33468 6360
rect 33514 6326 33548 6360
rect 33594 6326 33628 6360
rect 33674 6326 33708 6360
rect 33754 6326 33788 6360
rect 33834 6326 33868 6360
rect 33914 6326 33948 6360
rect 33994 6326 34028 6360
rect 34074 6326 34108 6360
rect 34154 6326 34188 6360
rect 34234 6326 34268 6360
rect 34314 6326 34348 6360
rect 34394 6326 34428 6360
rect 34474 6326 34508 6360
rect 34554 6326 34588 6360
rect 34634 6326 34668 6360
rect 34714 6326 34748 6360
rect 34794 6326 34828 6360
rect 34874 6326 34908 6360
rect 34954 6326 34988 6360
rect 35034 6326 35068 6360
rect 35114 6326 35148 6360
rect 35194 6326 35228 6360
rect 35274 6326 35308 6360
rect 35354 6326 35388 6360
rect 35434 6326 35468 6360
rect 35514 6326 35548 6360
rect -34905 4787 -34871 4821
rect -34825 4787 -34791 4821
rect -34745 4787 -34711 4821
rect -34665 4787 -34631 4821
rect -34585 4787 -34551 4821
rect -34505 4787 -34471 4821
rect -34425 4787 -34391 4821
rect -34345 4787 -34311 4821
rect -34265 4787 -34231 4821
rect -34185 4787 -34151 4821
rect -34105 4787 -34071 4821
rect -34025 4787 -33991 4821
rect -33945 4787 -33911 4821
rect -33865 4787 -33831 4821
rect -33785 4787 -33751 4821
rect -33705 4787 -33671 4821
rect -33625 4787 -33591 4821
rect -33545 4787 -33511 4821
rect -33465 4787 -33431 4821
rect -33385 4787 -33351 4821
rect -33305 4787 -33271 4821
rect -33225 4787 -33191 4821
rect -33145 4787 -33111 4821
rect -33065 4787 -33031 4821
rect -32985 4787 -32951 4821
rect -32905 4787 -32871 4821
rect -32825 4787 -32791 4821
rect -32745 4787 -32711 4821
rect -32665 4787 -32631 4821
rect -32585 4787 -32551 4821
rect -32505 4787 -32471 4821
rect -32425 4787 -32391 4821
rect -32345 4787 -32311 4821
rect -32265 4787 -32231 4821
rect -32185 4787 -32151 4821
rect -32105 4787 -32071 4821
rect -32025 4787 -31991 4821
rect -31945 4787 -31911 4821
rect -31865 4787 -31831 4821
rect -31785 4787 -31751 4821
rect -31705 4787 -31671 4821
rect -31625 4787 -31591 4821
rect -31545 4787 -31511 4821
rect -31465 4787 -31431 4821
rect -31385 4787 -31351 4821
rect -31305 4787 -31271 4821
rect -31225 4787 -31191 4821
rect -31145 4787 -31111 4821
rect -31065 4787 -31031 4821
rect -30985 4787 -30951 4821
rect -30905 4787 -30871 4821
rect -30825 4787 -30791 4821
rect -30745 4787 -30711 4821
rect -30665 4787 -30631 4821
rect -30585 4787 -30551 4821
rect -30505 4787 -30471 4821
rect -30425 4787 -30391 4821
rect -30345 4787 -30311 4821
rect -30265 4787 -30231 4821
rect -30185 4787 -30151 4821
rect -30105 4787 -30071 4821
rect -30025 4787 -29991 4821
rect -29945 4787 -29911 4821
rect -29865 4787 -29831 4821
rect -29785 4787 -29751 4821
rect -29705 4787 -29671 4821
rect -29625 4787 -29591 4821
rect -29545 4787 -29511 4821
rect -29465 4787 -29431 4821
rect -29385 4787 -29351 4821
rect -29305 4787 -29271 4821
rect -29225 4787 -29191 4821
rect -29145 4787 -29111 4821
rect -29065 4787 -29031 4821
rect -28985 4787 -28951 4821
rect -28905 4787 -28871 4821
rect -28825 4787 -28791 4821
rect -28745 4787 -28711 4821
rect -28665 4787 -28631 4821
rect -28585 4787 -28551 4821
rect -28505 4787 -28471 4821
rect -28425 4787 -28391 4821
rect -28345 4787 -28311 4821
rect -28265 4787 -28231 4821
rect -28185 4787 -28151 4821
rect -28105 4787 -28071 4821
rect -28025 4787 -27991 4821
rect -27945 4787 -27911 4821
rect -27865 4787 -27831 4821
rect -27785 4787 -27751 4821
rect -27705 4787 -27671 4821
rect -27625 4787 -27591 4821
rect -27545 4787 -27511 4821
rect -27465 4787 -27431 4821
rect -27385 4787 -27351 4821
rect -27305 4787 -27271 4821
rect -27225 4787 -27191 4821
rect -27145 4787 -27111 4821
rect -27065 4787 -27031 4821
rect -26985 4787 -26951 4821
rect -26905 4787 -26871 4821
rect -26825 4787 -26791 4821
rect -26745 4787 -26711 4821
rect -26665 4787 -26631 4821
rect -26585 4787 -26551 4821
rect -26505 4787 -26471 4821
rect -26425 4787 -26391 4821
rect -26345 4787 -26311 4821
rect -26265 4787 -26231 4821
rect -26185 4787 -26151 4821
rect -26105 4787 -26071 4821
rect -26025 4787 -25991 4821
rect -25945 4787 -25911 4821
rect -25865 4787 -25831 4821
rect -25785 4787 -25751 4821
rect -25705 4787 -25671 4821
rect -25625 4787 -25591 4821
rect -25545 4787 -25511 4821
rect -25465 4787 -25431 4821
rect -25385 4787 -25351 4821
rect -25305 4787 -25271 4821
rect -25225 4787 -25191 4821
rect -25145 4787 -25111 4821
rect -25065 4787 -25031 4821
rect -24985 4787 -24951 4821
rect -24905 4787 -24871 4821
rect -24825 4787 -24791 4821
rect -24745 4787 -24711 4821
rect -24665 4787 -24631 4821
rect -24585 4787 -24551 4821
rect -24505 4787 -24471 4821
rect -24425 4787 -24391 4821
rect -24345 4787 -24311 4821
rect -24265 4787 -24231 4821
rect -24185 4787 -24151 4821
rect -24105 4787 -24071 4821
rect -24025 4787 -23991 4821
rect -23945 4787 -23911 4821
rect -23865 4787 -23831 4821
rect -23785 4787 -23751 4821
rect -23705 4787 -23671 4821
rect -23625 4787 -23591 4821
rect -23545 4787 -23511 4821
rect -23465 4787 -23431 4821
rect -23385 4787 -23351 4821
rect -23305 4787 -23271 4821
rect -23225 4787 -23191 4821
rect -23145 4787 -23111 4821
rect -23065 4787 -23031 4821
rect -22985 4787 -22951 4821
rect -22905 4787 -22871 4821
rect -22825 4787 -22791 4821
rect -22745 4787 -22711 4821
rect -22665 4787 -22631 4821
rect -22585 4787 -22551 4821
rect -22505 4787 -22471 4821
rect -22425 4787 -22391 4821
rect -22345 4787 -22311 4821
rect -22265 4787 -22231 4821
rect -22185 4787 -22151 4821
rect -22105 4787 -22071 4821
rect -22025 4787 -21991 4821
rect -21944 4787 -21910 4821
rect -21864 4787 -21830 4821
rect -21784 4787 -21750 4821
rect -21704 4787 -21670 4821
rect -21624 4787 -21590 4821
rect -21544 4787 -21510 4821
rect -21464 4787 -21430 4821
rect -21384 4787 -21350 4821
rect -21304 4787 -21270 4821
rect -21224 4787 -21190 4821
rect -21144 4787 -21110 4821
rect -21064 4787 -21030 4821
rect -20984 4787 -20950 4821
rect -20904 4787 -20870 4821
rect -20824 4787 -20790 4821
rect -20744 4787 -20710 4821
rect -20664 4787 -20630 4821
rect -20584 4787 -20550 4821
rect -20504 4787 -20470 4821
rect -20424 4787 -20390 4821
rect -20344 4787 -20310 4821
rect -20264 4787 -20230 4821
rect -20184 4787 -20150 4821
rect -20104 4787 -20070 4821
rect -20024 4787 -19990 4821
rect -19944 4787 -19910 4821
rect -19864 4787 -19830 4821
rect -19784 4787 -19750 4821
rect -19704 4787 -19670 4821
rect -19624 4787 -19590 4821
rect -19544 4787 -19510 4821
rect -19464 4787 -19430 4821
rect -19384 4787 -19350 4821
rect -19304 4787 -19270 4821
rect -19224 4787 -19190 4821
rect -19144 4787 -19110 4821
rect -19064 4787 -19030 4821
rect -18984 4787 -18950 4821
rect -18904 4787 -18870 4821
rect -18824 4787 -18790 4821
rect -18744 4787 -18710 4821
rect -18664 4787 -18630 4821
rect -18584 4787 -18550 4821
rect -18504 4787 -18470 4821
rect -18424 4787 -18390 4821
rect -18344 4787 -18310 4821
rect -18264 4787 -18230 4821
rect -18184 4787 -18150 4821
rect -18104 4787 -18070 4821
rect -18024 4787 -17990 4821
rect -17944 4787 -17910 4821
rect -17864 4787 -17830 4821
rect -17784 4787 -17750 4821
rect -17704 4787 -17670 4821
rect -17624 4787 -17590 4821
rect -17544 4787 -17510 4821
rect -17464 4787 -17430 4821
rect -17384 4787 -17350 4821
rect -17304 4787 -17270 4821
rect -17224 4787 -17190 4821
rect -17144 4787 -17110 4821
rect -17064 4787 -17030 4821
rect -16984 4787 -16950 4821
rect -16904 4787 -16870 4821
rect -16824 4787 -16790 4821
rect -16744 4787 -16710 4821
rect -16664 4787 -16630 4821
rect -16584 4787 -16550 4821
rect -16504 4787 -16470 4821
rect -16424 4787 -16390 4821
rect -16344 4787 -16310 4821
rect -16264 4787 -16230 4821
rect -16184 4787 -16150 4821
rect -16104 4787 -16070 4821
rect -16024 4787 -15990 4821
rect -15944 4787 -15910 4821
rect -15864 4787 -15830 4821
rect -15784 4787 -15750 4821
rect -15704 4787 -15670 4821
rect -15624 4787 -15590 4821
rect -15544 4787 -15510 4821
rect -15464 4787 -15430 4821
rect -15384 4787 -15350 4821
rect -15304 4787 -15270 4821
rect -15224 4787 -15190 4821
rect -15144 4787 -15110 4821
rect -15064 4787 -15030 4821
rect -14984 4787 -14950 4821
rect -14904 4787 -14870 4821
rect -14824 4787 -14790 4821
rect -14744 4787 -14710 4821
rect -14664 4787 -14630 4821
rect -14584 4787 -14550 4821
rect -14504 4787 -14470 4821
rect -14424 4787 -14390 4821
rect -14344 4787 -14310 4821
rect -14264 4787 -14230 4821
rect -14184 4787 -14150 4821
rect -14104 4787 -14070 4821
rect -14024 4787 -13990 4821
rect -13944 4787 -13910 4821
rect -13864 4787 -13830 4821
rect -13784 4787 -13750 4821
rect -13704 4787 -13670 4821
rect -13624 4787 -13590 4821
rect -13544 4787 -13510 4821
rect -13464 4787 -13430 4821
rect -13384 4787 -13350 4821
rect -13304 4787 -13270 4821
rect -13224 4787 -13190 4821
rect -13144 4787 -13110 4821
rect -13064 4787 -13030 4821
rect -12984 4787 -12950 4821
rect -12904 4787 -12870 4821
rect -12824 4787 -12790 4821
rect -12744 4787 -12710 4821
rect -12664 4787 -12630 4821
rect -12584 4787 -12550 4821
rect -12504 4787 -12470 4821
rect -12424 4787 -12390 4821
rect -12344 4787 -12310 4821
rect -12264 4787 -12230 4821
rect -12184 4787 -12150 4821
rect -12104 4787 -12070 4821
rect -12024 4787 -11990 4821
rect -11944 4787 -11910 4821
rect -11864 4787 -11830 4821
rect -11784 4787 -11750 4821
rect -11704 4787 -11670 4821
rect -11624 4787 -11590 4821
rect -11544 4787 -11510 4821
rect -11464 4787 -11430 4821
rect -11384 4787 -11350 4821
rect -11304 4787 -11270 4821
rect -11224 4787 -11190 4821
rect -11144 4787 -11110 4821
rect -11064 4787 -11030 4821
rect -10984 4787 -10950 4821
rect -10904 4787 -10870 4821
rect -10824 4787 -10790 4821
rect -10744 4787 -10710 4821
rect -10664 4787 -10630 4821
rect -10584 4787 -10550 4821
rect -10504 4787 -10470 4821
rect -10424 4787 -10390 4821
rect -10344 4787 -10310 4821
rect -10264 4787 -10230 4821
rect -10184 4787 -10150 4821
rect -10104 4787 -10070 4821
rect -10024 4787 -9990 4821
rect -9944 4787 -9910 4821
rect -9864 4787 -9830 4821
rect -9784 4787 -9750 4821
rect -9704 4787 -9670 4821
rect -9624 4787 -9590 4821
rect -9544 4787 -9510 4821
rect -9464 4787 -9430 4821
rect -9384 4787 -9350 4821
rect -9304 4787 -9270 4821
rect -9224 4787 -9190 4821
rect -9144 4787 -9110 4821
rect -9064 4787 -9030 4821
rect -8983 4787 -8949 4821
rect -8903 4787 -8869 4821
rect -8823 4787 -8789 4821
rect -8743 4787 -8709 4821
rect -8663 4787 -8629 4821
rect -8583 4787 -8549 4821
rect -8503 4787 -8469 4821
rect -8423 4787 -8389 4821
rect -8343 4787 -8309 4821
rect -8263 4787 -8229 4821
rect -8183 4787 -8149 4821
rect -8103 4787 -8069 4821
rect -8023 4787 -7989 4821
rect -7943 4787 -7909 4821
rect -7863 4787 -7829 4821
rect -7783 4787 -7749 4821
rect -7703 4787 -7669 4821
rect -7623 4787 -7589 4821
rect -7543 4787 -7509 4821
rect -7463 4787 -7429 4821
rect -7383 4787 -7349 4821
rect -7303 4787 -7269 4821
rect -7223 4787 -7189 4821
rect -7143 4787 -7109 4821
rect -7063 4787 -7029 4821
rect -6983 4787 -6949 4821
rect -6903 4787 -6869 4821
rect -6823 4787 -6789 4821
rect -6743 4787 -6709 4821
rect -6663 4787 -6629 4821
rect -6583 4787 -6549 4821
rect -6503 4787 -6469 4821
rect -6423 4787 -6389 4821
rect -6343 4787 -6309 4821
rect -6263 4787 -6229 4821
rect -6183 4787 -6149 4821
rect -6103 4787 -6069 4821
rect -6023 4787 -5989 4821
rect -5943 4787 -5909 4821
rect -5863 4787 -5829 4821
rect -5783 4787 -5749 4821
rect -5703 4787 -5669 4821
rect -5623 4787 -5589 4821
rect -5543 4787 -5509 4821
rect -5463 4787 -5429 4821
rect -5383 4787 -5349 4821
rect -5303 4787 -5269 4821
rect -5223 4787 -5189 4821
rect -5143 4787 -5109 4821
rect -5063 4787 -5029 4821
rect -4983 4787 -4949 4821
rect -4903 4787 -4869 4821
rect -4823 4787 -4789 4821
rect -4743 4787 -4709 4821
rect -4663 4787 -4629 4821
rect -4583 4787 -4549 4821
rect -4503 4787 -4469 4821
rect -4423 4787 -4389 4821
rect -4343 4787 -4309 4821
rect -4263 4787 -4229 4821
rect -4183 4787 -4149 4821
rect -4103 4787 -4069 4821
rect -4023 4787 -3989 4821
rect -3943 4787 -3909 4821
rect -3863 4787 -3829 4821
rect -3783 4787 -3749 4821
rect -3703 4787 -3669 4821
rect -3623 4787 -3589 4821
rect -3543 4787 -3509 4821
rect -3463 4787 -3429 4821
rect -3383 4787 -3349 4821
rect -3303 4787 -3269 4821
rect -3223 4787 -3189 4821
rect -3143 4787 -3109 4821
rect -3063 4787 -3029 4821
rect -2983 4787 -2949 4821
rect -2903 4787 -2869 4821
rect -2823 4787 -2789 4821
rect -2743 4787 -2709 4821
rect -2663 4787 -2629 4821
rect -2583 4787 -2549 4821
rect -2503 4787 -2469 4821
rect -2423 4787 -2389 4821
rect -2343 4787 -2309 4821
rect -2263 4787 -2229 4821
rect -2183 4787 -2149 4821
rect -2103 4787 -2069 4821
rect -2023 4787 -1989 4821
rect -1943 4787 -1909 4821
rect -1863 4787 -1829 4821
rect -1783 4787 -1749 4821
rect -1703 4787 -1669 4821
rect -1623 4787 -1589 4821
rect -1543 4787 -1509 4821
rect -1463 4787 -1429 4821
rect -1383 4787 -1349 4821
rect -1303 4787 -1269 4821
rect -1223 4787 -1189 4821
rect -1143 4787 -1109 4821
rect -1063 4787 -1029 4821
rect -983 4787 -949 4821
rect -903 4787 -869 4821
rect -823 4787 -789 4821
rect -743 4787 -709 4821
rect -663 4787 -629 4821
rect -583 4787 -549 4821
rect -503 4787 -469 4821
rect -423 4787 -389 4821
rect 1681 4787 1715 4821
rect 1761 4787 1795 4821
rect 1841 4787 1875 4821
rect 1921 4787 1955 4821
rect 2001 4787 2035 4821
rect 2081 4787 2115 4821
rect 2161 4787 2195 4821
rect 2241 4787 2275 4821
rect 2321 4787 2355 4821
rect 2401 4787 2435 4821
rect 2481 4787 2515 4821
rect 2561 4787 2595 4821
rect 2641 4787 2675 4821
rect 2721 4787 2755 4821
rect 2801 4787 2835 4821
rect 2881 4787 2915 4821
rect 2961 4787 2995 4821
rect 3041 4787 3075 4821
rect 3121 4787 3155 4821
rect 3201 4787 3235 4821
rect 3281 4787 3315 4821
rect 3361 4787 3395 4821
rect 3441 4787 3475 4821
rect 3521 4787 3555 4821
rect 3601 4787 3635 4821
rect 3681 4787 3715 4821
rect 3761 4787 3795 4821
rect 3841 4787 3875 4821
rect 3921 4787 3955 4821
rect 4001 4787 4035 4821
rect 4081 4787 4115 4821
rect 4161 4787 4195 4821
rect 4241 4787 4275 4821
rect 4321 4787 4355 4821
rect 4401 4787 4435 4821
rect 4481 4787 4515 4821
rect 4561 4787 4595 4821
rect 4641 4787 4675 4821
rect 4721 4787 4755 4821
rect 4801 4787 4835 4821
rect 4881 4787 4915 4821
rect 4961 4787 4995 4821
rect 5041 4787 5075 4821
rect 5121 4787 5155 4821
rect 5201 4787 5235 4821
rect 5281 4787 5315 4821
rect 5361 4787 5395 4821
rect 5441 4787 5475 4821
rect 5521 4787 5555 4821
rect 5601 4787 5635 4821
rect 5681 4787 5715 4821
rect 5761 4787 5795 4821
rect 5841 4787 5875 4821
rect 5921 4787 5955 4821
rect 6001 4787 6035 4821
rect 6081 4787 6115 4821
rect 6161 4787 6195 4821
rect 6241 4787 6275 4821
rect 6321 4787 6355 4821
rect 6401 4787 6435 4821
rect 6481 4787 6515 4821
rect 6561 4787 6595 4821
rect 6641 4787 6675 4821
rect 6721 4787 6755 4821
rect 6801 4787 6835 4821
rect 6881 4787 6915 4821
rect 6961 4787 6995 4821
rect 7041 4787 7075 4821
rect 7121 4787 7155 4821
rect 7201 4787 7235 4821
rect 7281 4787 7315 4821
rect 7361 4787 7395 4821
rect 7441 4787 7475 4821
rect 7521 4787 7555 4821
rect 7601 4787 7635 4821
rect 7681 4787 7715 4821
rect 7761 4787 7795 4821
rect 7841 4787 7875 4821
rect 7921 4787 7955 4821
rect 8001 4787 8035 4821
rect 8081 4787 8115 4821
rect 8161 4787 8195 4821
rect 8241 4787 8275 4821
rect 8321 4787 8355 4821
rect 8401 4787 8435 4821
rect 8481 4787 8515 4821
rect 8561 4787 8595 4821
rect 8641 4787 8675 4821
rect 8721 4787 8755 4821
rect 8801 4787 8835 4821
rect 8881 4787 8915 4821
rect 8961 4787 8995 4821
rect 9041 4787 9075 4821
rect 9121 4787 9155 4821
rect 9201 4787 9235 4821
rect 9281 4787 9315 4821
rect 9361 4787 9395 4821
rect 9441 4787 9475 4821
rect 9521 4787 9555 4821
rect 9601 4787 9635 4821
rect 9681 4787 9715 4821
rect 9761 4787 9795 4821
rect 9841 4787 9875 4821
rect 9921 4787 9955 4821
rect 10001 4787 10035 4821
rect 10081 4787 10115 4821
rect 10161 4787 10195 4821
rect 10241 4787 10275 4821
rect 10321 4787 10355 4821
rect 10401 4787 10435 4821
rect 10481 4787 10515 4821
rect 10561 4787 10595 4821
rect 10641 4787 10675 4821
rect 10721 4787 10755 4821
rect 10801 4787 10835 4821
rect 10881 4787 10915 4821
rect 10961 4787 10995 4821
rect 11041 4787 11075 4821
rect 11121 4787 11155 4821
rect 11201 4787 11235 4821
rect 11281 4787 11315 4821
rect 11361 4787 11395 4821
rect 11441 4787 11475 4821
rect 11521 4787 11555 4821
rect 11601 4787 11635 4821
rect 11681 4787 11715 4821
rect 11761 4787 11795 4821
rect 11841 4787 11875 4821
rect 11921 4787 11955 4821
rect 12001 4787 12035 4821
rect 12081 4787 12115 4821
rect 12161 4787 12195 4821
rect 12241 4787 12275 4821
rect 12321 4787 12355 4821
rect 12401 4787 12435 4821
rect 12481 4787 12515 4821
rect 12561 4787 12595 4821
rect 12641 4787 12675 4821
rect 12721 4787 12755 4821
rect 12801 4787 12835 4821
rect 12881 4787 12915 4821
rect 12961 4787 12995 4821
rect 13041 4787 13075 4821
rect 13121 4787 13155 4821
rect 13201 4787 13235 4821
rect 13281 4787 13315 4821
rect 13361 4787 13395 4821
rect 13441 4787 13475 4821
rect 13521 4787 13555 4821
rect 13601 4787 13635 4821
rect 13681 4787 13715 4821
rect 13761 4787 13795 4821
rect 13841 4787 13875 4821
rect 13921 4787 13955 4821
rect 14001 4787 14035 4821
rect 14081 4787 14115 4821
rect 14161 4787 14195 4821
rect 14241 4787 14275 4821
rect 14321 4787 14355 4821
rect 14401 4787 14435 4821
rect 14481 4787 14515 4821
rect 14561 4787 14595 4821
rect 14642 4787 14676 4821
rect 14722 4787 14756 4821
rect 14802 4787 14836 4821
rect 14882 4787 14916 4821
rect 14962 4787 14996 4821
rect 15042 4787 15076 4821
rect 15122 4787 15156 4821
rect 15202 4787 15236 4821
rect 15282 4787 15316 4821
rect 15362 4787 15396 4821
rect 15442 4787 15476 4821
rect 15522 4787 15556 4821
rect 15602 4787 15636 4821
rect 15682 4787 15716 4821
rect 15762 4787 15796 4821
rect 15842 4787 15876 4821
rect 15922 4787 15956 4821
rect 16002 4787 16036 4821
rect 16082 4787 16116 4821
rect 16162 4787 16196 4821
rect 16242 4787 16276 4821
rect 16322 4787 16356 4821
rect 16402 4787 16436 4821
rect 16482 4787 16516 4821
rect 16562 4787 16596 4821
rect 16642 4787 16676 4821
rect 16722 4787 16756 4821
rect 16802 4787 16836 4821
rect 16882 4787 16916 4821
rect 16962 4787 16996 4821
rect 17042 4787 17076 4821
rect 17122 4787 17156 4821
rect 17202 4787 17236 4821
rect 17282 4787 17316 4821
rect 17362 4787 17396 4821
rect 17442 4787 17476 4821
rect 17522 4787 17556 4821
rect 17602 4787 17636 4821
rect 17682 4787 17716 4821
rect 17762 4787 17796 4821
rect 17842 4787 17876 4821
rect 17922 4787 17956 4821
rect 18002 4787 18036 4821
rect 18082 4787 18116 4821
rect 18162 4787 18196 4821
rect 18242 4787 18276 4821
rect 18322 4787 18356 4821
rect 18402 4787 18436 4821
rect 18482 4787 18516 4821
rect 18562 4787 18596 4821
rect 18642 4787 18676 4821
rect 18722 4787 18756 4821
rect 18802 4787 18836 4821
rect 18882 4787 18916 4821
rect 18962 4787 18996 4821
rect 19042 4787 19076 4821
rect 19122 4787 19156 4821
rect 19202 4787 19236 4821
rect 19282 4787 19316 4821
rect 19362 4787 19396 4821
rect 19442 4787 19476 4821
rect 19522 4787 19556 4821
rect 19602 4787 19636 4821
rect 19682 4787 19716 4821
rect 19762 4787 19796 4821
rect 19842 4787 19876 4821
rect 19922 4787 19956 4821
rect 20002 4787 20036 4821
rect 20082 4787 20116 4821
rect 20162 4787 20196 4821
rect 20242 4787 20276 4821
rect 20322 4787 20356 4821
rect 20402 4787 20436 4821
rect 20482 4787 20516 4821
rect 20562 4787 20596 4821
rect 20642 4787 20676 4821
rect 20722 4787 20756 4821
rect 20802 4787 20836 4821
rect 20882 4787 20916 4821
rect 20962 4787 20996 4821
rect 21042 4787 21076 4821
rect 21122 4787 21156 4821
rect 21202 4787 21236 4821
rect 21282 4787 21316 4821
rect 21362 4787 21396 4821
rect 21442 4787 21476 4821
rect 21522 4787 21556 4821
rect 21602 4787 21636 4821
rect 21682 4787 21716 4821
rect 21762 4787 21796 4821
rect 21842 4787 21876 4821
rect 21922 4787 21956 4821
rect 22002 4787 22036 4821
rect 22082 4787 22116 4821
rect 22162 4787 22196 4821
rect 22242 4787 22276 4821
rect 22322 4787 22356 4821
rect 22402 4787 22436 4821
rect 22482 4787 22516 4821
rect 22562 4787 22596 4821
rect 22642 4787 22676 4821
rect 22722 4787 22756 4821
rect 22802 4787 22836 4821
rect 22882 4787 22916 4821
rect 22962 4787 22996 4821
rect 23042 4787 23076 4821
rect 23122 4787 23156 4821
rect 23202 4787 23236 4821
rect 23282 4787 23316 4821
rect 23362 4787 23396 4821
rect 23442 4787 23476 4821
rect 23522 4787 23556 4821
rect 23602 4787 23636 4821
rect 23682 4787 23716 4821
rect 23762 4787 23796 4821
rect 23842 4787 23876 4821
rect 23922 4787 23956 4821
rect 24002 4787 24036 4821
rect 24082 4787 24116 4821
rect 24162 4787 24196 4821
rect 24242 4787 24276 4821
rect 24322 4787 24356 4821
rect 24402 4787 24436 4821
rect 24482 4787 24516 4821
rect 24562 4787 24596 4821
rect 24642 4787 24676 4821
rect 24722 4787 24756 4821
rect 24802 4787 24836 4821
rect 24882 4787 24916 4821
rect 24962 4787 24996 4821
rect 25042 4787 25076 4821
rect 25122 4787 25156 4821
rect 25202 4787 25236 4821
rect 25282 4787 25316 4821
rect 25362 4787 25396 4821
rect 25442 4787 25476 4821
rect 25522 4787 25556 4821
rect 25602 4787 25636 4821
rect 25682 4787 25716 4821
rect 25762 4787 25796 4821
rect 25842 4787 25876 4821
rect 25922 4787 25956 4821
rect 26002 4787 26036 4821
rect 26082 4787 26116 4821
rect 26162 4787 26196 4821
rect 26242 4787 26276 4821
rect 26322 4787 26356 4821
rect 26402 4787 26436 4821
rect 26482 4787 26516 4821
rect 26562 4787 26596 4821
rect 26642 4787 26676 4821
rect 26722 4787 26756 4821
rect 26802 4787 26836 4821
rect 26882 4787 26916 4821
rect 26962 4787 26996 4821
rect 27042 4787 27076 4821
rect 27122 4787 27156 4821
rect 27202 4787 27236 4821
rect 27282 4787 27316 4821
rect 27362 4787 27396 4821
rect 27442 4787 27476 4821
rect 27522 4787 27556 4821
rect 27603 4787 27637 4821
rect 27683 4787 27717 4821
rect 27763 4787 27797 4821
rect 27843 4787 27877 4821
rect 27923 4787 27957 4821
rect 28003 4787 28037 4821
rect 28083 4787 28117 4821
rect 28163 4787 28197 4821
rect 28243 4787 28277 4821
rect 28323 4787 28357 4821
rect 28403 4787 28437 4821
rect 28483 4787 28517 4821
rect 28563 4787 28597 4821
rect 28643 4787 28677 4821
rect 28723 4787 28757 4821
rect 28803 4787 28837 4821
rect 28883 4787 28917 4821
rect 28963 4787 28997 4821
rect 29043 4787 29077 4821
rect 29123 4787 29157 4821
rect 29203 4787 29237 4821
rect 29283 4787 29317 4821
rect 29363 4787 29397 4821
rect 29443 4787 29477 4821
rect 29523 4787 29557 4821
rect 29603 4787 29637 4821
rect 29683 4787 29717 4821
rect 29763 4787 29797 4821
rect 29843 4787 29877 4821
rect 29923 4787 29957 4821
rect 30003 4787 30037 4821
rect 30083 4787 30117 4821
rect 30163 4787 30197 4821
rect 30243 4787 30277 4821
rect 30323 4787 30357 4821
rect 30403 4787 30437 4821
rect 30483 4787 30517 4821
rect 30563 4787 30597 4821
rect 30643 4787 30677 4821
rect 30723 4787 30757 4821
rect 30803 4787 30837 4821
rect 30883 4787 30917 4821
rect 30963 4787 30997 4821
rect 31043 4787 31077 4821
rect 31123 4787 31157 4821
rect 31203 4787 31237 4821
rect 31283 4787 31317 4821
rect 31363 4787 31397 4821
rect 31443 4787 31477 4821
rect 31523 4787 31557 4821
rect 31603 4787 31637 4821
rect 31683 4787 31717 4821
rect 31763 4787 31797 4821
rect 31843 4787 31877 4821
rect 31923 4787 31957 4821
rect 32003 4787 32037 4821
rect 32083 4787 32117 4821
rect 32163 4787 32197 4821
rect 32243 4787 32277 4821
rect 32323 4787 32357 4821
rect 32403 4787 32437 4821
rect 32483 4787 32517 4821
rect 32563 4787 32597 4821
rect 32643 4787 32677 4821
rect 32723 4787 32757 4821
rect 32803 4787 32837 4821
rect 32883 4787 32917 4821
rect 32963 4787 32997 4821
rect 33043 4787 33077 4821
rect 33123 4787 33157 4821
rect 33203 4787 33237 4821
rect 33283 4787 33317 4821
rect 33363 4787 33397 4821
rect 33443 4787 33477 4821
rect 33523 4787 33557 4821
rect 33603 4787 33637 4821
rect 33683 4787 33717 4821
rect 33763 4787 33797 4821
rect 33843 4787 33877 4821
rect 33923 4787 33957 4821
rect 34003 4787 34037 4821
rect 34083 4787 34117 4821
rect 34163 4787 34197 4821
rect 34243 4787 34277 4821
rect 34323 4787 34357 4821
rect 34403 4787 34437 4821
rect 34483 4787 34517 4821
rect 34563 4787 34597 4821
rect 34643 4787 34677 4821
rect 34723 4787 34757 4821
rect 34803 4787 34837 4821
rect 34883 4787 34917 4821
rect 34963 4787 34997 4821
rect 35043 4787 35077 4821
rect 35123 4787 35157 4821
rect 35203 4787 35237 4821
rect 35283 4787 35317 4821
rect 35363 4787 35397 4821
rect 35443 4787 35477 4821
rect 35523 4787 35557 4821
rect 35603 4787 35637 4821
rect 35683 4787 35717 4821
rect 35763 4787 35797 4821
rect 35843 4787 35877 4821
rect 35923 4787 35957 4821
rect 36003 4787 36037 4821
rect 36083 4787 36117 4821
rect 36163 4787 36197 4821
<< metal1 >>
rect -37898 17197 -3290 17230
rect -37898 17163 -37852 17197
rect -37818 17163 -37772 17197
rect -37738 17163 -37692 17197
rect -37658 17163 -37612 17197
rect -37578 17163 -37532 17197
rect -37498 17163 -37452 17197
rect -37418 17163 -37372 17197
rect -37338 17163 -37292 17197
rect -37258 17163 -37212 17197
rect -37178 17163 -37132 17197
rect -37098 17163 -37052 17197
rect -37018 17163 -36972 17197
rect -36938 17163 -36892 17197
rect -36858 17163 -36812 17197
rect -36778 17163 -36732 17197
rect -36698 17163 -36652 17197
rect -36618 17163 -36572 17197
rect -36538 17163 -36492 17197
rect -36458 17163 -36412 17197
rect -36378 17163 -36332 17197
rect -36298 17163 -36252 17197
rect -36218 17163 -36172 17197
rect -36138 17163 -36092 17197
rect -36058 17163 -36012 17197
rect -35978 17163 -35932 17197
rect -35898 17163 -35852 17197
rect -35818 17163 -35772 17197
rect -35738 17163 -35692 17197
rect -35658 17163 -35612 17197
rect -35578 17163 -35532 17197
rect -35498 17163 -35452 17197
rect -35418 17163 -35372 17197
rect -35338 17163 -35292 17197
rect -35258 17163 -35212 17197
rect -35178 17163 -35132 17197
rect -35098 17163 -35052 17197
rect -35018 17163 -34972 17197
rect -34938 17163 -34892 17197
rect -34858 17163 -34812 17197
rect -34778 17163 -34732 17197
rect -34698 17163 -34652 17197
rect -34618 17163 -34572 17197
rect -34538 17163 -34492 17197
rect -34458 17163 -34412 17197
rect -34378 17163 -34332 17197
rect -34298 17163 -34252 17197
rect -34218 17163 -34172 17197
rect -34138 17163 -34092 17197
rect -34058 17163 -34012 17197
rect -33978 17163 -33932 17197
rect -33898 17163 -33852 17197
rect -33818 17163 -33772 17197
rect -33738 17163 -33692 17197
rect -33658 17163 -33612 17197
rect -33578 17163 -33532 17197
rect -33498 17163 -33452 17197
rect -33418 17163 -33372 17197
rect -33338 17163 -33292 17197
rect -33258 17163 -33212 17197
rect -33178 17163 -33132 17197
rect -33098 17163 -33052 17197
rect -33018 17163 -32972 17197
rect -32938 17163 -32892 17197
rect -32858 17163 -32812 17197
rect -32778 17163 -32732 17197
rect -32698 17163 -32652 17197
rect -32618 17163 -32572 17197
rect -32538 17163 -32492 17197
rect -32458 17163 -32412 17197
rect -32378 17163 -32332 17197
rect -32298 17163 -32252 17197
rect -32218 17163 -32172 17197
rect -32138 17163 -32092 17197
rect -32058 17163 -32012 17197
rect -31978 17163 -31932 17197
rect -31898 17163 -31852 17197
rect -31818 17163 -31772 17197
rect -31738 17163 -31692 17197
rect -31658 17163 -31612 17197
rect -31578 17163 -31532 17197
rect -31498 17163 -31452 17197
rect -31418 17163 -31372 17197
rect -31338 17163 -31292 17197
rect -31258 17163 -31212 17197
rect -31178 17163 -31132 17197
rect -31098 17163 -31052 17197
rect -31018 17163 -30972 17197
rect -30938 17163 -30892 17197
rect -30858 17163 -30812 17197
rect -30778 17163 -30732 17197
rect -30698 17163 -30652 17197
rect -30618 17163 -30572 17197
rect -30538 17163 -30492 17197
rect -30458 17163 -30412 17197
rect -30378 17163 -30332 17197
rect -30298 17163 -30252 17197
rect -30218 17163 -30172 17197
rect -30138 17163 -30092 17197
rect -30058 17163 -30012 17197
rect -29978 17163 -29932 17197
rect -29898 17163 -29852 17197
rect -29818 17163 -29772 17197
rect -29738 17163 -29692 17197
rect -29658 17163 -29612 17197
rect -29578 17163 -29532 17197
rect -29498 17163 -29452 17197
rect -29418 17163 -29372 17197
rect -29338 17163 -29292 17197
rect -29258 17163 -29212 17197
rect -29178 17163 -29132 17197
rect -29098 17163 -29052 17197
rect -29018 17163 -28972 17197
rect -28938 17163 -28892 17197
rect -28858 17163 -28812 17197
rect -28778 17163 -28732 17197
rect -28698 17163 -28652 17197
rect -28618 17163 -28572 17197
rect -28538 17163 -28492 17197
rect -28458 17163 -28412 17197
rect -28378 17163 -28332 17197
rect -28298 17163 -28252 17197
rect -28218 17163 -28172 17197
rect -28138 17163 -28092 17197
rect -28058 17163 -28012 17197
rect -27978 17163 -27932 17197
rect -27898 17163 -27852 17197
rect -27818 17163 -27772 17197
rect -27738 17163 -27692 17197
rect -27658 17163 -27612 17197
rect -27578 17163 -27532 17197
rect -27498 17163 -27452 17197
rect -27418 17163 -27372 17197
rect -27338 17163 -27292 17197
rect -27258 17163 -27212 17197
rect -27178 17163 -27132 17197
rect -27098 17163 -27052 17197
rect -27018 17163 -26972 17197
rect -26938 17163 -26892 17197
rect -26858 17163 -26812 17197
rect -26778 17163 -26732 17197
rect -26698 17163 -26652 17197
rect -26618 17163 -26572 17197
rect -26538 17163 -26492 17197
rect -26458 17163 -26412 17197
rect -26378 17163 -26332 17197
rect -26298 17163 -26252 17197
rect -26218 17163 -26172 17197
rect -26138 17163 -26092 17197
rect -26058 17163 -26012 17197
rect -25978 17163 -25932 17197
rect -25898 17163 -25852 17197
rect -25818 17163 -25772 17197
rect -25738 17163 -25692 17197
rect -25658 17163 -25612 17197
rect -25578 17163 -25532 17197
rect -25498 17163 -25452 17197
rect -25418 17163 -25372 17197
rect -25338 17163 -25292 17197
rect -25258 17163 -25212 17197
rect -25178 17163 -25132 17197
rect -25098 17163 -25052 17197
rect -25018 17163 -24972 17197
rect -24938 17163 -24891 17197
rect -24857 17163 -24811 17197
rect -24777 17163 -24731 17197
rect -24697 17163 -24651 17197
rect -24617 17163 -24571 17197
rect -24537 17163 -24491 17197
rect -24457 17163 -24411 17197
rect -24377 17163 -24331 17197
rect -24297 17163 -24251 17197
rect -24217 17163 -24171 17197
rect -24137 17163 -24091 17197
rect -24057 17163 -24011 17197
rect -23977 17163 -23931 17197
rect -23897 17163 -23851 17197
rect -23817 17163 -23771 17197
rect -23737 17163 -23691 17197
rect -23657 17163 -23611 17197
rect -23577 17163 -23531 17197
rect -23497 17163 -23451 17197
rect -23417 17163 -23371 17197
rect -23337 17163 -23291 17197
rect -23257 17163 -23211 17197
rect -23177 17163 -23131 17197
rect -23097 17163 -23051 17197
rect -23017 17163 -22971 17197
rect -22937 17163 -22891 17197
rect -22857 17163 -22811 17197
rect -22777 17163 -22731 17197
rect -22697 17163 -22651 17197
rect -22617 17163 -22571 17197
rect -22537 17163 -22491 17197
rect -22457 17163 -22411 17197
rect -22377 17163 -22331 17197
rect -22297 17163 -22251 17197
rect -22217 17163 -22171 17197
rect -22137 17163 -22091 17197
rect -22057 17163 -22011 17197
rect -21977 17163 -21931 17197
rect -21897 17163 -21851 17197
rect -21817 17163 -21771 17197
rect -21737 17163 -21691 17197
rect -21657 17163 -21611 17197
rect -21577 17163 -21531 17197
rect -21497 17163 -21451 17197
rect -21417 17163 -21371 17197
rect -21337 17163 -21291 17197
rect -21257 17163 -21211 17197
rect -21177 17163 -21131 17197
rect -21097 17163 -21051 17197
rect -21017 17163 -20971 17197
rect -20937 17163 -20891 17197
rect -20857 17163 -20811 17197
rect -20777 17163 -20731 17197
rect -20697 17163 -20651 17197
rect -20617 17163 -20571 17197
rect -20537 17163 -20491 17197
rect -20457 17163 -20411 17197
rect -20377 17163 -20331 17197
rect -20297 17163 -20251 17197
rect -20217 17163 -20171 17197
rect -20137 17163 -20091 17197
rect -20057 17163 -20011 17197
rect -19977 17163 -19931 17197
rect -19897 17163 -19851 17197
rect -19817 17163 -19771 17197
rect -19737 17163 -19691 17197
rect -19657 17163 -19611 17197
rect -19577 17163 -19531 17197
rect -19497 17163 -19451 17197
rect -19417 17163 -19371 17197
rect -19337 17163 -19291 17197
rect -19257 17163 -19211 17197
rect -19177 17163 -19131 17197
rect -19097 17163 -19051 17197
rect -19017 17163 -18971 17197
rect -18937 17163 -18891 17197
rect -18857 17163 -18811 17197
rect -18777 17163 -18731 17197
rect -18697 17163 -18651 17197
rect -18617 17163 -18571 17197
rect -18537 17163 -18491 17197
rect -18457 17163 -18411 17197
rect -18377 17163 -18331 17197
rect -18297 17163 -18251 17197
rect -18217 17163 -18171 17197
rect -18137 17163 -18091 17197
rect -18057 17163 -18011 17197
rect -17977 17163 -17931 17197
rect -17897 17163 -17851 17197
rect -17817 17163 -17771 17197
rect -17737 17163 -17691 17197
rect -17657 17163 -17611 17197
rect -17577 17163 -17531 17197
rect -17497 17163 -17451 17197
rect -17417 17163 -17371 17197
rect -17337 17163 -17291 17197
rect -17257 17163 -17211 17197
rect -17177 17163 -17131 17197
rect -17097 17163 -17051 17197
rect -17017 17163 -16971 17197
rect -16937 17163 -16891 17197
rect -16857 17163 -16811 17197
rect -16777 17163 -16731 17197
rect -16697 17163 -16651 17197
rect -16617 17163 -16571 17197
rect -16537 17163 -16491 17197
rect -16457 17163 -16411 17197
rect -16377 17163 -16331 17197
rect -16297 17163 -16251 17197
rect -16217 17163 -16171 17197
rect -16137 17163 -16091 17197
rect -16057 17163 -16011 17197
rect -15977 17163 -15931 17197
rect -15897 17163 -15851 17197
rect -15817 17163 -15771 17197
rect -15737 17163 -15691 17197
rect -15657 17163 -15611 17197
rect -15577 17163 -15531 17197
rect -15497 17163 -15451 17197
rect -15417 17163 -15371 17197
rect -15337 17163 -15291 17197
rect -15257 17163 -15211 17197
rect -15177 17163 -15131 17197
rect -15097 17163 -15051 17197
rect -15017 17163 -14971 17197
rect -14937 17163 -14891 17197
rect -14857 17163 -14811 17197
rect -14777 17163 -14731 17197
rect -14697 17163 -14651 17197
rect -14617 17163 -14571 17197
rect -14537 17163 -14491 17197
rect -14457 17163 -14411 17197
rect -14377 17163 -14331 17197
rect -14297 17163 -14251 17197
rect -14217 17163 -14171 17197
rect -14137 17163 -14091 17197
rect -14057 17163 -14011 17197
rect -13977 17163 -13931 17197
rect -13897 17163 -13851 17197
rect -13817 17163 -13771 17197
rect -13737 17163 -13691 17197
rect -13657 17163 -13611 17197
rect -13577 17163 -13531 17197
rect -13497 17163 -13451 17197
rect -13417 17163 -13371 17197
rect -13337 17163 -13291 17197
rect -13257 17163 -13211 17197
rect -13177 17163 -13131 17197
rect -13097 17163 -13051 17197
rect -13017 17163 -12971 17197
rect -12937 17163 -12891 17197
rect -12857 17163 -12811 17197
rect -12777 17163 -12731 17197
rect -12697 17163 -12651 17197
rect -12617 17163 -12571 17197
rect -12537 17163 -12491 17197
rect -12457 17163 -12411 17197
rect -12377 17163 -12331 17197
rect -12297 17163 -12251 17197
rect -12217 17163 -12171 17197
rect -12137 17163 -12091 17197
rect -12057 17163 -12011 17197
rect -11977 17163 -11930 17197
rect -11896 17163 -11850 17197
rect -11816 17163 -11770 17197
rect -11736 17163 -11690 17197
rect -11656 17163 -11610 17197
rect -11576 17163 -11530 17197
rect -11496 17163 -11450 17197
rect -11416 17163 -11370 17197
rect -11336 17163 -11290 17197
rect -11256 17163 -11210 17197
rect -11176 17163 -11130 17197
rect -11096 17163 -11050 17197
rect -11016 17163 -10970 17197
rect -10936 17163 -10890 17197
rect -10856 17163 -10810 17197
rect -10776 17163 -10730 17197
rect -10696 17163 -10650 17197
rect -10616 17163 -10570 17197
rect -10536 17163 -10490 17197
rect -10456 17163 -10410 17197
rect -10376 17163 -10330 17197
rect -10296 17163 -10250 17197
rect -10216 17163 -10170 17197
rect -10136 17163 -10090 17197
rect -10056 17163 -10010 17197
rect -9976 17163 -9930 17197
rect -9896 17163 -9850 17197
rect -9816 17163 -9770 17197
rect -9736 17163 -9690 17197
rect -9656 17163 -9610 17197
rect -9576 17163 -9530 17197
rect -9496 17163 -9450 17197
rect -9416 17163 -9370 17197
rect -9336 17163 -9290 17197
rect -9256 17163 -9210 17197
rect -9176 17163 -9130 17197
rect -9096 17163 -9050 17197
rect -9016 17163 -8970 17197
rect -8936 17163 -8890 17197
rect -8856 17163 -8810 17197
rect -8776 17163 -8730 17197
rect -8696 17163 -8650 17197
rect -8616 17163 -8570 17197
rect -8536 17163 -8490 17197
rect -8456 17163 -8410 17197
rect -8376 17163 -8330 17197
rect -8296 17163 -8250 17197
rect -8216 17163 -8170 17197
rect -8136 17163 -8090 17197
rect -8056 17163 -8010 17197
rect -7976 17163 -7930 17197
rect -7896 17163 -7850 17197
rect -7816 17163 -7770 17197
rect -7736 17163 -7690 17197
rect -7656 17163 -7610 17197
rect -7576 17163 -7530 17197
rect -7496 17163 -7450 17197
rect -7416 17163 -7370 17197
rect -7336 17163 -7290 17197
rect -7256 17163 -7210 17197
rect -7176 17163 -7130 17197
rect -7096 17163 -7050 17197
rect -7016 17163 -6970 17197
rect -6936 17163 -6890 17197
rect -6856 17163 -6810 17197
rect -6776 17163 -6730 17197
rect -6696 17163 -6650 17197
rect -6616 17163 -6570 17197
rect -6536 17163 -6490 17197
rect -6456 17163 -6410 17197
rect -6376 17163 -6330 17197
rect -6296 17163 -6250 17197
rect -6216 17163 -6170 17197
rect -6136 17163 -6090 17197
rect -6056 17163 -6010 17197
rect -5976 17163 -5930 17197
rect -5896 17163 -5850 17197
rect -5816 17163 -5770 17197
rect -5736 17163 -5690 17197
rect -5656 17163 -5610 17197
rect -5576 17163 -5530 17197
rect -5496 17163 -5450 17197
rect -5416 17163 -5370 17197
rect -5336 17163 -5290 17197
rect -5256 17163 -5210 17197
rect -5176 17163 -5130 17197
rect -5096 17163 -5050 17197
rect -5016 17163 -4970 17197
rect -4936 17163 -4890 17197
rect -4856 17163 -4810 17197
rect -4776 17163 -4730 17197
rect -4696 17163 -4650 17197
rect -4616 17163 -4570 17197
rect -4536 17163 -4490 17197
rect -4456 17163 -4410 17197
rect -4376 17163 -4330 17197
rect -4296 17163 -4250 17197
rect -4216 17163 -4170 17197
rect -4136 17163 -4090 17197
rect -4056 17163 -4010 17197
rect -3976 17163 -3930 17197
rect -3896 17163 -3850 17197
rect -3816 17163 -3770 17197
rect -3736 17163 -3690 17197
rect -3656 17163 -3610 17197
rect -3576 17163 -3530 17197
rect -3496 17163 -3450 17197
rect -3416 17163 -3370 17197
rect -3336 17163 -3290 17197
rect -37898 17130 -3290 17163
rect -1942 17197 2397 17230
rect -1942 17163 -1929 17197
rect -1895 17163 -1849 17197
rect -1815 17163 -1769 17197
rect -1735 17163 -1689 17197
rect -1655 17163 -1609 17197
rect -1575 17163 -1529 17197
rect -1495 17163 -1449 17197
rect -1415 17163 -1369 17197
rect -1335 17163 -1289 17197
rect -1255 17163 -1209 17197
rect -1175 17163 -1129 17197
rect -1095 17163 -1049 17197
rect -1015 17163 -969 17197
rect -935 17163 -889 17197
rect -855 17163 -809 17197
rect -775 17163 -729 17197
rect -695 17163 -649 17197
rect -615 17163 -569 17197
rect -535 17163 -489 17197
rect -455 17163 -409 17197
rect -375 17163 -329 17197
rect -295 17163 -249 17197
rect -215 17163 -169 17197
rect -135 17163 -89 17197
rect -55 17163 -9 17197
rect 25 17163 71 17197
rect 105 17163 151 17197
rect 185 17163 231 17197
rect 265 17163 311 17197
rect 345 17163 391 17197
rect 425 17163 471 17197
rect 505 17163 551 17197
rect 585 17163 631 17197
rect 665 17163 711 17197
rect 745 17163 791 17197
rect 825 17163 871 17197
rect 905 17163 951 17197
rect 985 17163 1031 17197
rect 1065 17163 1111 17197
rect 1145 17163 1191 17197
rect 1225 17163 1271 17197
rect 1305 17163 1351 17197
rect 1385 17163 1431 17197
rect 1465 17163 1511 17197
rect 1545 17163 1591 17197
rect 1625 17163 1671 17197
rect 1705 17163 1751 17197
rect 1785 17163 1831 17197
rect 1865 17163 1911 17197
rect 1945 17163 1991 17197
rect 2025 17163 2071 17197
rect 2105 17163 2151 17197
rect 2185 17163 2231 17197
rect 2265 17163 2311 17197
rect 2345 17163 2397 17197
rect -1942 17130 2397 17163
rect 3744 17197 38351 17230
rect 3744 17163 3790 17197
rect 3824 17163 3870 17197
rect 3904 17163 3950 17197
rect 3984 17163 4030 17197
rect 4064 17163 4110 17197
rect 4144 17163 4190 17197
rect 4224 17163 4270 17197
rect 4304 17163 4350 17197
rect 4384 17163 4430 17197
rect 4464 17163 4510 17197
rect 4544 17163 4590 17197
rect 4624 17163 4670 17197
rect 4704 17163 4750 17197
rect 4784 17163 4830 17197
rect 4864 17163 4910 17197
rect 4944 17163 4990 17197
rect 5024 17163 5070 17197
rect 5104 17163 5150 17197
rect 5184 17163 5230 17197
rect 5264 17163 5310 17197
rect 5344 17163 5390 17197
rect 5424 17163 5470 17197
rect 5504 17163 5550 17197
rect 5584 17163 5630 17197
rect 5664 17163 5710 17197
rect 5744 17163 5790 17197
rect 5824 17163 5870 17197
rect 5904 17163 5950 17197
rect 5984 17163 6030 17197
rect 6064 17163 6110 17197
rect 6144 17163 6190 17197
rect 6224 17163 6270 17197
rect 6304 17163 6350 17197
rect 6384 17163 6430 17197
rect 6464 17163 6510 17197
rect 6544 17163 6590 17197
rect 6624 17163 6670 17197
rect 6704 17163 6750 17197
rect 6784 17163 6830 17197
rect 6864 17163 6910 17197
rect 6944 17163 6990 17197
rect 7024 17163 7070 17197
rect 7104 17163 7150 17197
rect 7184 17163 7230 17197
rect 7264 17163 7310 17197
rect 7344 17163 7390 17197
rect 7424 17163 7470 17197
rect 7504 17163 7550 17197
rect 7584 17163 7630 17197
rect 7664 17163 7710 17197
rect 7744 17163 7790 17197
rect 7824 17163 7870 17197
rect 7904 17163 7950 17197
rect 7984 17163 8030 17197
rect 8064 17163 8110 17197
rect 8144 17163 8190 17197
rect 8224 17163 8270 17197
rect 8304 17163 8350 17197
rect 8384 17163 8430 17197
rect 8464 17163 8510 17197
rect 8544 17163 8590 17197
rect 8624 17163 8670 17197
rect 8704 17163 8750 17197
rect 8784 17163 8830 17197
rect 8864 17163 8910 17197
rect 8944 17163 8990 17197
rect 9024 17163 9070 17197
rect 9104 17163 9150 17197
rect 9184 17163 9230 17197
rect 9264 17163 9310 17197
rect 9344 17163 9390 17197
rect 9424 17163 9470 17197
rect 9504 17163 9550 17197
rect 9584 17163 9630 17197
rect 9664 17163 9710 17197
rect 9744 17163 9790 17197
rect 9824 17163 9870 17197
rect 9904 17163 9950 17197
rect 9984 17163 10030 17197
rect 10064 17163 10110 17197
rect 10144 17163 10190 17197
rect 10224 17163 10270 17197
rect 10304 17163 10350 17197
rect 10384 17163 10430 17197
rect 10464 17163 10510 17197
rect 10544 17163 10590 17197
rect 10624 17163 10670 17197
rect 10704 17163 10750 17197
rect 10784 17163 10830 17197
rect 10864 17163 10910 17197
rect 10944 17163 10990 17197
rect 11024 17163 11070 17197
rect 11104 17163 11150 17197
rect 11184 17163 11230 17197
rect 11264 17163 11310 17197
rect 11344 17163 11390 17197
rect 11424 17163 11470 17197
rect 11504 17163 11550 17197
rect 11584 17163 11630 17197
rect 11664 17163 11710 17197
rect 11744 17163 11790 17197
rect 11824 17163 11870 17197
rect 11904 17163 11950 17197
rect 11984 17163 12030 17197
rect 12064 17163 12110 17197
rect 12144 17163 12190 17197
rect 12224 17163 12270 17197
rect 12304 17163 12350 17197
rect 12384 17163 12430 17197
rect 12464 17163 12510 17197
rect 12544 17163 12590 17197
rect 12624 17163 12670 17197
rect 12704 17163 12750 17197
rect 12784 17163 12830 17197
rect 12864 17163 12910 17197
rect 12944 17163 12990 17197
rect 13024 17163 13070 17197
rect 13104 17163 13150 17197
rect 13184 17163 13230 17197
rect 13264 17163 13310 17197
rect 13344 17163 13390 17197
rect 13424 17163 13470 17197
rect 13504 17163 13550 17197
rect 13584 17163 13630 17197
rect 13664 17163 13710 17197
rect 13744 17163 13790 17197
rect 13824 17163 13870 17197
rect 13904 17163 13950 17197
rect 13984 17163 14030 17197
rect 14064 17163 14110 17197
rect 14144 17163 14190 17197
rect 14224 17163 14270 17197
rect 14304 17163 14350 17197
rect 14384 17163 14430 17197
rect 14464 17163 14510 17197
rect 14544 17163 14590 17197
rect 14624 17163 14670 17197
rect 14704 17163 14750 17197
rect 14784 17163 14830 17197
rect 14864 17163 14910 17197
rect 14944 17163 14990 17197
rect 15024 17163 15070 17197
rect 15104 17163 15150 17197
rect 15184 17163 15230 17197
rect 15264 17163 15310 17197
rect 15344 17163 15390 17197
rect 15424 17163 15470 17197
rect 15504 17163 15550 17197
rect 15584 17163 15630 17197
rect 15664 17163 15710 17197
rect 15744 17163 15790 17197
rect 15824 17163 15870 17197
rect 15904 17163 15950 17197
rect 15984 17163 16030 17197
rect 16064 17163 16110 17197
rect 16144 17163 16190 17197
rect 16224 17163 16270 17197
rect 16304 17163 16350 17197
rect 16384 17163 16430 17197
rect 16464 17163 16510 17197
rect 16544 17163 16590 17197
rect 16624 17163 16670 17197
rect 16704 17163 16751 17197
rect 16785 17163 16831 17197
rect 16865 17163 16911 17197
rect 16945 17163 16991 17197
rect 17025 17163 17071 17197
rect 17105 17163 17151 17197
rect 17185 17163 17231 17197
rect 17265 17163 17311 17197
rect 17345 17163 17391 17197
rect 17425 17163 17471 17197
rect 17505 17163 17551 17197
rect 17585 17163 17631 17197
rect 17665 17163 17711 17197
rect 17745 17163 17791 17197
rect 17825 17163 17871 17197
rect 17905 17163 17951 17197
rect 17985 17163 18031 17197
rect 18065 17163 18111 17197
rect 18145 17163 18191 17197
rect 18225 17163 18271 17197
rect 18305 17163 18351 17197
rect 18385 17163 18431 17197
rect 18465 17163 18511 17197
rect 18545 17163 18591 17197
rect 18625 17163 18671 17197
rect 18705 17163 18751 17197
rect 18785 17163 18831 17197
rect 18865 17163 18911 17197
rect 18945 17163 18991 17197
rect 19025 17163 19071 17197
rect 19105 17163 19151 17197
rect 19185 17163 19231 17197
rect 19265 17163 19311 17197
rect 19345 17163 19391 17197
rect 19425 17163 19471 17197
rect 19505 17163 19551 17197
rect 19585 17163 19631 17197
rect 19665 17163 19711 17197
rect 19745 17163 19791 17197
rect 19825 17163 19871 17197
rect 19905 17163 19951 17197
rect 19985 17163 20031 17197
rect 20065 17163 20111 17197
rect 20145 17163 20191 17197
rect 20225 17163 20271 17197
rect 20305 17163 20351 17197
rect 20385 17163 20431 17197
rect 20465 17163 20511 17197
rect 20545 17163 20591 17197
rect 20625 17163 20671 17197
rect 20705 17163 20751 17197
rect 20785 17163 20831 17197
rect 20865 17163 20911 17197
rect 20945 17163 20991 17197
rect 21025 17163 21071 17197
rect 21105 17163 21151 17197
rect 21185 17163 21231 17197
rect 21265 17163 21311 17197
rect 21345 17163 21391 17197
rect 21425 17163 21471 17197
rect 21505 17163 21551 17197
rect 21585 17163 21631 17197
rect 21665 17163 21711 17197
rect 21745 17163 21791 17197
rect 21825 17163 21871 17197
rect 21905 17163 21951 17197
rect 21985 17163 22031 17197
rect 22065 17163 22111 17197
rect 22145 17163 22191 17197
rect 22225 17163 22271 17197
rect 22305 17163 22351 17197
rect 22385 17163 22431 17197
rect 22465 17163 22511 17197
rect 22545 17163 22591 17197
rect 22625 17163 22671 17197
rect 22705 17163 22751 17197
rect 22785 17163 22831 17197
rect 22865 17163 22911 17197
rect 22945 17163 22991 17197
rect 23025 17163 23071 17197
rect 23105 17163 23151 17197
rect 23185 17163 23231 17197
rect 23265 17163 23311 17197
rect 23345 17163 23391 17197
rect 23425 17163 23471 17197
rect 23505 17163 23551 17197
rect 23585 17163 23631 17197
rect 23665 17163 23711 17197
rect 23745 17163 23791 17197
rect 23825 17163 23871 17197
rect 23905 17163 23951 17197
rect 23985 17163 24031 17197
rect 24065 17163 24111 17197
rect 24145 17163 24191 17197
rect 24225 17163 24271 17197
rect 24305 17163 24351 17197
rect 24385 17163 24431 17197
rect 24465 17163 24511 17197
rect 24545 17163 24591 17197
rect 24625 17163 24671 17197
rect 24705 17163 24751 17197
rect 24785 17163 24831 17197
rect 24865 17163 24911 17197
rect 24945 17163 24991 17197
rect 25025 17163 25071 17197
rect 25105 17163 25151 17197
rect 25185 17163 25231 17197
rect 25265 17163 25311 17197
rect 25345 17163 25391 17197
rect 25425 17163 25471 17197
rect 25505 17163 25551 17197
rect 25585 17163 25631 17197
rect 25665 17163 25711 17197
rect 25745 17163 25791 17197
rect 25825 17163 25871 17197
rect 25905 17163 25951 17197
rect 25985 17163 26031 17197
rect 26065 17163 26111 17197
rect 26145 17163 26191 17197
rect 26225 17163 26271 17197
rect 26305 17163 26351 17197
rect 26385 17163 26431 17197
rect 26465 17163 26511 17197
rect 26545 17163 26591 17197
rect 26625 17163 26671 17197
rect 26705 17163 26751 17197
rect 26785 17163 26831 17197
rect 26865 17163 26911 17197
rect 26945 17163 26991 17197
rect 27025 17163 27071 17197
rect 27105 17163 27151 17197
rect 27185 17163 27231 17197
rect 27265 17163 27311 17197
rect 27345 17163 27391 17197
rect 27425 17163 27471 17197
rect 27505 17163 27551 17197
rect 27585 17163 27631 17197
rect 27665 17163 27711 17197
rect 27745 17163 27791 17197
rect 27825 17163 27871 17197
rect 27905 17163 27951 17197
rect 27985 17163 28031 17197
rect 28065 17163 28111 17197
rect 28145 17163 28191 17197
rect 28225 17163 28271 17197
rect 28305 17163 28351 17197
rect 28385 17163 28431 17197
rect 28465 17163 28511 17197
rect 28545 17163 28591 17197
rect 28625 17163 28671 17197
rect 28705 17163 28751 17197
rect 28785 17163 28831 17197
rect 28865 17163 28911 17197
rect 28945 17163 28991 17197
rect 29025 17163 29071 17197
rect 29105 17163 29151 17197
rect 29185 17163 29231 17197
rect 29265 17163 29311 17197
rect 29345 17163 29391 17197
rect 29425 17163 29471 17197
rect 29505 17163 29551 17197
rect 29585 17163 29631 17197
rect 29665 17163 29711 17197
rect 29745 17163 29791 17197
rect 29825 17163 29871 17197
rect 29905 17163 29951 17197
rect 29985 17163 30031 17197
rect 30065 17163 30111 17197
rect 30145 17163 30191 17197
rect 30225 17163 30271 17197
rect 30305 17163 30351 17197
rect 30385 17163 30431 17197
rect 30465 17163 30511 17197
rect 30545 17163 30591 17197
rect 30625 17163 30671 17197
rect 30705 17163 30751 17197
rect 30785 17163 30831 17197
rect 30865 17163 30911 17197
rect 30945 17163 30991 17197
rect 31025 17163 31071 17197
rect 31105 17163 31151 17197
rect 31185 17163 31231 17197
rect 31265 17163 31311 17197
rect 31345 17163 31391 17197
rect 31425 17163 31471 17197
rect 31505 17163 31551 17197
rect 31585 17163 31631 17197
rect 31665 17163 31711 17197
rect 31745 17163 31791 17197
rect 31825 17163 31871 17197
rect 31905 17163 31951 17197
rect 31985 17163 32031 17197
rect 32065 17163 32111 17197
rect 32145 17163 32191 17197
rect 32225 17163 32271 17197
rect 32305 17163 32351 17197
rect 32385 17163 32431 17197
rect 32465 17163 32511 17197
rect 32545 17163 32591 17197
rect 32625 17163 32671 17197
rect 32705 17163 32751 17197
rect 32785 17163 32831 17197
rect 32865 17163 32911 17197
rect 32945 17163 32991 17197
rect 33025 17163 33071 17197
rect 33105 17163 33151 17197
rect 33185 17163 33231 17197
rect 33265 17163 33311 17197
rect 33345 17163 33391 17197
rect 33425 17163 33471 17197
rect 33505 17163 33551 17197
rect 33585 17163 33631 17197
rect 33665 17163 33711 17197
rect 33745 17163 33791 17197
rect 33825 17163 33871 17197
rect 33905 17163 33951 17197
rect 33985 17163 34031 17197
rect 34065 17163 34111 17197
rect 34145 17163 34191 17197
rect 34225 17163 34271 17197
rect 34305 17163 34351 17197
rect 34385 17163 34431 17197
rect 34465 17163 34511 17197
rect 34545 17163 34591 17197
rect 34625 17163 34671 17197
rect 34705 17163 34751 17197
rect 34785 17163 34831 17197
rect 34865 17163 34911 17197
rect 34945 17163 34991 17197
rect 35025 17163 35071 17197
rect 35105 17163 35151 17197
rect 35185 17163 35231 17197
rect 35265 17163 35311 17197
rect 35345 17163 35391 17197
rect 35425 17163 35471 17197
rect 35505 17163 35551 17197
rect 35585 17163 35631 17197
rect 35665 17163 35711 17197
rect 35745 17163 35791 17197
rect 35825 17163 35871 17197
rect 35905 17163 35951 17197
rect 35985 17163 36031 17197
rect 36065 17163 36111 17197
rect 36145 17163 36191 17197
rect 36225 17163 36271 17197
rect 36305 17163 36351 17197
rect 36385 17163 36431 17197
rect 36465 17163 36511 17197
rect 36545 17163 36591 17197
rect 36625 17163 36671 17197
rect 36705 17163 36751 17197
rect 36785 17163 36831 17197
rect 36865 17163 36911 17197
rect 36945 17163 36991 17197
rect 37025 17163 37071 17197
rect 37105 17163 37151 17197
rect 37185 17163 37231 17197
rect 37265 17163 37311 17197
rect 37345 17163 37391 17197
rect 37425 17163 37471 17197
rect 37505 17163 37551 17197
rect 37585 17163 37631 17197
rect 37665 17163 37711 17197
rect 37745 17163 37791 17197
rect 37825 17163 37871 17197
rect 37905 17163 37951 17197
rect 37985 17163 38031 17197
rect 38065 17163 38111 17197
rect 38145 17163 38191 17197
rect 38225 17163 38271 17197
rect 38305 17163 38351 17197
rect 3744 17130 38351 17163
rect 18621 17129 18881 17130
rect -37898 9338 -3290 9371
rect -37898 9304 -37852 9338
rect -37818 9304 -37772 9338
rect -37738 9304 -37692 9338
rect -37658 9304 -37612 9338
rect -37578 9304 -37532 9338
rect -37498 9304 -37452 9338
rect -37418 9304 -37372 9338
rect -37338 9304 -37292 9338
rect -37258 9304 -37212 9338
rect -37178 9304 -37132 9338
rect -37098 9304 -37052 9338
rect -37018 9304 -36972 9338
rect -36938 9304 -36892 9338
rect -36858 9304 -36812 9338
rect -36778 9304 -36732 9338
rect -36698 9304 -36652 9338
rect -36618 9304 -36572 9338
rect -36538 9304 -36492 9338
rect -36458 9304 -36412 9338
rect -36378 9304 -36332 9338
rect -36298 9304 -36252 9338
rect -36218 9304 -36172 9338
rect -36138 9304 -36092 9338
rect -36058 9304 -36012 9338
rect -35978 9304 -35932 9338
rect -35898 9304 -35852 9338
rect -35818 9304 -35772 9338
rect -35738 9304 -35692 9338
rect -35658 9304 -35612 9338
rect -35578 9304 -35532 9338
rect -35498 9304 -35452 9338
rect -35418 9304 -35372 9338
rect -35338 9304 -35292 9338
rect -35258 9304 -35212 9338
rect -35178 9304 -35132 9338
rect -35098 9304 -35052 9338
rect -35018 9304 -34972 9338
rect -34938 9304 -34892 9338
rect -34858 9304 -34812 9338
rect -34778 9304 -34732 9338
rect -34698 9304 -34652 9338
rect -34618 9304 -34572 9338
rect -34538 9304 -34492 9338
rect -34458 9304 -34412 9338
rect -34378 9304 -34332 9338
rect -34298 9304 -34252 9338
rect -34218 9304 -34172 9338
rect -34138 9304 -34092 9338
rect -34058 9304 -34012 9338
rect -33978 9304 -33932 9338
rect -33898 9304 -33852 9338
rect -33818 9304 -33772 9338
rect -33738 9304 -33692 9338
rect -33658 9304 -33612 9338
rect -33578 9304 -33532 9338
rect -33498 9304 -33452 9338
rect -33418 9304 -33372 9338
rect -33338 9304 -33292 9338
rect -33258 9304 -33212 9338
rect -33178 9304 -33132 9338
rect -33098 9304 -33052 9338
rect -33018 9304 -32972 9338
rect -32938 9304 -32892 9338
rect -32858 9304 -32812 9338
rect -32778 9304 -32732 9338
rect -32698 9304 -32652 9338
rect -32618 9304 -32572 9338
rect -32538 9304 -32492 9338
rect -32458 9304 -32412 9338
rect -32378 9304 -32332 9338
rect -32298 9304 -32252 9338
rect -32218 9304 -32172 9338
rect -32138 9304 -32092 9338
rect -32058 9304 -32012 9338
rect -31978 9304 -31932 9338
rect -31898 9304 -31852 9338
rect -31818 9304 -31772 9338
rect -31738 9304 -31692 9338
rect -31658 9304 -31612 9338
rect -31578 9304 -31532 9338
rect -31498 9304 -31452 9338
rect -31418 9304 -31372 9338
rect -31338 9304 -31292 9338
rect -31258 9304 -31212 9338
rect -31178 9304 -31132 9338
rect -31098 9304 -31052 9338
rect -31018 9304 -30972 9338
rect -30938 9304 -30892 9338
rect -30858 9304 -30812 9338
rect -30778 9304 -30732 9338
rect -30698 9304 -30652 9338
rect -30618 9304 -30572 9338
rect -30538 9304 -30492 9338
rect -30458 9304 -30412 9338
rect -30378 9304 -30332 9338
rect -30298 9304 -30252 9338
rect -30218 9304 -30172 9338
rect -30138 9304 -30092 9338
rect -30058 9304 -30012 9338
rect -29978 9304 -29932 9338
rect -29898 9304 -29852 9338
rect -29818 9304 -29772 9338
rect -29738 9304 -29692 9338
rect -29658 9304 -29612 9338
rect -29578 9304 -29532 9338
rect -29498 9304 -29452 9338
rect -29418 9304 -29372 9338
rect -29338 9304 -29292 9338
rect -29258 9304 -29212 9338
rect -29178 9304 -29132 9338
rect -29098 9304 -29052 9338
rect -29018 9304 -28972 9338
rect -28938 9304 -28892 9338
rect -28858 9304 -28812 9338
rect -28778 9304 -28732 9338
rect -28698 9304 -28652 9338
rect -28618 9304 -28572 9338
rect -28538 9304 -28492 9338
rect -28458 9304 -28412 9338
rect -28378 9304 -28332 9338
rect -28298 9304 -28252 9338
rect -28218 9304 -28172 9338
rect -28138 9304 -28092 9338
rect -28058 9304 -28012 9338
rect -27978 9304 -27932 9338
rect -27898 9304 -27852 9338
rect -27818 9304 -27772 9338
rect -27738 9304 -27692 9338
rect -27658 9304 -27612 9338
rect -27578 9304 -27532 9338
rect -27498 9304 -27452 9338
rect -27418 9304 -27372 9338
rect -27338 9304 -27292 9338
rect -27258 9304 -27212 9338
rect -27178 9304 -27132 9338
rect -27098 9304 -27052 9338
rect -27018 9304 -26972 9338
rect -26938 9304 -26892 9338
rect -26858 9304 -26812 9338
rect -26778 9304 -26732 9338
rect -26698 9304 -26652 9338
rect -26618 9304 -26572 9338
rect -26538 9304 -26492 9338
rect -26458 9304 -26412 9338
rect -26378 9304 -26332 9338
rect -26298 9304 -26252 9338
rect -26218 9304 -26172 9338
rect -26138 9304 -26092 9338
rect -26058 9304 -26012 9338
rect -25978 9304 -25932 9338
rect -25898 9304 -25852 9338
rect -25818 9304 -25772 9338
rect -25738 9304 -25692 9338
rect -25658 9304 -25612 9338
rect -25578 9304 -25532 9338
rect -25498 9304 -25452 9338
rect -25418 9304 -25372 9338
rect -25338 9304 -25292 9338
rect -25258 9304 -25212 9338
rect -25178 9304 -25132 9338
rect -25098 9304 -25052 9338
rect -25018 9304 -24972 9338
rect -24938 9304 -24891 9338
rect -24857 9304 -24811 9338
rect -24777 9304 -24731 9338
rect -24697 9304 -24651 9338
rect -24617 9304 -24571 9338
rect -24537 9304 -24491 9338
rect -24457 9304 -24411 9338
rect -24377 9304 -24331 9338
rect -24297 9304 -24251 9338
rect -24217 9304 -24171 9338
rect -24137 9304 -24091 9338
rect -24057 9304 -24011 9338
rect -23977 9304 -23931 9338
rect -23897 9304 -23851 9338
rect -23817 9304 -23771 9338
rect -23737 9304 -23691 9338
rect -23657 9304 -23611 9338
rect -23577 9304 -23531 9338
rect -23497 9304 -23451 9338
rect -23417 9304 -23371 9338
rect -23337 9304 -23291 9338
rect -23257 9304 -23211 9338
rect -23177 9304 -23131 9338
rect -23097 9304 -23051 9338
rect -23017 9304 -22971 9338
rect -22937 9304 -22891 9338
rect -22857 9304 -22811 9338
rect -22777 9304 -22731 9338
rect -22697 9304 -22651 9338
rect -22617 9304 -22571 9338
rect -22537 9304 -22491 9338
rect -22457 9304 -22411 9338
rect -22377 9304 -22331 9338
rect -22297 9304 -22251 9338
rect -22217 9304 -22171 9338
rect -22137 9304 -22091 9338
rect -22057 9304 -22011 9338
rect -21977 9304 -21931 9338
rect -21897 9304 -21851 9338
rect -21817 9304 -21771 9338
rect -21737 9304 -21691 9338
rect -21657 9304 -21611 9338
rect -21577 9304 -21531 9338
rect -21497 9304 -21451 9338
rect -21417 9304 -21371 9338
rect -21337 9304 -21291 9338
rect -21257 9304 -21211 9338
rect -21177 9304 -21131 9338
rect -21097 9304 -21051 9338
rect -21017 9304 -20971 9338
rect -20937 9304 -20891 9338
rect -20857 9304 -20811 9338
rect -20777 9304 -20731 9338
rect -20697 9304 -20651 9338
rect -20617 9304 -20571 9338
rect -20537 9304 -20491 9338
rect -20457 9304 -20411 9338
rect -20377 9304 -20331 9338
rect -20297 9304 -20251 9338
rect -20217 9304 -20171 9338
rect -20137 9304 -20091 9338
rect -20057 9304 -20011 9338
rect -19977 9304 -19931 9338
rect -19897 9304 -19851 9338
rect -19817 9304 -19771 9338
rect -19737 9304 -19691 9338
rect -19657 9304 -19611 9338
rect -19577 9304 -19531 9338
rect -19497 9304 -19451 9338
rect -19417 9304 -19371 9338
rect -19337 9304 -19291 9338
rect -19257 9304 -19211 9338
rect -19177 9304 -19131 9338
rect -19097 9304 -19051 9338
rect -19017 9304 -18971 9338
rect -18937 9304 -18891 9338
rect -18857 9304 -18811 9338
rect -18777 9304 -18731 9338
rect -18697 9304 -18651 9338
rect -18617 9304 -18571 9338
rect -18537 9304 -18491 9338
rect -18457 9304 -18411 9338
rect -18377 9304 -18331 9338
rect -18297 9304 -18251 9338
rect -18217 9304 -18171 9338
rect -18137 9304 -18091 9338
rect -18057 9304 -18011 9338
rect -17977 9304 -17931 9338
rect -17897 9304 -17851 9338
rect -17817 9304 -17771 9338
rect -17737 9304 -17691 9338
rect -17657 9304 -17611 9338
rect -17577 9304 -17531 9338
rect -17497 9304 -17451 9338
rect -17417 9304 -17371 9338
rect -17337 9304 -17291 9338
rect -17257 9304 -17211 9338
rect -17177 9304 -17131 9338
rect -17097 9304 -17051 9338
rect -17017 9304 -16971 9338
rect -16937 9304 -16891 9338
rect -16857 9304 -16811 9338
rect -16777 9304 -16731 9338
rect -16697 9304 -16651 9338
rect -16617 9304 -16571 9338
rect -16537 9304 -16491 9338
rect -16457 9304 -16411 9338
rect -16377 9304 -16331 9338
rect -16297 9304 -16251 9338
rect -16217 9304 -16171 9338
rect -16137 9304 -16091 9338
rect -16057 9304 -16011 9338
rect -15977 9304 -15931 9338
rect -15897 9304 -15851 9338
rect -15817 9304 -15771 9338
rect -15737 9304 -15691 9338
rect -15657 9304 -15611 9338
rect -15577 9304 -15531 9338
rect -15497 9304 -15451 9338
rect -15417 9304 -15371 9338
rect -15337 9304 -15291 9338
rect -15257 9304 -15211 9338
rect -15177 9304 -15131 9338
rect -15097 9304 -15051 9338
rect -15017 9304 -14971 9338
rect -14937 9304 -14891 9338
rect -14857 9304 -14811 9338
rect -14777 9304 -14731 9338
rect -14697 9304 -14651 9338
rect -14617 9304 -14571 9338
rect -14537 9304 -14491 9338
rect -14457 9304 -14411 9338
rect -14377 9304 -14331 9338
rect -14297 9304 -14251 9338
rect -14217 9304 -14171 9338
rect -14137 9304 -14091 9338
rect -14057 9304 -14011 9338
rect -13977 9304 -13931 9338
rect -13897 9304 -13851 9338
rect -13817 9304 -13771 9338
rect -13737 9304 -13691 9338
rect -13657 9304 -13611 9338
rect -13577 9304 -13531 9338
rect -13497 9304 -13451 9338
rect -13417 9304 -13371 9338
rect -13337 9304 -13291 9338
rect -13257 9304 -13211 9338
rect -13177 9304 -13131 9338
rect -13097 9304 -13051 9338
rect -13017 9304 -12971 9338
rect -12937 9304 -12891 9338
rect -12857 9304 -12811 9338
rect -12777 9304 -12731 9338
rect -12697 9304 -12651 9338
rect -12617 9304 -12571 9338
rect -12537 9304 -12491 9338
rect -12457 9304 -12411 9338
rect -12377 9304 -12331 9338
rect -12297 9304 -12251 9338
rect -12217 9304 -12171 9338
rect -12137 9304 -12091 9338
rect -12057 9304 -12011 9338
rect -11977 9304 -11930 9338
rect -11896 9304 -11850 9338
rect -11816 9304 -11770 9338
rect -11736 9304 -11690 9338
rect -11656 9304 -11610 9338
rect -11576 9304 -11530 9338
rect -11496 9304 -11450 9338
rect -11416 9304 -11370 9338
rect -11336 9304 -11290 9338
rect -11256 9304 -11210 9338
rect -11176 9304 -11130 9338
rect -11096 9304 -11050 9338
rect -11016 9304 -10970 9338
rect -10936 9304 -10890 9338
rect -10856 9304 -10810 9338
rect -10776 9304 -10730 9338
rect -10696 9304 -10650 9338
rect -10616 9304 -10570 9338
rect -10536 9304 -10490 9338
rect -10456 9304 -10410 9338
rect -10376 9304 -10330 9338
rect -10296 9304 -10250 9338
rect -10216 9304 -10170 9338
rect -10136 9304 -10090 9338
rect -10056 9304 -10010 9338
rect -9976 9304 -9930 9338
rect -9896 9304 -9850 9338
rect -9816 9304 -9770 9338
rect -9736 9304 -9690 9338
rect -9656 9304 -9610 9338
rect -9576 9304 -9530 9338
rect -9496 9304 -9450 9338
rect -9416 9304 -9370 9338
rect -9336 9304 -9290 9338
rect -9256 9304 -9210 9338
rect -9176 9304 -9130 9338
rect -9096 9304 -9050 9338
rect -9016 9304 -8970 9338
rect -8936 9304 -8890 9338
rect -8856 9304 -8810 9338
rect -8776 9304 -8730 9338
rect -8696 9304 -8650 9338
rect -8616 9304 -8570 9338
rect -8536 9304 -8490 9338
rect -8456 9304 -8410 9338
rect -8376 9304 -8330 9338
rect -8296 9304 -8250 9338
rect -8216 9304 -8170 9338
rect -8136 9304 -8090 9338
rect -8056 9304 -8010 9338
rect -7976 9304 -7930 9338
rect -7896 9304 -7850 9338
rect -7816 9304 -7770 9338
rect -7736 9304 -7690 9338
rect -7656 9304 -7610 9338
rect -7576 9304 -7530 9338
rect -7496 9304 -7450 9338
rect -7416 9304 -7370 9338
rect -7336 9304 -7290 9338
rect -7256 9304 -7210 9338
rect -7176 9304 -7130 9338
rect -7096 9304 -7050 9338
rect -7016 9304 -6970 9338
rect -6936 9304 -6890 9338
rect -6856 9304 -6810 9338
rect -6776 9304 -6730 9338
rect -6696 9304 -6650 9338
rect -6616 9304 -6570 9338
rect -6536 9304 -6490 9338
rect -6456 9304 -6410 9338
rect -6376 9304 -6330 9338
rect -6296 9304 -6250 9338
rect -6216 9304 -6170 9338
rect -6136 9304 -6090 9338
rect -6056 9304 -6010 9338
rect -5976 9304 -5930 9338
rect -5896 9304 -5850 9338
rect -5816 9304 -5770 9338
rect -5736 9304 -5690 9338
rect -5656 9304 -5610 9338
rect -5576 9304 -5530 9338
rect -5496 9304 -5450 9338
rect -5416 9304 -5370 9338
rect -5336 9304 -5290 9338
rect -5256 9304 -5210 9338
rect -5176 9304 -5130 9338
rect -5096 9304 -5050 9338
rect -5016 9304 -4970 9338
rect -4936 9304 -4890 9338
rect -4856 9304 -4810 9338
rect -4776 9304 -4730 9338
rect -4696 9304 -4650 9338
rect -4616 9304 -4570 9338
rect -4536 9304 -4490 9338
rect -4456 9304 -4410 9338
rect -4376 9304 -4330 9338
rect -4296 9304 -4250 9338
rect -4216 9304 -4170 9338
rect -4136 9304 -4090 9338
rect -4056 9304 -4010 9338
rect -3976 9304 -3930 9338
rect -3896 9304 -3850 9338
rect -3816 9304 -3770 9338
rect -3736 9304 -3690 9338
rect -3656 9304 -3610 9338
rect -3576 9304 -3530 9338
rect -3496 9304 -3450 9338
rect -3416 9304 -3370 9338
rect -3336 9304 -3290 9338
rect -37898 9271 -3290 9304
rect -1942 9338 2397 9371
rect -1942 9304 -1929 9338
rect -1895 9304 -1849 9338
rect -1815 9304 -1769 9338
rect -1735 9304 -1689 9338
rect -1655 9304 -1609 9338
rect -1575 9304 -1529 9338
rect -1495 9304 -1449 9338
rect -1415 9304 -1369 9338
rect -1335 9304 -1289 9338
rect -1255 9304 -1209 9338
rect -1175 9304 -1129 9338
rect -1095 9304 -1049 9338
rect -1015 9304 -969 9338
rect -935 9304 -889 9338
rect -855 9304 -809 9338
rect -775 9304 -729 9338
rect -695 9304 -649 9338
rect -615 9304 -569 9338
rect -535 9304 -489 9338
rect -455 9304 -409 9338
rect -375 9304 -329 9338
rect -295 9304 -249 9338
rect -215 9304 -169 9338
rect -135 9304 -89 9338
rect -55 9304 -9 9338
rect 25 9304 71 9338
rect 105 9304 151 9338
rect 185 9304 231 9338
rect 265 9304 311 9338
rect 345 9304 391 9338
rect 425 9304 471 9338
rect 505 9304 551 9338
rect 585 9304 631 9338
rect 665 9304 711 9338
rect 745 9304 791 9338
rect 825 9304 871 9338
rect 905 9304 951 9338
rect 985 9304 1031 9338
rect 1065 9304 1111 9338
rect 1145 9304 1191 9338
rect 1225 9304 1271 9338
rect 1305 9304 1351 9338
rect 1385 9304 1431 9338
rect 1465 9304 1511 9338
rect 1545 9304 1591 9338
rect 1625 9304 1671 9338
rect 1705 9304 1751 9338
rect 1785 9304 1831 9338
rect 1865 9304 1911 9338
rect 1945 9304 1991 9338
rect 2025 9304 2071 9338
rect 2105 9304 2151 9338
rect 2185 9304 2231 9338
rect 2265 9304 2311 9338
rect 2345 9304 2397 9338
rect -1942 9271 2397 9304
rect 3744 9338 38351 9371
rect 3744 9304 3790 9338
rect 3824 9304 3870 9338
rect 3904 9304 3950 9338
rect 3984 9304 4030 9338
rect 4064 9304 4110 9338
rect 4144 9304 4190 9338
rect 4224 9304 4270 9338
rect 4304 9304 4350 9338
rect 4384 9304 4430 9338
rect 4464 9304 4510 9338
rect 4544 9304 4590 9338
rect 4624 9304 4670 9338
rect 4704 9304 4750 9338
rect 4784 9304 4830 9338
rect 4864 9304 4910 9338
rect 4944 9304 4990 9338
rect 5024 9304 5070 9338
rect 5104 9304 5150 9338
rect 5184 9304 5230 9338
rect 5264 9304 5310 9338
rect 5344 9304 5390 9338
rect 5424 9304 5470 9338
rect 5504 9304 5550 9338
rect 5584 9304 5630 9338
rect 5664 9304 5710 9338
rect 5744 9304 5790 9338
rect 5824 9304 5870 9338
rect 5904 9304 5950 9338
rect 5984 9304 6030 9338
rect 6064 9304 6110 9338
rect 6144 9304 6190 9338
rect 6224 9304 6270 9338
rect 6304 9304 6350 9338
rect 6384 9304 6430 9338
rect 6464 9304 6510 9338
rect 6544 9304 6590 9338
rect 6624 9304 6670 9338
rect 6704 9304 6750 9338
rect 6784 9304 6830 9338
rect 6864 9304 6910 9338
rect 6944 9304 6990 9338
rect 7024 9304 7070 9338
rect 7104 9304 7150 9338
rect 7184 9304 7230 9338
rect 7264 9304 7310 9338
rect 7344 9304 7390 9338
rect 7424 9304 7470 9338
rect 7504 9304 7550 9338
rect 7584 9304 7630 9338
rect 7664 9304 7710 9338
rect 7744 9304 7790 9338
rect 7824 9304 7870 9338
rect 7904 9304 7950 9338
rect 7984 9304 8030 9338
rect 8064 9304 8110 9338
rect 8144 9304 8190 9338
rect 8224 9304 8270 9338
rect 8304 9304 8350 9338
rect 8384 9304 8430 9338
rect 8464 9304 8510 9338
rect 8544 9304 8590 9338
rect 8624 9304 8670 9338
rect 8704 9304 8750 9338
rect 8784 9304 8830 9338
rect 8864 9304 8910 9338
rect 8944 9304 8990 9338
rect 9024 9304 9070 9338
rect 9104 9304 9150 9338
rect 9184 9304 9230 9338
rect 9264 9304 9310 9338
rect 9344 9304 9390 9338
rect 9424 9304 9470 9338
rect 9504 9304 9550 9338
rect 9584 9304 9630 9338
rect 9664 9304 9710 9338
rect 9744 9304 9790 9338
rect 9824 9304 9870 9338
rect 9904 9304 9950 9338
rect 9984 9304 10030 9338
rect 10064 9304 10110 9338
rect 10144 9304 10190 9338
rect 10224 9304 10270 9338
rect 10304 9304 10350 9338
rect 10384 9304 10430 9338
rect 10464 9304 10510 9338
rect 10544 9304 10590 9338
rect 10624 9304 10670 9338
rect 10704 9304 10750 9338
rect 10784 9304 10830 9338
rect 10864 9304 10910 9338
rect 10944 9304 10990 9338
rect 11024 9304 11070 9338
rect 11104 9304 11150 9338
rect 11184 9304 11230 9338
rect 11264 9304 11310 9338
rect 11344 9304 11390 9338
rect 11424 9304 11470 9338
rect 11504 9304 11550 9338
rect 11584 9304 11630 9338
rect 11664 9304 11710 9338
rect 11744 9304 11790 9338
rect 11824 9304 11870 9338
rect 11904 9304 11950 9338
rect 11984 9304 12030 9338
rect 12064 9304 12110 9338
rect 12144 9304 12190 9338
rect 12224 9304 12270 9338
rect 12304 9304 12350 9338
rect 12384 9304 12430 9338
rect 12464 9304 12510 9338
rect 12544 9304 12590 9338
rect 12624 9304 12670 9338
rect 12704 9304 12750 9338
rect 12784 9304 12830 9338
rect 12864 9304 12910 9338
rect 12944 9304 12990 9338
rect 13024 9304 13070 9338
rect 13104 9304 13150 9338
rect 13184 9304 13230 9338
rect 13264 9304 13310 9338
rect 13344 9304 13390 9338
rect 13424 9304 13470 9338
rect 13504 9304 13550 9338
rect 13584 9304 13630 9338
rect 13664 9304 13710 9338
rect 13744 9304 13790 9338
rect 13824 9304 13870 9338
rect 13904 9304 13950 9338
rect 13984 9304 14030 9338
rect 14064 9304 14110 9338
rect 14144 9304 14190 9338
rect 14224 9304 14270 9338
rect 14304 9304 14350 9338
rect 14384 9304 14430 9338
rect 14464 9304 14510 9338
rect 14544 9304 14590 9338
rect 14624 9304 14670 9338
rect 14704 9304 14750 9338
rect 14784 9304 14830 9338
rect 14864 9304 14910 9338
rect 14944 9304 14990 9338
rect 15024 9304 15070 9338
rect 15104 9304 15150 9338
rect 15184 9304 15230 9338
rect 15264 9304 15310 9338
rect 15344 9304 15390 9338
rect 15424 9304 15470 9338
rect 15504 9304 15550 9338
rect 15584 9304 15630 9338
rect 15664 9304 15710 9338
rect 15744 9304 15790 9338
rect 15824 9304 15870 9338
rect 15904 9304 15950 9338
rect 15984 9304 16030 9338
rect 16064 9304 16110 9338
rect 16144 9304 16190 9338
rect 16224 9304 16270 9338
rect 16304 9304 16350 9338
rect 16384 9304 16430 9338
rect 16464 9304 16510 9338
rect 16544 9304 16590 9338
rect 16624 9304 16670 9338
rect 16704 9304 16751 9338
rect 16785 9304 16831 9338
rect 16865 9304 16911 9338
rect 16945 9304 16991 9338
rect 17025 9304 17071 9338
rect 17105 9304 17151 9338
rect 17185 9304 17231 9338
rect 17265 9304 17311 9338
rect 17345 9304 17391 9338
rect 17425 9304 17471 9338
rect 17505 9304 17551 9338
rect 17585 9304 17631 9338
rect 17665 9304 17711 9338
rect 17745 9304 17791 9338
rect 17825 9304 17871 9338
rect 17905 9304 17951 9338
rect 17985 9304 18031 9338
rect 18065 9304 18111 9338
rect 18145 9304 18191 9338
rect 18225 9304 18271 9338
rect 18305 9304 18351 9338
rect 18385 9304 18431 9338
rect 18465 9304 18511 9338
rect 18545 9304 18591 9338
rect 18625 9304 18671 9338
rect 18705 9304 18751 9338
rect 18785 9304 18831 9338
rect 18865 9304 18911 9338
rect 18945 9304 18991 9338
rect 19025 9304 19071 9338
rect 19105 9304 19151 9338
rect 19185 9304 19231 9338
rect 19265 9304 19311 9338
rect 19345 9304 19391 9338
rect 19425 9304 19471 9338
rect 19505 9304 19551 9338
rect 19585 9304 19631 9338
rect 19665 9304 19711 9338
rect 19745 9304 19791 9338
rect 19825 9304 19871 9338
rect 19905 9304 19951 9338
rect 19985 9304 20031 9338
rect 20065 9304 20111 9338
rect 20145 9304 20191 9338
rect 20225 9304 20271 9338
rect 20305 9304 20351 9338
rect 20385 9304 20431 9338
rect 20465 9304 20511 9338
rect 20545 9304 20591 9338
rect 20625 9304 20671 9338
rect 20705 9304 20751 9338
rect 20785 9304 20831 9338
rect 20865 9304 20911 9338
rect 20945 9304 20991 9338
rect 21025 9304 21071 9338
rect 21105 9304 21151 9338
rect 21185 9304 21231 9338
rect 21265 9304 21311 9338
rect 21345 9304 21391 9338
rect 21425 9304 21471 9338
rect 21505 9304 21551 9338
rect 21585 9304 21631 9338
rect 21665 9304 21711 9338
rect 21745 9304 21791 9338
rect 21825 9304 21871 9338
rect 21905 9304 21951 9338
rect 21985 9304 22031 9338
rect 22065 9304 22111 9338
rect 22145 9304 22191 9338
rect 22225 9304 22271 9338
rect 22305 9304 22351 9338
rect 22385 9304 22431 9338
rect 22465 9304 22511 9338
rect 22545 9304 22591 9338
rect 22625 9304 22671 9338
rect 22705 9304 22751 9338
rect 22785 9304 22831 9338
rect 22865 9304 22911 9338
rect 22945 9304 22991 9338
rect 23025 9304 23071 9338
rect 23105 9304 23151 9338
rect 23185 9304 23231 9338
rect 23265 9304 23311 9338
rect 23345 9304 23391 9338
rect 23425 9304 23471 9338
rect 23505 9304 23551 9338
rect 23585 9304 23631 9338
rect 23665 9304 23711 9338
rect 23745 9304 23791 9338
rect 23825 9304 23871 9338
rect 23905 9304 23951 9338
rect 23985 9304 24031 9338
rect 24065 9304 24111 9338
rect 24145 9304 24191 9338
rect 24225 9304 24271 9338
rect 24305 9304 24351 9338
rect 24385 9304 24431 9338
rect 24465 9304 24511 9338
rect 24545 9304 24591 9338
rect 24625 9304 24671 9338
rect 24705 9304 24751 9338
rect 24785 9304 24831 9338
rect 24865 9304 24911 9338
rect 24945 9304 24991 9338
rect 25025 9304 25071 9338
rect 25105 9304 25151 9338
rect 25185 9304 25231 9338
rect 25265 9304 25311 9338
rect 25345 9304 25391 9338
rect 25425 9304 25471 9338
rect 25505 9304 25551 9338
rect 25585 9304 25631 9338
rect 25665 9304 25711 9338
rect 25745 9304 25791 9338
rect 25825 9304 25871 9338
rect 25905 9304 25951 9338
rect 25985 9304 26031 9338
rect 26065 9304 26111 9338
rect 26145 9304 26191 9338
rect 26225 9304 26271 9338
rect 26305 9304 26351 9338
rect 26385 9304 26431 9338
rect 26465 9304 26511 9338
rect 26545 9304 26591 9338
rect 26625 9304 26671 9338
rect 26705 9304 26751 9338
rect 26785 9304 26831 9338
rect 26865 9304 26911 9338
rect 26945 9304 26991 9338
rect 27025 9304 27071 9338
rect 27105 9304 27151 9338
rect 27185 9304 27231 9338
rect 27265 9304 27311 9338
rect 27345 9304 27391 9338
rect 27425 9304 27471 9338
rect 27505 9304 27551 9338
rect 27585 9304 27631 9338
rect 27665 9304 27711 9338
rect 27745 9304 27791 9338
rect 27825 9304 27871 9338
rect 27905 9304 27951 9338
rect 27985 9304 28031 9338
rect 28065 9304 28111 9338
rect 28145 9304 28191 9338
rect 28225 9304 28271 9338
rect 28305 9304 28351 9338
rect 28385 9304 28431 9338
rect 28465 9304 28511 9338
rect 28545 9304 28591 9338
rect 28625 9304 28671 9338
rect 28705 9304 28751 9338
rect 28785 9304 28831 9338
rect 28865 9304 28911 9338
rect 28945 9304 28991 9338
rect 29025 9304 29071 9338
rect 29105 9304 29151 9338
rect 29185 9304 29231 9338
rect 29265 9304 29311 9338
rect 29345 9304 29391 9338
rect 29425 9304 29471 9338
rect 29505 9304 29551 9338
rect 29585 9304 29631 9338
rect 29665 9304 29711 9338
rect 29745 9304 29791 9338
rect 29825 9304 29871 9338
rect 29905 9304 29951 9338
rect 29985 9304 30031 9338
rect 30065 9304 30111 9338
rect 30145 9304 30191 9338
rect 30225 9304 30271 9338
rect 30305 9304 30351 9338
rect 30385 9304 30431 9338
rect 30465 9304 30511 9338
rect 30545 9304 30591 9338
rect 30625 9304 30671 9338
rect 30705 9304 30751 9338
rect 30785 9304 30831 9338
rect 30865 9304 30911 9338
rect 30945 9304 30991 9338
rect 31025 9304 31071 9338
rect 31105 9304 31151 9338
rect 31185 9304 31231 9338
rect 31265 9304 31311 9338
rect 31345 9304 31391 9338
rect 31425 9304 31471 9338
rect 31505 9304 31551 9338
rect 31585 9304 31631 9338
rect 31665 9304 31711 9338
rect 31745 9304 31791 9338
rect 31825 9304 31871 9338
rect 31905 9304 31951 9338
rect 31985 9304 32031 9338
rect 32065 9304 32111 9338
rect 32145 9304 32191 9338
rect 32225 9304 32271 9338
rect 32305 9304 32351 9338
rect 32385 9304 32431 9338
rect 32465 9304 32511 9338
rect 32545 9304 32591 9338
rect 32625 9304 32671 9338
rect 32705 9304 32751 9338
rect 32785 9304 32831 9338
rect 32865 9304 32911 9338
rect 32945 9304 32991 9338
rect 33025 9304 33071 9338
rect 33105 9304 33151 9338
rect 33185 9304 33231 9338
rect 33265 9304 33311 9338
rect 33345 9304 33391 9338
rect 33425 9304 33471 9338
rect 33505 9304 33551 9338
rect 33585 9304 33631 9338
rect 33665 9304 33711 9338
rect 33745 9304 33791 9338
rect 33825 9304 33871 9338
rect 33905 9304 33951 9338
rect 33985 9304 34031 9338
rect 34065 9304 34111 9338
rect 34145 9304 34191 9338
rect 34225 9304 34271 9338
rect 34305 9304 34351 9338
rect 34385 9304 34431 9338
rect 34465 9304 34511 9338
rect 34545 9304 34591 9338
rect 34625 9304 34671 9338
rect 34705 9304 34751 9338
rect 34785 9304 34831 9338
rect 34865 9304 34911 9338
rect 34945 9304 34991 9338
rect 35025 9304 35071 9338
rect 35105 9304 35151 9338
rect 35185 9304 35231 9338
rect 35265 9304 35311 9338
rect 35345 9304 35391 9338
rect 35425 9304 35471 9338
rect 35505 9304 35551 9338
rect 35585 9304 35631 9338
rect 35665 9304 35711 9338
rect 35745 9304 35791 9338
rect 35825 9304 35871 9338
rect 35905 9304 35951 9338
rect 35985 9304 36031 9338
rect 36065 9304 36111 9338
rect 36145 9304 36191 9338
rect 36225 9304 36271 9338
rect 36305 9304 36351 9338
rect 36385 9304 36431 9338
rect 36465 9304 36511 9338
rect 36545 9304 36591 9338
rect 36625 9304 36671 9338
rect 36705 9304 36751 9338
rect 36785 9304 36831 9338
rect 36865 9304 36911 9338
rect 36945 9304 36991 9338
rect 37025 9304 37071 9338
rect 37105 9304 37151 9338
rect 37185 9304 37231 9338
rect 37265 9304 37311 9338
rect 37345 9304 37391 9338
rect 37425 9304 37471 9338
rect 37505 9304 37551 9338
rect 37585 9304 37631 9338
rect 37665 9304 37711 9338
rect 37745 9304 37791 9338
rect 37825 9304 37871 9338
rect 37905 9304 37951 9338
rect 37985 9304 38031 9338
rect 38065 9304 38111 9338
rect 38145 9304 38191 9338
rect 38225 9304 38271 9338
rect 38305 9304 38351 9338
rect 3744 9271 38351 9304
rect -3640 7967 1316 7983
rect -3640 7933 1266 7967
rect 1300 7933 1316 7967
rect -3640 7917 1316 7933
rect -3650 6737 -1290 6753
rect -3650 6703 -1340 6737
rect -1306 6703 -1290 6737
rect -3650 6687 -1290 6703
rect -37897 6360 35594 6393
rect -37897 6326 -37851 6360
rect -37817 6326 -37771 6360
rect -37737 6326 -37691 6360
rect -37657 6326 -37611 6360
rect -37577 6326 -37531 6360
rect -37497 6326 -37451 6360
rect -37417 6326 -37371 6360
rect -37337 6326 -37291 6360
rect -37257 6326 -37211 6360
rect -37177 6326 -37131 6360
rect -37097 6326 -37051 6360
rect -37017 6326 -36971 6360
rect -36937 6326 -36891 6360
rect -36857 6326 -36811 6360
rect -36777 6326 -36731 6360
rect -36697 6326 -36651 6360
rect -36617 6326 -36571 6360
rect -36537 6326 -36491 6360
rect -36457 6326 -36411 6360
rect -36377 6326 -36331 6360
rect -36297 6326 -36251 6360
rect -36217 6326 -36171 6360
rect -36137 6326 -36091 6360
rect -36057 6326 -36011 6360
rect -35977 6326 -35931 6360
rect -35897 6326 -35851 6360
rect -35817 6326 -35771 6360
rect -35737 6326 -35691 6360
rect -35657 6326 -35611 6360
rect -35577 6326 -35531 6360
rect -35497 6326 -35451 6360
rect -35417 6326 -35371 6360
rect -35337 6326 -35291 6360
rect -35257 6326 -35211 6360
rect -35177 6326 -35131 6360
rect -35097 6326 -35051 6360
rect -35017 6326 -34971 6360
rect -34937 6326 -34891 6360
rect -34857 6326 -34811 6360
rect -34777 6326 -34731 6360
rect -34697 6326 -34651 6360
rect -34617 6326 -34571 6360
rect -34537 6326 -34491 6360
rect -34457 6326 -34411 6360
rect -34377 6326 -34331 6360
rect -34297 6326 -34251 6360
rect -34217 6326 -34171 6360
rect -34137 6326 -34091 6360
rect -34057 6326 -34011 6360
rect -33977 6326 -33931 6360
rect -33897 6326 -33851 6360
rect -33817 6326 -33771 6360
rect -33737 6326 -33691 6360
rect -33657 6326 -33611 6360
rect -33577 6326 -33531 6360
rect -33497 6326 -33451 6360
rect -33417 6326 -33371 6360
rect -33337 6326 -33291 6360
rect -33257 6326 -33211 6360
rect -33177 6326 -33131 6360
rect -33097 6326 -33051 6360
rect -33017 6326 -32971 6360
rect -32937 6326 -32891 6360
rect -32857 6326 -32811 6360
rect -32777 6326 -32731 6360
rect -32697 6326 -32651 6360
rect -32617 6326 -32571 6360
rect -32537 6326 -32491 6360
rect -32457 6326 -32411 6360
rect -32377 6326 -32331 6360
rect -32297 6326 -32251 6360
rect -32217 6326 -32171 6360
rect -32137 6326 -32091 6360
rect -32057 6326 -32011 6360
rect -31977 6326 -31931 6360
rect -31897 6326 -31851 6360
rect -31817 6326 -31771 6360
rect -31737 6326 -31691 6360
rect -31657 6326 -31611 6360
rect -31577 6326 -31531 6360
rect -31497 6326 -31451 6360
rect -31417 6326 -31371 6360
rect -31337 6326 -31291 6360
rect -31257 6326 -31211 6360
rect -31177 6326 -31131 6360
rect -31097 6326 -31051 6360
rect -31017 6326 -30971 6360
rect -30937 6326 -30891 6360
rect -30857 6326 -30811 6360
rect -30777 6326 -30731 6360
rect -30697 6326 -30651 6360
rect -30617 6326 -30571 6360
rect -30537 6326 -30491 6360
rect -30457 6326 -30411 6360
rect -30377 6326 -30331 6360
rect -30297 6326 -30251 6360
rect -30217 6326 -30171 6360
rect -30137 6326 -30091 6360
rect -30057 6326 -30011 6360
rect -29977 6326 -29931 6360
rect -29897 6326 -29851 6360
rect -29817 6326 -29771 6360
rect -29737 6326 -29691 6360
rect -29657 6326 -29611 6360
rect -29577 6326 -29531 6360
rect -29497 6326 -29451 6360
rect -29417 6326 -29371 6360
rect -29337 6326 -29291 6360
rect -29257 6326 -29211 6360
rect -29177 6326 -29131 6360
rect -29097 6326 -29051 6360
rect -29017 6326 -28971 6360
rect -28937 6326 -28891 6360
rect -28857 6326 -28811 6360
rect -28777 6326 -28731 6360
rect -28697 6326 -28651 6360
rect -28617 6326 -28571 6360
rect -28537 6326 -28491 6360
rect -28457 6326 -28411 6360
rect -28377 6326 -28331 6360
rect -28297 6326 -28251 6360
rect -28217 6326 -28171 6360
rect -28137 6326 -28091 6360
rect -28057 6326 -28011 6360
rect -27977 6326 -27931 6360
rect -27897 6326 -27851 6360
rect -27817 6326 -27771 6360
rect -27737 6326 -27691 6360
rect -27657 6326 -27611 6360
rect -27577 6326 -27531 6360
rect -27497 6326 -27451 6360
rect -27417 6326 -27371 6360
rect -27337 6326 -27291 6360
rect -27257 6326 -27211 6360
rect -27177 6326 -27131 6360
rect -27097 6326 -27051 6360
rect -27017 6326 -26971 6360
rect -26937 6326 -26891 6360
rect -26857 6326 -26811 6360
rect -26777 6326 -26731 6360
rect -26697 6326 -26651 6360
rect -26617 6326 -26571 6360
rect -26537 6326 -26491 6360
rect -26457 6326 -26411 6360
rect -26377 6326 -26331 6360
rect -26297 6326 -26251 6360
rect -26217 6326 -26171 6360
rect -26137 6326 -26091 6360
rect -26057 6326 -26011 6360
rect -25977 6326 -25931 6360
rect -25897 6326 -25851 6360
rect -25817 6326 -25771 6360
rect -25737 6326 -25691 6360
rect -25657 6326 -25611 6360
rect -25577 6326 -25531 6360
rect -25497 6326 -25451 6360
rect -25417 6326 -25371 6360
rect -25337 6326 -25291 6360
rect -25257 6326 -25211 6360
rect -25177 6326 -25131 6360
rect -25097 6326 -25051 6360
rect -25017 6326 -24971 6360
rect -24937 6326 -24890 6360
rect -24856 6326 -24810 6360
rect -24776 6326 -24730 6360
rect -24696 6326 -24650 6360
rect -24616 6326 -24570 6360
rect -24536 6326 -24490 6360
rect -24456 6326 -24410 6360
rect -24376 6326 -24330 6360
rect -24296 6326 -24250 6360
rect -24216 6326 -24170 6360
rect -24136 6326 -24090 6360
rect -24056 6326 -24010 6360
rect -23976 6326 -23930 6360
rect -23896 6326 -23850 6360
rect -23816 6326 -23770 6360
rect -23736 6326 -23690 6360
rect -23656 6326 -23610 6360
rect -23576 6326 -23530 6360
rect -23496 6326 -23450 6360
rect -23416 6326 -23370 6360
rect -23336 6326 -23290 6360
rect -23256 6326 -23210 6360
rect -23176 6326 -23130 6360
rect -23096 6326 -23050 6360
rect -23016 6326 -22970 6360
rect -22936 6326 -22890 6360
rect -22856 6326 -22810 6360
rect -22776 6326 -22730 6360
rect -22696 6326 -22650 6360
rect -22616 6326 -22570 6360
rect -22536 6326 -22490 6360
rect -22456 6326 -22410 6360
rect -22376 6326 -22330 6360
rect -22296 6326 -22250 6360
rect -22216 6326 -22170 6360
rect -22136 6326 -22090 6360
rect -22056 6326 -22010 6360
rect -21976 6326 -21930 6360
rect -21896 6326 -21850 6360
rect -21816 6326 -21770 6360
rect -21736 6326 -21690 6360
rect -21656 6326 -21610 6360
rect -21576 6326 -21530 6360
rect -21496 6326 -21450 6360
rect -21416 6326 -21370 6360
rect -21336 6326 -21290 6360
rect -21256 6326 -21210 6360
rect -21176 6326 -21130 6360
rect -21096 6326 -21050 6360
rect -21016 6326 -20970 6360
rect -20936 6326 -20890 6360
rect -20856 6326 -20810 6360
rect -20776 6326 -20730 6360
rect -20696 6326 -20650 6360
rect -20616 6326 -20570 6360
rect -20536 6326 -20490 6360
rect -20456 6326 -20410 6360
rect -20376 6326 -20330 6360
rect -20296 6326 -20250 6360
rect -20216 6326 -20170 6360
rect -20136 6326 -20090 6360
rect -20056 6326 -20010 6360
rect -19976 6326 -19930 6360
rect -19896 6326 -19850 6360
rect -19816 6326 -19770 6360
rect -19736 6326 -19690 6360
rect -19656 6326 -19610 6360
rect -19576 6326 -19530 6360
rect -19496 6326 -19450 6360
rect -19416 6326 -19370 6360
rect -19336 6326 -19290 6360
rect -19256 6326 -19210 6360
rect -19176 6326 -19130 6360
rect -19096 6326 -19050 6360
rect -19016 6326 -18970 6360
rect -18936 6326 -18890 6360
rect -18856 6326 -18810 6360
rect -18776 6326 -18730 6360
rect -18696 6326 -18650 6360
rect -18616 6326 -18570 6360
rect -18536 6326 -18490 6360
rect -18456 6326 -18410 6360
rect -18376 6326 -18330 6360
rect -18296 6326 -18250 6360
rect -18216 6326 -18170 6360
rect -18136 6326 -18090 6360
rect -18056 6326 -18010 6360
rect -17976 6326 -17930 6360
rect -17896 6326 -17850 6360
rect -17816 6326 -17770 6360
rect -17736 6326 -17690 6360
rect -17656 6326 -17610 6360
rect -17576 6326 -17530 6360
rect -17496 6326 -17450 6360
rect -17416 6326 -17370 6360
rect -17336 6326 -17290 6360
rect -17256 6326 -17210 6360
rect -17176 6326 -17130 6360
rect -17096 6326 -17050 6360
rect -17016 6326 -16970 6360
rect -16936 6326 -16890 6360
rect -16856 6326 -16810 6360
rect -16776 6326 -16730 6360
rect -16696 6326 -16650 6360
rect -16616 6326 -16570 6360
rect -16536 6326 -16490 6360
rect -16456 6326 -16410 6360
rect -16376 6326 -16330 6360
rect -16296 6326 -16250 6360
rect -16216 6326 -16170 6360
rect -16136 6326 -16090 6360
rect -16056 6326 -16010 6360
rect -15976 6326 -15930 6360
rect -15896 6326 -15850 6360
rect -15816 6326 -15770 6360
rect -15736 6326 -15690 6360
rect -15656 6326 -15610 6360
rect -15576 6326 -15530 6360
rect -15496 6326 -15450 6360
rect -15416 6326 -15370 6360
rect -15336 6326 -15290 6360
rect -15256 6326 -15210 6360
rect -15176 6326 -15130 6360
rect -15096 6326 -15050 6360
rect -15016 6326 -14970 6360
rect -14936 6326 -14890 6360
rect -14856 6326 -14810 6360
rect -14776 6326 -14730 6360
rect -14696 6326 -14650 6360
rect -14616 6326 -14570 6360
rect -14536 6326 -14490 6360
rect -14456 6326 -14410 6360
rect -14376 6326 -14330 6360
rect -14296 6326 -14250 6360
rect -14216 6326 -14170 6360
rect -14136 6326 -14090 6360
rect -14056 6326 -14010 6360
rect -13976 6326 -13930 6360
rect -13896 6326 -13850 6360
rect -13816 6326 -13770 6360
rect -13736 6326 -13690 6360
rect -13656 6326 -13610 6360
rect -13576 6326 -13530 6360
rect -13496 6326 -13450 6360
rect -13416 6326 -13370 6360
rect -13336 6326 -13290 6360
rect -13256 6326 -13210 6360
rect -13176 6326 -13130 6360
rect -13096 6326 -13050 6360
rect -13016 6326 -12970 6360
rect -12936 6326 -12890 6360
rect -12856 6326 -12810 6360
rect -12776 6326 -12730 6360
rect -12696 6326 -12650 6360
rect -12616 6326 -12570 6360
rect -12536 6326 -12490 6360
rect -12456 6326 -12410 6360
rect -12376 6326 -12330 6360
rect -12296 6326 -12250 6360
rect -12216 6326 -12170 6360
rect -12136 6326 -12090 6360
rect -12056 6326 -12010 6360
rect -11976 6326 -11929 6360
rect -11895 6326 -11849 6360
rect -11815 6326 -11769 6360
rect -11735 6326 -11689 6360
rect -11655 6326 -11609 6360
rect -11575 6326 -11529 6360
rect -11495 6326 -11449 6360
rect -11415 6326 -11369 6360
rect -11335 6326 -11289 6360
rect -11255 6326 -11209 6360
rect -11175 6326 -11129 6360
rect -11095 6326 -11049 6360
rect -11015 6326 -10969 6360
rect -10935 6326 -10889 6360
rect -10855 6326 -10809 6360
rect -10775 6326 -10729 6360
rect -10695 6326 -10649 6360
rect -10615 6326 -10569 6360
rect -10535 6326 -10489 6360
rect -10455 6326 -10409 6360
rect -10375 6326 -10329 6360
rect -10295 6326 -10249 6360
rect -10215 6326 -10169 6360
rect -10135 6326 -10089 6360
rect -10055 6326 -10009 6360
rect -9975 6326 -9929 6360
rect -9895 6326 -9849 6360
rect -9815 6326 -9769 6360
rect -9735 6326 -9689 6360
rect -9655 6326 -9609 6360
rect -9575 6326 -9529 6360
rect -9495 6326 -9449 6360
rect -9415 6326 -9369 6360
rect -9335 6326 -9289 6360
rect -9255 6326 -9209 6360
rect -9175 6326 -9129 6360
rect -9095 6326 -9049 6360
rect -9015 6326 -8969 6360
rect -8935 6326 -8889 6360
rect -8855 6326 -8809 6360
rect -8775 6326 -8729 6360
rect -8695 6326 -8649 6360
rect -8615 6326 -8569 6360
rect -8535 6326 -8489 6360
rect -8455 6326 -8409 6360
rect -8375 6326 -8329 6360
rect -8295 6326 -8249 6360
rect -8215 6326 -8169 6360
rect -8135 6326 -8089 6360
rect -8055 6326 -8009 6360
rect -7975 6326 -7929 6360
rect -7895 6326 -7849 6360
rect -7815 6326 -7769 6360
rect -7735 6326 -7689 6360
rect -7655 6326 -7609 6360
rect -7575 6326 -7529 6360
rect -7495 6326 -7449 6360
rect -7415 6326 -7369 6360
rect -7335 6326 -7289 6360
rect -7255 6326 -7209 6360
rect -7175 6326 -7129 6360
rect -7095 6326 -7049 6360
rect -7015 6326 -6969 6360
rect -6935 6326 -6889 6360
rect -6855 6326 -6809 6360
rect -6775 6326 -6729 6360
rect -6695 6326 -6649 6360
rect -6615 6326 -6569 6360
rect -6535 6326 -6489 6360
rect -6455 6326 -6409 6360
rect -6375 6326 -6329 6360
rect -6295 6326 -6249 6360
rect -6215 6326 -6169 6360
rect -6135 6326 -6089 6360
rect -6055 6326 -6009 6360
rect -5975 6326 -5929 6360
rect -5895 6326 -5849 6360
rect -5815 6326 -5769 6360
rect -5735 6326 -5689 6360
rect -5655 6326 -5609 6360
rect -5575 6326 -5529 6360
rect -5495 6326 -5449 6360
rect -5415 6326 -5369 6360
rect -5335 6326 -5289 6360
rect -5255 6326 -5209 6360
rect -5175 6326 -5129 6360
rect -5095 6326 -5049 6360
rect -5015 6326 -4969 6360
rect -4935 6326 -4889 6360
rect -4855 6326 -4809 6360
rect -4775 6326 -4729 6360
rect -4695 6326 -4649 6360
rect -4615 6326 -4569 6360
rect -4535 6326 -4489 6360
rect -4455 6326 -4409 6360
rect -4375 6326 -4329 6360
rect -4295 6326 -4249 6360
rect -4215 6326 -4169 6360
rect -4135 6326 -4089 6360
rect -4055 6326 -4009 6360
rect -3975 6326 -3929 6360
rect -3895 6326 -3849 6360
rect -3815 6326 -3769 6360
rect -3735 6326 -3689 6360
rect -3655 6326 -3609 6360
rect -3575 6326 -3529 6360
rect -3495 6326 -3449 6360
rect -3415 6326 -3369 6360
rect -3335 6326 -3289 6360
rect -3255 6326 -3209 6360
rect -3175 6326 -3129 6360
rect -3095 6326 -3049 6360
rect -3015 6326 -2969 6360
rect -2935 6326 -2889 6360
rect -2855 6326 -2809 6360
rect -2775 6326 -2729 6360
rect -2695 6326 -2649 6360
rect -2615 6326 -2569 6360
rect -2535 6326 -2489 6360
rect -2455 6326 -2409 6360
rect -2375 6326 -2329 6360
rect -2295 6326 -2249 6360
rect -2215 6326 -2169 6360
rect -2135 6326 -2089 6360
rect -2055 6326 -2009 6360
rect -1975 6326 -1929 6360
rect -1895 6326 -1849 6360
rect -1815 6326 -1769 6360
rect -1735 6326 -1689 6360
rect -1655 6326 -1609 6360
rect -1575 6326 -1529 6360
rect -1495 6326 -1449 6360
rect -1415 6326 -1369 6360
rect -1335 6326 -1289 6360
rect -1255 6326 -1209 6360
rect -1175 6326 -1129 6360
rect -1095 6326 -1049 6360
rect -1015 6326 -969 6360
rect -935 6326 -889 6360
rect -855 6326 -809 6360
rect -775 6326 -729 6360
rect -695 6326 -649 6360
rect -615 6326 -569 6360
rect -535 6326 -489 6360
rect -455 6326 -409 6360
rect -375 6326 -329 6360
rect -295 6326 -249 6360
rect -215 6326 -169 6360
rect -135 6326 -89 6360
rect -55 6326 -9 6360
rect 25 6326 71 6360
rect 105 6326 151 6360
rect 185 6326 231 6360
rect 265 6326 311 6360
rect 345 6326 391 6360
rect 425 6326 471 6360
rect 505 6326 551 6360
rect 585 6326 631 6360
rect 665 6326 711 6360
rect 745 6326 791 6360
rect 825 6326 871 6360
rect 905 6326 951 6360
rect 985 6326 1031 6360
rect 1065 6326 1111 6360
rect 1145 6326 1191 6360
rect 1225 6326 1271 6360
rect 1305 6326 1351 6360
rect 1385 6326 1431 6360
rect 1465 6326 1511 6360
rect 1545 6326 1591 6360
rect 1625 6326 1671 6360
rect 1705 6326 1751 6360
rect 1785 6326 1831 6360
rect 1865 6326 1911 6360
rect 1945 6326 1991 6360
rect 2025 6326 2071 6360
rect 2105 6326 2151 6360
rect 2185 6326 2231 6360
rect 2265 6326 2311 6360
rect 2345 6326 2391 6360
rect 2425 6326 2471 6360
rect 2505 6326 2551 6360
rect 2585 6326 2631 6360
rect 2665 6326 2711 6360
rect 2745 6326 2791 6360
rect 2825 6326 2871 6360
rect 2905 6326 2951 6360
rect 2985 6326 3031 6360
rect 3065 6326 3111 6360
rect 3145 6326 3191 6360
rect 3225 6326 3271 6360
rect 3305 6326 3351 6360
rect 3385 6326 3431 6360
rect 3465 6326 3511 6360
rect 3545 6326 3591 6360
rect 3625 6326 3671 6360
rect 3705 6326 3751 6360
rect 3785 6326 3831 6360
rect 3865 6326 3911 6360
rect 3945 6326 3991 6360
rect 4025 6326 4071 6360
rect 4105 6326 4151 6360
rect 4185 6326 4231 6360
rect 4265 6326 4311 6360
rect 4345 6326 4391 6360
rect 4425 6326 4471 6360
rect 4505 6326 4551 6360
rect 4585 6326 4631 6360
rect 4665 6326 4711 6360
rect 4745 6326 4791 6360
rect 4825 6326 4871 6360
rect 4905 6326 4951 6360
rect 4985 6326 5031 6360
rect 5065 6326 5111 6360
rect 5145 6326 5191 6360
rect 5225 6326 5271 6360
rect 5305 6326 5351 6360
rect 5385 6326 5431 6360
rect 5465 6326 5511 6360
rect 5545 6326 5591 6360
rect 5625 6326 5671 6360
rect 5705 6326 5751 6360
rect 5785 6326 5831 6360
rect 5865 6326 5911 6360
rect 5945 6326 5991 6360
rect 6025 6326 6071 6360
rect 6105 6326 6151 6360
rect 6185 6326 6231 6360
rect 6265 6326 6311 6360
rect 6345 6326 6391 6360
rect 6425 6326 6471 6360
rect 6505 6326 6551 6360
rect 6585 6326 6631 6360
rect 6665 6326 6711 6360
rect 6745 6326 6791 6360
rect 6825 6326 6871 6360
rect 6905 6326 6951 6360
rect 6985 6326 7031 6360
rect 7065 6326 7111 6360
rect 7145 6326 7191 6360
rect 7225 6326 7271 6360
rect 7305 6326 7351 6360
rect 7385 6326 7431 6360
rect 7465 6326 7511 6360
rect 7545 6326 7591 6360
rect 7625 6326 7671 6360
rect 7705 6326 7751 6360
rect 7785 6326 7831 6360
rect 7865 6326 7911 6360
rect 7945 6326 7991 6360
rect 8025 6326 8071 6360
rect 8105 6326 8151 6360
rect 8185 6326 8231 6360
rect 8265 6326 8311 6360
rect 8345 6326 8391 6360
rect 8425 6326 8471 6360
rect 8505 6326 8551 6360
rect 8585 6326 8631 6360
rect 8665 6326 8711 6360
rect 8745 6326 8791 6360
rect 8825 6326 8871 6360
rect 8905 6326 8951 6360
rect 8985 6326 9031 6360
rect 9065 6326 9111 6360
rect 9145 6326 9191 6360
rect 9225 6326 9271 6360
rect 9305 6326 9351 6360
rect 9385 6326 9431 6360
rect 9465 6326 9511 6360
rect 9545 6326 9591 6360
rect 9625 6326 9672 6360
rect 9706 6326 9752 6360
rect 9786 6326 9832 6360
rect 9866 6326 9912 6360
rect 9946 6326 9992 6360
rect 10026 6326 10072 6360
rect 10106 6326 10152 6360
rect 10186 6326 10232 6360
rect 10266 6326 10312 6360
rect 10346 6326 10392 6360
rect 10426 6326 10472 6360
rect 10506 6326 10552 6360
rect 10586 6326 10632 6360
rect 10666 6326 10712 6360
rect 10746 6326 10792 6360
rect 10826 6326 10872 6360
rect 10906 6326 10952 6360
rect 10986 6326 11032 6360
rect 11066 6326 11112 6360
rect 11146 6326 11192 6360
rect 11226 6326 11272 6360
rect 11306 6326 11352 6360
rect 11386 6326 11432 6360
rect 11466 6326 11512 6360
rect 11546 6326 11592 6360
rect 11626 6326 11672 6360
rect 11706 6326 11752 6360
rect 11786 6326 11832 6360
rect 11866 6326 11912 6360
rect 11946 6326 11992 6360
rect 12026 6326 12072 6360
rect 12106 6326 12152 6360
rect 12186 6326 12232 6360
rect 12266 6326 12312 6360
rect 12346 6326 12392 6360
rect 12426 6326 12472 6360
rect 12506 6326 12552 6360
rect 12586 6326 12632 6360
rect 12666 6326 12712 6360
rect 12746 6326 12792 6360
rect 12826 6326 12872 6360
rect 12906 6326 12952 6360
rect 12986 6326 13032 6360
rect 13066 6326 13112 6360
rect 13146 6326 13192 6360
rect 13226 6326 13272 6360
rect 13306 6326 13352 6360
rect 13386 6326 13432 6360
rect 13466 6326 13512 6360
rect 13546 6326 13592 6360
rect 13626 6326 13672 6360
rect 13706 6326 13752 6360
rect 13786 6326 13832 6360
rect 13866 6326 13912 6360
rect 13946 6326 13992 6360
rect 14026 6326 14072 6360
rect 14106 6326 14152 6360
rect 14186 6326 14232 6360
rect 14266 6326 14312 6360
rect 14346 6326 14392 6360
rect 14426 6326 14472 6360
rect 14506 6326 14552 6360
rect 14586 6326 14632 6360
rect 14666 6326 14712 6360
rect 14746 6326 14792 6360
rect 14826 6326 14872 6360
rect 14906 6326 14952 6360
rect 14986 6326 15032 6360
rect 15066 6326 15112 6360
rect 15146 6326 15192 6360
rect 15226 6326 15272 6360
rect 15306 6326 15352 6360
rect 15386 6326 15432 6360
rect 15466 6326 15512 6360
rect 15546 6326 15592 6360
rect 15626 6326 15672 6360
rect 15706 6326 15752 6360
rect 15786 6326 15832 6360
rect 15866 6326 15912 6360
rect 15946 6326 15992 6360
rect 16026 6326 16072 6360
rect 16106 6326 16152 6360
rect 16186 6326 16232 6360
rect 16266 6326 16312 6360
rect 16346 6326 16392 6360
rect 16426 6326 16472 6360
rect 16506 6326 16552 6360
rect 16586 6326 16632 6360
rect 16666 6326 16712 6360
rect 16746 6326 16792 6360
rect 16826 6326 16872 6360
rect 16906 6326 16952 6360
rect 16986 6326 17032 6360
rect 17066 6326 17112 6360
rect 17146 6326 17192 6360
rect 17226 6326 17272 6360
rect 17306 6326 17352 6360
rect 17386 6326 17432 6360
rect 17466 6326 17512 6360
rect 17546 6326 17592 6360
rect 17626 6326 17672 6360
rect 17706 6326 17752 6360
rect 17786 6326 17832 6360
rect 17866 6326 17912 6360
rect 17946 6326 17992 6360
rect 18026 6326 18072 6360
rect 18106 6326 18152 6360
rect 18186 6326 18232 6360
rect 18266 6326 18312 6360
rect 18346 6326 18392 6360
rect 18426 6326 18472 6360
rect 18506 6326 18552 6360
rect 18586 6326 18632 6360
rect 18666 6326 18712 6360
rect 18746 6326 18792 6360
rect 18826 6326 18872 6360
rect 18906 6326 18952 6360
rect 18986 6326 19032 6360
rect 19066 6326 19112 6360
rect 19146 6326 19192 6360
rect 19226 6326 19272 6360
rect 19306 6326 19352 6360
rect 19386 6326 19432 6360
rect 19466 6326 19512 6360
rect 19546 6326 19592 6360
rect 19626 6326 19672 6360
rect 19706 6326 19752 6360
rect 19786 6326 19832 6360
rect 19866 6326 19912 6360
rect 19946 6326 19992 6360
rect 20026 6326 20072 6360
rect 20106 6326 20152 6360
rect 20186 6326 20232 6360
rect 20266 6326 20312 6360
rect 20346 6326 20392 6360
rect 20426 6326 20472 6360
rect 20506 6326 20552 6360
rect 20586 6326 20632 6360
rect 20666 6326 20712 6360
rect 20746 6326 20792 6360
rect 20826 6326 20872 6360
rect 20906 6326 20952 6360
rect 20986 6326 21032 6360
rect 21066 6326 21112 6360
rect 21146 6326 21192 6360
rect 21226 6326 21272 6360
rect 21306 6326 21352 6360
rect 21386 6326 21432 6360
rect 21466 6326 21512 6360
rect 21546 6326 21592 6360
rect 21626 6326 21672 6360
rect 21706 6326 21752 6360
rect 21786 6326 21832 6360
rect 21866 6326 21912 6360
rect 21946 6326 21992 6360
rect 22026 6326 22072 6360
rect 22106 6326 22152 6360
rect 22186 6326 22232 6360
rect 22266 6326 22312 6360
rect 22346 6326 22392 6360
rect 22426 6326 22472 6360
rect 22506 6326 22552 6360
rect 22586 6326 22633 6360
rect 22667 6326 22713 6360
rect 22747 6326 22793 6360
rect 22827 6326 22873 6360
rect 22907 6326 22953 6360
rect 22987 6326 23033 6360
rect 23067 6326 23113 6360
rect 23147 6326 23193 6360
rect 23227 6326 23273 6360
rect 23307 6326 23353 6360
rect 23387 6326 23433 6360
rect 23467 6326 23513 6360
rect 23547 6326 23593 6360
rect 23627 6326 23673 6360
rect 23707 6326 23753 6360
rect 23787 6326 23833 6360
rect 23867 6326 23913 6360
rect 23947 6326 23993 6360
rect 24027 6326 24073 6360
rect 24107 6326 24153 6360
rect 24187 6326 24233 6360
rect 24267 6326 24313 6360
rect 24347 6326 24393 6360
rect 24427 6326 24473 6360
rect 24507 6326 24553 6360
rect 24587 6326 24633 6360
rect 24667 6326 24713 6360
rect 24747 6326 24793 6360
rect 24827 6326 24873 6360
rect 24907 6326 24953 6360
rect 24987 6326 25033 6360
rect 25067 6326 25113 6360
rect 25147 6326 25193 6360
rect 25227 6326 25273 6360
rect 25307 6326 25353 6360
rect 25387 6326 25433 6360
rect 25467 6326 25513 6360
rect 25547 6326 25593 6360
rect 25627 6326 25673 6360
rect 25707 6326 25753 6360
rect 25787 6326 25833 6360
rect 25867 6326 25913 6360
rect 25947 6326 25993 6360
rect 26027 6326 26073 6360
rect 26107 6326 26153 6360
rect 26187 6326 26233 6360
rect 26267 6326 26313 6360
rect 26347 6326 26393 6360
rect 26427 6326 26473 6360
rect 26507 6326 26553 6360
rect 26587 6326 26633 6360
rect 26667 6326 26713 6360
rect 26747 6326 26793 6360
rect 26827 6326 26873 6360
rect 26907 6326 26953 6360
rect 26987 6326 27033 6360
rect 27067 6326 27113 6360
rect 27147 6326 27193 6360
rect 27227 6326 27273 6360
rect 27307 6326 27353 6360
rect 27387 6326 27433 6360
rect 27467 6326 27513 6360
rect 27547 6326 27593 6360
rect 27627 6326 27673 6360
rect 27707 6326 27753 6360
rect 27787 6326 27833 6360
rect 27867 6326 27913 6360
rect 27947 6326 27993 6360
rect 28027 6326 28073 6360
rect 28107 6326 28153 6360
rect 28187 6326 28233 6360
rect 28267 6326 28313 6360
rect 28347 6326 28393 6360
rect 28427 6326 28473 6360
rect 28507 6326 28553 6360
rect 28587 6326 28633 6360
rect 28667 6326 28713 6360
rect 28747 6326 28793 6360
rect 28827 6326 28873 6360
rect 28907 6326 28953 6360
rect 28987 6326 29033 6360
rect 29067 6326 29113 6360
rect 29147 6326 29193 6360
rect 29227 6326 29273 6360
rect 29307 6326 29353 6360
rect 29387 6326 29433 6360
rect 29467 6326 29513 6360
rect 29547 6326 29593 6360
rect 29627 6326 29673 6360
rect 29707 6326 29753 6360
rect 29787 6326 29833 6360
rect 29867 6326 29913 6360
rect 29947 6326 29993 6360
rect 30027 6326 30073 6360
rect 30107 6326 30153 6360
rect 30187 6326 30233 6360
rect 30267 6326 30313 6360
rect 30347 6326 30393 6360
rect 30427 6326 30473 6360
rect 30507 6326 30553 6360
rect 30587 6326 30633 6360
rect 30667 6326 30713 6360
rect 30747 6326 30793 6360
rect 30827 6326 30873 6360
rect 30907 6326 30953 6360
rect 30987 6326 31033 6360
rect 31067 6326 31113 6360
rect 31147 6326 31193 6360
rect 31227 6326 31274 6360
rect 31308 6326 31354 6360
rect 31388 6326 31434 6360
rect 31468 6326 31514 6360
rect 31548 6326 31594 6360
rect 31628 6326 31674 6360
rect 31708 6326 31754 6360
rect 31788 6326 31834 6360
rect 31868 6326 31914 6360
rect 31948 6326 31994 6360
rect 32028 6326 32074 6360
rect 32108 6326 32154 6360
rect 32188 6326 32234 6360
rect 32268 6326 32314 6360
rect 32348 6326 32394 6360
rect 32428 6326 32474 6360
rect 32508 6326 32554 6360
rect 32588 6326 32634 6360
rect 32668 6326 32714 6360
rect 32748 6326 32794 6360
rect 32828 6326 32874 6360
rect 32908 6326 32954 6360
rect 32988 6326 33034 6360
rect 33068 6326 33114 6360
rect 33148 6326 33194 6360
rect 33228 6326 33274 6360
rect 33308 6326 33354 6360
rect 33388 6326 33434 6360
rect 33468 6326 33514 6360
rect 33548 6326 33594 6360
rect 33628 6326 33674 6360
rect 33708 6326 33754 6360
rect 33788 6326 33834 6360
rect 33868 6326 33914 6360
rect 33948 6326 33994 6360
rect 34028 6326 34074 6360
rect 34108 6326 34154 6360
rect 34188 6326 34234 6360
rect 34268 6326 34314 6360
rect 34348 6326 34394 6360
rect 34428 6326 34474 6360
rect 34508 6326 34554 6360
rect 34588 6326 34634 6360
rect 34668 6326 34714 6360
rect 34748 6326 34794 6360
rect 34828 6326 34874 6360
rect 34908 6326 34954 6360
rect 34988 6326 35034 6360
rect 35068 6326 35114 6360
rect 35148 6326 35194 6360
rect 35228 6326 35274 6360
rect 35308 6326 35354 6360
rect 35388 6326 35434 6360
rect 35468 6326 35514 6360
rect 35548 6326 35594 6360
rect -37897 6293 35594 6326
rect -34951 4821 -343 4854
rect -34951 4787 -34905 4821
rect -34871 4787 -34825 4821
rect -34791 4787 -34745 4821
rect -34711 4787 -34665 4821
rect -34631 4787 -34585 4821
rect -34551 4787 -34505 4821
rect -34471 4787 -34425 4821
rect -34391 4787 -34345 4821
rect -34311 4787 -34265 4821
rect -34231 4787 -34185 4821
rect -34151 4787 -34105 4821
rect -34071 4787 -34025 4821
rect -33991 4787 -33945 4821
rect -33911 4787 -33865 4821
rect -33831 4787 -33785 4821
rect -33751 4787 -33705 4821
rect -33671 4787 -33625 4821
rect -33591 4787 -33545 4821
rect -33511 4787 -33465 4821
rect -33431 4787 -33385 4821
rect -33351 4787 -33305 4821
rect -33271 4787 -33225 4821
rect -33191 4787 -33145 4821
rect -33111 4787 -33065 4821
rect -33031 4787 -32985 4821
rect -32951 4787 -32905 4821
rect -32871 4787 -32825 4821
rect -32791 4787 -32745 4821
rect -32711 4787 -32665 4821
rect -32631 4787 -32585 4821
rect -32551 4787 -32505 4821
rect -32471 4787 -32425 4821
rect -32391 4787 -32345 4821
rect -32311 4787 -32265 4821
rect -32231 4787 -32185 4821
rect -32151 4787 -32105 4821
rect -32071 4787 -32025 4821
rect -31991 4787 -31945 4821
rect -31911 4787 -31865 4821
rect -31831 4787 -31785 4821
rect -31751 4787 -31705 4821
rect -31671 4787 -31625 4821
rect -31591 4787 -31545 4821
rect -31511 4787 -31465 4821
rect -31431 4787 -31385 4821
rect -31351 4787 -31305 4821
rect -31271 4787 -31225 4821
rect -31191 4787 -31145 4821
rect -31111 4787 -31065 4821
rect -31031 4787 -30985 4821
rect -30951 4787 -30905 4821
rect -30871 4787 -30825 4821
rect -30791 4787 -30745 4821
rect -30711 4787 -30665 4821
rect -30631 4787 -30585 4821
rect -30551 4787 -30505 4821
rect -30471 4787 -30425 4821
rect -30391 4787 -30345 4821
rect -30311 4787 -30265 4821
rect -30231 4787 -30185 4821
rect -30151 4787 -30105 4821
rect -30071 4787 -30025 4821
rect -29991 4787 -29945 4821
rect -29911 4787 -29865 4821
rect -29831 4787 -29785 4821
rect -29751 4787 -29705 4821
rect -29671 4787 -29625 4821
rect -29591 4787 -29545 4821
rect -29511 4787 -29465 4821
rect -29431 4787 -29385 4821
rect -29351 4787 -29305 4821
rect -29271 4787 -29225 4821
rect -29191 4787 -29145 4821
rect -29111 4787 -29065 4821
rect -29031 4787 -28985 4821
rect -28951 4787 -28905 4821
rect -28871 4787 -28825 4821
rect -28791 4787 -28745 4821
rect -28711 4787 -28665 4821
rect -28631 4787 -28585 4821
rect -28551 4787 -28505 4821
rect -28471 4787 -28425 4821
rect -28391 4787 -28345 4821
rect -28311 4787 -28265 4821
rect -28231 4787 -28185 4821
rect -28151 4787 -28105 4821
rect -28071 4787 -28025 4821
rect -27991 4787 -27945 4821
rect -27911 4787 -27865 4821
rect -27831 4787 -27785 4821
rect -27751 4787 -27705 4821
rect -27671 4787 -27625 4821
rect -27591 4787 -27545 4821
rect -27511 4787 -27465 4821
rect -27431 4787 -27385 4821
rect -27351 4787 -27305 4821
rect -27271 4787 -27225 4821
rect -27191 4787 -27145 4821
rect -27111 4787 -27065 4821
rect -27031 4787 -26985 4821
rect -26951 4787 -26905 4821
rect -26871 4787 -26825 4821
rect -26791 4787 -26745 4821
rect -26711 4787 -26665 4821
rect -26631 4787 -26585 4821
rect -26551 4787 -26505 4821
rect -26471 4787 -26425 4821
rect -26391 4787 -26345 4821
rect -26311 4787 -26265 4821
rect -26231 4787 -26185 4821
rect -26151 4787 -26105 4821
rect -26071 4787 -26025 4821
rect -25991 4787 -25945 4821
rect -25911 4787 -25865 4821
rect -25831 4787 -25785 4821
rect -25751 4787 -25705 4821
rect -25671 4787 -25625 4821
rect -25591 4787 -25545 4821
rect -25511 4787 -25465 4821
rect -25431 4787 -25385 4821
rect -25351 4787 -25305 4821
rect -25271 4787 -25225 4821
rect -25191 4787 -25145 4821
rect -25111 4787 -25065 4821
rect -25031 4787 -24985 4821
rect -24951 4787 -24905 4821
rect -24871 4787 -24825 4821
rect -24791 4787 -24745 4821
rect -24711 4787 -24665 4821
rect -24631 4787 -24585 4821
rect -24551 4787 -24505 4821
rect -24471 4787 -24425 4821
rect -24391 4787 -24345 4821
rect -24311 4787 -24265 4821
rect -24231 4787 -24185 4821
rect -24151 4787 -24105 4821
rect -24071 4787 -24025 4821
rect -23991 4787 -23945 4821
rect -23911 4787 -23865 4821
rect -23831 4787 -23785 4821
rect -23751 4787 -23705 4821
rect -23671 4787 -23625 4821
rect -23591 4787 -23545 4821
rect -23511 4787 -23465 4821
rect -23431 4787 -23385 4821
rect -23351 4787 -23305 4821
rect -23271 4787 -23225 4821
rect -23191 4787 -23145 4821
rect -23111 4787 -23065 4821
rect -23031 4787 -22985 4821
rect -22951 4787 -22905 4821
rect -22871 4787 -22825 4821
rect -22791 4787 -22745 4821
rect -22711 4787 -22665 4821
rect -22631 4787 -22585 4821
rect -22551 4787 -22505 4821
rect -22471 4787 -22425 4821
rect -22391 4787 -22345 4821
rect -22311 4787 -22265 4821
rect -22231 4787 -22185 4821
rect -22151 4787 -22105 4821
rect -22071 4787 -22025 4821
rect -21991 4787 -21944 4821
rect -21910 4787 -21864 4821
rect -21830 4787 -21784 4821
rect -21750 4787 -21704 4821
rect -21670 4787 -21624 4821
rect -21590 4787 -21544 4821
rect -21510 4787 -21464 4821
rect -21430 4787 -21384 4821
rect -21350 4787 -21304 4821
rect -21270 4787 -21224 4821
rect -21190 4787 -21144 4821
rect -21110 4787 -21064 4821
rect -21030 4787 -20984 4821
rect -20950 4787 -20904 4821
rect -20870 4787 -20824 4821
rect -20790 4787 -20744 4821
rect -20710 4787 -20664 4821
rect -20630 4787 -20584 4821
rect -20550 4787 -20504 4821
rect -20470 4787 -20424 4821
rect -20390 4787 -20344 4821
rect -20310 4787 -20264 4821
rect -20230 4787 -20184 4821
rect -20150 4787 -20104 4821
rect -20070 4787 -20024 4821
rect -19990 4787 -19944 4821
rect -19910 4787 -19864 4821
rect -19830 4787 -19784 4821
rect -19750 4787 -19704 4821
rect -19670 4787 -19624 4821
rect -19590 4787 -19544 4821
rect -19510 4787 -19464 4821
rect -19430 4787 -19384 4821
rect -19350 4787 -19304 4821
rect -19270 4787 -19224 4821
rect -19190 4787 -19144 4821
rect -19110 4787 -19064 4821
rect -19030 4787 -18984 4821
rect -18950 4787 -18904 4821
rect -18870 4787 -18824 4821
rect -18790 4787 -18744 4821
rect -18710 4787 -18664 4821
rect -18630 4787 -18584 4821
rect -18550 4787 -18504 4821
rect -18470 4787 -18424 4821
rect -18390 4787 -18344 4821
rect -18310 4787 -18264 4821
rect -18230 4787 -18184 4821
rect -18150 4787 -18104 4821
rect -18070 4787 -18024 4821
rect -17990 4787 -17944 4821
rect -17910 4787 -17864 4821
rect -17830 4787 -17784 4821
rect -17750 4787 -17704 4821
rect -17670 4787 -17624 4821
rect -17590 4787 -17544 4821
rect -17510 4787 -17464 4821
rect -17430 4787 -17384 4821
rect -17350 4787 -17304 4821
rect -17270 4787 -17224 4821
rect -17190 4787 -17144 4821
rect -17110 4787 -17064 4821
rect -17030 4787 -16984 4821
rect -16950 4787 -16904 4821
rect -16870 4787 -16824 4821
rect -16790 4787 -16744 4821
rect -16710 4787 -16664 4821
rect -16630 4787 -16584 4821
rect -16550 4787 -16504 4821
rect -16470 4787 -16424 4821
rect -16390 4787 -16344 4821
rect -16310 4787 -16264 4821
rect -16230 4787 -16184 4821
rect -16150 4787 -16104 4821
rect -16070 4787 -16024 4821
rect -15990 4787 -15944 4821
rect -15910 4787 -15864 4821
rect -15830 4787 -15784 4821
rect -15750 4787 -15704 4821
rect -15670 4787 -15624 4821
rect -15590 4787 -15544 4821
rect -15510 4787 -15464 4821
rect -15430 4787 -15384 4821
rect -15350 4787 -15304 4821
rect -15270 4787 -15224 4821
rect -15190 4787 -15144 4821
rect -15110 4787 -15064 4821
rect -15030 4787 -14984 4821
rect -14950 4787 -14904 4821
rect -14870 4787 -14824 4821
rect -14790 4787 -14744 4821
rect -14710 4787 -14664 4821
rect -14630 4787 -14584 4821
rect -14550 4787 -14504 4821
rect -14470 4787 -14424 4821
rect -14390 4787 -14344 4821
rect -14310 4787 -14264 4821
rect -14230 4787 -14184 4821
rect -14150 4787 -14104 4821
rect -14070 4787 -14024 4821
rect -13990 4787 -13944 4821
rect -13910 4787 -13864 4821
rect -13830 4787 -13784 4821
rect -13750 4787 -13704 4821
rect -13670 4787 -13624 4821
rect -13590 4787 -13544 4821
rect -13510 4787 -13464 4821
rect -13430 4787 -13384 4821
rect -13350 4787 -13304 4821
rect -13270 4787 -13224 4821
rect -13190 4787 -13144 4821
rect -13110 4787 -13064 4821
rect -13030 4787 -12984 4821
rect -12950 4787 -12904 4821
rect -12870 4787 -12824 4821
rect -12790 4787 -12744 4821
rect -12710 4787 -12664 4821
rect -12630 4787 -12584 4821
rect -12550 4787 -12504 4821
rect -12470 4787 -12424 4821
rect -12390 4787 -12344 4821
rect -12310 4787 -12264 4821
rect -12230 4787 -12184 4821
rect -12150 4787 -12104 4821
rect -12070 4787 -12024 4821
rect -11990 4787 -11944 4821
rect -11910 4787 -11864 4821
rect -11830 4787 -11784 4821
rect -11750 4787 -11704 4821
rect -11670 4787 -11624 4821
rect -11590 4787 -11544 4821
rect -11510 4787 -11464 4821
rect -11430 4787 -11384 4821
rect -11350 4787 -11304 4821
rect -11270 4787 -11224 4821
rect -11190 4787 -11144 4821
rect -11110 4787 -11064 4821
rect -11030 4787 -10984 4821
rect -10950 4787 -10904 4821
rect -10870 4787 -10824 4821
rect -10790 4787 -10744 4821
rect -10710 4787 -10664 4821
rect -10630 4787 -10584 4821
rect -10550 4787 -10504 4821
rect -10470 4787 -10424 4821
rect -10390 4787 -10344 4821
rect -10310 4787 -10264 4821
rect -10230 4787 -10184 4821
rect -10150 4787 -10104 4821
rect -10070 4787 -10024 4821
rect -9990 4787 -9944 4821
rect -9910 4787 -9864 4821
rect -9830 4787 -9784 4821
rect -9750 4787 -9704 4821
rect -9670 4787 -9624 4821
rect -9590 4787 -9544 4821
rect -9510 4787 -9464 4821
rect -9430 4787 -9384 4821
rect -9350 4787 -9304 4821
rect -9270 4787 -9224 4821
rect -9190 4787 -9144 4821
rect -9110 4787 -9064 4821
rect -9030 4787 -8983 4821
rect -8949 4787 -8903 4821
rect -8869 4787 -8823 4821
rect -8789 4787 -8743 4821
rect -8709 4787 -8663 4821
rect -8629 4787 -8583 4821
rect -8549 4787 -8503 4821
rect -8469 4787 -8423 4821
rect -8389 4787 -8343 4821
rect -8309 4787 -8263 4821
rect -8229 4787 -8183 4821
rect -8149 4787 -8103 4821
rect -8069 4787 -8023 4821
rect -7989 4787 -7943 4821
rect -7909 4787 -7863 4821
rect -7829 4787 -7783 4821
rect -7749 4787 -7703 4821
rect -7669 4787 -7623 4821
rect -7589 4787 -7543 4821
rect -7509 4787 -7463 4821
rect -7429 4787 -7383 4821
rect -7349 4787 -7303 4821
rect -7269 4787 -7223 4821
rect -7189 4787 -7143 4821
rect -7109 4787 -7063 4821
rect -7029 4787 -6983 4821
rect -6949 4787 -6903 4821
rect -6869 4787 -6823 4821
rect -6789 4787 -6743 4821
rect -6709 4787 -6663 4821
rect -6629 4787 -6583 4821
rect -6549 4787 -6503 4821
rect -6469 4787 -6423 4821
rect -6389 4787 -6343 4821
rect -6309 4787 -6263 4821
rect -6229 4787 -6183 4821
rect -6149 4787 -6103 4821
rect -6069 4787 -6023 4821
rect -5989 4787 -5943 4821
rect -5909 4787 -5863 4821
rect -5829 4787 -5783 4821
rect -5749 4787 -5703 4821
rect -5669 4787 -5623 4821
rect -5589 4787 -5543 4821
rect -5509 4787 -5463 4821
rect -5429 4787 -5383 4821
rect -5349 4787 -5303 4821
rect -5269 4787 -5223 4821
rect -5189 4787 -5143 4821
rect -5109 4787 -5063 4821
rect -5029 4787 -4983 4821
rect -4949 4787 -4903 4821
rect -4869 4787 -4823 4821
rect -4789 4787 -4743 4821
rect -4709 4787 -4663 4821
rect -4629 4787 -4583 4821
rect -4549 4787 -4503 4821
rect -4469 4787 -4423 4821
rect -4389 4787 -4343 4821
rect -4309 4787 -4263 4821
rect -4229 4787 -4183 4821
rect -4149 4787 -4103 4821
rect -4069 4787 -4023 4821
rect -3989 4787 -3943 4821
rect -3909 4787 -3863 4821
rect -3829 4787 -3783 4821
rect -3749 4787 -3703 4821
rect -3669 4787 -3623 4821
rect -3589 4787 -3543 4821
rect -3509 4787 -3463 4821
rect -3429 4787 -3383 4821
rect -3349 4787 -3303 4821
rect -3269 4787 -3223 4821
rect -3189 4787 -3143 4821
rect -3109 4787 -3063 4821
rect -3029 4787 -2983 4821
rect -2949 4787 -2903 4821
rect -2869 4787 -2823 4821
rect -2789 4787 -2743 4821
rect -2709 4787 -2663 4821
rect -2629 4787 -2583 4821
rect -2549 4787 -2503 4821
rect -2469 4787 -2423 4821
rect -2389 4787 -2343 4821
rect -2309 4787 -2263 4821
rect -2229 4787 -2183 4821
rect -2149 4787 -2103 4821
rect -2069 4787 -2023 4821
rect -1989 4787 -1943 4821
rect -1909 4787 -1863 4821
rect -1829 4787 -1783 4821
rect -1749 4787 -1703 4821
rect -1669 4787 -1623 4821
rect -1589 4787 -1543 4821
rect -1509 4787 -1463 4821
rect -1429 4787 -1383 4821
rect -1349 4787 -1303 4821
rect -1269 4787 -1223 4821
rect -1189 4787 -1143 4821
rect -1109 4787 -1063 4821
rect -1029 4787 -983 4821
rect -949 4787 -903 4821
rect -869 4787 -823 4821
rect -789 4787 -743 4821
rect -709 4787 -663 4821
rect -629 4787 -583 4821
rect -549 4787 -503 4821
rect -469 4787 -423 4821
rect -389 4787 -343 4821
rect -34951 4754 -343 4787
rect 1635 4821 36243 4854
rect 1635 4787 1681 4821
rect 1715 4787 1761 4821
rect 1795 4787 1841 4821
rect 1875 4787 1921 4821
rect 1955 4787 2001 4821
rect 2035 4787 2081 4821
rect 2115 4787 2161 4821
rect 2195 4787 2241 4821
rect 2275 4787 2321 4821
rect 2355 4787 2401 4821
rect 2435 4787 2481 4821
rect 2515 4787 2561 4821
rect 2595 4787 2641 4821
rect 2675 4787 2721 4821
rect 2755 4787 2801 4821
rect 2835 4787 2881 4821
rect 2915 4787 2961 4821
rect 2995 4787 3041 4821
rect 3075 4787 3121 4821
rect 3155 4787 3201 4821
rect 3235 4787 3281 4821
rect 3315 4787 3361 4821
rect 3395 4787 3441 4821
rect 3475 4787 3521 4821
rect 3555 4787 3601 4821
rect 3635 4787 3681 4821
rect 3715 4787 3761 4821
rect 3795 4787 3841 4821
rect 3875 4787 3921 4821
rect 3955 4787 4001 4821
rect 4035 4787 4081 4821
rect 4115 4787 4161 4821
rect 4195 4787 4241 4821
rect 4275 4787 4321 4821
rect 4355 4787 4401 4821
rect 4435 4787 4481 4821
rect 4515 4787 4561 4821
rect 4595 4787 4641 4821
rect 4675 4787 4721 4821
rect 4755 4787 4801 4821
rect 4835 4787 4881 4821
rect 4915 4787 4961 4821
rect 4995 4787 5041 4821
rect 5075 4787 5121 4821
rect 5155 4787 5201 4821
rect 5235 4787 5281 4821
rect 5315 4787 5361 4821
rect 5395 4787 5441 4821
rect 5475 4787 5521 4821
rect 5555 4787 5601 4821
rect 5635 4787 5681 4821
rect 5715 4787 5761 4821
rect 5795 4787 5841 4821
rect 5875 4787 5921 4821
rect 5955 4787 6001 4821
rect 6035 4787 6081 4821
rect 6115 4787 6161 4821
rect 6195 4787 6241 4821
rect 6275 4787 6321 4821
rect 6355 4787 6401 4821
rect 6435 4787 6481 4821
rect 6515 4787 6561 4821
rect 6595 4787 6641 4821
rect 6675 4787 6721 4821
rect 6755 4787 6801 4821
rect 6835 4787 6881 4821
rect 6915 4787 6961 4821
rect 6995 4787 7041 4821
rect 7075 4787 7121 4821
rect 7155 4787 7201 4821
rect 7235 4787 7281 4821
rect 7315 4787 7361 4821
rect 7395 4787 7441 4821
rect 7475 4787 7521 4821
rect 7555 4787 7601 4821
rect 7635 4787 7681 4821
rect 7715 4787 7761 4821
rect 7795 4787 7841 4821
rect 7875 4787 7921 4821
rect 7955 4787 8001 4821
rect 8035 4787 8081 4821
rect 8115 4787 8161 4821
rect 8195 4787 8241 4821
rect 8275 4787 8321 4821
rect 8355 4787 8401 4821
rect 8435 4787 8481 4821
rect 8515 4787 8561 4821
rect 8595 4787 8641 4821
rect 8675 4787 8721 4821
rect 8755 4787 8801 4821
rect 8835 4787 8881 4821
rect 8915 4787 8961 4821
rect 8995 4787 9041 4821
rect 9075 4787 9121 4821
rect 9155 4787 9201 4821
rect 9235 4787 9281 4821
rect 9315 4787 9361 4821
rect 9395 4787 9441 4821
rect 9475 4787 9521 4821
rect 9555 4787 9601 4821
rect 9635 4787 9681 4821
rect 9715 4787 9761 4821
rect 9795 4787 9841 4821
rect 9875 4787 9921 4821
rect 9955 4787 10001 4821
rect 10035 4787 10081 4821
rect 10115 4787 10161 4821
rect 10195 4787 10241 4821
rect 10275 4787 10321 4821
rect 10355 4787 10401 4821
rect 10435 4787 10481 4821
rect 10515 4787 10561 4821
rect 10595 4787 10641 4821
rect 10675 4787 10721 4821
rect 10755 4787 10801 4821
rect 10835 4787 10881 4821
rect 10915 4787 10961 4821
rect 10995 4787 11041 4821
rect 11075 4787 11121 4821
rect 11155 4787 11201 4821
rect 11235 4787 11281 4821
rect 11315 4787 11361 4821
rect 11395 4787 11441 4821
rect 11475 4787 11521 4821
rect 11555 4787 11601 4821
rect 11635 4787 11681 4821
rect 11715 4787 11761 4821
rect 11795 4787 11841 4821
rect 11875 4787 11921 4821
rect 11955 4787 12001 4821
rect 12035 4787 12081 4821
rect 12115 4787 12161 4821
rect 12195 4787 12241 4821
rect 12275 4787 12321 4821
rect 12355 4787 12401 4821
rect 12435 4787 12481 4821
rect 12515 4787 12561 4821
rect 12595 4787 12641 4821
rect 12675 4787 12721 4821
rect 12755 4787 12801 4821
rect 12835 4787 12881 4821
rect 12915 4787 12961 4821
rect 12995 4787 13041 4821
rect 13075 4787 13121 4821
rect 13155 4787 13201 4821
rect 13235 4787 13281 4821
rect 13315 4787 13361 4821
rect 13395 4787 13441 4821
rect 13475 4787 13521 4821
rect 13555 4787 13601 4821
rect 13635 4787 13681 4821
rect 13715 4787 13761 4821
rect 13795 4787 13841 4821
rect 13875 4787 13921 4821
rect 13955 4787 14001 4821
rect 14035 4787 14081 4821
rect 14115 4787 14161 4821
rect 14195 4787 14241 4821
rect 14275 4787 14321 4821
rect 14355 4787 14401 4821
rect 14435 4787 14481 4821
rect 14515 4787 14561 4821
rect 14595 4787 14642 4821
rect 14676 4787 14722 4821
rect 14756 4787 14802 4821
rect 14836 4787 14882 4821
rect 14916 4787 14962 4821
rect 14996 4787 15042 4821
rect 15076 4787 15122 4821
rect 15156 4787 15202 4821
rect 15236 4787 15282 4821
rect 15316 4787 15362 4821
rect 15396 4787 15442 4821
rect 15476 4787 15522 4821
rect 15556 4787 15602 4821
rect 15636 4787 15682 4821
rect 15716 4787 15762 4821
rect 15796 4787 15842 4821
rect 15876 4787 15922 4821
rect 15956 4787 16002 4821
rect 16036 4787 16082 4821
rect 16116 4787 16162 4821
rect 16196 4787 16242 4821
rect 16276 4787 16322 4821
rect 16356 4787 16402 4821
rect 16436 4787 16482 4821
rect 16516 4787 16562 4821
rect 16596 4787 16642 4821
rect 16676 4787 16722 4821
rect 16756 4787 16802 4821
rect 16836 4787 16882 4821
rect 16916 4787 16962 4821
rect 16996 4787 17042 4821
rect 17076 4787 17122 4821
rect 17156 4787 17202 4821
rect 17236 4787 17282 4821
rect 17316 4787 17362 4821
rect 17396 4787 17442 4821
rect 17476 4787 17522 4821
rect 17556 4787 17602 4821
rect 17636 4787 17682 4821
rect 17716 4787 17762 4821
rect 17796 4787 17842 4821
rect 17876 4787 17922 4821
rect 17956 4787 18002 4821
rect 18036 4787 18082 4821
rect 18116 4787 18162 4821
rect 18196 4787 18242 4821
rect 18276 4787 18322 4821
rect 18356 4787 18402 4821
rect 18436 4787 18482 4821
rect 18516 4787 18562 4821
rect 18596 4787 18642 4821
rect 18676 4787 18722 4821
rect 18756 4787 18802 4821
rect 18836 4787 18882 4821
rect 18916 4787 18962 4821
rect 18996 4787 19042 4821
rect 19076 4787 19122 4821
rect 19156 4787 19202 4821
rect 19236 4787 19282 4821
rect 19316 4787 19362 4821
rect 19396 4787 19442 4821
rect 19476 4787 19522 4821
rect 19556 4787 19602 4821
rect 19636 4787 19682 4821
rect 19716 4787 19762 4821
rect 19796 4787 19842 4821
rect 19876 4787 19922 4821
rect 19956 4787 20002 4821
rect 20036 4787 20082 4821
rect 20116 4787 20162 4821
rect 20196 4787 20242 4821
rect 20276 4787 20322 4821
rect 20356 4787 20402 4821
rect 20436 4787 20482 4821
rect 20516 4787 20562 4821
rect 20596 4787 20642 4821
rect 20676 4787 20722 4821
rect 20756 4787 20802 4821
rect 20836 4787 20882 4821
rect 20916 4787 20962 4821
rect 20996 4787 21042 4821
rect 21076 4787 21122 4821
rect 21156 4787 21202 4821
rect 21236 4787 21282 4821
rect 21316 4787 21362 4821
rect 21396 4787 21442 4821
rect 21476 4787 21522 4821
rect 21556 4787 21602 4821
rect 21636 4787 21682 4821
rect 21716 4787 21762 4821
rect 21796 4787 21842 4821
rect 21876 4787 21922 4821
rect 21956 4787 22002 4821
rect 22036 4787 22082 4821
rect 22116 4787 22162 4821
rect 22196 4787 22242 4821
rect 22276 4787 22322 4821
rect 22356 4787 22402 4821
rect 22436 4787 22482 4821
rect 22516 4787 22562 4821
rect 22596 4787 22642 4821
rect 22676 4787 22722 4821
rect 22756 4787 22802 4821
rect 22836 4787 22882 4821
rect 22916 4787 22962 4821
rect 22996 4787 23042 4821
rect 23076 4787 23122 4821
rect 23156 4787 23202 4821
rect 23236 4787 23282 4821
rect 23316 4787 23362 4821
rect 23396 4787 23442 4821
rect 23476 4787 23522 4821
rect 23556 4787 23602 4821
rect 23636 4787 23682 4821
rect 23716 4787 23762 4821
rect 23796 4787 23842 4821
rect 23876 4787 23922 4821
rect 23956 4787 24002 4821
rect 24036 4787 24082 4821
rect 24116 4787 24162 4821
rect 24196 4787 24242 4821
rect 24276 4787 24322 4821
rect 24356 4787 24402 4821
rect 24436 4787 24482 4821
rect 24516 4787 24562 4821
rect 24596 4787 24642 4821
rect 24676 4787 24722 4821
rect 24756 4787 24802 4821
rect 24836 4787 24882 4821
rect 24916 4787 24962 4821
rect 24996 4787 25042 4821
rect 25076 4787 25122 4821
rect 25156 4787 25202 4821
rect 25236 4787 25282 4821
rect 25316 4787 25362 4821
rect 25396 4787 25442 4821
rect 25476 4787 25522 4821
rect 25556 4787 25602 4821
rect 25636 4787 25682 4821
rect 25716 4787 25762 4821
rect 25796 4787 25842 4821
rect 25876 4787 25922 4821
rect 25956 4787 26002 4821
rect 26036 4787 26082 4821
rect 26116 4787 26162 4821
rect 26196 4787 26242 4821
rect 26276 4787 26322 4821
rect 26356 4787 26402 4821
rect 26436 4787 26482 4821
rect 26516 4787 26562 4821
rect 26596 4787 26642 4821
rect 26676 4787 26722 4821
rect 26756 4787 26802 4821
rect 26836 4787 26882 4821
rect 26916 4787 26962 4821
rect 26996 4787 27042 4821
rect 27076 4787 27122 4821
rect 27156 4787 27202 4821
rect 27236 4787 27282 4821
rect 27316 4787 27362 4821
rect 27396 4787 27442 4821
rect 27476 4787 27522 4821
rect 27556 4787 27603 4821
rect 27637 4787 27683 4821
rect 27717 4787 27763 4821
rect 27797 4787 27843 4821
rect 27877 4787 27923 4821
rect 27957 4787 28003 4821
rect 28037 4787 28083 4821
rect 28117 4787 28163 4821
rect 28197 4787 28243 4821
rect 28277 4787 28323 4821
rect 28357 4787 28403 4821
rect 28437 4787 28483 4821
rect 28517 4787 28563 4821
rect 28597 4787 28643 4821
rect 28677 4787 28723 4821
rect 28757 4787 28803 4821
rect 28837 4787 28883 4821
rect 28917 4787 28963 4821
rect 28997 4787 29043 4821
rect 29077 4787 29123 4821
rect 29157 4787 29203 4821
rect 29237 4787 29283 4821
rect 29317 4787 29363 4821
rect 29397 4787 29443 4821
rect 29477 4787 29523 4821
rect 29557 4787 29603 4821
rect 29637 4787 29683 4821
rect 29717 4787 29763 4821
rect 29797 4787 29843 4821
rect 29877 4787 29923 4821
rect 29957 4787 30003 4821
rect 30037 4787 30083 4821
rect 30117 4787 30163 4821
rect 30197 4787 30243 4821
rect 30277 4787 30323 4821
rect 30357 4787 30403 4821
rect 30437 4787 30483 4821
rect 30517 4787 30563 4821
rect 30597 4787 30643 4821
rect 30677 4787 30723 4821
rect 30757 4787 30803 4821
rect 30837 4787 30883 4821
rect 30917 4787 30963 4821
rect 30997 4787 31043 4821
rect 31077 4787 31123 4821
rect 31157 4787 31203 4821
rect 31237 4787 31283 4821
rect 31317 4787 31363 4821
rect 31397 4787 31443 4821
rect 31477 4787 31523 4821
rect 31557 4787 31603 4821
rect 31637 4787 31683 4821
rect 31717 4787 31763 4821
rect 31797 4787 31843 4821
rect 31877 4787 31923 4821
rect 31957 4787 32003 4821
rect 32037 4787 32083 4821
rect 32117 4787 32163 4821
rect 32197 4787 32243 4821
rect 32277 4787 32323 4821
rect 32357 4787 32403 4821
rect 32437 4787 32483 4821
rect 32517 4787 32563 4821
rect 32597 4787 32643 4821
rect 32677 4787 32723 4821
rect 32757 4787 32803 4821
rect 32837 4787 32883 4821
rect 32917 4787 32963 4821
rect 32997 4787 33043 4821
rect 33077 4787 33123 4821
rect 33157 4787 33203 4821
rect 33237 4787 33283 4821
rect 33317 4787 33363 4821
rect 33397 4787 33443 4821
rect 33477 4787 33523 4821
rect 33557 4787 33603 4821
rect 33637 4787 33683 4821
rect 33717 4787 33763 4821
rect 33797 4787 33843 4821
rect 33877 4787 33923 4821
rect 33957 4787 34003 4821
rect 34037 4787 34083 4821
rect 34117 4787 34163 4821
rect 34197 4787 34243 4821
rect 34277 4787 34323 4821
rect 34357 4787 34403 4821
rect 34437 4787 34483 4821
rect 34517 4787 34563 4821
rect 34597 4787 34643 4821
rect 34677 4787 34723 4821
rect 34757 4787 34803 4821
rect 34837 4787 34883 4821
rect 34917 4787 34963 4821
rect 34997 4787 35043 4821
rect 35077 4787 35123 4821
rect 35157 4787 35203 4821
rect 35237 4787 35283 4821
rect 35317 4787 35363 4821
rect 35397 4787 35443 4821
rect 35477 4787 35523 4821
rect 35557 4787 35603 4821
rect 35637 4787 35683 4821
rect 35717 4787 35763 4821
rect 35797 4787 35843 4821
rect 35877 4787 35923 4821
rect 35957 4787 36003 4821
rect 36037 4787 36083 4821
rect 36117 4787 36163 4821
rect 36197 4787 36243 4821
rect 1635 4754 36243 4787
<< metal2 >>
rect -1505 8709 38335 8743
rect 4101 8601 38333 8635
rect -25 5631 1341 5891
rect 1601 5631 1694 5891
rect 1614 4700 1694 5631
<< metal3 >>
rect -285 5891 -25 6493
rect 1341 5891 1601 6493
<< metal4 >>
rect -20677 11271 -20455 11471
rect -20677 10191 -20477 11271
rect 3394 11270 18881 11470
rect -20677 9991 -1983 10191
rect -2183 8362 -1983 9991
rect 3394 8362 3594 11270
<< via4 >>
rect -3848 7838 -3612 8074
rect -3848 6600 -3612 6836
rect -276 6505 -40 6741
rect 1350 6505 1586 6741
rect -273 5643 -37 5879
rect 1353 5643 1589 5879
<< metal5 >>
rect -3941 8074 -3520 8166
rect -3941 7838 -3848 8074
rect -3612 7838 -3520 8074
rect -3941 7746 -3520 7838
rect -3941 6836 -3520 6928
rect -3941 6600 -3848 6836
rect -3612 6600 -3520 6836
rect -3941 6508 -3520 6600
rect -369 6741 52 6833
rect -369 6505 -276 6741
rect -40 6505 52 6741
rect -369 6413 52 6505
rect 1257 6741 1678 6833
rect 1257 6505 1350 6741
rect 1586 6505 1678 6741
rect 1257 6413 1678 6505
rect -366 5879 55 5971
rect -366 5643 -273 5879
rect -37 5643 55 5879
rect -366 5551 55 5643
rect 1260 5879 1681 5971
rect 1260 5643 1353 5879
rect 1589 5643 1681 5879
rect 1260 5551 1681 5643
<< glass >>
rect -3940 7746 -3520 8166
rect -3940 6508 -3520 6928
rect -368 6413 52 6833
rect 1258 6413 1678 6833
rect -365 5551 55 5971
rect 1261 5551 1681 5971
use CASCODED_nmos_1v8_lvt_4p5_10finger  CASCODED_nmos_1v8_lvt_4p5_10finger_0
timestamp 1670967604
transform -1 0 824 0 1 6615
box -3590 209 -298 1270
use CASCODED_nmos_1v8_lvt_4p5_10finger  CASCODED_nmos_1v8_lvt_4p5_10finger_1
timestamp 1670967604
transform 1 0 486 0 1 6615
box -3590 209 -298 1270
use Li_via_M2  Li_via_M2_0
timestamp 1670967604
transform 1 0 4041 0 1 8598
box -20 -20 60 60
use Li_via_M2  Li_via_M2_1
timestamp 1670967604
transform 1 0 -1565 0 1 8706
box -20 -20 60 60
use Li_via_M2  Li_via_M2_2
timestamp 1670967604
transform 1 0 1634 0 1 4640
box -20 -20 60 60
use M1_vias_M4  M1_vias_M4_0
timestamp 1670967604
transform 1 0 -3380 0 1 7996
box -480 -170 -220 90
use M1_vias_M4  M1_vias_M4_1
timestamp 1670967604
transform 1 0 -3380 0 1 6758
box -480 -170 -220 90
use M1_vias_M4  M1_vias_M4_2
timestamp 1670967604
transform 1 0 1821 0 1 5801
box -480 -170 -220 90
use M1_vias_M4  M1_vias_M4_3
timestamp 1670967604
transform 1 0 195 0 1 5801
box -480 -170 -220 90
use M1_vias_M4  M1_vias_M4_4
timestamp 1670967604
transform 1 0 1818 0 1 6663
box -480 -170 -220 90
use M1_vias_M4  M1_vias_M4_5
timestamp 1670967604
transform 1 0 192 0 1 6663
box -480 -170 -220 90
use M1_vias_M4  M1_vias_M4_6
timestamp 1670967604
transform 1 0 -1738 0 1 8272
box -480 -170 -220 90
use M1_vias_M4  M1_vias_M4_7
timestamp 1670967604
transform 1 0 3843 0 1 8272
box -480 -170 -220 90
use M1_vias_M4  M1_vias_M4_8
timestamp 1670967604
transform 1 0 19101 0 1 17039
box -480 -170 -220 90
use M1_vias_M4  M1_vias_M4_9
timestamp 1670967604
transform 1 0 -20234 0 1 17040
box -480 -170 -220 90
use Resistor_20k  Resistor_20k_0
timestamp 1670967604
transform 1 0 3134 0 1 7413
box 1122 690 2146 1692
use Resistor_20k  Resistor_20k_1
timestamp 1670967604
transform 1 0 -2411 0 1 7414
box 1122 690 2146 1692
use Square_Inductor_10t_2s_1w_180dout  Square_Inductor_10t_2s_1w_180dout_0
timestamp 1670967604
transform 1 0 6541 0 1 16650
box -5060 -5380 30140 29820
use Square_Inductor_10t_2s_1w_180dout  Square_Inductor_10t_2s_1w_180dout_1
timestamp 1670967604
transform 1 0 -32795 0 1 16651
box -5060 -5380 30140 29820
use Vdd_power_rail  Vdd_power_rail_0
timestamp 1670967604
transform 1 0 4027 0 1 15970
box -1630 1160 -250 1260
use Vdd_power_rail  Vdd_power_rail_1
timestamp 1670967604
transform 1 0 -1692 0 1 15970
box -1630 1160 -250 1260
use Vdd_power_rail  Vdd_power_rail_2
timestamp 1670967604
transform 1 0 4027 0 1 8111
box -1630 1160 -250 1260
use Vdd_power_rail  Vdd_power_rail_3
timestamp 1670967604
transform 1 0 -1692 0 1 8111
box -1630 1160 -250 1260
use Vdd_power_rail  Vdd_power_rail_4
timestamp 1670967604
transform 1 0 4027 0 1 8111
box -1630 1160 -250 1260
use Vdd_power_rail  Vdd_power_rail_5
timestamp 1670967604
transform 1 0 -1692 0 1 8111
box -1630 1160 -250 1260
use Via_P_Licon_Li  Via_P_Licon_Li_0
timestamp 1670967604
transform 1 0 882 0 1 6813
box 368 1104 434 1170
use Via_P_Licon_Li  Via_P_Licon_Li_1
timestamp 1670967604
transform 1 0 -1724 0 1 5583
box 368 1104 434 1170
use Via_P_Licon_Li  Via_P_Licon_Li_2
timestamp 1670967604
transform 1 0 -3218 0 1 6800
box 368 1104 434 1170
use Via_P_Licon_Li  Via_P_Licon_Li_3
timestamp 1670967604
transform 1 0 2388 0 1 6800
box 368 1104 434 1170
use simple_current_mirror  simple_current_mirror_0
timestamp 1670967989
transform 1 0 -105 0 1 3560
box -299 -197 1778 1294
<< labels >>
flabel metal1 s -3460 7929 -3409 7972 2 FreeSans 100000 0 0 0 IN1
port 1 nsew
flabel metal1 s -3460 6699 -3419 6738 2 FreeSans 100000 0 0 0 IN2
port 2 nsew
flabel metal1 s 551 6326 665 6360 2 FreeSans 100000 0 0 0 Ground
port 3 nsew
flabel metal1 s 471 9304 1145 9338 2 FreeSans 100000 0 0 0 VDD
port 4 nsew
flabel metal1 s -570 17162 104 17196 2 FreeSans 100000 0 0 0 VDD
port 4 nsew
flabel metal2 s 5489 8714 5514 8737 2 FreeSans 100000 0 0 0 OUT1
port 5 nsew
flabel metal2 s 5490 8607 5517 8627 2 FreeSans 100000 0 0 0 OUT2
port 6 nsew
<< properties >>
string path 7.355 30.225 7.355 32.465 
<< end >>
