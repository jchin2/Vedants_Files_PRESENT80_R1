magic
tech sky130A
timestamp 1662731941
<< nwell >>
rect -75 130 160 500
<< nmos >>
rect 65 -55 80 95
<< pmos >>
rect 65 165 80 465
<< ndiff >>
rect 5 80 65 95
rect 5 50 20 80
rect 50 50 65 80
rect 5 -10 65 50
rect 5 -40 20 -10
rect 50 -40 65 -10
rect 5 -55 65 -40
rect 80 80 140 95
rect 80 50 95 80
rect 125 50 140 80
rect 80 -10 140 50
rect 80 -40 95 -10
rect 125 -40 140 -10
rect 80 -55 140 -40
<< pdiff >>
rect 5 450 65 465
rect 5 420 20 450
rect 50 420 65 450
rect 5 360 65 420
rect 5 330 20 360
rect 50 330 65 360
rect 5 300 65 330
rect 5 270 20 300
rect 50 270 65 300
rect 5 210 65 270
rect 5 180 20 210
rect 50 180 65 210
rect 5 165 65 180
rect 80 450 140 465
rect 80 420 95 450
rect 125 420 140 450
rect 80 360 140 420
rect 80 330 95 360
rect 125 330 140 360
rect 80 300 140 330
rect 80 270 95 300
rect 125 270 140 300
rect 80 210 140 270
rect 80 180 95 210
rect 125 180 140 210
rect 80 165 140 180
<< ndiffc >>
rect 20 50 50 80
rect 20 -40 50 -10
rect 95 50 125 80
rect 95 -40 125 -10
<< pdiffc >>
rect 20 420 50 450
rect 20 330 50 360
rect 20 270 50 300
rect 20 180 50 210
rect 95 420 125 450
rect 95 330 125 360
rect 95 270 125 300
rect 95 180 125 210
<< psubdiff >>
rect -55 80 5 95
rect -55 50 -40 80
rect -10 50 5 80
rect -55 -10 5 50
rect -55 -40 -40 -10
rect -10 -40 5 -10
rect -55 -55 5 -40
<< nsubdiff >>
rect -55 450 5 465
rect -55 420 -40 450
rect -10 420 5 450
rect -55 360 5 420
rect -55 330 -40 360
rect -10 330 5 360
rect -55 300 5 330
rect -55 270 -40 300
rect -10 270 5 300
rect -55 210 5 270
rect -55 180 -40 210
rect -10 180 5 210
rect -55 165 5 180
<< psubdiffcont >>
rect -40 50 -10 80
rect -40 -40 -10 -10
<< nsubdiffcont >>
rect -40 420 -10 450
rect -40 330 -10 360
rect -40 270 -10 300
rect -40 180 -10 210
<< poly >>
rect 65 465 80 480
rect 65 150 80 165
rect 25 140 80 150
rect 25 120 35 140
rect 55 120 80 140
rect 25 110 80 120
rect 65 95 80 110
rect 65 -70 80 -55
<< polycont >>
rect 35 120 55 140
<< locali >>
rect -75 515 160 525
rect -75 495 -65 515
rect -45 495 -25 515
rect -5 495 15 515
rect 35 495 55 515
rect 75 495 95 515
rect 115 495 135 515
rect 155 495 160 515
rect -75 485 160 495
rect -50 460 5 485
rect -50 450 60 460
rect -50 420 -40 450
rect -10 420 20 450
rect 50 420 60 450
rect -50 360 60 420
rect -50 330 -40 360
rect -10 330 20 360
rect 50 330 60 360
rect -50 300 60 330
rect -50 270 -40 300
rect -10 270 20 300
rect 50 270 60 300
rect -50 210 60 270
rect -50 180 -40 210
rect -10 180 20 210
rect 50 180 60 210
rect -50 170 60 180
rect 85 450 135 460
rect 85 420 95 450
rect 125 420 135 450
rect 85 360 135 420
rect 85 330 95 360
rect 125 330 135 360
rect 85 300 135 330
rect 85 270 95 300
rect 125 270 135 300
rect 85 210 135 270
rect 85 180 95 210
rect 125 180 135 210
rect 85 170 135 180
rect 25 140 65 150
rect -75 120 35 140
rect 55 120 65 140
rect 25 110 65 120
rect 110 140 135 170
rect 110 120 160 140
rect 110 90 135 120
rect -50 80 60 90
rect -50 50 -40 80
rect -10 50 20 80
rect 50 50 60 80
rect -50 -10 60 50
rect -50 -40 -40 -10
rect -10 -40 20 -10
rect 50 -40 60 -10
rect -50 -50 60 -40
rect 85 80 135 90
rect 85 50 95 80
rect 125 50 135 80
rect 85 -10 135 50
rect 85 -40 95 -10
rect 125 -40 135 -10
rect 85 -50 135 -40
rect -50 -75 5 -50
rect -75 -85 160 -75
rect -75 -105 -65 -85
rect -45 -105 -25 -85
rect -5 -105 15 -85
rect 35 -105 55 -85
rect 75 -105 95 -85
rect 115 -105 135 -85
rect 155 -105 160 -85
rect -75 -115 160 -105
<< viali >>
rect -65 495 -45 515
rect -25 495 -5 515
rect 15 495 35 515
rect 55 495 75 515
rect 95 495 115 515
rect 135 495 155 515
rect -65 -105 -45 -85
rect -25 -105 -5 -85
rect 15 -105 35 -85
rect 55 -105 75 -85
rect 95 -105 115 -85
rect 135 -105 155 -85
<< metal1 >>
rect -75 515 160 545
rect -75 495 -65 515
rect -45 495 -25 515
rect -5 495 15 515
rect 35 495 55 515
rect 75 495 95 515
rect 115 495 135 515
rect 155 495 160 515
rect -75 465 160 495
rect -75 -85 160 -55
rect -75 -105 -65 -85
rect -45 -105 -25 -85
rect -5 -105 15 -85
rect 35 -105 55 -85
rect 75 -105 95 -85
rect 115 -105 135 -85
rect 155 -105 160 -85
rect -75 -135 160 -105
<< labels >>
rlabel metal1 -65 495 -45 515 7 A
port 1 w
rlabel locali -75 120 -55 140 7 B
port 2 w
rlabel metal1 -65 -105 -45 -85 7 D
port 4 w
rlabel locali 140 120 160 140 7 C
port 3 w
<< end >>
