* NGSPICE file created from CMOS_PRESENT80_R1_flat.ext - technology: sky130A

.subckt CMOS_PRESENT80_R1_flat GND k0 k0_bar x0 x0_bar x1_bar x1 k1_bar k1 k2 k2_bar
+ x2 x2_bar x3_bar x3 k3_bar k3 s3 s2 s1 s0 VDD
X0 a_n2290_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t4 GND.t160 GND.t159 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n787_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t2 GND.t39 GND.t38 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n732_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t4 GND.t101 GND.t100 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X3 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR a_n2140_n2118# GND.t25 GND.t24 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n4395_n1508# x2_bar.t0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t3 VDD.t23 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X5 a_275_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t2 a_575_n3696# VDD.t57 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X6 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A a_425_1648# GND.t125 GND.t1 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n2290_370# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t4 GND.t80 GND.t79 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_425_n1508# VDD.t143 VDD.t4 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X9 a_n432_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t3 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A GND.t67 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X10 GND.t41 x0_bar.t0 a_n4395_1038# GND.t40 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X11 a_n732_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t2 VDD.t169 VDD.t168 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X12 a_n4395_1038# k0_bar.t0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t2 GND.t59 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t5 a_n732_n2118# GND.t137 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X14 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t1 x1.t0 a_n4695_n540# VDD.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X15 GND.t77 x2_bar.t1 a_n4395_n2118# GND.t76 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X16 a_n4695_n540# k1_bar.t0 VDD.t68 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X17 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND a_n787_n10008# GND.t123 GND.t122 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X18 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t0 a_n2345_n6852# VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X19 s2.t1 a_275_n5942# GND.t115 GND.t114 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X20 a_n4395_370# k1_bar.t1 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t2 GND.t59 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X21 a_n2140_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t4 a_n2290_n7820# VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X22 a_n4395_n2118# k2_bar.t0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t1 GND.t46 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X23 a_425_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t2 VDD.t46 VDD.t8 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X24 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_425_n1508# GND.t140 GND.t139 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X25 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t2 k3.t0 a_n4695_n2786# GND.t65 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X26 VDD.t39 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t3 a_n2495_n3696# VDD.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X27 a_n2290_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t4 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X28 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t1 a_n2495_n10008# GND.t64 GND.t63 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X29 a_n732_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t5 GND.t88 GND.t87 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X30 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t5 a_n2290_1648# VDD.t182 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X31 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n2140_n8430# VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X32 a_n2290_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t4 VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X33 VDD.t170 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A a_425_n1508# VDD.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X34 a_n4695_n2786# x3.t0 GND.t147 GND.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X35 a_n787_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t3 a_n787_1648# VDD.t69 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X36 VDD.t71 k3.t1 a_n4395_n3696# VDD.t70 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X37 a_n787_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t6 VDD.t167 VDD.t166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X38 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t1 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t6 GND.t136 GND.t135 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X39 a_275_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t2 a_575_n6852# VDD.t20 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X40 a_n1990_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t5 a_n2140_n2118# VDD.t101 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X41 a_n432_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t4 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A VDD.t58 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X42 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR a_n787_1038# GND.t99 GND.t98 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X43 a_n2140_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t6 a_n2290_n8430# GND.t158 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X44 a_n2345_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t5 a_n2045_n5942# GND.t42 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X45 a_425_n540# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A a_425_370# GND.t81 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X46 a_n4695_370# x1.t1 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X47 a_425_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t5 GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X48 a_n4395_n3696# x3_bar.t0 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t0 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X49 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t5 a_n732_n7820# VDD.t154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X50 a_n2290_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t7 GND.t34 GND.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X51 s3.t1 a_275_n9098# GND.t97 GND.t96 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X52 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n2140_n8430# GND.t111 GND.t110 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X53 a_n1990_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t6 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A GND.t0 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X54 a_n2140_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t7 a_n2290_n540# VDD.t142 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X55 a_425_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A a_425_n2118# GND.t22 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X56 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B a_425_n540# GND.t2 GND.t1 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X57 VDD.t141 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t8 a_n432_n1508# VDD.t140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X58 a_575_n10008# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND a_425_n10008# VDD.t54 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X59 a_n2290_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t6 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X60 VDD.t153 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t6 a_n1990_n1508# VDD.t152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X61 GND.t30 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t3 a_275_n2786# GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X62 a_n2140_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t9 a_n2290_n4664# VDD.t139 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X63 s0.t0 a_1637_1038# VDD.t66 VDD.t65 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X64 VDD.t151 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t7 a_n787_n540# VDD.t150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X65 a_n1990_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t6 a_n2140_n2118# GND.t148 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X66 a_n432_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t7 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A GND.t89 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X67 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND a_425_n7820# VDD.t64 VDD.t63 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X68 a_n2345_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t8 VDD.t149 VDD.t148 sky130_fd_pr__pfet_01v8 ad=3.6e+12p pd=1.44e+07u as=0p ps=0u w=3e+06u l=150000u
X69 a_n787_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t2 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X70 a_n2495_n10008# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t7 VDD.t181 VDD.t180 sky130_fd_pr__pfet_01v8 ad=3.6e+12p pd=1.44e+07u as=0p ps=0u w=3e+06u l=150000u
X71 a_n2290_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t7 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X72 a_425_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X73 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t10 a_n732_n8430# GND.t134 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X74 a_n787_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t3 GND.t120 GND.t6 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X75 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t1 a_n2345_n6852# GND.t48 GND.t47 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X76 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n2140_n5274# VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X77 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t3 k0.t0 a_n4695_1038# GND.t138 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X78 a_n432_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t4 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A VDD.t42 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X79 a_n4695_1038# x0.t0 GND.t43 GND.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X80 GND.t106 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t5 a_n432_n2118# GND.t105 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X81 a_575_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_425_n3696# VDD.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X82 a_425_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X83 a_1637_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A VDD.t118 VDD.t117 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X84 GND.t15 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t7 a_n1990_n2118# GND.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X85 a_n2140_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t9 a_n2290_n5274# GND.t104 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X86 VDD.t60 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_425_1648# VDD.t59 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X87 a_n2140_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t8 a_n2290_370# GND.t131 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X88 a_n2345_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t8 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X89 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND a_425_n7820# GND.t84 GND.t83 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X90 a_425_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t8 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X91 a_n787_n10008# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t8 VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X92 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t9 a_n732_n4664# VDD.t156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X93 a_n2290_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t11 GND.t133 GND.t132 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X94 VDD.t81 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_425_n7820# VDD.t80 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X95 VDD.t110 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t9 a_n2495_n3696# VDD.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X96 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n2140_n5274# GND.t62 GND.t61 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X97 GND.t163 x3_bar.t1 a_n4395_n2786# GND.t76 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X98 GND.t91 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t3 a_275_n5942# GND.t90 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X99 a_n1990_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t6 a_n2140_n8430# VDD.t21 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X100 GND.t51 x1_bar.t0 a_n4395_370# GND.t40 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X101 a_n432_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t9 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A GND.t149 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X102 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_425_n4664# VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X103 a_n4395_n2786# k3_bar.t0 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t3 GND.t46 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X104 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t10 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X105 a_425_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t11 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X106 a_425_n540# CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X107 VDD.t122 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR a_n787_n3696# VDD.t121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X108 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t0 a_n2495_n10008# VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X109 a_425_n6852# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND VDD.t163 VDD.t162 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X110 VDD.t75 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A a_425_n540# VDD.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X111 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t9 a_n732_n5274# GND.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X112 a_425_n7820# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_425_n8430# GND.t68 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X113 a_n787_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t12 VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X114 a_575_n6852# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_425_n6852# VDD.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X115 VDD.t136 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t13 a_n432_n7820# VDD.t135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X116 a_n1990_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t10 a_n2140_n8430# GND.t66 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X117 VDD.t179 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t10 a_n1990_n7820# VDD.t178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X118 a_n2345_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t10 GND.t45 GND.t44 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X119 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t14 a_n2290_1038# GND.t131 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X120 GND.t36 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t10 a_n1990_370# GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X121 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_425_n4664# GND.t55 GND.t54 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X122 a_n2290_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t11 GND.t156 GND.t79 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X123 a_425_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t8 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X124 GND.t13 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t9 a_n787_1038# GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X125 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t3 k1.t0 a_n4695_370# GND.t138 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X126 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n2140_n540# GND.t73 GND.t72 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X127 a_425_370# CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X128 a_n787_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t12 GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X129 GND.t82 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND a_275_n2786# GND.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X130 VDD.t134 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t15 a_n1990_1648# VDD.t133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X131 GND.t95 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t2 a_275_n9098# GND.t94 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X132 a_n2345_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t13 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X133 VDD.t79 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A a_425_n4664# VDD.t78 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X134 a_275_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X135 a_n1990_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t11 a_n2140_n5274# VDD.t108 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X136 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A a_n787_n540# GND.t128 GND.t98 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X137 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND a_n787_n3696# VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X138 GND.t58 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t10 a_n432_n8430# GND.t57 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X139 VDD.t177 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t12 a_n2345_n6852# VDD.t176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X140 GND.t93 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t7 a_n1990_n8430# GND.t92 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X141 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t13 VDD.t175 VDD.t174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X142 VDD.t48 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n787_n6852# VDD.t47 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X143 a_425_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t11 GND.t162 GND.t143 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X144 a_1637_1038# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B a_1637_1648# VDD.t55 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X145 s0.t1 a_1637_1038# GND.t86 GND.t85 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X146 a_n787_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t11 a_n787_370# GND.t12 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X147 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t12 a_n2195_n2786# GND.t78 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X148 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t0 a_n2495_n3696# VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X149 a_n787_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t8 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X150 a_425_n4664# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A a_425_n5274# GND.t52 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X151 VDD.t173 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t14 a_n1990_n540# VDD.t152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X152 a_n2345_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t16 GND.t130 GND.t129 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X153 VDD.t172 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t15 a_n432_n4664# VDD.t171 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X154 VDD.t147 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t12 a_n1990_n4664# VDD.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X155 a_n1990_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t12 a_n2140_n5274# GND.t56 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X156 a_n2195_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t14 a_n2345_n2786# GND.t121 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X157 a_n732_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t13 VDD.t107 VDD.t106 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X158 a_n787_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR a_n787_n2786# GND.t124 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X159 GND.t144 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND a_275_n5942# GND.t143 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X160 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A a_425_1648# VDD.t124 VDD.t123 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X161 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t1 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t15 GND.t146 GND.t145 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X162 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t0 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t16 VDD.t165 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X163 a_425_1038# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR GND.t117 GND.t4 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X164 a_1637_1038# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A GND.t119 GND.t118 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X165 VDD.t158 k0.t1 a_n4395_1648# VDD.t157 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X166 a_275_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND GND.t53 GND.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X167 a_n4395_1648# x0_bar.t1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t1 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X168 a_425_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_425_1038# GND.t81 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X169 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t0 x2.t0 a_n4695_n1508# VDD.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X170 a_n787_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t17 GND.t75 GND.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X171 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND a_n787_n6852# VDD.t161 VDD.t160 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X172 s1.t0 a_275_n2786# VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X173 GND.t50 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t9 a_n432_n5274# GND.t49 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X174 GND.t11 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t14 a_n1990_n5274# GND.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X175 a_n4695_n1508# k2_bar.t1 VDD.t164 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X176 a_n732_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t17 GND.t32 GND.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X177 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t13 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X178 a_275_n9098# CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t3 a_575_n10008# VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X179 a_n2045_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t18 a_n2195_n5942# GND.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X180 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B a_425_n540# VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X181 VDD.t36 k1.t1 a_n4395_n540# VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X182 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t2 k2.t0 a_n4695_n2118# GND.t65 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X183 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND a_n787_n3696# GND.t109 GND.t108 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X184 a_n2195_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t16 a_n2345_n5942# GND.t155 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X185 VDD.t132 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t18 a_n2495_n10008# VDD.t131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X186 a_n4395_n540# x1_bar.t1 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t0 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X187 GND.t116 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND a_275_n9098# GND.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X188 a_n787_n6852# CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n787_n5942# GND.t60 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X189 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR a_n787_1038# VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X190 a_n4695_n2118# x2.t1 GND.t19 GND.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X191 a_425_n10008# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND VDD.t100 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X192 a_275_n9098# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND GND.t69 GND.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X193 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t14 GND.t113 GND.t112 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X194 a_n787_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t10 GND.t151 GND.t150 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X195 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t1 a_n2495_n3696# GND.t103 GND.t102 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X196 s2.t0 a_275_n5942# VDD.t98 VDD.t97 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X197 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n2140_n540# VDD.t56 VDD.t18 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X198 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t17 a_n2290_n1508# VDD.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X199 VDD.t27 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t13 a_n2495_n10008# VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X200 a_n1990_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t11 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A VDD.t159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X201 GND.t107 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t12 a_n1990_1038# GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X202 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t1 x3.t1 a_n4695_n3696# VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X203 a_n2290_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t14 VDD.t51 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X204 a_n2495_n10008# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t15 a_n2195_n9098# GND.t26 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X205 a_n732_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t15 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X206 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR a_n2140_n2118# VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X207 a_n1990_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t13 a_n2140_n540# GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X208 a_n4695_n3696# k3_bar.t1 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X209 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A a_n787_n540# VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X210 a_n2195_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t18 a_n2345_n9098# GND.t154 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X211 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND a_n787_n6852# GND.t142 GND.t141 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X212 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t19 GND.t153 GND.t152 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X213 a_n432_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t11 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X214 s1.t1 a_275_n2786# GND.t127 GND.t126 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X215 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t0 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t19 VDD.t130 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X216 GND.t71 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B a_1637_1038# GND.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X217 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t15 a_n2290_n2118# GND.t161 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X218 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND a_n787_n10008# VDD.t120 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X219 VDD.t7 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n787_n10008# VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X220 a_n787_n10008# CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n787_n9098# GND.t3 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X221 VDD.t103 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t16 a_n2345_n6852# VDD.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X222 s3.t0 a_275_n9098# VDD.t73 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X223 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t0 x0.t1 a_n4695_1648# VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X224 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t19 a_n732_n1508# VDD.t155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X225 a_n4695_1648# k0_bar.t1 VDD.t87 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X226 a_n1990_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t17 a_n2140_n540# VDD.t101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X227 VDD.t94 k2.t1 a_n4395_n1508# VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
R0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t18 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t7 1221.07
R1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n10 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t17 993.097
R2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n13 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t5 993.097
R3 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t10 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t6 924.95
R4 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t15 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t9 924.95
R5 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t14 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t8 923.343
R6 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t10 633.02
R7 CMOS_sbox_0/CMOS_s2_0/CMOS_XOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t15 633.02
R8 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t14 633.02
R9 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t19 579.86
R10 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t16 570.366
R11 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t12 570.366
R12 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t13 547.727
R13 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n6 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/B 539.692
R14 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n12 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/B 539.692
R15 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n6 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/B 427.962
R16 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n8 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/C 422.28
R17 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t18 392.02
R18 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n11 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 391.88
R19 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n14 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/A 391.88
R20 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n10 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t4 356.59
R21 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n13 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t11 356.59
R22 CMOS_4in_XOR_0/CMOS_INV_2/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n5 78.72
R23 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n7 78.72
R24 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n10 78.72
R25 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n13 78.72
R26 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n16 CMOS_4in_XOR_0/CMOS_INV_2/A 57.376
R27 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n9 CMOS_sbox_0/CMOS_s2_0/CMOS_XOR_0/B 45.03
R28 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n18 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t2 24
R29 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n18 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t3 24
R30 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n43 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t1 19.7
R31 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n43 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t0 19.7
R32 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n19 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n18 8.472
R33 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n25 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n23 5.44
R34 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n25 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n24 5.44
R35 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n42 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n41 4.61
R36 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n30 4.609
R37 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n28 4.5
R38 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n17 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n21 4.5
R39 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n42 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n47 4.5
R40 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n37 4.5
R41 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n48 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n52 4.5
R42 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n4 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n54 4.302
R43 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n45 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n44 3.472
R44 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n9 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n8 3.393
R45 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n11 CMOS_sbox_0/CMOS_s2_0/x0 3.332
R46 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n25 3.144
R47 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n14 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n12 3.064
R48 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n38 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n29 3.018
R49 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n44 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n43 2.773
R50 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n41 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n39 2.56
R51 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n47 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n46 2.56
R52 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n21 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n19 2.4
R53 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n28 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n27 2.4
R54 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n30 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n31 2.24
R55 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n37 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n34 1.92
R56 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n52 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n51 1.92
R57 CMOS_sbox_0/CMOS_s1_0/x0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n11 1.597
R58 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n38 1.383
R59 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n8 CMOS_sbox_0/CMOS_s3_0/x0 1.374
R60 CMOS_4in_XOR_0/XOR0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n15 1.253
R61 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n15 CMOS_sbox_0/CMOS_s0_0/x0 1.252
R62 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n17 1.125
R63 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n4 1.125
R64 CMOS_4in_XOR_0/CMOS_XOR_3/XOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n55 1.062
R65 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n3 1.159
R66 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n37 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n36 0.8
R67 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n52 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n50 0.8
R68 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n16 CMOS_4in_XOR_0/XOR0 0.796
R69 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n55 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n1 0.538
R70 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n55 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n0 0.53
R71 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n30 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n33 0.48
R72 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n15 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n14 0.335
R73 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n21 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n20 0.32
R74 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n28 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n26 0.32
R75 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n12 CMOS_sbox_0/CMOS_s1_0/x0 0.267
R76 CMOS_sbox_0/CMOS_s3_0/x0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n6 0.217
R77 CMOS_4in_XOR_0/CMOS_XOR_3/XOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n16 0.215
R78 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n41 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n40 0.16
R79 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n47 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n45 0.16
R80 CMOS_sbox_0/CMOS_s2_0/x0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n9 0.156
R81 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n4 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n48 0.114
R82 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n48 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n42 0.221
R83 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n38 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n2 0.092
R84 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n17 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n22 0.079
R85 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n54 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n53 0.059
R86 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n50 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n49 0.055
R87 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n36 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n35 0.055
R88 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n33 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n32 0.05
R89 GND.n792 GND.t152 4563.98
R90 GND.n792 GND.t145 4563.98
R91 GND.n808 GND.t112 4563.98
R92 GND.n808 GND.t135 4563.98
R93 GND.n125 GND.t110 2383.33
R94 GND.n476 GND.t24 2383.33
R95 GND.n698 GND.t72 1283.79
R96 GND.n699 GND.n698 284.705
R97 GND.n572 GND.t118 180.204
R98 GND.n801 GND.n800 164.96
R99 GND.n810 GND.n804 164.96
R100 GND.n162 GND.t158 159.607
R101 GND.n93 GND.t134 159.607
R102 GND.n336 GND.t104 159.607
R103 GND.n269 GND.t157 159.607
R104 GND.n722 GND.t131 159.607
R105 GND.n753 GND.t138 159.607
R106 GND.n444 GND.t137 159.607
R107 GND.n513 GND.t161 159.607
R108 GND.n126 GND.n125 150.98
R109 GND.n477 GND.n476 150.98
R110 GND.n4 GND.t65 150.98
R111 GND.n564 GND.t70 135.153
R112 GND.n170 GND.t33 133.725
R113 GND.n101 GND.t100 133.725
R114 GND.n344 GND.t132 133.725
R115 GND.n277 GND.t87 133.725
R116 GND.n730 GND.t79 133.725
R117 GND.n744 GND.t8 133.725
R118 GND.n452 GND.t31 133.725
R119 GND.n521 GND.t159 133.725
R120 GND.n857 GND.t18 133.725
R121 GND.n152 GND.t66 125.098
R122 GND.n81 GND.t89 125.098
R123 GND.n326 GND.t56 125.098
R124 GND.n257 GND.t149 125.098
R125 GND.n712 GND.t0 125.098
R126 GND.n764 GND.t59 125.098
R127 GND.n432 GND.t67 125.098
R128 GND.n503 GND.t148 125.098
R129 GND.n839 GND.t46 125.098
R130 GND.n170 GND.t129 103.529
R131 GND.n101 GND.t38 103.529
R132 GND.n54 GND.t20 103.529
R133 GND.n300 GND.t47 103.529
R134 GND.n344 GND.t44 103.529
R135 GND.n277 GND.t150 103.529
R136 GND.n230 GND.t143 103.529
R137 GND.n665 GND.t6 103.529
R138 GND.n618 GND.t4 103.529
R139 GND.n452 GND.t74 103.529
R140 GND.n405 GND.t27 103.529
R141 GND.n521 GND.t16 103.529
R142 GND.n144 GND.t92 99.215
R143 GND.n72 GND.t57 99.215
R144 GND.n318 GND.t10 99.215
R145 GND.n248 GND.t49 99.215
R146 GND.n704 GND.t35 99.215
R147 GND.n772 GND.t40 99.215
R148 GND.n423 GND.t105 99.215
R149 GND.n495 GND.t14 99.215
R150 GND.n831 GND.t76 99.215
R151 GND.n542 GND.t85 90.102
R152 GND.n134 GND.t63 77.647
R153 GND.n162 GND.t154 77.647
R154 GND.n93 GND.t3 77.647
R155 GND.n14 GND.t96 77.647
R156 GND.n45 GND.t68 77.647
R157 GND.n295 GND.t61 77.647
R158 GND.n336 GND.t155 77.647
R159 GND.n269 GND.t60 77.647
R160 GND.n190 GND.t114 77.647
R161 GND.n221 GND.t52 77.647
R162 GND.n657 GND.t12 77.647
R163 GND.n610 GND.t81 77.647
R164 GND.n444 GND.t124 77.647
R165 GND.n365 GND.t126 77.647
R166 GND.n396 GND.t22 77.647
R167 GND.n485 GND.t102 77.647
R168 GND.n513 GND.t121 77.647
R169 GND.n156 GND.t26 51.764
R170 GND.n72 GND.t122 51.764
R171 GND.n23 GND.t83 51.764
R172 GND.n37 GND.t94 51.764
R173 GND.n330 GND.t37 51.764
R174 GND.n248 GND.t141 51.764
R175 GND.n199 GND.t54 51.764
R176 GND.n213 GND.t90 51.764
R177 GND.n635 GND.t98 51.764
R178 GND.n589 GND.t1 51.764
R179 GND.n423 GND.t108 51.764
R180 GND.n374 GND.t139 51.764
R181 GND.n388 GND.t29 51.764
R182 GND.n507 GND.t78 51.764
R183 GND GND.n863 45.074
R184 CMOS_4in_XOR_0/GND GND.n0 40.19
R185 GND.n181 GND.n180 37.883
R186 GND.n355 GND.n354 35.52
R187 GND.n801 GND.n736 35.52
R188 GND.n804 GND.n531 35.52
R189 GND.n743 GND.t43 30.21
R190 GND.n6 GND.t136 30.21
R191 GND.n830 GND.t163 30.21
R192 GND.n861 GND.t147 30.21
R193 GND.n179 GND.t130 30.21
R194 GND.n138 GND.t64 30.21
R195 GND.n110 GND.t39 30.21
R196 GND.n76 GND.t123 30.21
R197 GND.n36 GND.t95 30.21
R198 GND.n18 GND.t97 30.21
R199 GND.n353 GND.t45 30.21
R200 GND.n304 GND.t48 30.21
R201 GND.n286 GND.t151 30.21
R202 GND.n252 GND.t142 30.21
R203 GND.n212 GND.t91 30.21
R204 GND.n194 GND.t115 30.21
R205 GND.n593 GND.t2 30.21
R206 GND.n626 GND.t5 30.21
R207 GND.n639 GND.t128 30.21
R208 GND.n673 GND.t120 30.21
R209 GND.n703 GND.t36 30.21
R210 GND.n734 GND.t80 30.21
R211 GND.n685 GND.t73 30.21
R212 GND.n738 GND.t146 30.21
R213 GND.n776 GND.t51 30.21
R214 GND.n743 GND.t9 30.21
R215 GND.n530 GND.t17 30.21
R216 GND.n489 GND.t103 30.21
R217 GND.n461 GND.t75 30.21
R218 GND.n427 GND.t109 30.21
R219 GND.n387 GND.t30 30.21
R220 GND.n369 GND.t127 30.21
R221 GND.n6 GND.t113 30.21
R222 GND.n830 GND.t77 30.21
R223 GND.n861 GND.t19 30.21
R224 GND.n27 GND.t84 30.21
R225 GND.n62 GND.t21 30.21
R226 GND.n71 GND.t58 30.21
R227 GND.n105 GND.t101 30.21
R228 GND.n124 GND.t111 30.21
R229 GND.n143 GND.t93 30.21
R230 GND.n174 GND.t34 30.21
R231 GND.n203 GND.t55 30.21
R232 GND.n238 GND.t162 30.21
R233 GND.n247 GND.t50 30.21
R234 GND.n281 GND.t88 30.21
R235 GND.n299 GND.t62 30.21
R236 GND.n317 GND.t11 30.21
R237 GND.n348 GND.t133 30.21
R238 GND.n546 GND.t86 30.21
R239 GND.n559 GND.t71 30.21
R240 GND.n580 GND.t119 30.21
R241 GND.n593 GND.t125 30.21
R242 GND.n626 GND.t117 30.21
R243 GND.n639 GND.t99 30.21
R244 GND.n652 GND.t13 30.21
R245 GND.n673 GND.t7 30.21
R246 GND.n703 GND.t107 30.21
R247 GND.n734 GND.t156 30.21
R248 GND.n738 GND.t153 30.21
R249 GND.n776 GND.t41 30.21
R250 GND.n378 GND.t140 30.21
R251 GND.n413 GND.t28 30.21
R252 GND.n422 GND.t106 30.21
R253 GND.n456 GND.t32 30.21
R254 GND.n475 GND.t25 30.21
R255 GND.n494 GND.t15 30.21
R256 GND.n525 GND.t160 30.21
R257 GND.n808 GND.n807 28.947
R258 GND.n322 GND.t42 25.882
R259 GND.n9 GND.t69 24
R260 GND.n9 GND.t116 24
R261 GND.n185 GND.t53 24
R262 GND.n185 GND.t144 24
R263 GND.n360 GND.t23 24
R264 GND.n360 GND.t82 24
R265 GND.n810 GND.n809 17.263
R266 GND.n95 GND.n92 11.52
R267 GND.n47 GND.n44 11.52
R268 GND.n164 GND.n161 11.52
R269 GND.n271 GND.n268 11.52
R270 GND.n223 GND.n220 11.52
R271 GND.n338 GND.n335 11.52
R272 GND.n659 GND.n656 11.52
R273 GND.n612 GND.n609 11.52
R274 GND.n566 GND.n563 11.52
R275 GND.n724 GND.n721 11.52
R276 GND.n797 GND.n795 11.52
R277 GND.n758 GND.n755 11.52
R278 GND.n446 GND.n443 11.52
R279 GND.n398 GND.n395 11.52
R280 GND.n515 GND.n512 11.52
R281 GND.n817 GND.n816 11.52
R282 GND.n851 GND.n848 11.52
R283 GND.n355 GND.n182 9.77
R284 GND.n804 GND.n357 9.77
R285 GND.n802 GND.n801 9.77
R286 GND.n12 GND.n11 9.154
R287 GND.n16 GND.n15 9.154
R288 GND.n15 GND.n14 9.154
R289 GND.n21 GND.n20 9.154
R290 GND.n20 GND.n19 9.154
R291 GND.n25 GND.n24 9.154
R292 GND.n24 GND.n23 9.154
R293 GND.n30 GND.n29 9.154
R294 GND.n29 GND.n28 9.154
R295 GND.n34 GND.n33 9.154
R296 GND.n33 GND.n32 9.154
R297 GND.n39 GND.n38 9.154
R298 GND.n38 GND.n37 9.154
R299 GND.n44 GND.n43 9.154
R300 GND.n43 GND.n42 9.154
R301 GND.n47 GND.n46 9.154
R302 GND.n46 GND.n45 9.154
R303 GND.n51 GND.n50 9.154
R304 GND.n50 GND.n49 9.154
R305 GND.n56 GND.n55 9.154
R306 GND.n55 GND.n54 9.154
R307 GND.n60 GND.n59 9.154
R308 GND.n69 GND.n68 9.154
R309 GND.n74 GND.n73 9.154
R310 GND.n73 GND.n72 9.154
R311 GND.n79 GND.n78 9.154
R312 GND.n78 GND.n77 9.154
R313 GND.n83 GND.n82 9.154
R314 GND.n82 GND.n81 9.154
R315 GND.n87 GND.n86 9.154
R316 GND.n86 GND.n85 9.154
R317 GND.n92 GND.n91 9.154
R318 GND.n91 GND.n90 9.154
R319 GND.n95 GND.n94 9.154
R320 GND.n94 GND.n93 9.154
R321 GND.n99 GND.n98 9.154
R322 GND.n98 GND.n97 9.154
R323 GND.n103 GND.n102 9.154
R324 GND.n102 GND.n101 9.154
R325 GND.n108 GND.n107 9.154
R326 GND.n114 GND.n113 9.154
R327 GND.n117 GND.n116 9.154
R328 GND.n122 GND.n121 9.154
R329 GND.n128 GND.n127 9.154
R330 GND.n127 GND.n126 9.154
R331 GND.n132 GND.n131 9.154
R332 GND.n131 GND.n130 9.154
R333 GND.n136 GND.n135 9.154
R334 GND.n135 GND.n134 9.154
R335 GND.n141 GND.n140 9.154
R336 GND.n140 GND.n139 9.154
R337 GND.n146 GND.n145 9.154
R338 GND.n145 GND.n144 9.154
R339 GND.n150 GND.n149 9.154
R340 GND.n149 GND.n148 9.154
R341 GND.n154 GND.n153 9.154
R342 GND.n153 GND.n152 9.154
R343 GND.n158 GND.n157 9.154
R344 GND.n157 GND.n156 9.154
R345 GND.n161 GND.n8 9.154
R346 GND.n8 GND.n7 9.154
R347 GND.n164 GND.n163 9.154
R348 GND.n163 GND.n162 9.154
R349 GND.n168 GND.n167 9.154
R350 GND.n167 GND.n166 9.154
R351 GND.n172 GND.n171 9.154
R352 GND.n171 GND.n170 9.154
R353 GND.n177 GND.n176 9.154
R354 GND.n188 GND.n187 9.154
R355 GND.n192 GND.n191 9.154
R356 GND.n191 GND.n190 9.154
R357 GND.n197 GND.n196 9.154
R358 GND.n196 GND.n195 9.154
R359 GND.n201 GND.n200 9.154
R360 GND.n200 GND.n199 9.154
R361 GND.n206 GND.n205 9.154
R362 GND.n205 GND.n204 9.154
R363 GND.n210 GND.n209 9.154
R364 GND.n209 GND.n208 9.154
R365 GND.n215 GND.n214 9.154
R366 GND.n214 GND.n213 9.154
R367 GND.n220 GND.n219 9.154
R368 GND.n219 GND.n218 9.154
R369 GND.n223 GND.n222 9.154
R370 GND.n222 GND.n221 9.154
R371 GND.n227 GND.n226 9.154
R372 GND.n226 GND.n225 9.154
R373 GND.n232 GND.n231 9.154
R374 GND.n231 GND.n230 9.154
R375 GND.n236 GND.n235 9.154
R376 GND.n245 GND.n244 9.154
R377 GND.n250 GND.n249 9.154
R378 GND.n249 GND.n248 9.154
R379 GND.n255 GND.n254 9.154
R380 GND.n254 GND.n253 9.154
R381 GND.n259 GND.n258 9.154
R382 GND.n258 GND.n257 9.154
R383 GND.n263 GND.n262 9.154
R384 GND.n262 GND.n261 9.154
R385 GND.n268 GND.n267 9.154
R386 GND.n267 GND.n266 9.154
R387 GND.n271 GND.n270 9.154
R388 GND.n270 GND.n269 9.154
R389 GND.n275 GND.n274 9.154
R390 GND.n274 GND.n273 9.154
R391 GND.n279 GND.n278 9.154
R392 GND.n278 GND.n277 9.154
R393 GND.n284 GND.n283 9.154
R394 GND.n293 GND.n292 9.154
R395 GND.n297 GND.n296 9.154
R396 GND.n296 GND.n295 9.154
R397 GND.n302 GND.n301 9.154
R398 GND.n301 GND.n300 9.154
R399 GND.n307 GND.n306 9.154
R400 GND.n306 GND.n305 9.154
R401 GND.n311 GND.n310 9.154
R402 GND.n310 GND.n309 9.154
R403 GND.n315 GND.n314 9.154
R404 GND.n314 GND.n313 9.154
R405 GND.n320 GND.n319 9.154
R406 GND.n319 GND.n318 9.154
R407 GND.n324 GND.n323 9.154
R408 GND.n323 GND.n322 9.154
R409 GND.n328 GND.n327 9.154
R410 GND.n327 GND.n326 9.154
R411 GND.n332 GND.n331 9.154
R412 GND.n331 GND.n330 9.154
R413 GND.n335 GND.n184 9.154
R414 GND.n184 GND.n183 9.154
R415 GND.n338 GND.n337 9.154
R416 GND.n337 GND.n336 9.154
R417 GND.n342 GND.n341 9.154
R418 GND.n341 GND.n340 9.154
R419 GND.n346 GND.n345 9.154
R420 GND.n345 GND.n344 9.154
R421 GND.n351 GND.n350 9.154
R422 GND.n540 GND.n539 9.154
R423 GND.n544 GND.n543 9.154
R424 GND.n543 GND.n542 9.154
R425 GND.n549 GND.n548 9.154
R426 GND.n548 GND.n547 9.154
R427 GND.n553 GND.n552 9.154
R428 GND.n552 GND.n551 9.154
R429 GND.n557 GND.n556 9.154
R430 GND.n556 GND.n555 9.154
R431 GND.n563 GND.n562 9.154
R432 GND.n562 GND.n561 9.154
R433 GND.n566 GND.n565 9.154
R434 GND.n565 GND.n564 9.154
R435 GND.n570 GND.n569 9.154
R436 GND.n569 GND.n568 9.154
R437 GND.n574 GND.n573 9.154
R438 GND.n573 GND.n572 9.154
R439 GND.n578 GND.n577 9.154
R440 GND.n587 GND.n586 9.154
R441 GND.n591 GND.n590 9.154
R442 GND.n590 GND.n589 9.154
R443 GND.n596 GND.n595 9.154
R444 GND.n595 GND.n594 9.154
R445 GND.n600 GND.n599 9.154
R446 GND.n599 GND.n598 9.154
R447 GND.n604 GND.n603 9.154
R448 GND.n603 GND.n602 9.154
R449 GND.n609 GND.n608 9.154
R450 GND.n608 GND.n607 9.154
R451 GND.n612 GND.n611 9.154
R452 GND.n611 GND.n610 9.154
R453 GND.n616 GND.n615 9.154
R454 GND.n615 GND.n614 9.154
R455 GND.n620 GND.n619 9.154
R456 GND.n619 GND.n618 9.154
R457 GND.n624 GND.n623 9.154
R458 GND.n633 GND.n632 9.154
R459 GND.n637 GND.n636 9.154
R460 GND.n636 GND.n635 9.154
R461 GND.n642 GND.n641 9.154
R462 GND.n641 GND.n640 9.154
R463 GND.n646 GND.n645 9.154
R464 GND.n645 GND.n644 9.154
R465 GND.n650 GND.n649 9.154
R466 GND.n649 GND.n648 9.154
R467 GND.n656 GND.n655 9.154
R468 GND.n655 GND.n654 9.154
R469 GND.n659 GND.n658 9.154
R470 GND.n658 GND.n657 9.154
R471 GND.n663 GND.n662 9.154
R472 GND.n662 GND.n661 9.154
R473 GND.n667 GND.n666 9.154
R474 GND.n666 GND.n665 9.154
R475 GND.n671 GND.n670 9.154
R476 GND.n680 GND.n679 9.154
R477 GND.n683 GND.n682 9.154
R478 GND.n688 GND.n687 9.154
R479 GND.n691 GND.n690 9.154
R480 GND.n696 GND.n695 9.154
R481 GND.n701 GND.n700 9.154
R482 GND.n700 GND.n699 9.154
R483 GND.n706 GND.n705 9.154
R484 GND.n705 GND.n704 9.154
R485 GND.n710 GND.n709 9.154
R486 GND.n709 GND.n708 9.154
R487 GND.n714 GND.n713 9.154
R488 GND.n713 GND.n712 9.154
R489 GND.n718 GND.n717 9.154
R490 GND.n717 GND.n716 9.154
R491 GND.n721 GND.n537 9.154
R492 GND.n537 GND.n536 9.154
R493 GND.n724 GND.n723 9.154
R494 GND.n723 GND.n722 9.154
R495 GND.n728 GND.n727 9.154
R496 GND.n727 GND.n726 9.154
R497 GND.n732 GND.n731 9.154
R498 GND.n731 GND.n730 9.154
R499 GND.n535 GND.n534 9.154
R500 GND.n797 GND.n796 9.154
R501 GND.n795 GND.n794 9.154
R502 GND.n787 GND.n786 9.154
R503 GND.n786 GND.n785 9.154
R504 GND.n783 GND.n782 9.154
R505 GND.n782 GND.n781 9.154
R506 GND.n779 GND.n778 9.154
R507 GND.n778 GND.n777 9.154
R508 GND.n774 GND.n773 9.154
R509 GND.n773 GND.n772 9.154
R510 GND.n770 GND.n769 9.154
R511 GND.n769 GND.n768 9.154
R512 GND.n766 GND.n765 9.154
R513 GND.n765 GND.n764 9.154
R514 GND.n762 GND.n761 9.154
R515 GND.n761 GND.n760 9.154
R516 GND.n758 GND.n757 9.154
R517 GND.n757 GND.n756 9.154
R518 GND.n755 GND.n754 9.154
R519 GND.n754 GND.n753 9.154
R520 GND.n750 GND.n749 9.154
R521 GND.n749 GND.n748 9.154
R522 GND.n746 GND.n745 9.154
R523 GND.n745 GND.n744 9.154
R524 GND.n741 GND.n740 9.154
R525 GND.n363 GND.n362 9.154
R526 GND.n367 GND.n366 9.154
R527 GND.n366 GND.n365 9.154
R528 GND.n372 GND.n371 9.154
R529 GND.n371 GND.n370 9.154
R530 GND.n376 GND.n375 9.154
R531 GND.n375 GND.n374 9.154
R532 GND.n381 GND.n380 9.154
R533 GND.n380 GND.n379 9.154
R534 GND.n385 GND.n384 9.154
R535 GND.n384 GND.n383 9.154
R536 GND.n390 GND.n389 9.154
R537 GND.n389 GND.n388 9.154
R538 GND.n395 GND.n394 9.154
R539 GND.n394 GND.n393 9.154
R540 GND.n398 GND.n397 9.154
R541 GND.n397 GND.n396 9.154
R542 GND.n402 GND.n401 9.154
R543 GND.n401 GND.n400 9.154
R544 GND.n407 GND.n406 9.154
R545 GND.n406 GND.n405 9.154
R546 GND.n411 GND.n410 9.154
R547 GND.n420 GND.n419 9.154
R548 GND.n425 GND.n424 9.154
R549 GND.n424 GND.n423 9.154
R550 GND.n430 GND.n429 9.154
R551 GND.n429 GND.n428 9.154
R552 GND.n434 GND.n433 9.154
R553 GND.n433 GND.n432 9.154
R554 GND.n438 GND.n437 9.154
R555 GND.n437 GND.n436 9.154
R556 GND.n443 GND.n442 9.154
R557 GND.n442 GND.n441 9.154
R558 GND.n446 GND.n445 9.154
R559 GND.n445 GND.n444 9.154
R560 GND.n450 GND.n449 9.154
R561 GND.n449 GND.n448 9.154
R562 GND.n454 GND.n453 9.154
R563 GND.n453 GND.n452 9.154
R564 GND.n459 GND.n458 9.154
R565 GND.n465 GND.n464 9.154
R566 GND.n468 GND.n467 9.154
R567 GND.n473 GND.n472 9.154
R568 GND.n479 GND.n478 9.154
R569 GND.n478 GND.n477 9.154
R570 GND.n483 GND.n482 9.154
R571 GND.n482 GND.n481 9.154
R572 GND.n487 GND.n486 9.154
R573 GND.n486 GND.n485 9.154
R574 GND.n492 GND.n491 9.154
R575 GND.n491 GND.n490 9.154
R576 GND.n497 GND.n496 9.154
R577 GND.n496 GND.n495 9.154
R578 GND.n501 GND.n500 9.154
R579 GND.n500 GND.n499 9.154
R580 GND.n505 GND.n504 9.154
R581 GND.n504 GND.n503 9.154
R582 GND.n509 GND.n508 9.154
R583 GND.n508 GND.n507 9.154
R584 GND.n512 GND.n359 9.154
R585 GND.n359 GND.n358 9.154
R586 GND.n515 GND.n514 9.154
R587 GND.n514 GND.n513 9.154
R588 GND.n519 GND.n518 9.154
R589 GND.n518 GND.n517 9.154
R590 GND.n523 GND.n522 9.154
R591 GND.n522 GND.n521 9.154
R592 GND.n528 GND.n527 9.154
R593 GND.n812 GND.n811 9.154
R594 GND.n816 GND.n815 9.154
R595 GND.n820 GND.n819 9.154
R596 GND.n824 GND.n823 9.154
R597 GND.n823 GND.n822 9.154
R598 GND.n828 GND.n827 9.154
R599 GND.n827 GND.n826 9.154
R600 GND.n833 GND.n832 9.154
R601 GND.n832 GND.n831 9.154
R602 GND.n837 GND.n836 9.154
R603 GND.n836 GND.n835 9.154
R604 GND.n841 GND.n840 9.154
R605 GND.n840 GND.n839 9.154
R606 GND.n845 GND.n844 9.154
R607 GND.n844 GND.n843 9.154
R608 GND.n848 GND.n5 9.154
R609 GND.n5 GND.n4 9.154
R610 GND.n851 GND.n850 9.154
R611 GND.n850 GND.n849 9.154
R612 GND.n855 GND.n854 9.154
R613 GND.n854 GND.n853 9.154
R614 GND.n859 GND.n858 9.154
R615 GND.n858 GND.n857 9.154
R616 GND.n3 GND.n2 9.154
R617 GND.n121 GND.n120 8.108
R618 GND.n11 GND.n10 8.108
R619 GND.n187 GND.n186 8.108
R620 GND.n679 GND.n678 8.108
R621 GND.n687 GND.n686 8.108
R622 GND.n695 GND.n694 8.108
R623 GND.n794 GND.n793 8.108
R624 GND.n791 GND.n790 8.108
R625 GND.n362 GND.n361 8.108
R626 GND.n472 GND.n471 8.108
R627 GND.n806 GND.n805 8.108
R628 GND.n53 GND.n9 6.21
R629 GND.n229 GND.n185 6.21
R630 GND.n404 GND.n360 6.21
R631 GND.n182 GND.n181 4.797
R632 GND.n803 GND.n802 4.782
R633 GND.n357 GND.n356 4.782
R634 GND.n180 GND.n179 4.706
R635 GND.n354 GND.n353 4.706
R636 GND.n531 GND.n530 4.706
R637 GND.n17 GND.n16 4.65
R638 GND.n22 GND.n21 4.65
R639 GND.n26 GND.n25 4.65
R640 GND.n31 GND.n30 4.65
R641 GND.n35 GND.n34 4.65
R642 GND.n40 GND.n39 4.65
R643 GND.n44 GND.n41 4.65
R644 GND.n48 GND.n47 4.65
R645 GND.n52 GND.n51 4.65
R646 GND.n57 GND.n56 4.65
R647 GND.n61 GND.n60 4.65
R648 GND.n64 GND.n63 4.65
R649 GND.n66 GND.n65 4.65
R650 GND.n70 GND.n69 4.65
R651 GND.n75 GND.n74 4.65
R652 GND.n80 GND.n79 4.65
R653 GND.n84 GND.n83 4.65
R654 GND.n88 GND.n87 4.65
R655 GND.n92 GND.n89 4.65
R656 GND.n96 GND.n95 4.65
R657 GND.n100 GND.n99 4.65
R658 GND.n104 GND.n103 4.65
R659 GND.n109 GND.n108 4.65
R660 GND.n112 GND.n111 4.65
R661 GND.n115 GND.n114 4.65
R662 GND.n118 GND.n117 4.65
R663 GND.n123 GND.n122 4.65
R664 GND.n129 GND.n128 4.65
R665 GND.n133 GND.n132 4.65
R666 GND.n137 GND.n136 4.65
R667 GND.n142 GND.n141 4.65
R668 GND.n147 GND.n146 4.65
R669 GND.n151 GND.n150 4.65
R670 GND.n155 GND.n154 4.65
R671 GND.n159 GND.n158 4.65
R672 GND.n161 GND.n160 4.65
R673 GND.n165 GND.n164 4.65
R674 GND.n169 GND.n168 4.65
R675 GND.n173 GND.n172 4.65
R676 GND.n178 GND.n177 4.65
R677 GND.n193 GND.n192 4.65
R678 GND.n198 GND.n197 4.65
R679 GND.n202 GND.n201 4.65
R680 GND.n207 GND.n206 4.65
R681 GND.n211 GND.n210 4.65
R682 GND.n216 GND.n215 4.65
R683 GND.n220 GND.n217 4.65
R684 GND.n224 GND.n223 4.65
R685 GND.n228 GND.n227 4.65
R686 GND.n233 GND.n232 4.65
R687 GND.n237 GND.n236 4.65
R688 GND.n240 GND.n239 4.65
R689 GND.n242 GND.n241 4.65
R690 GND.n246 GND.n245 4.65
R691 GND.n251 GND.n250 4.65
R692 GND.n256 GND.n255 4.65
R693 GND.n260 GND.n259 4.65
R694 GND.n264 GND.n263 4.65
R695 GND.n268 GND.n265 4.65
R696 GND.n272 GND.n271 4.65
R697 GND.n276 GND.n275 4.65
R698 GND.n280 GND.n279 4.65
R699 GND.n285 GND.n284 4.65
R700 GND.n288 GND.n287 4.65
R701 GND.n290 GND.n289 4.65
R702 GND.n294 GND.n293 4.65
R703 GND.n298 GND.n297 4.65
R704 GND.n303 GND.n302 4.65
R705 GND.n308 GND.n307 4.65
R706 GND.n312 GND.n311 4.65
R707 GND.n316 GND.n315 4.65
R708 GND.n321 GND.n320 4.65
R709 GND.n325 GND.n324 4.65
R710 GND.n329 GND.n328 4.65
R711 GND.n333 GND.n332 4.65
R712 GND.n335 GND.n334 4.65
R713 GND.n339 GND.n338 4.65
R714 GND.n343 GND.n342 4.65
R715 GND.n347 GND.n346 4.65
R716 GND.n352 GND.n351 4.65
R717 GND.n545 GND.n544 4.65
R718 GND.n550 GND.n549 4.65
R719 GND.n554 GND.n553 4.65
R720 GND.n558 GND.n557 4.65
R721 GND.n563 GND.n560 4.65
R722 GND.n567 GND.n566 4.65
R723 GND.n571 GND.n570 4.65
R724 GND.n575 GND.n574 4.65
R725 GND.n579 GND.n578 4.65
R726 GND.n582 GND.n581 4.65
R727 GND.n584 GND.n583 4.65
R728 GND.n588 GND.n587 4.65
R729 GND.n592 GND.n591 4.65
R730 GND.n597 GND.n596 4.65
R731 GND.n601 GND.n600 4.65
R732 GND.n605 GND.n604 4.65
R733 GND.n609 GND.n606 4.65
R734 GND.n613 GND.n612 4.65
R735 GND.n617 GND.n616 4.65
R736 GND.n621 GND.n620 4.65
R737 GND.n625 GND.n624 4.65
R738 GND.n628 GND.n627 4.65
R739 GND.n630 GND.n629 4.65
R740 GND.n634 GND.n633 4.65
R741 GND.n638 GND.n637 4.65
R742 GND.n643 GND.n642 4.65
R743 GND.n647 GND.n646 4.65
R744 GND.n651 GND.n650 4.65
R745 GND.n656 GND.n653 4.65
R746 GND.n660 GND.n659 4.65
R747 GND.n664 GND.n663 4.65
R748 GND.n668 GND.n667 4.65
R749 GND.n672 GND.n671 4.65
R750 GND.n675 GND.n674 4.65
R751 GND.n677 GND.n676 4.65
R752 GND.n681 GND.n680 4.65
R753 GND.n684 GND.n683 4.65
R754 GND.n689 GND.n688 4.65
R755 GND.n692 GND.n691 4.65
R756 GND.n697 GND.n696 4.65
R757 GND.n702 GND.n701 4.65
R758 GND.n707 GND.n706 4.65
R759 GND.n711 GND.n710 4.65
R760 GND.n715 GND.n714 4.65
R761 GND.n719 GND.n718 4.65
R762 GND.n721 GND.n720 4.65
R763 GND.n725 GND.n724 4.65
R764 GND.n729 GND.n728 4.65
R765 GND.n733 GND.n732 4.65
R766 GND.n798 GND.n797 4.65
R767 GND.n795 GND.n789 4.65
R768 GND.n788 GND.n787 4.65
R769 GND.n784 GND.n783 4.65
R770 GND.n780 GND.n779 4.65
R771 GND.n775 GND.n774 4.65
R772 GND.n771 GND.n770 4.65
R773 GND.n767 GND.n766 4.65
R774 GND.n763 GND.n762 4.65
R775 GND.n759 GND.n758 4.65
R776 GND.n755 GND.n752 4.65
R777 GND.n751 GND.n750 4.65
R778 GND.n747 GND.n746 4.65
R779 GND.n368 GND.n367 4.65
R780 GND.n373 GND.n372 4.65
R781 GND.n377 GND.n376 4.65
R782 GND.n382 GND.n381 4.65
R783 GND.n386 GND.n385 4.65
R784 GND.n391 GND.n390 4.65
R785 GND.n395 GND.n392 4.65
R786 GND.n399 GND.n398 4.65
R787 GND.n403 GND.n402 4.65
R788 GND.n408 GND.n407 4.65
R789 GND.n412 GND.n411 4.65
R790 GND.n415 GND.n414 4.65
R791 GND.n417 GND.n416 4.65
R792 GND.n421 GND.n420 4.65
R793 GND.n426 GND.n425 4.65
R794 GND.n431 GND.n430 4.65
R795 GND.n435 GND.n434 4.65
R796 GND.n439 GND.n438 4.65
R797 GND.n443 GND.n440 4.65
R798 GND.n447 GND.n446 4.65
R799 GND.n451 GND.n450 4.65
R800 GND.n455 GND.n454 4.65
R801 GND.n460 GND.n459 4.65
R802 GND.n463 GND.n462 4.65
R803 GND.n466 GND.n465 4.65
R804 GND.n469 GND.n468 4.65
R805 GND.n474 GND.n473 4.65
R806 GND.n480 GND.n479 4.65
R807 GND.n484 GND.n483 4.65
R808 GND.n488 GND.n487 4.65
R809 GND.n493 GND.n492 4.65
R810 GND.n498 GND.n497 4.65
R811 GND.n502 GND.n501 4.65
R812 GND.n506 GND.n505 4.65
R813 GND.n510 GND.n509 4.65
R814 GND.n512 GND.n511 4.65
R815 GND.n516 GND.n515 4.65
R816 GND.n520 GND.n519 4.65
R817 GND.n524 GND.n523 4.65
R818 GND.n529 GND.n528 4.65
R819 GND.n816 GND.n814 4.65
R820 GND.n818 GND.n817 4.65
R821 GND.n821 GND.n820 4.65
R822 GND.n825 GND.n824 4.65
R823 GND.n829 GND.n828 4.65
R824 GND.n834 GND.n833 4.65
R825 GND.n838 GND.n837 4.65
R826 GND.n842 GND.n841 4.65
R827 GND.n846 GND.n845 4.65
R828 GND.n848 GND.n847 4.65
R829 GND.n852 GND.n851 4.65
R830 GND.n856 GND.n855 4.65
R831 GND.n860 GND.n859 4.65
R832 GND.n804 GND.n803 3.127
R833 GND.n801 GND.n532 3.127
R834 GND.n356 GND.n355 3.127
R835 GND.n586 GND.n585 2.759
R836 GND.n632 GND.n631 2.759
R837 GND.n59 GND.n58 2.759
R838 GND.n235 GND.n234 2.759
R839 GND.n623 GND.n622 2.759
R840 GND.n670 GND.n669 2.759
R841 GND.n410 GND.n409 2.759
R842 GND.n813 GND.n810 2.613
R843 GND.n736 GND.n735 2.612
R844 GND.n800 GND.n799 2.612
R845 GND.n742 GND.n0 2.612
R846 GND.n863 GND.n862 2.612
R847 GND.n13 GND.n12 2.562
R848 GND.n189 GND.n188 2.562
R849 GND.n541 GND.n540 2.562
R850 GND.n364 GND.n363 2.562
R851 GND.n813 GND.n812 2.562
R852 GND.n735 GND.n535 2.562
R853 GND.n799 GND.n737 2.562
R854 GND.n742 GND.n741 2.562
R855 GND.n862 GND.n3 2.562
R856 GND.n532 CMOS_sbox_0/GND 2.379
R857 GND.n539 GND.n538 1.853
R858 GND.n577 GND.n576 1.853
R859 GND.n534 GND.n533 1.593
R860 GND.n2 GND.n1 1.593
R861 GND.n740 GND.n739 1.593
R862 GND.n814 GND.n813 1.145
R863 GND.n17 GND.n13 1.145
R864 GND.n193 GND.n189 1.145
R865 GND.n545 GND.n541 1.145
R866 GND.n368 GND.n364 1.145
R867 GND.n799 GND.n798 1.145
R868 GND.n862 GND.n861 1.09
R869 GND.n735 GND.n734 1.09
R870 GND.n743 GND.n742 1.09
R871 GND.n66 GND.n64 0.525
R872 GND.n242 GND.n240 0.525
R873 GND.n584 GND.n582 0.525
R874 GND.n630 GND.n628 0.525
R875 GND.n417 GND.n415 0.525
R876 GND.n120 GND.n119 0.524
R877 GND.n793 GND.n792 0.524
R878 GND.n694 GND.n693 0.524
R879 GND.n792 GND.n791 0.524
R880 GND.n471 GND.n470 0.524
R881 GND.n809 GND.n808 0.524
R882 GND.n808 GND.n806 0.524
R883 GND.n115 GND.n112 0.507
R884 GND.n290 GND.n288 0.507
R885 GND.n677 GND.n675 0.507
R886 GND.n466 GND.n463 0.507
R887 GND.n821 GND.n818 0.09
R888 GND.n825 GND.n821 0.09
R889 GND.n829 GND.n825 0.09
R890 GND.n838 GND.n834 0.09
R891 GND.n842 GND.n838 0.09
R892 GND.n846 GND.n842 0.09
R893 GND.n847 GND.n846 0.09
R894 GND.n856 GND.n852 0.09
R895 GND.n860 GND.n856 0.09
R896 GND.n26 GND.n22 0.09
R897 GND.n35 GND.n31 0.09
R898 GND.n41 GND.n40 0.09
R899 GND.n52 GND.n48 0.09
R900 GND.n61 GND.n57 0.09
R901 GND.n70 GND.n66 0.09
R902 GND.n84 GND.n80 0.09
R903 GND.n88 GND.n84 0.09
R904 GND.n89 GND.n88 0.09
R905 GND.n100 GND.n96 0.09
R906 GND.n104 GND.n100 0.09
R907 GND.n118 GND.n115 0.09
R908 GND.n123 GND.n118 0.09
R909 GND.n133 GND.n129 0.09
R910 GND.n137 GND.n133 0.09
R911 GND.n151 GND.n147 0.09
R912 GND.n155 GND.n151 0.09
R913 GND.n159 GND.n155 0.09
R914 GND.n160 GND.n159 0.09
R915 GND.n169 GND.n165 0.09
R916 GND.n173 GND.n169 0.09
R917 GND.n202 GND.n198 0.09
R918 GND.n211 GND.n207 0.09
R919 GND.n217 GND.n216 0.09
R920 GND.n228 GND.n224 0.09
R921 GND.n237 GND.n233 0.09
R922 GND.n246 GND.n242 0.09
R923 GND.n260 GND.n256 0.09
R924 GND.n264 GND.n260 0.09
R925 GND.n265 GND.n264 0.09
R926 GND.n276 GND.n272 0.09
R927 GND.n280 GND.n276 0.09
R928 GND.n294 GND.n290 0.09
R929 GND.n298 GND.n294 0.09
R930 GND.n312 GND.n308 0.09
R931 GND.n316 GND.n312 0.09
R932 GND.n325 GND.n321 0.09
R933 GND.n329 GND.n325 0.09
R934 GND.n333 GND.n329 0.09
R935 GND.n334 GND.n333 0.09
R936 GND.n343 GND.n339 0.09
R937 GND.n347 GND.n343 0.09
R938 GND.n554 GND.n550 0.09
R939 GND.n558 GND.n554 0.09
R940 GND.n560 GND.n558 0.09
R941 GND.n571 GND.n567 0.09
R942 GND.n575 GND.n571 0.09
R943 GND.n579 GND.n575 0.09
R944 GND.n588 GND.n584 0.09
R945 GND.n592 GND.n588 0.09
R946 GND.n601 GND.n597 0.09
R947 GND.n605 GND.n601 0.09
R948 GND.n606 GND.n605 0.09
R949 GND.n617 GND.n613 0.09
R950 GND.n621 GND.n617 0.09
R951 GND.n625 GND.n621 0.09
R952 GND.n634 GND.n630 0.09
R953 GND.n638 GND.n634 0.09
R954 GND.n647 GND.n643 0.09
R955 GND.n651 GND.n647 0.09
R956 GND.n653 GND.n651 0.09
R957 GND.n664 GND.n660 0.09
R958 GND.n668 GND.n664 0.09
R959 GND.n672 GND.n668 0.09
R960 GND.n681 GND.n677 0.09
R961 GND.n684 GND.n681 0.09
R962 GND.n692 GND.n689 0.09
R963 GND.n697 GND.n692 0.09
R964 GND.n702 GND.n697 0.09
R965 GND.n711 GND.n707 0.09
R966 GND.n715 GND.n711 0.09
R967 GND.n719 GND.n715 0.09
R968 GND.n720 GND.n719 0.09
R969 GND.n729 GND.n725 0.09
R970 GND.n733 GND.n729 0.09
R971 GND.n789 GND.n788 0.09
R972 GND.n788 GND.n784 0.09
R973 GND.n784 GND.n780 0.09
R974 GND.n775 GND.n771 0.09
R975 GND.n771 GND.n767 0.09
R976 GND.n767 GND.n763 0.09
R977 GND.n763 GND.n759 0.09
R978 GND.n752 GND.n751 0.09
R979 GND.n751 GND.n747 0.09
R980 GND.n377 GND.n373 0.09
R981 GND.n386 GND.n382 0.09
R982 GND.n392 GND.n391 0.09
R983 GND.n403 GND.n399 0.09
R984 GND.n412 GND.n408 0.09
R985 GND.n421 GND.n417 0.09
R986 GND.n435 GND.n431 0.09
R987 GND.n439 GND.n435 0.09
R988 GND.n440 GND.n439 0.09
R989 GND.n451 GND.n447 0.09
R990 GND.n455 GND.n451 0.09
R991 GND.n469 GND.n466 0.09
R992 GND.n474 GND.n469 0.09
R993 GND.n484 GND.n480 0.09
R994 GND.n488 GND.n484 0.09
R995 GND.n502 GND.n498 0.09
R996 GND.n506 GND.n502 0.09
R997 GND.n510 GND.n506 0.09
R998 GND.n511 GND.n510 0.09
R999 GND.n520 GND.n516 0.09
R1000 GND.n524 GND.n520 0.09
R1001 GND.n292 GND.n291 0.089
R1002 GND.n802 CMOS_sbox_0/CMOS_s0_0/GND 0.085
R1003 CMOS_sbox_0/CMOS_s1_0/GND GND.n357 0.085
R1004 GND.n182 CMOS_sbox_0/CMOS_s2_0/GND 0.085
R1005 GND.n27 GND.n26 0.078
R1006 GND.n40 GND.n36 0.078
R1007 GND.n76 GND.n75 0.078
R1008 GND.n203 GND.n202 0.078
R1009 GND.n216 GND.n212 0.078
R1010 GND.n252 GND.n251 0.078
R1011 GND.n546 GND.n545 0.078
R1012 GND.n593 GND.n592 0.078
R1013 GND.n639 GND.n638 0.078
R1014 GND.n378 GND.n377 0.078
R1015 GND.n391 GND.n387 0.078
R1016 GND.n427 GND.n426 0.078
R1017 GND.n527 GND.n526 0.074
R1018 GND.n107 GND.n106 0.074
R1019 GND.n176 GND.n175 0.074
R1020 GND.n283 GND.n282 0.074
R1021 GND.n350 GND.n349 0.074
R1022 GND.n458 GND.n457 0.074
R1023 GND.n18 GND.n17 0.072
R1024 GND.n194 GND.n193 0.072
R1025 GND.n369 GND.n368 0.072
R1026 GND.n124 GND.n123 0.071
R1027 GND.n138 GND.n137 0.071
R1028 GND.n299 GND.n298 0.071
R1029 GND.n685 GND.n684 0.071
R1030 GND.n475 GND.n474 0.071
R1031 GND.n489 GND.n488 0.071
R1032 GND.n834 GND.n830 0.065
R1033 GND.n852 CMOS_4in_XOR_0/CMOS_XOR_0/GND 0.065
R1034 GND.n48 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/GND 0.065
R1035 GND.n75 GND.n71 0.065
R1036 GND.n96 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/GND 0.065
R1037 GND.n147 GND.n143 0.065
R1038 GND.n165 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/GND 0.065
R1039 GND.n224 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/GND 0.065
R1040 GND.n251 GND.n247 0.065
R1041 GND.n272 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/GND 0.065
R1042 GND.n321 GND.n317 0.065
R1043 GND.n339 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/GND 0.065
R1044 GND.n567 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/GND 0.065
R1045 GND.n613 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/GND 0.065
R1046 GND.n660 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/GND 0.065
R1047 GND.n707 GND.n703 0.065
R1048 GND.n725 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/GND 0.065
R1049 GND.n776 GND.n775 0.065
R1050 GND.n752 CMOS_4in_XOR_0/CMOS_XOR_2/GND 0.065
R1051 GND.n399 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/GND 0.065
R1052 GND.n426 GND.n422 0.065
R1053 GND.n447 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/GND 0.065
R1054 GND.n498 GND.n494 0.065
R1055 GND.n516 GND 0.065
R1056 GND.n57 GND.n53 0.063
R1057 GND.n233 GND.n229 0.063
R1058 GND.n304 GND.n303 0.063
R1059 GND.n408 GND.n404 0.063
R1060 GND.n803 CMOS_sbox_0/CMOS_s1_0/GND 0.063
R1061 GND.n356 CMOS_sbox_0/CMOS_s2_0/GND 0.062
R1062 GND.n532 CMOS_sbox_0/CMOS_s0_0/GND 0.062
R1063 GND.n64 GND.n62 0.056
R1064 GND.n112 GND.n110 0.056
R1065 GND.n240 GND.n238 0.056
R1066 GND.n288 GND.n286 0.056
R1067 GND.n582 GND.n580 0.056
R1068 GND.n628 GND.n626 0.056
R1069 GND.n675 GND.n673 0.056
R1070 GND.n415 GND.n413 0.056
R1071 GND.n463 GND.n461 0.056
R1072 GND.n861 GND.n860 0.055
R1073 GND.n105 GND.n104 0.055
R1074 GND.n174 GND.n173 0.055
R1075 GND.n281 GND.n280 0.055
R1076 GND.n348 GND.n347 0.055
R1077 GND.n734 GND.n733 0.055
R1078 GND.n747 GND.n743 0.055
R1079 GND.n456 GND.n455 0.055
R1080 GND.n525 GND.n524 0.055
R1081 CMOS_4in_XOR_0/CMOS_INV_0/GND GND.n6 0.05
R1082 GND.n738 CMOS_4in_XOR_0/CMOS_INV_1/GND 0.05
R1083 GND.n181 CMOS_sbox_0/CMOS_s3_0/GND 0.048
R1084 GND.n68 GND.n67 0.047
R1085 GND.n244 GND.n243 0.047
R1086 GND.n419 GND.n418 0.047
R1087 GND.n109 GND.n105 0.035
R1088 GND.n178 GND.n174 0.035
R1089 GND.n285 GND.n281 0.035
R1090 GND.n352 GND.n348 0.035
R1091 GND.n460 GND.n456 0.035
R1092 GND.n529 GND.n525 0.035
R1093 GND.n62 GND.n61 0.033
R1094 GND.n110 GND.n109 0.033
R1095 GND.n179 GND.n178 0.033
R1096 GND.n238 GND.n237 0.033
R1097 GND.n286 GND.n285 0.033
R1098 GND.n353 GND.n352 0.033
R1099 GND.n580 GND.n579 0.033
R1100 GND.n626 GND.n625 0.033
R1101 GND.n673 GND.n672 0.033
R1102 GND.n413 GND.n412 0.033
R1103 GND.n461 GND.n460 0.033
R1104 GND.n530 GND.n529 0.033
R1105 GND.n53 GND.n52 0.026
R1106 GND.n229 GND.n228 0.026
R1107 GND.n308 GND.n304 0.026
R1108 GND.n404 GND.n403 0.026
R1109 GND.n830 GND.n829 0.025
R1110 GND.n847 CMOS_4in_XOR_0/CMOS_XOR_0/GND 0.025
R1111 GND.n41 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/GND 0.025
R1112 GND.n71 GND.n70 0.025
R1113 GND.n89 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/GND 0.025
R1114 GND.n143 GND.n142 0.025
R1115 GND.n160 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/GND 0.025
R1116 GND.n217 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/GND 0.025
R1117 GND.n247 GND.n246 0.025
R1118 GND.n265 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/GND 0.025
R1119 GND.n317 GND.n316 0.025
R1120 GND.n334 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/GND 0.025
R1121 GND.n606 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/GND 0.025
R1122 GND.n703 GND.n702 0.025
R1123 GND.n720 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/GND 0.025
R1124 GND.n780 GND.n776 0.025
R1125 GND.n759 CMOS_4in_XOR_0/CMOS_XOR_2/GND 0.025
R1126 GND.n392 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/GND 0.025
R1127 GND.n422 GND.n421 0.025
R1128 GND.n440 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/GND 0.025
R1129 GND.n494 GND.n493 0.025
R1130 GND.n511 GND 0.025
R1131 GND.n814 CMOS_4in_XOR_0/CMOS_INV_0/GND 0.021
R1132 GND.n798 CMOS_4in_XOR_0/CMOS_INV_1/GND 0.021
R1133 GND.n818 GND.n6 0.018
R1134 GND.n129 GND.n124 0.018
R1135 GND.n142 GND.n138 0.018
R1136 GND.n303 GND.n299 0.018
R1137 GND.n560 GND.n559 0.018
R1138 GND.n653 GND.n652 0.018
R1139 GND.n689 GND.n685 0.018
R1140 GND.n789 GND.n738 0.018
R1141 GND.n480 GND.n475 0.018
R1142 GND.n493 GND.n489 0.018
R1143 GND.n22 GND.n18 0.017
R1144 GND.n198 GND.n194 0.017
R1145 GND.n373 GND.n369 0.017
R1146 GND.n31 GND.n27 0.011
R1147 GND.n36 GND.n35 0.011
R1148 GND.n80 GND.n76 0.011
R1149 GND.n207 GND.n203 0.011
R1150 GND.n212 GND.n211 0.011
R1151 GND.n256 GND.n252 0.011
R1152 GND.n550 GND.n546 0.011
R1153 GND.n597 GND.n593 0.011
R1154 GND.n643 GND.n639 0.011
R1155 GND.n382 GND.n378 0.011
R1156 GND.n387 GND.n386 0.011
R1157 GND.n431 GND.n427 0.011
R1158 GND.n559 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/GND 0.006
R1159 GND.n652 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/GND 0.006
R1160 CMOS_4in_XOR_0/GND GND 0.006
R1161 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t14 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t11 1345.61
R1162 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t10 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t17 1345.61
R1163 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t9 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t12 1221.07
R1164 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n9 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t16 811.366
R1165 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t4 683.32
R1166 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n12 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t9 630.3
R1167 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t15 616.084
R1168 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t13 616.084
R1169 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t2 579.86
R1170 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t8 547.727
R1171 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t7 528.72
R1172 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t3 528.72
R1173 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t6 528.72
R1174 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t14 392.02
R1175 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t10 392.02
R1176 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n9 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t5 329.366
R1177 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n11 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/A_bar 286.14
R1178 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n2 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/A_bar 285.868
R1179 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n15 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n14 280.68
R1180 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n10 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/A 264.208
R1181 CMOS_4in_XOR_0/CMOS_INV_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t0 136.873
R1182 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n1 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/B_bar 125.96
R1183 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n9 78.72
R1184 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n15 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t1 76.998
R1185 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n13 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n12 38.547
R1186 CMOS_4in_XOR_0/CMOS_INV_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n15 28.16
R1187 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n8 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n7 12.409
R1188 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n4 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n3 12.409
R1189 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n8 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n6 11.74
R1190 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n6 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n5 8.764
R1191 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n15 CMOS_4in_XOR_0/XOR3_bar 3.805
R1192 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n7 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/B_bar 3.68
R1193 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 3.68
R1194 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n0 3.68
R1195 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n6 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/B 2.72
R1196 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n12 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/A 2.72
R1197 CMOS_sbox_0/CMOS_s1_0/x3_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n2 2.313
R1198 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n4 CMOS_sbox_0/CMOS_s1_0/x3_bar 2.167
R1199 CMOS_sbox_0/CMOS_s3_0/x3_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n8 2.167
R1200 CMOS_sbox_0/CMOS_s2_0/x3_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n11 2.112
R1201 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n10 CMOS_sbox_0/CMOS_s3_0/x3_bar 1.708
R1202 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n14 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n13 1.443
R1203 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n1 1.408
R1204 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n1 CMOS_sbox_0/CMOS_s0_0/x3_bar 1.202
R1205 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n11 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n10 1.109
R1206 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n14 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n4 1.015
R1207 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n13 CMOS_sbox_0/CMOS_s2_0/x3_bar 0.291
R1208 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t8 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t10 1221.07
R1209 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t11 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t7 1221.07
R1210 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n6 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t5 993.097
R1211 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t12 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t9 924.95
R1212 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t6 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t15 924.95
R1213 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/D CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t8 633.02
R1214 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t12 633.02
R1215 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t6 633.02
R1216 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t14 579.86
R1217 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t13 547.727
R1218 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n9 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/B 393.772
R1219 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n11 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 393.772
R1220 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_2/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t11 392.02
R1221 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n6 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t4 356.59
R1222 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n8 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/D 232.012
R1223 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n10 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_2/A 214.75
R1224 CMOS_4in_XOR_0/CMOS_INV_3/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n5 78.72
R1225 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n13 CMOS_4in_XOR_0/CMOS_INV_3/A 57.376
R1226 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n15 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t1 24
R1227 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n15 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t2 24
R1228 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n40 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t3 19.7
R1229 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n40 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t0 19.7
R1230 CMOS_sbox_0/CMOS_s3_0/x2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n7 16.257
R1231 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n6 8.764
R1232 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n16 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n15 8.472
R1233 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n22 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n20 5.44
R1234 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n22 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n21 5.44
R1235 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n39 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n38 4.61
R1236 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n27 4.609
R1237 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n25 4.5
R1238 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n14 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n18 4.5
R1239 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n34 4.5
R1240 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n39 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n44 4.5
R1241 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n45 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n49 4.5
R1242 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n9 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n8 4.448
R1243 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n4 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n51 4.302
R1244 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n12 CMOS_sbox_0/CMOS_s2_0/x2 3.602
R1245 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n42 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n41 3.472
R1246 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n22 3.144
R1247 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n35 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n26 3.02
R1248 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n41 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n40 2.773
R1249 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n7 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/A 2.72
R1250 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n10 CMOS_sbox_0/CMOS_s0_0/x2 2.618
R1251 CMOS_4in_XOR_0/XOR2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n12 2.614
R1252 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n38 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n36 2.56
R1253 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n44 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n43 2.56
R1254 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n18 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n16 2.4
R1255 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n25 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n24 2.4
R1256 CMOS_sbox_0/CMOS_s1_0/x2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n10 2.3
R1257 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n27 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n28 2.24
R1258 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n34 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n31 1.92
R1259 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n49 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n48 1.92
R1260 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n35 1.382
R1261 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n14 1.125
R1262 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n4 1.125
R1263 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n12 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n11 1.103
R1264 CMOS_4in_XOR_0/CMOS_XOR_0/XOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n52 1.062
R1265 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n3 1.159
R1266 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n34 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n33 0.8
R1267 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n49 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n47 0.8
R1268 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n13 CMOS_4in_XOR_0/XOR2 0.796
R1269 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n52 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n1 0.538
R1270 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n52 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n0 0.53
R1271 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n27 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n30 0.48
R1272 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n18 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n17 0.32
R1273 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n25 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n23 0.32
R1274 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n8 CMOS_sbox_0/CMOS_s3_0/x2 0.264
R1275 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n11 CMOS_sbox_0/CMOS_s1_0/x2 0.218
R1276 CMOS_sbox_0/CMOS_s2_0/x2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n9 0.218
R1277 CMOS_4in_XOR_0/CMOS_XOR_0/XOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n13 0.215
R1278 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n38 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n37 0.16
R1279 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n44 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n42 0.16
R1280 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n4 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n45 0.114
R1281 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n45 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n39 0.221
R1282 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n35 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n2 0.092
R1283 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n14 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n19 0.079
R1284 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n51 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n50 0.06
R1285 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n33 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n32 0.055
R1286 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n47 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n46 0.054
R1287 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n30 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n29 0.05
R1288 x2_bar.t1 x2_bar.t0 1345.61
R1289 x2_bar x2_bar.t1 392.02
R1290 x2_bar CMOS_4in_XOR_0/x2_bar 264.8
R1291 VDD.n626 VDD.n625 1822.05
R1292 VDD.t178 VDD.t95 552.101
R1293 VDD.n625 VDD.t49 535.897
R1294 VDD.n368 VDD.t63 371.739
R1295 VDD.n550 VDD.t44 371.739
R1296 VDD.t32 VDD.t140 206.521
R1297 VDD.t155 VDD.t106 206.521
R1298 VDD.t80 VDD.t24 206.521
R1299 VDD.t58 VDD.t135 206.521
R1300 VDD.t154 VDD.t104 206.521
R1301 VDD.t21 VDD.t2 206.521
R1302 VDD.t2 VDD.t14 206.521
R1303 VDD.t78 VDD.t12 206.521
R1304 VDD.t42 VDD.t171 206.521
R1305 VDD.t156 VDD.t168 206.521
R1306 VDD.t108 VDD.t139 206.521
R1307 VDD.t139 VDD.t28 206.521
R1308 VDD.n862 VDD.n861 200.48
R1309 VDD.n661 VDD.t146 196.884
R1310 VDD.n368 VDD.t80 165.217
R1311 VDD.n550 VDD.t78 165.217
R1312 VDD.n477 VDD.t21 112.898
R1313 VDD.n761 VDD.t155 110.144
R1314 VDD.n411 VDD.t154 110.144
R1315 VDD.n593 VDD.t156 110.144
R1316 VDD.n761 VDD.t32 96.376
R1317 VDD.n411 VDD.t58 96.376
R1318 VDD.n593 VDD.t42 96.376
R1319 VDD.n477 VDD.t178 93.623
R1320 VDD.n920 VDD.t11 38.206
R1321 VDD.n164 VDD.t182 38.206
R1322 VDD.n871 VDD.t16 36.141
R1323 VDD.n928 VDD.t90 32.01
R1324 VDD.n1014 VDD.t86 32.01
R1325 VDD.n172 VDD.t113 32.01
R1326 VDD.n908 VDD.t10 29.945
R1327 VDD.n1032 VDD.t22 29.945
R1328 VDD.n154 VDD.t159 29.945
R1329 VDD.n369 VDD.n368 29.141
R1330 VDD.n551 VDD.n550 29.141
R1331 VDD.n762 VDD.n761 26.226
R1332 VDD.n412 VDD.n411 26.226
R1333 VDD.n594 VDD.n593 26.226
R1334 VDD.n223 VDD.t99 24.782
R1335 VDD.n270 VDD.t111 24.782
R1336 VDD.n326 VDD.t131 24.782
R1337 VDD.n128 VDD.t166 24.782
R1338 VDD.n82 VDD.t115 24.782
R1339 VDD.n35 VDD.t117 24.782
R1340 VDD.n900 VDD.t70 23.75
R1341 VDD.n1040 VDD.t157 23.75
R1342 VDD.n146 VDD.t133 23.75
R1343 VDD.n779 VDD.t88 23.312
R1344 VDD.n380 VDD.t162 23.312
R1345 VDD.n429 VDD.t33 23.312
R1346 VDD.n454 VDD.t40 23.312
R1347 VDD.n504 VDD.t148 23.312
R1348 VDD.n562 VDD.t61 23.312
R1349 VDD.n611 VDD.t137 23.312
R1350 VDD.n684 VDD.t38 23.312
R1351 VDD.n704 VDD.t143 22.029
R1352 VDD.n717 VDD.t170 22.029
R1353 VDD.n738 VDD.t46 22.029
R1354 VDD.n801 VDD.t19 22.029
R1355 VDD.n818 VDD.t153 22.029
R1356 VDD.n851 VDD.t51 22.029
R1357 VDD.n388 VDD.t25 22.029
R1358 VDD.n508 VDD.t15 22.029
R1359 VDD.n471 VDD.t179 22.029
R1360 VDD.n453 VDD.t96 22.029
R1361 VDD.n433 VDD.t105 22.029
R1362 VDD.n397 VDD.t136 22.029
R1363 VDD.n366 VDD.t81 22.029
R1364 VDD.n353 VDD.t64 22.029
R1365 VDD.n570 VDD.t13 22.029
R1366 VDD.n688 VDD.t29 22.029
R1367 VDD.n652 VDD.t147 22.029
R1368 VDD.n634 VDD.t50 22.029
R1369 VDD.n615 VDD.t169 22.029
R1370 VDD.n579 VDD.t172 22.029
R1371 VDD.n548 VDD.t79 22.029
R1372 VDD.n535 VDD.t45 22.029
R1373 VDD.n176 VDD.t114 22.029
R1374 VDD.n145 VDD.t134 22.029
R1375 VDD.n136 VDD.t167 22.029
R1376 VDD.n103 VDD.t77 22.029
R1377 VDD.n90 VDD.t116 22.029
R1378 VDD.n69 VDD.t60 22.029
R1379 VDD.n56 VDD.t124 22.029
R1380 VDD.n43 VDD.t118 22.029
R1381 VDD.n10 VDD.t66 22.029
R1382 VDD.n783 VDD.t107 22.029
R1383 VDD.n747 VDD.t141 22.029
R1384 VDD.n939 VDD.t145 22.029
R1385 VDD.n965 VDD.t94 22.029
R1386 VDD.n998 VDD.t164 22.029
R1387 VDD.n1013 VDD.t87 22.029
R1388 VDD.n1044 VDD.t158 22.029
R1389 VDD.n1061 VDD.t175 22.029
R1390 VDD.n704 VDD.t5 22.029
R1391 VDD.n717 VDD.t75 22.029
R1392 VDD.n738 VDD.t9 22.029
R1393 VDD.n752 VDD.t128 22.029
R1394 VDD.n766 VDD.t151 22.029
R1395 VDD.n788 VDD.t89 22.029
R1396 VDD.n801 VDD.t56 22.029
R1397 VDD.n818 VDD.t173 22.029
R1398 VDD.n851 VDD.t31 22.029
R1399 VDD.n190 VDD.t73 22.029
R1400 VDD.n231 VDD.t100 22.029
R1401 VDD.n244 VDD.t120 22.029
R1402 VDD.n257 VDD.t7 22.029
R1403 VDD.n278 VDD.t112 22.029
R1404 VDD.n291 VDD.t53 22.029
R1405 VDD.n308 VDD.t27 22.029
R1406 VDD.n344 VDD.t98 22.029
R1407 VDD.n388 VDD.t163 22.029
R1408 VDD.n402 VDD.t161 22.029
R1409 VDD.n416 VDD.t48 22.029
R1410 VDD.n438 VDD.t34 22.029
R1411 VDD.n458 VDD.t41 22.029
R1412 VDD.n476 VDD.t103 22.029
R1413 VDD.n513 VDD.t149 22.029
R1414 VDD.n873 VDD.t130 22.029
R1415 VDD.n899 VDD.t71 22.029
R1416 VDD.n932 VDD.t91 22.029
R1417 VDD.n526 VDD.t126 22.029
R1418 VDD.n570 VDD.t62 22.029
R1419 VDD.n584 VDD.t93 22.029
R1420 VDD.n598 VDD.t122 22.029
R1421 VDD.n620 VDD.t138 22.029
R1422 VDD.n647 VDD.t83 22.029
R1423 VDD.n666 VDD.t110 22.029
R1424 VDD.n939 VDD.t165 22.029
R1425 VDD.n965 VDD.t36 22.029
R1426 VDD.n998 VDD.t68 22.029
R1427 VDD.n662 VDD.n661 21.37
R1428 VDD.n986 VDD.t37 21.073
R1429 VDD.n839 VDD.t142 21.073
R1430 VDD.n181 VDD.t181 19.7
R1431 VDD.n181 VDD.t132 19.7
R1432 VDD.n490 VDD.t85 19.7
R1433 VDD.n490 VDD.t177 19.7
R1434 VDD.n517 VDD.t1 19.7
R1435 VDD.n517 VDD.t39 19.7
R1436 VDD.n186 VDD.t72 18.586
R1437 VDD.n215 VDD.t54 18.586
R1438 VDD.n262 VDD.t6 18.586
R1439 VDD.n287 VDD.t52 18.586
R1440 VDD.n317 VDD.t180 18.586
R1441 VDD.n880 VDD.t129 18.586
R1442 VDD.n867 VDD.t174 18.586
R1443 VDD.n120 VDD.t69 18.586
R1444 VDD.n74 VDD.t59 18.586
R1445 VDD.n27 VDD.t55 18.586
R1446 VDD.n994 VDD.t67 17.655
R1447 VDD.n847 VDD.t30 17.655
R1448 VDD.n771 VDD.t150 17.484
R1449 VDD.n340 VDD.t97 17.484
R1450 VDD.n372 VDD.t43 17.484
R1451 VDD.n421 VDD.t47 17.484
R1452 VDD.n496 VDD.t176 17.484
R1453 VDD.n522 VDD.t125 17.484
R1454 VDD.n554 VDD.t17 17.484
R1455 VDD.n603 VDD.t121 17.484
R1456 VDD.n643 VDD.t82 17.484
R1457 VDD.n675 VDD.t0 17.484
R1458 VDD.n974 VDD.t23 16.516
R1459 VDD.n827 VDD.t101 16.516
R1460 VDD.n730 VDD.t8 13.669
R1461 VDD.n966 VDD.t35 13.099
R1462 VDD.n819 VDD.t152 13.099
R1463 VDD.t102 VDD.n477 12.627
R1464 VDD.n207 VDD.t3 12.391
R1465 VDD.n240 VDD.t119 12.391
R1466 VDD.n309 VDD.t26 12.391
R1467 VDD.n99 VDD.t76 12.391
R1468 VDD.n52 VDD.t123 12.391
R1469 VDD.n6 VDD.t65 12.391
R1470 VDD.n748 VDD.t127 11.656
R1471 VDD.n362 VDD.t20 11.656
R1472 VDD.n398 VDD.t160 11.656
R1473 VDD.n486 VDD.t84 11.656
R1474 VDD.n544 VDD.t57 11.656
R1475 VDD.n580 VDD.t92 11.656
R1476 VDD.n667 VDD.t109 11.656
R1477 VDD.n724 VDD.n721 11.52
R1478 VDD.n773 VDD.n770 11.52
R1479 VDD.n217 VDD.n214 11.52
R1480 VDD.n264 VDD.n261 11.52
R1481 VDD.n319 VDD.n316 11.52
R1482 VDD.n374 VDD.n371 11.52
R1483 VDD.n423 VDD.n420 11.52
R1484 VDD.n498 VDD.n495 11.52
R1485 VDD.n556 VDD.n553 11.52
R1486 VDD.n605 VDD.n602 11.52
R1487 VDD.n677 VDD.n674 11.52
R1488 VDD.n885 VDD.n882 11.52
R1489 VDD.n922 VDD.n919 11.52
R1490 VDD.n166 VDD.n163 11.52
R1491 VDD.n1026 VDD.n1025 11.52
R1492 VDD.n122 VDD.n119 11.52
R1493 VDD.n76 VDD.n73 11.52
R1494 VDD.n29 VDD.n26 11.52
R1495 VDD.n841 VDD.n838 11.52
R1496 VDD.n951 VDD.n948 11.52
R1497 VDD.n988 VDD.n985 11.52
R1498 VDD.n946 VDD.t144 10.251
R1499 VDD.n797 VDD.t18 10.251
R1500 VDD.n722 VDD.t74 10.251
R1501 VDD.n661 VDD.t108 9.637
R1502 VDD.n698 VDD.n697 8.855
R1503 VDD.n745 VDD.n744 8.855
R1504 VDD.n184 VDD.n183 8.855
R1505 VDD.n238 VDD.n237 8.855
R1506 VDD.n285 VDD.n284 8.855
R1507 VDD.n289 VDD.n288 8.855
R1508 VDD.n288 VDD.n287 8.855
R1509 VDD.n294 VDD.n293 8.855
R1510 VDD.n293 VDD.n292 8.855
R1511 VDD.n298 VDD.n297 8.855
R1512 VDD.n297 VDD.n296 8.855
R1513 VDD.n302 VDD.n301 8.855
R1514 VDD.n301 VDD.n300 8.855
R1515 VDD.n306 VDD.n305 8.855
R1516 VDD.n305 VDD.n304 8.855
R1517 VDD.n311 VDD.n310 8.855
R1518 VDD.n310 VDD.n309 8.855
R1519 VDD.n316 VDD.n315 8.855
R1520 VDD.n315 VDD.n314 8.855
R1521 VDD.n319 VDD.n318 8.855
R1522 VDD.n318 VDD.n317 8.855
R1523 VDD.n323 VDD.n322 8.855
R1524 VDD.n322 VDD.n321 8.855
R1525 VDD.n328 VDD.n327 8.855
R1526 VDD.n327 VDD.n326 8.855
R1527 VDD.n332 VDD.n331 8.855
R1528 VDD.n242 VDD.n241 8.855
R1529 VDD.n241 VDD.n240 8.855
R1530 VDD.n247 VDD.n246 8.855
R1531 VDD.n246 VDD.n245 8.855
R1532 VDD.n251 VDD.n250 8.855
R1533 VDD.n250 VDD.n249 8.855
R1534 VDD.n255 VDD.n254 8.855
R1535 VDD.n254 VDD.n253 8.855
R1536 VDD.n261 VDD.n260 8.855
R1537 VDD.n260 VDD.n259 8.855
R1538 VDD.n264 VDD.n263 8.855
R1539 VDD.n263 VDD.n262 8.855
R1540 VDD.n268 VDD.n267 8.855
R1541 VDD.n267 VDD.n266 8.855
R1542 VDD.n272 VDD.n271 8.855
R1543 VDD.n271 VDD.n270 8.855
R1544 VDD.n276 VDD.n275 8.855
R1545 VDD.n188 VDD.n187 8.855
R1546 VDD.n187 VDD.n186 8.855
R1547 VDD.n193 VDD.n192 8.855
R1548 VDD.n192 VDD.n191 8.855
R1549 VDD.n197 VDD.n196 8.855
R1550 VDD.n196 VDD.n195 8.855
R1551 VDD.n201 VDD.n200 8.855
R1552 VDD.n200 VDD.n199 8.855
R1553 VDD.n205 VDD.n204 8.855
R1554 VDD.n204 VDD.n203 8.855
R1555 VDD.n209 VDD.n208 8.855
R1556 VDD.n208 VDD.n207 8.855
R1557 VDD.n214 VDD.n213 8.855
R1558 VDD.n213 VDD.n212 8.855
R1559 VDD.n217 VDD.n216 8.855
R1560 VDD.n216 VDD.n215 8.855
R1561 VDD.n221 VDD.n220 8.855
R1562 VDD.n220 VDD.n219 8.855
R1563 VDD.n225 VDD.n224 8.855
R1564 VDD.n224 VDD.n223 8.855
R1565 VDD.n229 VDD.n228 8.855
R1566 VDD.n338 VDD.n337 8.855
R1567 VDD.n395 VDD.n394 8.855
R1568 VDD.n447 VDD.n446 8.855
R1569 VDD.n446 VDD.n445 8.855
R1570 VDD.n451 VDD.n450 8.855
R1571 VDD.n450 VDD.n449 8.855
R1572 VDD.n456 VDD.n455 8.855
R1573 VDD.n455 VDD.n454 8.855
R1574 VDD.n461 VDD.n460 8.855
R1575 VDD.n460 VDD.n459 8.855
R1576 VDD.n465 VDD.n464 8.855
R1577 VDD.n464 VDD.n463 8.855
R1578 VDD.n469 VDD.n468 8.855
R1579 VDD.n468 VDD.n467 8.855
R1580 VDD.n474 VDD.n473 8.855
R1581 VDD.n473 VDD.n472 8.855
R1582 VDD.n480 VDD.n479 8.855
R1583 VDD.n479 VDD.n478 8.855
R1584 VDD.n484 VDD.n483 8.855
R1585 VDD.n483 VDD.n482 8.855
R1586 VDD.n488 VDD.n487 8.855
R1587 VDD.n487 VDD.n486 8.855
R1588 VDD.n495 VDD.n494 8.855
R1589 VDD.n494 VDD.n493 8.855
R1590 VDD.n498 VDD.n497 8.855
R1591 VDD.n497 VDD.n496 8.855
R1592 VDD.n502 VDD.n501 8.855
R1593 VDD.n501 VDD.n500 8.855
R1594 VDD.n506 VDD.n505 8.855
R1595 VDD.n505 VDD.n504 8.855
R1596 VDD.n511 VDD.n510 8.855
R1597 VDD.n443 VDD.n442 8.855
R1598 VDD.n442 VDD.n441 8.855
R1599 VDD.n400 VDD.n399 8.855
R1600 VDD.n399 VDD.n398 8.855
R1601 VDD.n405 VDD.n404 8.855
R1602 VDD.n404 VDD.n403 8.855
R1603 VDD.n409 VDD.n408 8.855
R1604 VDD.n408 VDD.n407 8.855
R1605 VDD.n414 VDD.n413 8.855
R1606 VDD.n413 VDD.n412 8.855
R1607 VDD.n420 VDD.n419 8.855
R1608 VDD.n419 VDD.n418 8.855
R1609 VDD.n423 VDD.n422 8.855
R1610 VDD.n422 VDD.n421 8.855
R1611 VDD.n427 VDD.n426 8.855
R1612 VDD.n426 VDD.n425 8.855
R1613 VDD.n431 VDD.n430 8.855
R1614 VDD.n430 VDD.n429 8.855
R1615 VDD.n436 VDD.n435 8.855
R1616 VDD.n342 VDD.n341 8.855
R1617 VDD.n341 VDD.n340 8.855
R1618 VDD.n347 VDD.n346 8.855
R1619 VDD.n346 VDD.n345 8.855
R1620 VDD.n351 VDD.n350 8.855
R1621 VDD.n350 VDD.n349 8.855
R1622 VDD.n356 VDD.n355 8.855
R1623 VDD.n355 VDD.n354 8.855
R1624 VDD.n360 VDD.n359 8.855
R1625 VDD.n359 VDD.n358 8.855
R1626 VDD.n364 VDD.n363 8.855
R1627 VDD.n363 VDD.n362 8.855
R1628 VDD.n371 VDD.n370 8.855
R1629 VDD.n370 VDD.n369 8.855
R1630 VDD.n374 VDD.n373 8.855
R1631 VDD.n373 VDD.n372 8.855
R1632 VDD.n378 VDD.n377 8.855
R1633 VDD.n377 VDD.n376 8.855
R1634 VDD.n382 VDD.n381 8.855
R1635 VDD.n381 VDD.n380 8.855
R1636 VDD.n386 VDD.n385 8.855
R1637 VDD.n520 VDD.n519 8.855
R1638 VDD.n577 VDD.n576 8.855
R1639 VDD.n629 VDD.n628 8.855
R1640 VDD.n877 VDD.n876 8.855
R1641 VDD.n882 VDD.n881 8.855
R1642 VDD.n881 VDD.n880 8.855
R1643 VDD.n885 VDD.n884 8.855
R1644 VDD.n884 VDD.n883 8.855
R1645 VDD.n889 VDD.n888 8.855
R1646 VDD.n888 VDD.n887 8.855
R1647 VDD.n893 VDD.n892 8.855
R1648 VDD.n892 VDD.n891 8.855
R1649 VDD.n897 VDD.n896 8.855
R1650 VDD.n896 VDD.n895 8.855
R1651 VDD.n902 VDD.n901 8.855
R1652 VDD.n901 VDD.n900 8.855
R1653 VDD.n906 VDD.n905 8.855
R1654 VDD.n905 VDD.n904 8.855
R1655 VDD.n910 VDD.n909 8.855
R1656 VDD.n909 VDD.n908 8.855
R1657 VDD.n914 VDD.n913 8.855
R1658 VDD.n913 VDD.n912 8.855
R1659 VDD.n919 VDD.n918 8.855
R1660 VDD.n918 VDD.n917 8.855
R1661 VDD.n922 VDD.n921 8.855
R1662 VDD.n921 VDD.n920 8.855
R1663 VDD.n926 VDD.n925 8.855
R1664 VDD.n925 VDD.n924 8.855
R1665 VDD.n930 VDD.n929 8.855
R1666 VDD.n929 VDD.n928 8.855
R1667 VDD.n935 VDD.n934 8.855
R1668 VDD.n632 VDD.n631 8.855
R1669 VDD.n637 VDD.n636 8.855
R1670 VDD.n636 VDD.n635 8.855
R1671 VDD.n641 VDD.n640 8.855
R1672 VDD.n640 VDD.n639 8.855
R1673 VDD.n645 VDD.n644 8.855
R1674 VDD.n644 VDD.n643 8.855
R1675 VDD.n650 VDD.n649 8.855
R1676 VDD.n649 VDD.n648 8.855
R1677 VDD.n655 VDD.n654 8.855
R1678 VDD.n654 VDD.n653 8.855
R1679 VDD.n659 VDD.n658 8.855
R1680 VDD.n658 VDD.n657 8.855
R1681 VDD.n664 VDD.n663 8.855
R1682 VDD.n663 VDD.n662 8.855
R1683 VDD.n669 VDD.n668 8.855
R1684 VDD.n668 VDD.n667 8.855
R1685 VDD.n674 VDD.n673 8.855
R1686 VDD.n673 VDD.n672 8.855
R1687 VDD.n677 VDD.n676 8.855
R1688 VDD.n676 VDD.n675 8.855
R1689 VDD.n681 VDD.n680 8.855
R1690 VDD.n680 VDD.n679 8.855
R1691 VDD.n686 VDD.n685 8.855
R1692 VDD.n685 VDD.n684 8.855
R1693 VDD.n691 VDD.n690 8.855
R1694 VDD.n582 VDD.n581 8.855
R1695 VDD.n581 VDD.n580 8.855
R1696 VDD.n587 VDD.n586 8.855
R1697 VDD.n586 VDD.n585 8.855
R1698 VDD.n591 VDD.n590 8.855
R1699 VDD.n590 VDD.n589 8.855
R1700 VDD.n596 VDD.n595 8.855
R1701 VDD.n595 VDD.n594 8.855
R1702 VDD.n602 VDD.n601 8.855
R1703 VDD.n601 VDD.n600 8.855
R1704 VDD.n605 VDD.n604 8.855
R1705 VDD.n604 VDD.n603 8.855
R1706 VDD.n609 VDD.n608 8.855
R1707 VDD.n608 VDD.n607 8.855
R1708 VDD.n613 VDD.n612 8.855
R1709 VDD.n612 VDD.n611 8.855
R1710 VDD.n618 VDD.n617 8.855
R1711 VDD.n524 VDD.n523 8.855
R1712 VDD.n523 VDD.n522 8.855
R1713 VDD.n529 VDD.n528 8.855
R1714 VDD.n528 VDD.n527 8.855
R1715 VDD.n533 VDD.n532 8.855
R1716 VDD.n532 VDD.n531 8.855
R1717 VDD.n538 VDD.n537 8.855
R1718 VDD.n537 VDD.n536 8.855
R1719 VDD.n542 VDD.n541 8.855
R1720 VDD.n541 VDD.n540 8.855
R1721 VDD.n546 VDD.n545 8.855
R1722 VDD.n545 VDD.n544 8.855
R1723 VDD.n553 VDD.n552 8.855
R1724 VDD.n552 VDD.n551 8.855
R1725 VDD.n556 VDD.n555 8.855
R1726 VDD.n555 VDD.n554 8.855
R1727 VDD.n560 VDD.n559 8.855
R1728 VDD.n559 VDD.n558 8.855
R1729 VDD.n564 VDD.n563 8.855
R1730 VDD.n563 VDD.n562 8.855
R1731 VDD.n568 VDD.n567 8.855
R1732 VDD.n4 VDD.n3 8.855
R1733 VDD.n8 VDD.n7 8.855
R1734 VDD.n7 VDD.n6 8.855
R1735 VDD.n13 VDD.n12 8.855
R1736 VDD.n12 VDD.n11 8.855
R1737 VDD.n17 VDD.n16 8.855
R1738 VDD.n16 VDD.n15 8.855
R1739 VDD.n21 VDD.n20 8.855
R1740 VDD.n20 VDD.n19 8.855
R1741 VDD.n26 VDD.n25 8.855
R1742 VDD.n25 VDD.n24 8.855
R1743 VDD.n29 VDD.n28 8.855
R1744 VDD.n28 VDD.n27 8.855
R1745 VDD.n33 VDD.n32 8.855
R1746 VDD.n32 VDD.n31 8.855
R1747 VDD.n37 VDD.n36 8.855
R1748 VDD.n36 VDD.n35 8.855
R1749 VDD.n41 VDD.n40 8.855
R1750 VDD.n50 VDD.n49 8.855
R1751 VDD.n54 VDD.n53 8.855
R1752 VDD.n53 VDD.n52 8.855
R1753 VDD.n59 VDD.n58 8.855
R1754 VDD.n58 VDD.n57 8.855
R1755 VDD.n63 VDD.n62 8.855
R1756 VDD.n62 VDD.n61 8.855
R1757 VDD.n67 VDD.n66 8.855
R1758 VDD.n66 VDD.n65 8.855
R1759 VDD.n73 VDD.n72 8.855
R1760 VDD.n72 VDD.n71 8.855
R1761 VDD.n76 VDD.n75 8.855
R1762 VDD.n75 VDD.n74 8.855
R1763 VDD.n80 VDD.n79 8.855
R1764 VDD.n79 VDD.n78 8.855
R1765 VDD.n84 VDD.n83 8.855
R1766 VDD.n83 VDD.n82 8.855
R1767 VDD.n88 VDD.n87 8.855
R1768 VDD.n97 VDD.n96 8.855
R1769 VDD.n101 VDD.n100 8.855
R1770 VDD.n100 VDD.n99 8.855
R1771 VDD.n106 VDD.n105 8.855
R1772 VDD.n105 VDD.n104 8.855
R1773 VDD.n110 VDD.n109 8.855
R1774 VDD.n109 VDD.n108 8.855
R1775 VDD.n114 VDD.n113 8.855
R1776 VDD.n113 VDD.n112 8.855
R1777 VDD.n119 VDD.n118 8.855
R1778 VDD.n118 VDD.n117 8.855
R1779 VDD.n122 VDD.n121 8.855
R1780 VDD.n121 VDD.n120 8.855
R1781 VDD.n126 VDD.n125 8.855
R1782 VDD.n125 VDD.n124 8.855
R1783 VDD.n130 VDD.n129 8.855
R1784 VDD.n129 VDD.n128 8.855
R1785 VDD.n134 VDD.n133 8.855
R1786 VDD.n143 VDD.n142 8.855
R1787 VDD.n148 VDD.n147 8.855
R1788 VDD.n147 VDD.n146 8.855
R1789 VDD.n152 VDD.n151 8.855
R1790 VDD.n151 VDD.n150 8.855
R1791 VDD.n156 VDD.n155 8.855
R1792 VDD.n155 VDD.n154 8.855
R1793 VDD.n160 VDD.n159 8.855
R1794 VDD.n159 VDD.n158 8.855
R1795 VDD.n163 VDD.n1 8.855
R1796 VDD.n1 VDD.n0 8.855
R1797 VDD.n166 VDD.n165 8.855
R1798 VDD.n165 VDD.n164 8.855
R1799 VDD.n170 VDD.n169 8.855
R1800 VDD.n169 VDD.n168 8.855
R1801 VDD.n174 VDD.n173 8.855
R1802 VDD.n173 VDD.n172 8.855
R1803 VDD.n179 VDD.n178 8.855
R1804 VDD.n750 VDD.n749 8.855
R1805 VDD.n749 VDD.n748 8.855
R1806 VDD.n755 VDD.n754 8.855
R1807 VDD.n754 VDD.n753 8.855
R1808 VDD.n759 VDD.n758 8.855
R1809 VDD.n758 VDD.n757 8.855
R1810 VDD.n764 VDD.n763 8.855
R1811 VDD.n763 VDD.n762 8.855
R1812 VDD.n770 VDD.n769 8.855
R1813 VDD.n769 VDD.n768 8.855
R1814 VDD.n773 VDD.n772 8.855
R1815 VDD.n772 VDD.n771 8.855
R1816 VDD.n777 VDD.n776 8.855
R1817 VDD.n776 VDD.n775 8.855
R1818 VDD.n781 VDD.n780 8.855
R1819 VDD.n780 VDD.n779 8.855
R1820 VDD.n786 VDD.n785 8.855
R1821 VDD.n702 VDD.n701 8.855
R1822 VDD.n701 VDD.n700 8.855
R1823 VDD.n707 VDD.n706 8.855
R1824 VDD.n706 VDD.n705 8.855
R1825 VDD.n711 VDD.n710 8.855
R1826 VDD.n710 VDD.n709 8.855
R1827 VDD.n715 VDD.n714 8.855
R1828 VDD.n714 VDD.n713 8.855
R1829 VDD.n721 VDD.n720 8.855
R1830 VDD.n720 VDD.n719 8.855
R1831 VDD.n724 VDD.n723 8.855
R1832 VDD.n723 VDD.n722 8.855
R1833 VDD.n728 VDD.n727 8.855
R1834 VDD.n727 VDD.n726 8.855
R1835 VDD.n732 VDD.n731 8.855
R1836 VDD.n731 VDD.n730 8.855
R1837 VDD.n736 VDD.n735 8.855
R1838 VDD.n795 VDD.n794 8.855
R1839 VDD.n799 VDD.n798 8.855
R1840 VDD.n798 VDD.n797 8.855
R1841 VDD.n804 VDD.n803 8.855
R1842 VDD.n803 VDD.n802 8.855
R1843 VDD.n808 VDD.n807 8.855
R1844 VDD.n807 VDD.n806 8.855
R1845 VDD.n812 VDD.n811 8.855
R1846 VDD.n811 VDD.n810 8.855
R1847 VDD.n816 VDD.n815 8.855
R1848 VDD.n815 VDD.n814 8.855
R1849 VDD.n821 VDD.n820 8.855
R1850 VDD.n820 VDD.n819 8.855
R1851 VDD.n825 VDD.n824 8.855
R1852 VDD.n824 VDD.n823 8.855
R1853 VDD.n829 VDD.n828 8.855
R1854 VDD.n828 VDD.n827 8.855
R1855 VDD.n833 VDD.n832 8.855
R1856 VDD.n832 VDD.n831 8.855
R1857 VDD.n838 VDD.n837 8.855
R1858 VDD.n837 VDD.n836 8.855
R1859 VDD.n841 VDD.n840 8.855
R1860 VDD.n840 VDD.n839 8.855
R1861 VDD.n845 VDD.n844 8.855
R1862 VDD.n844 VDD.n843 8.855
R1863 VDD.n849 VDD.n848 8.855
R1864 VDD.n848 VDD.n847 8.855
R1865 VDD.n854 VDD.n853 8.855
R1866 VDD.n943 VDD.n942 8.855
R1867 VDD.n948 VDD.n947 8.855
R1868 VDD.n947 VDD.n946 8.855
R1869 VDD.n951 VDD.n950 8.855
R1870 VDD.n950 VDD.n949 8.855
R1871 VDD.n955 VDD.n954 8.855
R1872 VDD.n954 VDD.n953 8.855
R1873 VDD.n959 VDD.n958 8.855
R1874 VDD.n958 VDD.n957 8.855
R1875 VDD.n963 VDD.n962 8.855
R1876 VDD.n962 VDD.n961 8.855
R1877 VDD.n968 VDD.n967 8.855
R1878 VDD.n967 VDD.n966 8.855
R1879 VDD.n972 VDD.n971 8.855
R1880 VDD.n971 VDD.n970 8.855
R1881 VDD.n976 VDD.n975 8.855
R1882 VDD.n975 VDD.n974 8.855
R1883 VDD.n980 VDD.n979 8.855
R1884 VDD.n979 VDD.n978 8.855
R1885 VDD.n985 VDD.n984 8.855
R1886 VDD.n984 VDD.n983 8.855
R1887 VDD.n988 VDD.n987 8.855
R1888 VDD.n987 VDD.n986 8.855
R1889 VDD.n992 VDD.n991 8.855
R1890 VDD.n991 VDD.n990 8.855
R1891 VDD.n996 VDD.n995 8.855
R1892 VDD.n995 VDD.n994 8.855
R1893 VDD.n1001 VDD.n1000 8.855
R1894 VDD.n865 VDD.n864 8.855
R1895 VDD.n869 VDD.n868 8.855
R1896 VDD.n868 VDD.n867 8.855
R1897 VDD.n1059 VDD.n1058 8.855
R1898 VDD.n1058 VDD.n1057 8.855
R1899 VDD.n1055 VDD.n1054 8.855
R1900 VDD.n1054 VDD.n1053 8.855
R1901 VDD.n1051 VDD.n1050 8.855
R1902 VDD.n1050 VDD.n1049 8.855
R1903 VDD.n1047 VDD.n1046 8.855
R1904 VDD.n1046 VDD.n1045 8.855
R1905 VDD.n1042 VDD.n1041 8.855
R1906 VDD.n1041 VDD.n1040 8.855
R1907 VDD.n1038 VDD.n1037 8.855
R1908 VDD.n1037 VDD.n1036 8.855
R1909 VDD.n1034 VDD.n1033 8.855
R1910 VDD.n1033 VDD.n1032 8.855
R1911 VDD.n1030 VDD.n1029 8.855
R1912 VDD.n1029 VDD.n1028 8.855
R1913 VDD.n1026 VDD.n872 8.855
R1914 VDD.n872 VDD.n871 8.855
R1915 VDD.n1025 VDD.n1024 8.855
R1916 VDD.n1024 VDD.n1023 8.855
R1917 VDD.n1020 VDD.n1019 8.855
R1918 VDD.n1019 VDD.n1018 8.855
R1919 VDD.n1016 VDD.n1015 8.855
R1920 VDD.n1015 VDD.n1014 8.855
R1921 VDD.n1011 VDD.n1010 8.855
R1922 VDD.n628 VDD.n627 7.349
R1923 VDD.n700 VDD.t4 6.834
R1924 VDD.n478 VDD.t102 5.828
R1925 VDD.n794 VDD.n793 5.273
R1926 VDD.n697 VDD.n696 5.273
R1927 VDD.n735 VDD.n734 5.273
R1928 VDD.n853 VDD.n852 5.273
R1929 VDD.n1000 VDD.n999 5.273
R1930 VDD.n942 VDD.n941 5.273
R1931 VDD.n516 VDD.n335 4.91
R1932 VDD.n1005 VDD.n938 4.91
R1933 VDD.n695 VDD.n516 4.775
R1934 VDD.n859 VDD.n858 4.775
R1935 VDD.n858 VDD.n695 4.775
R1936 VDD.n1006 VDD.n1005 4.775
R1937 VDD.n335 VDD.n334 4.65
R1938 VDD.n286 VDD.n285 4.65
R1939 VDD.n290 VDD.n289 4.65
R1940 VDD.n295 VDD.n294 4.65
R1941 VDD.n299 VDD.n298 4.65
R1942 VDD.n303 VDD.n302 4.65
R1943 VDD.n307 VDD.n306 4.65
R1944 VDD.n312 VDD.n311 4.65
R1945 VDD.n316 VDD.n313 4.65
R1946 VDD.n320 VDD.n319 4.65
R1947 VDD.n324 VDD.n323 4.65
R1948 VDD.n329 VDD.n328 4.65
R1949 VDD.n333 VDD.n332 4.65
R1950 VDD.n282 VDD.n281 4.65
R1951 VDD.n280 VDD.n279 4.65
R1952 VDD.n239 VDD.n238 4.65
R1953 VDD.n243 VDD.n242 4.65
R1954 VDD.n248 VDD.n247 4.65
R1955 VDD.n252 VDD.n251 4.65
R1956 VDD.n256 VDD.n255 4.65
R1957 VDD.n261 VDD.n258 4.65
R1958 VDD.n265 VDD.n264 4.65
R1959 VDD.n269 VDD.n268 4.65
R1960 VDD.n273 VDD.n272 4.65
R1961 VDD.n277 VDD.n276 4.65
R1962 VDD.n235 VDD.n234 4.65
R1963 VDD.n233 VDD.n232 4.65
R1964 VDD.n189 VDD.n188 4.65
R1965 VDD.n194 VDD.n193 4.65
R1966 VDD.n198 VDD.n197 4.65
R1967 VDD.n202 VDD.n201 4.65
R1968 VDD.n206 VDD.n205 4.65
R1969 VDD.n210 VDD.n209 4.65
R1970 VDD.n214 VDD.n211 4.65
R1971 VDD.n218 VDD.n217 4.65
R1972 VDD.n222 VDD.n221 4.65
R1973 VDD.n226 VDD.n225 4.65
R1974 VDD.n230 VDD.n229 4.65
R1975 VDD.n515 VDD.n514 4.65
R1976 VDD.n448 VDD.n447 4.65
R1977 VDD.n452 VDD.n451 4.65
R1978 VDD.n457 VDD.n456 4.65
R1979 VDD.n462 VDD.n461 4.65
R1980 VDD.n466 VDD.n465 4.65
R1981 VDD.n470 VDD.n469 4.65
R1982 VDD.n475 VDD.n474 4.65
R1983 VDD.n481 VDD.n480 4.65
R1984 VDD.n485 VDD.n484 4.65
R1985 VDD.n489 VDD.n488 4.65
R1986 VDD.n495 VDD.n492 4.65
R1987 VDD.n499 VDD.n498 4.65
R1988 VDD.n503 VDD.n502 4.65
R1989 VDD.n507 VDD.n506 4.65
R1990 VDD.n512 VDD.n511 4.65
R1991 VDD.n444 VDD.n443 4.65
R1992 VDD.n440 VDD.n439 4.65
R1993 VDD.n396 VDD.n395 4.65
R1994 VDD.n401 VDD.n400 4.65
R1995 VDD.n406 VDD.n405 4.65
R1996 VDD.n410 VDD.n409 4.65
R1997 VDD.n415 VDD.n414 4.65
R1998 VDD.n420 VDD.n417 4.65
R1999 VDD.n424 VDD.n423 4.65
R2000 VDD.n428 VDD.n427 4.65
R2001 VDD.n432 VDD.n431 4.65
R2002 VDD.n437 VDD.n436 4.65
R2003 VDD.n392 VDD.n391 4.65
R2004 VDD.n390 VDD.n389 4.65
R2005 VDD.n343 VDD.n342 4.65
R2006 VDD.n348 VDD.n347 4.65
R2007 VDD.n352 VDD.n351 4.65
R2008 VDD.n357 VDD.n356 4.65
R2009 VDD.n361 VDD.n360 4.65
R2010 VDD.n365 VDD.n364 4.65
R2011 VDD.n371 VDD.n367 4.65
R2012 VDD.n375 VDD.n374 4.65
R2013 VDD.n379 VDD.n378 4.65
R2014 VDD.n383 VDD.n382 4.65
R2015 VDD.n387 VDD.n386 4.65
R2016 VDD.n882 VDD.n879 4.65
R2017 VDD.n886 VDD.n885 4.65
R2018 VDD.n890 VDD.n889 4.65
R2019 VDD.n894 VDD.n893 4.65
R2020 VDD.n898 VDD.n897 4.65
R2021 VDD.n903 VDD.n902 4.65
R2022 VDD.n907 VDD.n906 4.65
R2023 VDD.n911 VDD.n910 4.65
R2024 VDD.n915 VDD.n914 4.65
R2025 VDD.n919 VDD.n916 4.65
R2026 VDD.n923 VDD.n922 4.65
R2027 VDD.n927 VDD.n926 4.65
R2028 VDD.n931 VDD.n930 4.65
R2029 VDD.n936 VDD.n935 4.65
R2030 VDD.n938 VDD.n937 4.65
R2031 VDD.n694 VDD.n693 4.65
R2032 VDD.n630 VDD.n629 4.65
R2033 VDD.n633 VDD.n632 4.65
R2034 VDD.n638 VDD.n637 4.65
R2035 VDD.n642 VDD.n641 4.65
R2036 VDD.n646 VDD.n645 4.65
R2037 VDD.n651 VDD.n650 4.65
R2038 VDD.n656 VDD.n655 4.65
R2039 VDD.n660 VDD.n659 4.65
R2040 VDD.n665 VDD.n664 4.65
R2041 VDD.n670 VDD.n669 4.65
R2042 VDD.n674 VDD.n671 4.65
R2043 VDD.n678 VDD.n677 4.65
R2044 VDD.n682 VDD.n681 4.65
R2045 VDD.n687 VDD.n686 4.65
R2046 VDD.n692 VDD.n691 4.65
R2047 VDD.n624 VDD.n623 4.65
R2048 VDD.n622 VDD.n621 4.65
R2049 VDD.n578 VDD.n577 4.65
R2050 VDD.n583 VDD.n582 4.65
R2051 VDD.n588 VDD.n587 4.65
R2052 VDD.n592 VDD.n591 4.65
R2053 VDD.n597 VDD.n596 4.65
R2054 VDD.n602 VDD.n599 4.65
R2055 VDD.n606 VDD.n605 4.65
R2056 VDD.n610 VDD.n609 4.65
R2057 VDD.n614 VDD.n613 4.65
R2058 VDD.n619 VDD.n618 4.65
R2059 VDD.n574 VDD.n573 4.65
R2060 VDD.n572 VDD.n571 4.65
R2061 VDD.n525 VDD.n524 4.65
R2062 VDD.n530 VDD.n529 4.65
R2063 VDD.n534 VDD.n533 4.65
R2064 VDD.n539 VDD.n538 4.65
R2065 VDD.n543 VDD.n542 4.65
R2066 VDD.n547 VDD.n546 4.65
R2067 VDD.n553 VDD.n549 4.65
R2068 VDD.n557 VDD.n556 4.65
R2069 VDD.n561 VDD.n560 4.65
R2070 VDD.n565 VDD.n564 4.65
R2071 VDD.n569 VDD.n568 4.65
R2072 VDD.n9 VDD.n8 4.65
R2073 VDD.n14 VDD.n13 4.65
R2074 VDD.n18 VDD.n17 4.65
R2075 VDD.n22 VDD.n21 4.65
R2076 VDD.n26 VDD.n23 4.65
R2077 VDD.n30 VDD.n29 4.65
R2078 VDD.n34 VDD.n33 4.65
R2079 VDD.n38 VDD.n37 4.65
R2080 VDD.n42 VDD.n41 4.65
R2081 VDD.n45 VDD.n44 4.65
R2082 VDD.n47 VDD.n46 4.65
R2083 VDD.n51 VDD.n50 4.65
R2084 VDD.n55 VDD.n54 4.65
R2085 VDD.n60 VDD.n59 4.65
R2086 VDD.n64 VDD.n63 4.65
R2087 VDD.n68 VDD.n67 4.65
R2088 VDD.n73 VDD.n70 4.65
R2089 VDD.n77 VDD.n76 4.65
R2090 VDD.n81 VDD.n80 4.65
R2091 VDD.n85 VDD.n84 4.65
R2092 VDD.n89 VDD.n88 4.65
R2093 VDD.n92 VDD.n91 4.65
R2094 VDD.n94 VDD.n93 4.65
R2095 VDD.n98 VDD.n97 4.65
R2096 VDD.n102 VDD.n101 4.65
R2097 VDD.n107 VDD.n106 4.65
R2098 VDD.n111 VDD.n110 4.65
R2099 VDD.n115 VDD.n114 4.65
R2100 VDD.n119 VDD.n116 4.65
R2101 VDD.n123 VDD.n122 4.65
R2102 VDD.n127 VDD.n126 4.65
R2103 VDD.n131 VDD.n130 4.65
R2104 VDD.n135 VDD.n134 4.65
R2105 VDD.n138 VDD.n137 4.65
R2106 VDD.n140 VDD.n139 4.65
R2107 VDD.n144 VDD.n143 4.65
R2108 VDD.n149 VDD.n148 4.65
R2109 VDD.n153 VDD.n152 4.65
R2110 VDD.n157 VDD.n156 4.65
R2111 VDD.n161 VDD.n160 4.65
R2112 VDD.n163 VDD.n162 4.65
R2113 VDD.n167 VDD.n166 4.65
R2114 VDD.n171 VDD.n170 4.65
R2115 VDD.n175 VDD.n174 4.65
R2116 VDD.n180 VDD.n179 4.65
R2117 VDD.n861 VDD.n860 4.65
R2118 VDD.n790 VDD.n789 4.65
R2119 VDD.n746 VDD.n745 4.65
R2120 VDD.n751 VDD.n750 4.65
R2121 VDD.n756 VDD.n755 4.65
R2122 VDD.n760 VDD.n759 4.65
R2123 VDD.n765 VDD.n764 4.65
R2124 VDD.n770 VDD.n767 4.65
R2125 VDD.n774 VDD.n773 4.65
R2126 VDD.n778 VDD.n777 4.65
R2127 VDD.n782 VDD.n781 4.65
R2128 VDD.n787 VDD.n786 4.65
R2129 VDD.n742 VDD.n741 4.65
R2130 VDD.n740 VDD.n739 4.65
R2131 VDD.n703 VDD.n702 4.65
R2132 VDD.n708 VDD.n707 4.65
R2133 VDD.n712 VDD.n711 4.65
R2134 VDD.n716 VDD.n715 4.65
R2135 VDD.n721 VDD.n718 4.65
R2136 VDD.n725 VDD.n724 4.65
R2137 VDD.n729 VDD.n728 4.65
R2138 VDD.n733 VDD.n732 4.65
R2139 VDD.n737 VDD.n736 4.65
R2140 VDD.n857 VDD.n856 4.65
R2141 VDD.n792 VDD.n791 4.65
R2142 VDD.n796 VDD.n795 4.65
R2143 VDD.n800 VDD.n799 4.65
R2144 VDD.n805 VDD.n804 4.65
R2145 VDD.n809 VDD.n808 4.65
R2146 VDD.n813 VDD.n812 4.65
R2147 VDD.n817 VDD.n816 4.65
R2148 VDD.n822 VDD.n821 4.65
R2149 VDD.n826 VDD.n825 4.65
R2150 VDD.n830 VDD.n829 4.65
R2151 VDD.n834 VDD.n833 4.65
R2152 VDD.n838 VDD.n835 4.65
R2153 VDD.n842 VDD.n841 4.65
R2154 VDD.n846 VDD.n845 4.65
R2155 VDD.n850 VDD.n849 4.65
R2156 VDD.n855 VDD.n854 4.65
R2157 VDD.n948 VDD.n945 4.65
R2158 VDD.n952 VDD.n951 4.65
R2159 VDD.n956 VDD.n955 4.65
R2160 VDD.n960 VDD.n959 4.65
R2161 VDD.n964 VDD.n963 4.65
R2162 VDD.n969 VDD.n968 4.65
R2163 VDD.n973 VDD.n972 4.65
R2164 VDD.n977 VDD.n976 4.65
R2165 VDD.n981 VDD.n980 4.65
R2166 VDD.n985 VDD.n982 4.65
R2167 VDD.n989 VDD.n988 4.65
R2168 VDD.n993 VDD.n992 4.65
R2169 VDD.n997 VDD.n996 4.65
R2170 VDD.n1002 VDD.n1001 4.65
R2171 VDD.n1004 VDD.n1003 4.65
R2172 VDD.n870 VDD.n869 4.65
R2173 VDD.n1060 VDD.n1059 4.65
R2174 VDD.n1056 VDD.n1055 4.65
R2175 VDD.n1052 VDD.n1051 4.65
R2176 VDD.n1048 VDD.n1047 4.65
R2177 VDD.n1043 VDD.n1042 4.65
R2178 VDD.n1039 VDD.n1038 4.65
R2179 VDD.n1035 VDD.n1034 4.65
R2180 VDD.n1031 VDD.n1030 4.65
R2181 VDD.n1027 VDD.n1026 4.65
R2182 VDD.n1025 VDD.n1022 4.65
R2183 VDD.n1021 VDD.n1020 4.65
R2184 VDD.n1017 VDD.n1016 4.65
R2185 VDD.n1012 VDD.n1011 4.65
R2186 VDD.n1008 VDD.n1007 4.65
R2187 VDD.n744 VDD.n743 4.396
R2188 VDD.n394 VDD.n393 4.396
R2189 VDD.n510 VDD.n509 4.396
R2190 VDD.n435 VDD.n434 4.396
R2191 VDD.n385 VDD.n384 4.396
R2192 VDD.n576 VDD.n575 4.396
R2193 VDD.n690 VDD.n689 4.396
R2194 VDD.n617 VDD.n616 4.396
R2195 VDD.n567 VDD.n566 4.396
R2196 VDD.n785 VDD.n784 4.396
R2197 VDD.n876 VDD.n875 4.288
R2198 VDD.n3 VDD.n2 4.288
R2199 VDD.n49 VDD.n48 4.288
R2200 VDD.n96 VDD.n95 4.288
R2201 VDD.n178 VDD.n177 4.288
R2202 VDD.n864 VDD.n863 4.288
R2203 VDD.n183 VDD.n182 4.288
R2204 VDD.n237 VDD.n236 4.288
R2205 VDD.n284 VDD.n283 4.288
R2206 VDD.n331 VDD.n330 4.288
R2207 VDD.n275 VDD.n274 4.288
R2208 VDD.n228 VDD.n227 4.288
R2209 VDD.n934 VDD.n933 4.288
R2210 VDD.n142 VDD.n141 4.288
R2211 VDD.n40 VDD.n39 4.288
R2212 VDD.n87 VDD.n86 4.288
R2213 VDD.n133 VDD.n132 4.288
R2214 VDD.n1010 VDD.n1009 4.288
R2215 VDD.n944 VDD.n940 2.613
R2216 VDD.n866 VDD.n862 2.613
R2217 VDD.n878 VDD.n874 2.612
R2218 VDD.n5 VDD.n4 2.562
R2219 VDD.n944 VDD.n943 2.562
R2220 VDD.n866 VDD.n865 2.562
R2221 VDD.n185 VDD.n184 2.562
R2222 VDD.n339 VDD.n338 2.562
R2223 VDD.n878 VDD.n877 2.562
R2224 VDD.n521 VDD.n520 2.562
R2225 VDD.n699 VDD.n698 2.562
R2226 VDD.n325 VDD.n181 2.329
R2227 VDD.n491 VDD.n490 2.329
R2228 VDD.n683 VDD.n517 2.329
R2229 VDD.n9 VDD.n5 1.145
R2230 VDD.n945 VDD.n944 1.145
R2231 VDD.n870 VDD.n866 1.145
R2232 VDD.n189 VDD.n185 1.145
R2233 VDD.n343 VDD.n339 1.145
R2234 VDD.n879 VDD.n878 1.145
R2235 VDD.n525 VDD.n521 1.145
R2236 VDD.n703 VDD.n699 1.145
R2237 VDD.n140 VDD.n138 0.957
R2238 VDD.n282 VDD.n280 0.777
R2239 VDD.n627 VDD.n626 0.754
R2240 VDD.n235 VDD.n233 0.525
R2241 VDD.n392 VDD.n390 0.525
R2242 VDD.n574 VDD.n572 0.525
R2243 VDD.n47 VDD.n45 0.525
R2244 VDD.n94 VDD.n92 0.525
R2245 VDD.n742 VDD.n740 0.525
R2246 VDD.n444 VDD.n440 0.507
R2247 VDD.n624 VDD.n622 0.507
R2248 VDD.n792 VDD.n790 0.507
R2249 VDD.n337 VDD.n336 0.227
R2250 VDD.n519 VDD.n518 0.227
R2251 VDD.n516 VDD.n515 0.135
R2252 VDD.n695 VDD.n694 0.135
R2253 VDD.n860 VDD.n859 0.135
R2254 VDD.n858 VDD.n857 0.135
R2255 VDD.n1005 VDD.n1004 0.135
R2256 VDD.n1008 VDD.n1006 0.135
R2257 VDD.n198 VDD.n194 0.09
R2258 VDD.n202 VDD.n198 0.09
R2259 VDD.n206 VDD.n202 0.09
R2260 VDD.n210 VDD.n206 0.09
R2261 VDD.n211 VDD.n210 0.09
R2262 VDD.n222 VDD.n218 0.09
R2263 VDD.n226 VDD.n222 0.09
R2264 VDD.n230 VDD.n226 0.09
R2265 VDD.n239 VDD.n235 0.09
R2266 VDD.n243 VDD.n239 0.09
R2267 VDD.n252 VDD.n248 0.09
R2268 VDD.n256 VDD.n252 0.09
R2269 VDD.n258 VDD.n256 0.09
R2270 VDD.n269 VDD.n265 0.09
R2271 VDD.n273 VDD.n269 0.09
R2272 VDD.n277 VDD.n273 0.09
R2273 VDD.n286 VDD.n282 0.09
R2274 VDD.n290 VDD.n286 0.09
R2275 VDD.n299 VDD.n295 0.09
R2276 VDD.n303 VDD.n299 0.09
R2277 VDD.n307 VDD.n303 0.09
R2278 VDD.n313 VDD.n312 0.09
R2279 VDD.n324 VDD.n320 0.09
R2280 VDD.n333 VDD.n329 0.09
R2281 VDD.n335 VDD.n333 0.09
R2282 VDD.n352 VDD.n348 0.09
R2283 VDD.n361 VDD.n357 0.09
R2284 VDD.n365 VDD.n361 0.09
R2285 VDD.n367 VDD.n365 0.09
R2286 VDD.n379 VDD.n375 0.09
R2287 VDD.n383 VDD.n379 0.09
R2288 VDD.n387 VDD.n383 0.09
R2289 VDD.n396 VDD.n392 0.09
R2290 VDD.n410 VDD.n406 0.09
R2291 VDD.n415 VDD.n410 0.09
R2292 VDD.n417 VDD.n415 0.09
R2293 VDD.n428 VDD.n424 0.09
R2294 VDD.n432 VDD.n428 0.09
R2295 VDD.n448 VDD.n444 0.09
R2296 VDD.n452 VDD.n448 0.09
R2297 VDD.n466 VDD.n462 0.09
R2298 VDD.n470 VDD.n466 0.09
R2299 VDD.n485 VDD.n481 0.09
R2300 VDD.n489 VDD.n485 0.09
R2301 VDD.n492 VDD.n489 0.09
R2302 VDD.n503 VDD.n499 0.09
R2303 VDD.n507 VDD.n503 0.09
R2304 VDD.n890 VDD.n886 0.09
R2305 VDD.n894 VDD.n890 0.09
R2306 VDD.n898 VDD.n894 0.09
R2307 VDD.n907 VDD.n903 0.09
R2308 VDD.n911 VDD.n907 0.09
R2309 VDD.n915 VDD.n911 0.09
R2310 VDD.n916 VDD.n915 0.09
R2311 VDD.n927 VDD.n923 0.09
R2312 VDD.n931 VDD.n927 0.09
R2313 VDD.n938 VDD.n936 0.09
R2314 VDD.n534 VDD.n530 0.09
R2315 VDD.n543 VDD.n539 0.09
R2316 VDD.n547 VDD.n543 0.09
R2317 VDD.n549 VDD.n547 0.09
R2318 VDD.n561 VDD.n557 0.09
R2319 VDD.n565 VDD.n561 0.09
R2320 VDD.n569 VDD.n565 0.09
R2321 VDD.n578 VDD.n574 0.09
R2322 VDD.n592 VDD.n588 0.09
R2323 VDD.n597 VDD.n592 0.09
R2324 VDD.n599 VDD.n597 0.09
R2325 VDD.n610 VDD.n606 0.09
R2326 VDD.n614 VDD.n610 0.09
R2327 VDD.n630 VDD.n624 0.09
R2328 VDD.n633 VDD.n630 0.09
R2329 VDD.n642 VDD.n638 0.09
R2330 VDD.n646 VDD.n642 0.09
R2331 VDD.n660 VDD.n656 0.09
R2332 VDD.n665 VDD.n660 0.09
R2333 VDD.n671 VDD.n670 0.09
R2334 VDD.n682 VDD.n678 0.09
R2335 VDD.n694 VDD.n692 0.09
R2336 VDD.n18 VDD.n14 0.09
R2337 VDD.n22 VDD.n18 0.09
R2338 VDD.n23 VDD.n22 0.09
R2339 VDD.n34 VDD.n30 0.09
R2340 VDD.n38 VDD.n34 0.09
R2341 VDD.n42 VDD.n38 0.09
R2342 VDD.n51 VDD.n47 0.09
R2343 VDD.n55 VDD.n51 0.09
R2344 VDD.n64 VDD.n60 0.09
R2345 VDD.n68 VDD.n64 0.09
R2346 VDD.n70 VDD.n68 0.09
R2347 VDD.n81 VDD.n77 0.09
R2348 VDD.n85 VDD.n81 0.09
R2349 VDD.n89 VDD.n85 0.09
R2350 VDD.n98 VDD.n94 0.09
R2351 VDD.n102 VDD.n98 0.09
R2352 VDD.n111 VDD.n107 0.09
R2353 VDD.n115 VDD.n111 0.09
R2354 VDD.n116 VDD.n115 0.09
R2355 VDD.n127 VDD.n123 0.09
R2356 VDD.n131 VDD.n127 0.09
R2357 VDD.n135 VDD.n131 0.09
R2358 VDD.n144 VDD.n140 0.09
R2359 VDD.n153 VDD.n149 0.09
R2360 VDD.n157 VDD.n153 0.09
R2361 VDD.n161 VDD.n157 0.09
R2362 VDD.n162 VDD.n161 0.09
R2363 VDD.n171 VDD.n167 0.09
R2364 VDD.n175 VDD.n171 0.09
R2365 VDD.n860 VDD.n180 0.09
R2366 VDD.n712 VDD.n708 0.09
R2367 VDD.n716 VDD.n712 0.09
R2368 VDD.n718 VDD.n716 0.09
R2369 VDD.n729 VDD.n725 0.09
R2370 VDD.n733 VDD.n729 0.09
R2371 VDD.n737 VDD.n733 0.09
R2372 VDD.n746 VDD.n742 0.09
R2373 VDD.n760 VDD.n756 0.09
R2374 VDD.n765 VDD.n760 0.09
R2375 VDD.n767 VDD.n765 0.09
R2376 VDD.n778 VDD.n774 0.09
R2377 VDD.n782 VDD.n778 0.09
R2378 VDD.n796 VDD.n792 0.09
R2379 VDD.n800 VDD.n796 0.09
R2380 VDD.n809 VDD.n805 0.09
R2381 VDD.n813 VDD.n809 0.09
R2382 VDD.n817 VDD.n813 0.09
R2383 VDD.n826 VDD.n822 0.09
R2384 VDD.n830 VDD.n826 0.09
R2385 VDD.n834 VDD.n830 0.09
R2386 VDD.n835 VDD.n834 0.09
R2387 VDD.n846 VDD.n842 0.09
R2388 VDD.n850 VDD.n846 0.09
R2389 VDD.n857 VDD.n855 0.09
R2390 VDD.n956 VDD.n952 0.09
R2391 VDD.n960 VDD.n956 0.09
R2392 VDD.n964 VDD.n960 0.09
R2393 VDD.n973 VDD.n969 0.09
R2394 VDD.n977 VDD.n973 0.09
R2395 VDD.n981 VDD.n977 0.09
R2396 VDD.n982 VDD.n981 0.09
R2397 VDD.n993 VDD.n989 0.09
R2398 VDD.n997 VDD.n993 0.09
R2399 VDD.n1004 VDD.n1002 0.09
R2400 VDD.n1060 VDD.n1056 0.09
R2401 VDD.n1056 VDD.n1052 0.09
R2402 VDD.n1052 VDD.n1048 0.09
R2403 VDD.n1043 VDD.n1039 0.09
R2404 VDD.n1039 VDD.n1035 0.09
R2405 VDD.n1035 VDD.n1031 0.09
R2406 VDD.n1031 VDD.n1027 0.09
R2407 VDD.n1022 VDD.n1021 0.09
R2408 VDD.n1021 VDD.n1017 0.09
R2409 VDD.n1012 VDD.n1008 0.09
R2410 VDD.n481 VDD.n476 0.086
R2411 VDD.n244 VDD.n243 0.078
R2412 VDD.n312 VDD.n308 0.078
R2413 VDD.n353 VDD.n352 0.078
R2414 VDD.n402 VDD.n401 0.078
R2415 VDD.n535 VDD.n534 0.078
R2416 VDD.n584 VDD.n583 0.078
R2417 VDD.n670 VDD.n666 0.078
R2418 VDD.n10 VDD.n9 0.078
R2419 VDD.n56 VDD.n55 0.078
R2420 VDD.n103 VDD.n102 0.078
R2421 VDD.n704 VDD.n703 0.078
R2422 VDD.n752 VDD.n751 0.078
R2423 VDD.n291 VDD.n290 0.071
R2424 VDD.n453 VDD.n452 0.071
R2425 VDD.n634 VDD.n633 0.071
R2426 VDD.n647 VDD.n646 0.071
R2427 VDD.n801 VDD.n800 0.071
R2428 VDD.n190 VDD.n189 0.07
R2429 VDD.n344 VDD.n343 0.07
R2430 VDD.n526 VDD.n525 0.07
R2431 VDD.n218 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_OR_0/VDD 0.065
R2432 VDD.n265 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/VDD 0.065
R2433 VDD.n320 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/VDD 0.065
R2434 VDD.n375 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/VDD 0.065
R2435 VDD.n401 VDD.n397 0.065
R2436 VDD.n424 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/VDD 0.065
R2437 VDD.n475 VDD.n471 0.065
R2438 VDD.n499 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/VDD 0.065
R2439 VDD.n903 VDD.n899 0.065
R2440 VDD.n923 CMOS_4in_XOR_0/CMOS_XOR_1/VDD 0.065
R2441 VDD.n557 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_OR_0/VDD 0.065
R2442 VDD.n583 VDD.n579 0.065
R2443 VDD.n606 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/VDD 0.065
R2444 VDD.n656 VDD.n652 0.065
R2445 VDD.n678 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/VDD 0.065
R2446 VDD.n30 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/VDD 0.065
R2447 VDD.n77 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/VDD 0.065
R2448 VDD.n123 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/VDD 0.065
R2449 VDD.n149 VDD.n145 0.065
R2450 VDD.n167 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/VDD 0.065
R2451 VDD.n725 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/VDD 0.065
R2452 VDD.n751 VDD.n747 0.065
R2453 VDD.n774 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/VDD 0.065
R2454 VDD.n822 VDD.n818 0.065
R2455 VDD.n842 VDD 0.065
R2456 VDD.n969 VDD.n965 0.065
R2457 VDD.n989 CMOS_4in_XOR_0/CMOS_XOR_0/VDD 0.065
R2458 VDD.n1044 VDD.n1043 0.065
R2459 VDD.n1022 CMOS_4in_XOR_0/CMOS_XOR_3/VDD 0.065
R2460 VDD.n329 VDD.n325 0.063
R2461 VDD.n458 VDD.n457 0.063
R2462 VDD.n687 VDD.n683 0.063
R2463 VDD.n233 VDD.n231 0.056
R2464 VDD.n280 VDD.n278 0.056
R2465 VDD.n390 VDD.n388 0.056
R2466 VDD.n440 VDD.n438 0.056
R2467 VDD.n515 VDD.n513 0.056
R2468 VDD.n572 VDD.n570 0.056
R2469 VDD.n622 VDD.n620 0.056
R2470 VDD.n45 VDD.n43 0.056
R2471 VDD.n92 VDD.n90 0.056
R2472 VDD.n138 VDD.n136 0.056
R2473 VDD.n740 VDD.n738 0.056
R2474 VDD.n790 VDD.n788 0.056
R2475 VDD.n433 VDD.n432 0.055
R2476 VDD.n508 VDD.n507 0.055
R2477 VDD.n932 VDD.n931 0.055
R2478 VDD.n615 VDD.n614 0.055
R2479 VDD.n688 VDD.n687 0.055
R2480 VDD.n176 VDD.n175 0.055
R2481 VDD.n783 VDD.n782 0.055
R2482 VDD.n851 VDD.n850 0.055
R2483 VDD.n998 VDD.n997 0.055
R2484 VDD.n1017 VDD.n1013 0.055
R2485 CMOS_4in_XOR_0/CMOS_INV_0/VDD VDD.n873 0.05
R2486 CMOS_4in_XOR_0/CMOS_INV_1/VDD VDD.n939 0.05
R2487 CMOS_4in_XOR_0/CMOS_INV_2/VDD VDD.n1061 0.05
R2488 VDD.n437 VDD.n433 0.035
R2489 VDD.n512 VDD.n508 0.035
R2490 VDD.n936 VDD.n932 0.035
R2491 VDD.n619 VDD.n615 0.035
R2492 VDD.n692 VDD.n688 0.035
R2493 VDD.n180 VDD.n176 0.035
R2494 VDD.n787 VDD.n783 0.035
R2495 VDD.n855 VDD.n851 0.035
R2496 VDD.n1002 VDD.n998 0.035
R2497 VDD.n1013 VDD.n1012 0.035
R2498 VDD.n231 VDD.n230 0.033
R2499 VDD.n278 VDD.n277 0.033
R2500 VDD.n388 VDD.n387 0.033
R2501 VDD.n438 VDD.n437 0.033
R2502 VDD.n513 VDD.n512 0.033
R2503 VDD.n570 VDD.n569 0.033
R2504 VDD.n620 VDD.n619 0.033
R2505 VDD.n43 VDD.n42 0.033
R2506 VDD.n90 VDD.n89 0.033
R2507 VDD.n136 VDD.n135 0.033
R2508 VDD.n738 VDD.n737 0.033
R2509 VDD.n788 VDD.n787 0.033
R2510 VDD.n516 CMOS_sbox_0/CMOS_s3_0/VDD 0.027
R2511 VDD.n695 CMOS_sbox_0/CMOS_s2_0/VDD 0.027
R2512 VDD.n859 CMOS_sbox_0/CMOS_s0_0/VDD 0.027
R2513 VDD.n858 CMOS_sbox_0/CMOS_s1_0/VDD 0.027
R2514 VDD.n325 VDD.n324 0.026
R2515 VDD.n462 VDD.n458 0.026
R2516 VDD.n683 VDD.n682 0.026
R2517 VDD.n211 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_OR_0/VDD 0.025
R2518 VDD.n313 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/VDD 0.025
R2519 VDD.n397 VDD.n396 0.025
R2520 VDD.n471 VDD.n470 0.025
R2521 VDD.n899 VDD.n898 0.025
R2522 VDD.n916 CMOS_4in_XOR_0/CMOS_XOR_1/VDD 0.025
R2523 VDD.n579 VDD.n578 0.025
R2524 VDD.n652 VDD.n651 0.025
R2525 VDD.n671 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/VDD 0.025
R2526 VDD.n23 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/VDD 0.025
R2527 VDD.n116 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/VDD 0.025
R2528 VDD.n145 VDD.n144 0.025
R2529 VDD.n162 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/VDD 0.025
R2530 VDD.n747 VDD.n746 0.025
R2531 VDD.n818 VDD.n817 0.025
R2532 VDD.n835 VDD 0.025
R2533 VDD.n965 VDD.n964 0.025
R2534 VDD.n982 CMOS_4in_XOR_0/CMOS_XOR_0/VDD 0.025
R2535 VDD.n1048 VDD.n1044 0.025
R2536 VDD.n1027 CMOS_4in_XOR_0/CMOS_XOR_3/VDD 0.025
R2537 VDD.n1006 CMOS_4in_XOR_0/VDD 0.022
R2538 VDD.n879 CMOS_4in_XOR_0/CMOS_INV_0/VDD 0.021
R2539 VDD.n945 CMOS_4in_XOR_0/CMOS_INV_1/VDD 0.021
R2540 CMOS_4in_XOR_0/CMOS_INV_2/VDD VDD.n870 0.021
R2541 VDD.n194 VDD.n190 0.02
R2542 VDD.n348 VDD.n344 0.02
R2543 VDD.n530 VDD.n526 0.02
R2544 VDD.n295 VDD.n291 0.018
R2545 VDD.n457 VDD.n453 0.018
R2546 VDD.n492 VDD.n491 0.018
R2547 VDD.n886 VDD.n873 0.018
R2548 VDD.n638 VDD.n634 0.018
R2549 VDD.n651 VDD.n647 0.018
R2550 VDD.n805 VDD.n801 0.018
R2551 VDD.n952 VDD.n939 0.018
R2552 VDD.n1061 VDD.n1060 0.018
R2553 VDD.n258 VDD.n257 0.017
R2554 VDD.n367 VDD.n366 0.017
R2555 VDD.n417 VDD.n416 0.017
R2556 VDD.n549 VDD.n548 0.017
R2557 VDD.n599 VDD.n598 0.017
R2558 VDD.n70 VDD.n69 0.017
R2559 VDD.n718 VDD.n717 0.017
R2560 VDD.n767 VDD.n766 0.017
R2561 VDD.n248 VDD.n244 0.011
R2562 VDD.n308 VDD.n307 0.011
R2563 VDD.n357 VDD.n353 0.011
R2564 VDD.n406 VDD.n402 0.011
R2565 VDD.n539 VDD.n535 0.011
R2566 VDD.n588 VDD.n584 0.011
R2567 VDD.n666 VDD.n665 0.011
R2568 VDD.n14 VDD.n10 0.011
R2569 VDD.n60 VDD.n56 0.011
R2570 VDD.n107 VDD.n103 0.011
R2571 VDD.n708 VDD.n704 0.011
R2572 VDD.n756 VDD.n752 0.011
R2573 CMOS_sbox_0/CMOS_s0_0/VDD CMOS_sbox_0/VDD 0.01
R2574 VDD.n257 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/VDD 0.007
R2575 VDD.n366 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/VDD 0.007
R2576 VDD.n416 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/VDD 0.007
R2577 VDD.n548 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_OR_0/VDD 0.007
R2578 VDD.n598 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/VDD 0.007
R2579 VDD.n69 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/VDD 0.007
R2580 VDD.n717 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/VDD 0.007
R2581 VDD.n766 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/VDD 0.007
R2582 VDD.n491 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/VDD 0.006
R2583 VDD.n476 VDD.n475 0.003
R2584 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t2 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t3 1221.07
R2585 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.n0 787.238
R2586 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t2 633.02
R2587 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t1 117.958
R2588 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT 91.717
R2589 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t0 45.156
R2590 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n13 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t9 993.097
R2591 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t7 993.097
R2592 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t13 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t10 924.95
R2593 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t8 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t5 924.95
R2594 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t15 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t14 924.95
R2595 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t13 633.02
R2596 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t8 633.02
R2597 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t15 633.02
R2598 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t6 579.86
R2599 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n9 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t17 579.86
R2600 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n11 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t16 570.366
R2601 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n11 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t18 570.366
R2602 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t19 547.727
R2603 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n9 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t12 547.727
R2604 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n13 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t11 356.59
R2605 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t4 356.59
R2606 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n4 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/B 317.612
R2607 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n14 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/A 173
R2608 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n6 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/A 173
R2609 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n12 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/C 158.792
R2610 CMOS_4in_XOR_0/CMOS_INV_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n3 78.72
R2611 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n11 78.72
R2612 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n13 78.72
R2613 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n5 78.72
R2614 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n18 CMOS_4in_XOR_0/CMOS_INV_0/A 57.376
R2615 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n12 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/B 42.892
R2616 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B 42.892
R2617 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n29 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t3 24
R2618 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n29 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t2 24
R2619 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n46 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t0 19.7
R2620 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n46 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t1 19.7
R2621 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n16 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n10 10.065
R2622 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n10 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n9 8.764
R2623 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n30 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n29 8.472
R2624 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n26 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n24 5.44
R2625 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n26 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n25 5.44
R2626 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n41 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n42 4.61
R2627 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n20 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n23 4.5
R2628 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n27 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n31 4.5
R2629 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n39 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n57 4.5
R2630 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n40 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n53 4.5
R2631 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n41 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n49 4.5
R2632 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n38 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n37 4.592
R2633 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n59 4.302
R2634 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n48 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n47 3.472
R2635 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n14 CMOS_sbox_0/CMOS_s3_0/x3 3.33
R2636 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n8 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n7 3.303
R2637 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n27 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n26 3.144
R2638 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n6 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n4 3.096
R2639 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n38 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n33 3.019
R2640 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n47 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n46 2.773
R2641 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n10 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 2.72
R2642 CMOS_4in_XOR_0/XOR3 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n17 2.576
R2643 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n49 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n45 2.56
R2644 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n42 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n44 2.56
R2645 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n23 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n21 2.4
R2646 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n31 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n30 2.4
R2647 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n17 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n8 2.25
R2648 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n53 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n50 2.24
R2649 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n57 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n54 1.92
R2650 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n37 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n36 1.92
R2651 CMOS_sbox_0/CMOS_s1_0/x3 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n6 1.646
R2652 CMOS_sbox_0/CMOS_s2_0/x3 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n14 1.599
R2653 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n15 CMOS_sbox_0/CMOS_s2_0/x3 1.304
R2654 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n20 1.127
R2655 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n16 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n15 1.126
R2656 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n27 1.125
R2657 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n2 1.125
R2658 CMOS_4in_XOR_0/CMOS_XOR_1/XOR CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n60 1.062
R2659 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n57 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n56 0.8
R2660 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n37 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n35 0.8
R2661 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n18 CMOS_4in_XOR_0/XOR3 0.796
R2662 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n32 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n38 0.718
R2663 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n32 0.666
R2664 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n60 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n0 0.571
R2665 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n60 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n1 0.529
R2666 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n53 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n52 0.48
R2667 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n23 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n22 0.32
R2668 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n31 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n28 0.32
R2669 CMOS_4in_XOR_0/CMOS_XOR_1/XOR CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n18 0.215
R2670 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n4 CMOS_sbox_0/CMOS_s0_0/x3 0.181
R2671 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n49 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n48 0.16
R2672 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n42 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n43 0.16
R2673 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n15 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n8 0.157
R2674 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n7 CMOS_sbox_0/CMOS_s1_0/x3 0.157
R2675 CMOS_sbox_0/CMOS_s3_0/x3 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n12 0.157
R2676 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n39 0.115
R2677 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n40 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n41 0.11
R2678 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n39 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n40 0.109
R2679 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n17 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n16 0.106
R2680 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n20 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n19 0.079
R2681 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n59 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n58 0.06
R2682 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n35 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n34 0.055
R2683 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n56 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n55 0.055
R2684 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n52 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n51 0.05
R2685 x0_bar.t0 x0_bar.t1 1345.61
R2686 x0_bar x0_bar.t0 392.02
R2687 x0_bar CMOS_4in_XOR_0/x0_bar 263.2
R2688 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t7 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t5 1345.61
R2689 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t12 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t11 1345.61
R2690 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t4 683.32
R2691 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n6 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t6 681.713
R2692 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t2 616.084
R2693 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t8 570.366
R2694 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t3 570.366
R2695 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t10 528.72
R2696 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t9 528.72
R2697 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n6 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t13 528.72
R2698 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 510.892
R2699 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n8 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/A_bar 505.226
R2700 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t7 392.02
R2701 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t12 392.02
R2702 CMOS_sbox_0/CMOS_s3_0/x0_bar CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/B_bar 346.044
R2703 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n7 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/B_bar 344.84
R2704 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n4 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/C 337.8
R2705 CMOS_4in_XOR_0/CMOS_INV_2/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t0 147.753
R2706 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n3 78.72
R2707 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n10 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t1 76.998
R2708 CMOS_4in_XOR_0/CMOS_INV_2/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n10 17.28
R2709 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n1 14.546
R2710 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n10 CMOS_4in_XOR_0/XOR0_bar 3.777
R2711 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n0 3.68
R2712 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n1 CMOS_sbox_0/CMOS_s2_0/CMOS_XOR_0/B_bar 3.68
R2713 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n6 3.68
R2714 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n2 CMOS_sbox_0/CMOS_s3_0/x0_bar 2.759
R2715 CMOS_sbox_0/CMOS_s2_0/x0_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n2 2.163
R2716 CMOS_sbox_0/CMOS_s1_0/x0_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n5 2.102
R2717 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n9 CMOS_sbox_0/CMOS_s0_0/x0_bar 1.501
R2718 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n4 CMOS_sbox_0/CMOS_s2_0/x0_bar 1.469
R2719 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n7 CMOS_sbox_0/CMOS_s1_0/x0_bar 1.444
R2720 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n8 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n7 1.417
R2721 CMOS_4in_XOR_0/XOR0_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n9 1.365
R2722 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n4 1.357
R2723 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n9 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n8 0.559
R2724 k0_bar.n0 k0_bar.t1 683.32
R2725 k0_bar.n0 k0_bar.t0 528.72
R2726 k0_bar CMOS_4in_XOR_0/k0_bar 108.96
R2727 k0_bar k0_bar.n0 3.68
R2728 x1.n0 x1.t0 993.097
R2729 x1.n0 x1.t1 356.59
R2730 x1 CMOS_4in_XOR_0/x1 119.2
R2731 x1 x1.n0 78.72
R2732 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t18 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t13 1221.07
R2733 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t14 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t10 1221.07
R2734 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n9 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t4 993.097
R2735 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n11 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t9 993.097
R2736 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n4 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t19 993.097
R2737 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t15 579.86
R2738 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t11 579.86
R2739 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n16 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t12 579.86
R2740 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t16 547.727
R2741 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t8 547.727
R2742 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n16 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t6 547.727
R2743 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n17 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/A 451.88
R2744 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n14 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/B 400.52
R2745 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n13 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t18 389.3
R2746 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n6 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t14 389.3
R2747 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n9 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t7 356.59
R2748 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n11 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t5 356.59
R2749 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n4 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t17 356.59
R2750 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n15 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/B 356.332
R2751 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n10 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/A 318.92
R2752 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n6 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n5 211.594
R2753 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n13 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n12 183.874
R2754 CMOS_4in_XOR_0/CMOS_INV_1/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n3 78.72
R2755 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n9 78.72
R2756 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n16 78.72
R2757 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n19 CMOS_4in_XOR_0/CMOS_INV_1/A 57.376
R2758 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n30 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t2 24
R2759 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n30 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t3 24
R2760 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n10 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n8 20.982
R2761 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n47 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t0 19.7
R2762 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n47 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t1 19.7
R2763 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n8 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n7 8.764
R2764 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n12 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n11 8.764
R2765 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n4 8.764
R2766 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n31 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n30 8.472
R2767 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n27 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n25 5.44
R2768 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n27 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n26 5.44
R2769 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n42 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n43 4.61
R2770 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n21 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n24 4.5
R2771 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n28 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n32 4.5
R2772 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n40 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n58 4.5
R2773 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n41 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n54 4.5
R2774 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n42 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n50 4.5
R2775 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n39 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n38 4.592
R2776 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n60 4.302
R2777 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n49 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n48 3.472
R2778 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n18 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n17 3.39
R2779 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n28 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n27 3.144
R2780 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n39 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n34 3.019
R2781 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n48 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n47 2.773
R2782 CMOS_sbox_0/CMOS_s1_0/x1 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n15 2.764
R2783 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n8 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/B 2.72
R2784 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n12 CMOS_sbox_0/CMOS_s2_0/CMOS_XOR_0/A 2.72
R2785 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n13 2.72
R2786 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 2.72
R2787 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n6 2.72
R2788 CMOS_sbox_0/CMOS_s2_0/x1 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n14 2.699
R2789 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n50 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n46 2.56
R2790 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n43 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n45 2.56
R2791 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n24 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n22 2.4
R2792 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n32 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n31 2.4
R2793 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n54 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n51 2.24
R2794 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n14 CMOS_sbox_0/CMOS_s3_0/x1 2.23
R2795 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n15 CMOS_sbox_0/CMOS_s2_0/x1 2.167
R2796 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n58 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n55 1.92
R2797 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n38 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n37 1.92
R2798 CMOS_4in_XOR_0/XOR1 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n18 1.902
R2799 CMOS_sbox_0/CMOS_s3_0/x1 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n10 1.597
R2800 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n18 CMOS_sbox_0/CMOS_s1_0/x1 1.369
R2801 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n21 1.127
R2802 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n28 1.125
R2803 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n2 1.125
R2804 CMOS_4in_XOR_0/CMOS_XOR_2/XOR CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n61 1.062
R2805 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n58 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n57 0.8
R2806 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n38 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n36 0.8
R2807 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n19 CMOS_4in_XOR_0/XOR1 0.796
R2808 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n33 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n39 0.718
R2809 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n33 0.666
R2810 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n61 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n0 0.571
R2811 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n61 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n1 0.529
R2812 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n54 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n53 0.48
R2813 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n24 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n23 0.32
R2814 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n32 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n29 0.32
R2815 CMOS_4in_XOR_0/CMOS_XOR_2/XOR CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n19 0.215
R2816 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n50 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n49 0.16
R2817 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n43 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n44 0.16
R2818 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n17 CMOS_sbox_0/CMOS_s0_0/x1 0.151
R2819 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n40 0.115
R2820 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n41 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n42 0.11
R2821 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n40 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n41 0.109
R2822 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n21 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n20 0.079
R2823 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n60 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n59 0.06
R2824 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n36 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n35 0.055
R2825 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n57 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n56 0.055
R2826 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n53 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n52 0.05
R2827 k1_bar.n0 k1_bar.t0 681.713
R2828 k1_bar.n0 k1_bar.t1 528.72
R2829 k1_bar CMOS_4in_XOR_0/k1_bar 109.28
R2830 k1_bar k1_bar.n0 3.68
R2831 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t2 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t3 1221.07
R2832 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.n0 739.238
R2833 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t2 633.02
R2834 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/OUT CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t1 114.438
R2835 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.n0 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/OUT 95.237
R2836 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.n0 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t0 45.156
R2837 s2.n2 s2.t0 120.552
R2838 s2.n1 s2.t1 98.438
R2839 s2 s2.n2 7.84
R2840 s2 s2.n1 3.68
R2841 s2.n1 s2.n0 3.084
R2842 s2.n0 CMOS_sbox_0/CMOS_s2_0/s2 0.374
R2843 k2_bar.n0 k2_bar.t1 683.32
R2844 k2_bar.n0 k2_bar.t0 528.72
R2845 k2_bar CMOS_4in_XOR_0/k2_bar 109.92
R2846 k2_bar k2_bar.n0 3.68
R2847 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t10 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t4 1345.61
R2848 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t13 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t15 1221.07
R2849 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t9 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t3 1221.07
R2850 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t7 683.32
R2851 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n11 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t14 683.32
R2852 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n4 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t13 630.3
R2853 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t11 579.86
R2854 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t5 579.86
R2855 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t8 547.727
R2856 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t2 547.727
R2857 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t12 528.72
R2858 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n11 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t6 528.72
R2859 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t10 392.02
R2860 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t9 392.02
R2861 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n10 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/B 285.69
R2862 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n8 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/B_bar 198.92
R2863 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n12 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 198.92
R2864 CMOS_4in_XOR_0/CMOS_INV_3/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t0 147.753
R2865 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n15 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t1 76.998
R2866 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n5 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/A_bar 44.234
R2867 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n4 41.121
R2868 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n6 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n3 17.994
R2869 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n9 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n1 17.994
R2870 CMOS_4in_XOR_0/CMOS_INV_3/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n15 17.28
R2871 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n2 8.764
R2872 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n0 8.764
R2873 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n14 CMOS_4in_XOR_0/XOR2_bar 4.541
R2874 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n7 3.68
R2875 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n11 3.68
R2876 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n15 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n14 3.033
R2877 CMOS_4in_XOR_0/XOR2_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n13 2.867
R2878 CMOS_sbox_0/CMOS_s1_0/x2_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n10 2.764
R2879 CMOS_sbox_0/CMOS_s3_0/x2_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n5 2.762
R2880 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n4 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/A 2.72
R2881 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n3 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/B 2.72
R2882 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/B 2.72
R2883 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n10 CMOS_sbox_0/CMOS_s0_0/x2_bar 2.157
R2884 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n9 CMOS_sbox_0/CMOS_s2_0/x2_bar 2.019
R2885 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n6 CMOS_sbox_0/CMOS_s3_0/x2_bar 2.019
R2886 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n8 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n6 1.697
R2887 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n13 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n9 1.242
R2888 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n12 CMOS_sbox_0/CMOS_s1_0/x2_bar 1.205
R2889 CMOS_sbox_0/CMOS_s2_0/x2_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n8 1.205
R2890 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n14 CMOS_4in_XOR_0/XOR2_bar 0.93
R2891 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n13 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n12 0.447
R2892 k3.t1 k3.t0 923.343
R2893 k3 k3.t1 633.02
R2894 k3 CMOS_4in_XOR_0/k3 264.8
R2895 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t3 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t2 1221.07
R2896 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.n0 787.238
R2897 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t3 633.02
R2898 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t1 117.958
R2899 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.n0 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT 91.717
R2900 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.n0 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t0 45.156
R2901 x3.n0 x3.t1 993.097
R2902 x3.n0 x3.t0 356.59
R2903 x3 CMOS_4in_XOR_0/x3 119.52
R2904 x3 x3.n0 78.72
R2905 x3_bar.t1 x3_bar.t0 1345.61
R2906 x3_bar x3_bar.t1 392.02
R2907 x3_bar CMOS_4in_XOR_0/x3_bar 263.52
R2908 s3.n2 s3.t0 120.552
R2909 s3.n1 s3.t1 98.438
R2910 s3 s3.n2 7.84
R2911 s3 s3.n1 3.68
R2912 s3.n1 s3.n0 3.084
R2913 s3.n0 CMOS_sbox_0/CMOS_s3_0/s3 0.374
R2914 s0 s0.t0 117.353
R2915 s0.n0 s0.t1 95.65
R2916 s0 s0.n0 10.009
R2917 s0.n0 CMOS_sbox_0/CMOS_s0_0/s0 0.913
R2918 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t7 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t6 1345.61
R2919 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t9 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t4 1345.61
R2920 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t5 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t11 1345.61
R2921 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t10 579.86
R2922 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t3 579.86
R2923 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n0 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t8 547.727
R2924 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n5 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t2 547.727
R2925 CMOS_sbox_0/CMOS_s3_0/x1_bar CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/A_bar 436.286
R2926 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t7 392.02
R2927 CMOS_sbox_0/CMOS_s2_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t9 392.02
R2928 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t5 392.02
R2929 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n6 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_2/B 380.227
R2930 CMOS_4in_XOR_0/CMOS_INV_1/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t0 136.873
R2931 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_2/B CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n5 78.72
R2932 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n8 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t1 76.998
R2933 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n3 CMOS_sbox_0/CMOS_s2_0/CMOS_XOR_0/A_bar 44.915
R2934 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n4 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 44.915
R2935 CMOS_4in_XOR_0/CMOS_INV_1/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n8 28.16
R2936 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n2 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n1 11.862
R2937 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n1 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n0 8.764
R2938 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n8 CMOS_4in_XOR_0/XOR1_bar 3.777
R2939 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n7 CMOS_sbox_0/CMOS_s0_0/x1_bar 3.078
R2940 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n1 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/B 2.72
R2941 CMOS_sbox_0/CMOS_s1_0/x1_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n4 2.663
R2942 CMOS_sbox_0/CMOS_s2_0/x1_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n3 2.663
R2943 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n4 CMOS_sbox_0/CMOS_s2_0/x1_bar 2.259
R2944 CMOS_4in_XOR_0/XOR1_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n7 2.11
R2945 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n7 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n6 1.54
R2946 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n2 CMOS_sbox_0/CMOS_s3_0/x1_bar 1.448
R2947 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n3 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n2 0.803
R2948 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n6 CMOS_sbox_0/CMOS_s1_0/x1_bar 0.294
R2949 k0.t1 k0.t0 924.95
R2950 k0 k0.t1 633.02
R2951 k0 CMOS_4in_XOR_0/k0 263.52
R2952 x0.n0 x0.t1 993.097
R2953 x0.n0 x0.t0 356.59
R2954 x0 CMOS_4in_XOR_0/x0 118.88
R2955 x0 x0.n0 78.72
R2956 x1_bar.t0 x1_bar.t1 1345.61
R2957 x1_bar x1_bar.t0 392.02
R2958 x1_bar CMOS_4in_XOR_0/x1_bar 263.52
R2959 k3_bar.n0 k3_bar.t1 681.713
R2960 k3_bar.n0 k3_bar.t0 528.72
R2961 k3_bar CMOS_4in_XOR_0/k3_bar 109.6
R2962 k3_bar k3_bar.n0 3.68
R2963 k1.t1 k1.t0 923.343
R2964 k1 k1.t1 633.02
R2965 k1 CMOS_4in_XOR_0/k1 265.44
R2966 x2.n0 x2.t0 993.097
R2967 x2.n0 x2.t1 356.59
R2968 x2 CMOS_4in_XOR_0/x2 119.2
R2969 x2 x2.n0 78.72
R2970 s1.n2 s1.t0 120.552
R2971 s1.n1 s1.t1 98.438
R2972 s1 s1.n2 7.84
R2973 s1 s1.n1 3.68
R2974 s1.n1 s1.n0 3.084
R2975 s1.n0 CMOS_sbox_0/CMOS_s1_0/s1 0.374
R2976 k2.t1 k2.t0 924.95
R2977 k2 k2.t1 633.02
R2978 k2 CMOS_4in_XOR_0/k2 264.8
C0 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND 0.00fF
C1 a_425_n7820# a_n432_n7820# 0.00fF
C2 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n2290_n2118# 0.01fF
C3 a_n1990_n540# a_n2140_n2118# 0.00fF
C4 a_425_n4664# a_575_n3696# 0.00fF
C5 a_n2290_n540# a_n2140_n540# 0.02fF
C6 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C7 a_n4395_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C8 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n432_n7820# 0.00fF
C9 a_n432_n4664# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND 0.00fF
C10 a_n2495_n10008# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.04fF
C11 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_n732_n7820# 0.01fF
C12 a_n2290_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.02fF
C13 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n1990_n5274# 0.00fF
C14 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.76fF
C15 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND 0.00fF
C16 a_n2290_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C17 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n2290_n8430# 0.01fF
C18 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.35fF
C19 a_n2195_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C20 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR a_n787_1038# 0.07fF
C21 a_425_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C22 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.21fF
C23 a_n2345_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.02fF
C24 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.00fF
C25 a_275_n5942# a_425_n5274# 0.00fF
C26 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2140_n540# 0.07fF
C27 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR 0.01fF
C28 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n2140_n8430# 0.06fF
C29 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n4695_n2786# 0.01fF
C30 a_n4395_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C31 a_n787_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C32 a_n2290_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C33 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_n2140_n2118# 0.01fF
C34 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_n1990_370# 0.00fF
C35 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n4395_1038# 0.00fF
C36 a_n2195_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C37 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_425_n2118# 0.01fF
C38 a_425_n7820# a_n732_n8430# 0.00fF
C39 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_275_n2786# 0.05fF
C40 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.03fF
C41 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT 0.10fF
C42 a_n2045_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C43 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.15fF
C44 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n4695_1038# 0.00fF
C45 a_n4395_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C46 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.01fF
C47 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar a_n732_n1508# 0.01fF
C48 a_n2345_n6852# a_n2290_n5274# 0.00fF
C49 a_n2290_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C50 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n732_n8430# 0.01fF
C51 a_425_n10008# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.00fF
C52 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A a_425_n1508# 0.09fF
C53 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_425_n4664# 0.08fF
C54 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.84fF
C55 a_425_n540# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A 0.00fF
C56 a_n432_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C57 a_275_n9098# a_425_n7820# 0.01fF
C58 a_n787_n10008# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.00fF
C59 a_n787_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C60 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n2290_n8430# 0.00fF
C61 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2290_n4664# 0.00fF
C62 a_n4395_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C63 a_275_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.04fF
C64 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n1990_n1508# 0.03fF
C65 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n4395_1648# 0.00fF
C66 a_n2345_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C67 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A a_n787_n3696# 0.01fF
C68 a_n1990_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C69 a_n787_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C70 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.08fF
C71 a_n787_n9098# a_n787_n10008# 0.01fF
C72 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A a_n1990_n1508# 0.00fF
C73 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.04fF
C74 a_275_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.10fF
C75 a_n2140_n540# a_n1990_n1508# 0.00fF
C76 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n4695_1648# 0.00fF
C77 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2290_370# 0.00fF
C78 a_n2140_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.15fF
C79 a_275_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.00fF
C80 a_n2195_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.00fF
C81 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C82 a_n787_n6852# a_575_n6852# 0.00fF
C83 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n4695_1038# 0.00fF
C84 a_n787_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C85 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND a_n2495_n10008# 0.00fF
C86 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n2495_n10008# 0.02fF
C87 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.35fF
C88 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n732_n1508# 0.01fF
C89 a_n1990_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C90 a_n432_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C91 a_n4395_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C92 a_n4695_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C93 a_n2290_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C94 a_n787_1038# a_n2290_1038# 0.00fF
C95 a_275_n5942# a_425_n7820# 0.01fF
C96 a_n432_n8430# a_n787_n10008# 0.00fF
C97 a_n787_n6852# a_425_n6852# 0.00fF
C98 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C99 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n787_n6852# 0.03fF
C100 a_275_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C101 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR a_1637_1038# 0.00fF
C102 a_425_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A 0.07fF
C103 a_275_n9098# a_575_n10008# 0.02fF
C104 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B 0.01fF
C105 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C106 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.09fF
C107 a_n1990_n4664# a_n2495_n3696# 0.00fF
C108 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n2290_n8430# 0.00fF
C109 a_n2345_n5942# a_n2345_n6852# 0.00fF
C110 a_n732_n7820# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.00fF
C111 a_425_n540# a_425_1038# 0.00fF
C112 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2345_n2786# 0.00fF
C113 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_n732_n5274# 0.00fF
C114 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n4695_1648# 0.00fF
C115 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.00fF
C116 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n1990_n7820# 0.01fF
C117 a_425_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C118 a_425_n1508# a_425_n3696# 0.00fF
C119 a_425_n1508# a_n732_n1508# 0.00fF
C120 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.03fF
C121 a_n787_n2786# a_n2495_n3696# 0.00fF
C122 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n1990_n5274# 0.00fF
C123 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.39fF
C124 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.03fF
C125 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.15fF
C126 a_n732_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.01fF
C127 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.09fF
C128 a_n1990_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C129 a_n787_n5942# a_275_n5942# 0.00fF
C130 a_n2345_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C131 a_425_n3696# a_n787_n3696# 0.00fF
C132 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n2140_n540# 0.02fF
C133 a_n4695_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C134 a_n787_n3696# a_n732_n1508# 0.00fF
C135 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_n432_n8430# 0.00fF
C136 a_n2345_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.13fF
C137 a_n2195_n9098# a_n2140_n8430# 0.00fF
C138 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_n787_370# 0.00fF
C139 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_n1990_1038# 0.01fF
C140 a_n732_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT 0.01fF
C141 a_n2290_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C142 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n787_n540# 0.04fF
C143 a_n2140_n5274# a_n1990_n5274# 0.01fF
C144 a_n2140_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.35fF
C145 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR 0.01fF
C146 a_n1990_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A 0.03fF
C147 a_425_n4664# a_575_n6852# 0.00fF
C148 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.17fF
C149 a_n1990_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C150 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C151 a_n4395_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C152 a_n2195_n2786# a_n2495_n3696# 0.01fF
C153 a_n2045_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C154 a_275_n2786# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.00fF
C155 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.01fF
C156 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n2290_1648# 0.00fF
C157 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_n432_n5274# 0.00fF
C158 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.04fF
C159 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.06fF
C160 a_n4395_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C161 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n4695_n540# 0.00fF
C162 a_n2195_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C163 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n2140_n540# 0.12fF
C164 a_n732_n8430# a_n2140_n8430# 0.00fF
C165 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.16fF
C166 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND a_575_n10008# 0.00fF
C167 a_425_n4664# a_425_n6852# 0.00fF
C168 a_n2140_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.33fF
C169 a_n2290_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C170 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.04fF
C171 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.07fF
C172 a_n1990_n4664# a_n2345_n6852# 0.00fF
C173 a_n2345_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.08fF
C174 a_n787_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT 0.01fF
C175 a_n432_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C176 a_n432_n4664# a_n787_n3696# 0.00fF
C177 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_575_n3696# 0.01fF
C178 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n787_n540# 0.00fF
C179 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n2290_370# 0.00fF
C180 a_n4695_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C181 a_n1990_n7820# a_n2495_n10008# 0.00fF
C182 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_425_n7820# 0.09fF
C183 a_n4395_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C184 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2290_n2118# 0.00fF
C185 a_n2195_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C186 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.05fF
C187 a_n2345_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.00fF
C188 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.23fF
C189 a_n2290_n4664# a_n2140_n5274# 0.02fF
C190 a_n787_n540# a_n1990_370# 0.00fF
C191 a_n2045_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C192 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.04fF
C193 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n2290_1648# 0.00fF
C194 a_n2290_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C195 a_425_n5274# a_425_n4664# 0.01fF
C196 a_n4395_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C197 a_n787_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.00fF
C198 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_n2195_n2786# 0.00fF
C199 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n2290_n7820# 0.01fF
C200 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A 0.32fF
C201 a_n787_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C202 a_425_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.01fF
C203 a_n2195_n5942# a_n2140_n5274# 0.00fF
C204 a_n787_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.01fF
C205 a_425_n540# a_n787_n540# 0.01fF
C206 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n2290_370# 0.00fF
C207 a_n432_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C208 a_n2345_n6852# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND 0.00fF
C209 a_575_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.00fF
C210 a_n432_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C211 a_n2345_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C212 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n787_n10008# 0.02fF
C213 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n1990_n7820# 0.00fF
C214 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.07fF
C215 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n787_1038# 0.08fF
C216 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A a_425_1038# 0.00fF
C217 a_n432_n8430# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.00fF
C218 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n732_n1508# 0.00fF
C219 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A a_n732_n5274# 0.01fF
C220 a_n4395_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.00fF
C221 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar a_n2290_n5274# 0.01fF
C222 a_n2495_n3696# a_n1990_n2118# 0.00fF
C223 a_n787_n5942# a_n787_n6852# 0.01fF
C224 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n732_n7820# 0.00fF
C225 a_n2195_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C226 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.12fF
C227 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_425_n3696# 0.00fF
C228 a_n2290_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C229 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n2140_n8430# 0.05fF
C230 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.14fF
C231 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_n732_n1508# 0.00fF
C232 a_n2345_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C233 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n2290_n7820# 0.00fF
C234 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2290_n8430# 0.00fF
C235 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_425_370# 0.00fF
C236 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.16fF
C237 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n4395_n1508# 0.00fF
C238 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.08fF
C239 a_n432_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C240 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.05fF
C241 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n732_n8430# 0.00fF
C242 a_n732_n4664# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.02fF
C243 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.86fF
C244 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A a_n1990_n5274# 0.00fF
C245 a_n787_n540# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B 0.00fF
C246 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n787_n10008# 0.05fF
C247 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C248 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n1990_n8430# 0.01fF
C249 a_n1990_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C250 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n732_n7820# 0.00fF
C251 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n4395_370# 0.00fF
C252 a_n2140_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.37fF
C253 a_n4695_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C254 a_425_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C255 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND a_275_n9098# 0.10fF
C256 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.24fF
C257 a_425_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C258 a_n1990_n4664# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.00fF
C259 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n2140_n5274# 0.08fF
C260 a_n787_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR 0.01fF
C261 a_n2345_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C262 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_n432_n7820# 0.03fF
C263 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n2290_n2118# 0.00fF
C264 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n2290_n7820# 0.00fF
C265 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2495_n3696# 0.11fF
C266 a_n2345_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C267 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.10fF
C268 a_n4695_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C269 a_n787_n540# a_n787_370# 0.01fF
C270 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.03fF
C271 a_n2195_n5942# a_n2140_n8430# 0.00fF
C272 a_n787_n6852# a_n432_n7820# 0.00fF
C273 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n1990_n8430# 0.00fF
C274 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n4395_370# 0.00fF
C275 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR 0.02fF
C276 a_n2290_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C277 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_n2140_n8430# 0.04fF
C278 a_n1990_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.00fF
C279 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar a_n732_n5274# 0.01fF
C280 a_n2495_n10008# a_n2290_n8430# 0.00fF
C281 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.02fF
C282 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.21fF
C283 a_n2345_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.14fF
C284 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C285 a_n1990_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.00fF
C286 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_425_n4664# 0.00fF
C287 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n732_n7820# 0.01fF
C288 a_n2290_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C289 a_n787_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C290 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.85fF
C291 a_n4395_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C292 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.06fF
C293 a_n2195_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C294 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_n732_n8430# 0.01fF
C295 a_n787_n540# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.05fF
C296 a_n4695_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C297 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C298 a_n787_1038# a_n787_370# 0.00fF
C299 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n1990_n5274# 0.01fF
C300 a_n2045_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C301 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.07fF
C302 a_n787_1038# a_n1990_1038# 0.00fF
C303 a_n2290_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C304 a_n1990_n7820# a_n2140_n8430# 0.03fF
C305 a_n4395_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.02fF
C306 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C307 a_n2495_n3696# a_n787_n3696# 0.00fF
C308 a_n2495_n3696# a_n1990_n1508# 0.00fF
C309 a_n732_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C310 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.04fF
C311 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n2290_n5274# 0.01fF
C312 a_n2140_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.21fF
C313 a_n787_n6852# a_n732_n8430# 0.00fF
C314 a_n1990_1648# a_n787_1038# 0.00fF
C315 a_n4695_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C316 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT 0.06fF
C317 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A 0.01fF
C318 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.05fF
C319 a_275_n9098# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.01fF
C320 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n2290_1038# 0.00fF
C321 a_n787_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.02fF
C322 a_n2290_n540# a_n787_n540# 0.00fF
C323 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.00fF
C324 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n2290_n8430# 0.01fF
C325 a_n432_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C326 a_275_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C327 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n1990_n8430# 0.00fF
C328 a_n4395_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C329 a_n787_n10008# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.05fF
C330 a_n2345_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C331 a_n787_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C332 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2345_n6852# 0.06fF
C333 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.58fF
C334 a_n1990_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C335 a_n1990_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.02fF
C336 a_n787_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C337 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n787_n540# 0.01fF
C338 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_425_n5274# 0.00fF
C339 a_n1990_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C340 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_425_n1508# 0.00fF
C341 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n4695_1038# 0.00fF
C342 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.02fF
C343 a_n432_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.03fF
C344 a_n787_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C345 a_n2045_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.00fF
C346 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.09fF
C347 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n2290_n5274# 0.01fF
C348 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2290_1648# 0.02fF
C349 a_n2290_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.02fF
C350 a_n2290_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.00fF
C351 a_n432_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C352 a_n2290_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C353 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B a_1637_1038# 0.08fF
C354 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.19fF
C355 a_275_n5942# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.00fF
C356 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n2290_1038# 0.00fF
C357 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n432_n8430# 0.01fF
C358 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_n787_n3696# 0.10fF
C359 a_275_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.02fF
C360 a_n432_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C361 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.03fF
C362 a_n2290_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.01fF
C363 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A 0.00fF
C364 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B 0.00fF
C365 a_n432_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.03fF
C366 a_n2195_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C367 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.02fF
C368 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.01fF
C369 a_275_n5942# a_n787_n6852# 0.01fF
C370 a_n4395_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C371 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.12fF
C372 a_n4695_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C373 a_n2140_n540# a_n2290_370# 0.01fF
C374 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n787_n10008# 0.02fF
C375 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n4695_1648# 0.00fF
C376 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n787_1038# 0.01fF
C377 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.09fF
C378 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.02fF
C379 a_n787_n540# a_425_370# 0.00fF
C380 a_n2195_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C381 a_n787_n2786# a_275_n2786# 0.00fF
C382 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A a_425_n3696# 0.00fF
C383 a_n787_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR 0.00fF
C384 a_n2345_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C385 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C386 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A a_n732_n1508# 0.02fF
C387 a_n732_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C388 a_n787_n9098# CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR 0.01fF
C389 a_275_n2786# a_575_n3696# 0.02fF
C390 a_425_n7820# a_425_n8430# 0.01fF
C391 a_425_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C392 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C393 a_n1990_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C394 a_n787_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C395 a_n787_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.07fF
C396 a_n2345_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C397 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT a_425_n10008# 0.01fF
C398 a_n2140_n5274# a_n2495_n3696# 0.01fF
C399 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_575_n6852# 0.01fF
C400 a_n787_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.05fF
C401 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_425_n8430# 0.01fF
C402 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_425_1648# 0.06fF
C403 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C404 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n732_n5274# 0.00fF
C405 a_n2345_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C406 a_n432_n1508# a_425_n1508# 0.00fF
C407 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT a_n787_n10008# 0.10fF
C408 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2290_n7820# 0.01fF
C409 a_n1990_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.00fF
C410 a_n1990_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C411 a_n2140_n2118# a_n2195_n2786# 0.00fF
C412 a_n2290_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C413 a_n4395_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C414 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n432_n2118# 0.01fF
C415 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n432_n8430# 0.00fF
C416 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_425_n6852# 0.01fF
C417 a_n432_n1508# a_n787_n3696# 0.00fF
C418 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.05fF
C419 a_n2345_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C420 a_275_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR 0.00fF
C421 a_n1990_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C422 a_n4395_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C423 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n1990_n540# 0.00fF
C424 a_425_1038# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A 0.00fF
C425 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.10fF
C426 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.03fF
C427 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n732_n7820# 0.01fF
C428 a_n732_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C429 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_275_n2786# 0.01fF
C430 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A a_425_n6852# 0.00fF
C431 a_n4695_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C432 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.01fF
C433 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.00fF
C434 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n1990_n5274# 0.00fF
C435 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.01fF
C436 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n732_n5274# 0.01fF
C437 a_n2345_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.10fF
C438 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2345_n9098# 0.00fF
C439 a_n2140_n8430# a_n2290_n8430# 0.01fF
C440 a_n432_n2118# a_425_n1508# 0.00fF
C441 a_275_n5942# a_425_n4664# 0.01fF
C442 a_n1990_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C443 a_n2495_n10008# a_n787_n10008# 0.00fF
C444 a_n732_n2118# a_n787_n540# 0.00fF
C445 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n787_n540# 0.00fF
C446 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_n2140_n5274# 0.01fF
C447 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 8.11fF
C448 a_n4695_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C449 a_n4395_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C450 a_n4395_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C451 a_n1990_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C452 a_425_1648# a_425_1038# 0.01fF
C453 a_n2195_n5942# a_n787_n6852# 0.00fF
C454 a_n1990_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C455 a_n432_n2118# a_n787_n3696# 0.00fF
C456 a_n1990_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C457 a_n2045_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C458 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n1990_370# 0.00fF
C459 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n2290_1648# 0.01fF
C460 a_n732_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.00fF
C461 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.08fF
C462 a_n787_1648# a_425_1648# 0.00fF
C463 a_n787_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C464 a_425_n5274# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.01fF
C465 a_n2345_n6852# a_n2140_n5274# 0.01fF
C466 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C467 a_n787_n6852# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.01fF
C468 a_n787_n5942# a_n2345_n6852# 0.00fF
C469 a_n2290_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C470 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n1990_n8430# 0.00fF
C471 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT a_n2345_n9098# 0.00fF
C472 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n4395_370# 0.00fF
C473 a_425_n7820# a_425_n10008# 0.00fF
C474 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT 0.06fF
C475 a_n732_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C476 a_n4395_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C477 a_n4695_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C478 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.94fF
C479 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR 0.00fF
C480 a_n1990_n7820# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.00fF
C481 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n2290_n2118# 0.01fF
C482 a_n787_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C483 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n787_n540# 0.09fF
C484 a_425_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C485 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A a_n787_n3696# 0.01fF
C486 a_n2140_n2118# a_n1990_n2118# 0.01fF
C487 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n787_n10008# 0.03fF
C488 a_1637_1648# a_1637_1038# 0.01fF
C489 a_n2045_n5942# a_n2140_n5274# 0.00fF
C490 a_n1990_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C491 a_n2290_n4664# CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR 0.00fF
C492 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n787_1038# 0.04fF
C493 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C494 a_n4695_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C495 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n4395_n2118# 0.00fF
C496 a_n4695_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C497 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.01fF
C498 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n4695_n3696# 0.02fF
C499 a_n2195_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C500 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar a_n2290_n5274# 0.01fF
C501 a_n432_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C502 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR 0.01fF
C503 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n1990_370# 0.00fF
C504 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.05fF
C505 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.04fF
C506 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.25fF
C507 a_n2290_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C508 a_n2290_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C509 a_n787_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C510 a_n432_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C511 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.01fF
C512 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_n732_n5274# 0.00fF
C513 a_n432_n4664# a_n787_n6852# 0.00fF
C514 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_n2140_n540# 0.03fF
C515 a_n432_n1508# CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR 0.00fF
C516 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n2290_n7820# 0.00fF
C517 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.00fF
C518 a_n2345_n9098# a_n2495_n10008# 0.01fF
C519 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.06fF
C520 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_425_n7820# 0.02fF
C521 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C522 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n787_1038# 0.01fF
C523 a_n432_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C524 a_n4695_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.02fF
C525 a_n2290_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C526 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.69fF
C527 a_n4395_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C528 a_n432_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND 0.00fF
C529 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.04fF
C530 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.04fF
C531 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n787_n6852# 0.05fF
C532 a_575_n10008# a_n787_n10008# 0.00fF
C533 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n4395_n2118# 0.00fF
C534 a_n732_n7820# a_425_n7820# 0.00fF
C535 a_n4695_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C536 a_425_n4664# a_425_n3696# 0.00fF
C537 a_n2195_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C538 a_n1990_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.02fF
C539 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.06fF
C540 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n2290_n8430# 0.00fF
C541 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR 0.04fF
C542 a_n732_n4664# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND 0.00fF
C543 a_n1990_n8430# a_n2495_n10008# 0.00fF
C544 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n732_n7820# 0.00fF
C545 a_n4395_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C546 a_n4395_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.02fF
C547 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2290_n5274# 0.00fF
C548 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.09fF
C549 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2140_n2118# 0.17fF
C550 a_n2345_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C551 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2290_1038# 0.01fF
C552 a_n2140_n2118# a_n2290_n1508# 0.02fF
C553 a_425_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C554 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_n2140_n5274# 0.01fF
C555 a_n787_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.01fF
C556 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n432_n8430# 0.01fF
C557 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT a_n787_n9098# 0.01fF
C558 a_n4695_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C559 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_275_n2786# 0.00fF
C560 a_275_n9098# a_425_n8430# 0.00fF
C561 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.06fF
C562 a_n432_n4664# CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR 0.00fF
C563 a_n2345_n6852# a_n2140_n8430# 0.01fF
C564 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n4695_1038# 0.00fF
C565 a_n2345_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C566 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_n432_n2118# 0.00fF
C567 a_n787_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C568 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n1990_1038# 0.00fF
C569 a_n787_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C570 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.06fF
C571 a_n2140_n5274# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.04fF
C572 a_n787_1038# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A 0.00fF
C573 a_n4395_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C574 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar a_n1990_n1508# 0.01fF
C575 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n1990_n2118# 0.00fF
C576 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n1990_n8430# 0.00fF
C577 a_n1990_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C578 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n4395_370# 0.02fF
C579 a_n432_n4664# a_425_n4664# 0.00fF
C580 a_n2045_n5942# a_n2140_n8430# 0.00fF
C581 a_n787_n10008# a_n432_n7820# 0.00fF
C582 a_n2345_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.08fF
C583 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C584 a_275_n2786# a_425_n1508# 0.01fF
C585 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.03fF
C586 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.00fF
C587 a_n4695_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C588 a_n4695_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C589 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.71fF
C590 a_n787_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C591 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n4695_1648# 0.00fF
C592 a_n4395_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C593 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND 0.04fF
C594 a_n2495_n10008# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C595 a_n787_n9098# a_n2495_n10008# 0.00fF
C596 a_n2140_n2118# a_n1990_n1508# 0.03fF
C597 a_n2195_n9098# a_n787_n10008# 0.00fF
C598 a_425_1648# a_n787_1038# 0.01fF
C599 a_275_n2786# a_n787_n3696# 0.01fF
C600 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.00fF
C601 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C602 a_425_n540# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B 0.05fF
C603 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n787_370# 0.00fF
C604 a_n4695_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C605 a_n2045_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C606 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.01fF
C607 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n1990_1038# 0.00fF
C608 a_n2290_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C609 a_n1990_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.01fF
C610 a_n2345_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.00fF
C611 a_425_n7820# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.08fF
C612 a_n1990_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C613 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n1990_n2118# 0.01fF
C614 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_425_n8430# 0.00fF
C615 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR 0.01fF
C616 a_n1990_n540# a_n2140_n540# 0.03fF
C617 a_n2290_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C618 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.06fF
C619 a_n732_n8430# a_n787_n10008# 0.00fF
C620 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_n432_n7820# 0.01fF
C621 a_n787_n10008# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C622 a_n4695_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C623 a_n1990_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C624 a_n2290_n7820# a_n2140_n8430# 0.02fF
C625 a_n787_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C626 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 10.11fF
C627 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.82fF
C628 a_n787_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C629 a_275_n9098# a_425_n10008# 0.02fF
C630 a_425_n540# a_n787_370# 0.00fF
C631 a_n2290_n4664# a_n2495_n3696# 0.00fF
C632 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.00fF
C633 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.97fF
C634 a_n2290_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C635 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n4395_n2786# 0.02fF
C636 a_275_n9098# a_n787_n10008# 0.01fF
C637 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C638 a_n1990_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C639 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_n2140_n8430# 0.01fF
C640 a_n787_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C641 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.00fF
C642 a_425_n7820# a_n432_n8430# 0.00fF
C643 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n2290_n5274# 0.00fF
C644 a_n2140_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.22fF
C645 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A a_1637_1038# 0.05fF
C646 a_n787_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C647 a_n2290_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.02fF
C648 a_n2345_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.03fF
C649 a_n732_n2118# a_n2140_n2118# 0.00fF
C650 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.04fF
C651 a_n732_n7820# a_n2140_n8430# 0.00fF
C652 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n2290_1038# 0.00fF
C653 a_n2290_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C654 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n4395_1038# 0.00fF
C655 a_n2345_n6852# a_n1990_n5274# 0.00fF
C656 a_n432_n5274# a_n787_n6852# 0.00fF
C657 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n432_n8430# 0.01fF
C658 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C659 a_575_n10008# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.00fF
C660 a_n787_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.05fF
C661 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C662 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_n732_n8430# 0.00fF
C663 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A a_n787_n540# 0.01fF
C664 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A 0.01fF
C665 a_425_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C666 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C667 a_425_n540# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.07fF
C668 a_n4395_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C669 a_n4695_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C670 a_n4395_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C671 a_n787_n3696# a_n732_n5274# 0.00fF
C672 a_n2140_n540# a_n787_n540# 0.02fF
C673 a_n2140_n5274# a_n2290_n5274# 0.01fF
C674 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n1990_n4664# 0.00fF
C675 a_n2045_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C676 a_n2290_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C677 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 10.47fF
C678 a_n2195_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C679 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.01fF
C680 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.02fF
C681 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n2290_1648# 0.00fF
C682 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.12fF
C683 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.05fF
C684 a_n787_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.02fF
C685 a_425_1648# a_1637_1038# 0.01fF
C686 a_n2345_n2786# a_n2495_n3696# 0.01fF
C687 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n1990_n1508# 0.00fF
C688 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n4395_1648# 0.00fF
C689 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.35fF
C690 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_425_n8430# 0.01fF
C691 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n1990_370# 0.00fF
C692 a_n2345_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C693 a_n1990_n8430# a_n2140_n8430# 0.01fF
C694 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND a_425_n10008# 0.01fF
C695 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n4395_1038# 0.00fF
C696 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND a_575_n6852# 0.00fF
C697 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR a_425_1648# 0.04fF
C698 a_n432_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.03fF
C699 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n787_n10008# 0.00fF
C700 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND a_n787_n10008# 0.07fF
C701 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.03fF
C702 a_n787_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C703 a_425_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C704 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n432_n5274# 0.00fF
C705 a_n732_n4664# a_n787_n3696# 0.00fF
C706 a_425_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.05fF
C707 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_275_n2786# 0.12fF
C708 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n2495_n10008# 0.01fF
C709 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_425_n3696# 0.01fF
C710 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND a_425_n6852# 0.01fF
C711 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND 0.00fF
C712 a_n2345_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C713 a_n432_n7820# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.00fF
C714 a_n1990_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C715 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n4395_n2118# 0.00fF
C716 a_n4395_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C717 a_n2195_n5942# a_n2345_n6852# 0.01fF
C718 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B 0.01fF
C719 a_n787_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.05fF
C720 a_275_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.05fF
C721 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2195_n2786# 0.00fF
C722 a_n787_n540# a_n2290_370# 0.00fF
C723 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_575_n6852# 0.00fF
C724 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n1990_n1508# 0.01fF
C725 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n4395_1648# 0.00fF
C726 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR 0.03fF
C727 a_n2290_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C728 a_n432_n5274# a_425_n4664# 0.00fF
C729 a_425_n1508# a_575_n3696# 0.00fF
C730 a_n787_n2786# a_n787_n3696# 0.01fF
C731 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_n2345_n2786# 0.00fF
C732 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n732_n5274# 0.00fF
C733 a_425_n540# a_425_n1508# 0.01fF
C734 a_n787_n540# a_n732_n1508# 0.00fF
C735 a_n432_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.01fF
C736 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.01fF
C737 a_275_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.01fF
C738 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_425_n6852# 0.00fF
C739 a_n2195_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C740 a_n2345_n6852# a_n787_n6852# 0.01fF
C741 a_425_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.01fF
C742 a_575_n3696# a_n787_n3696# 0.00fF
C743 a_425_n540# a_425_370# 0.01fF
C744 a_n732_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C745 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 13.27fF
C746 a_275_n2786# a_425_n2118# 0.00fF
C747 a_n4695_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C748 a_n4395_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C749 a_n2140_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.14fF
C750 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n2495_n10008# 0.15fF
C751 a_n1990_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C752 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR a_n732_n1508# 0.01fF
C753 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_425_1038# 0.01fF
C754 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR 0.02fF
C755 a_n2345_n6852# a_n1990_n7820# 0.00fF
C756 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A a_n787_370# 0.00fF
C757 a_n1990_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C758 a_n1990_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C759 a_n432_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT 0.01fF
C760 a_n732_n8430# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.00fF
C761 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A a_n1990_n5274# 0.00fF
C762 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C763 a_n2140_n5274# a_n732_n5274# 0.00fF
C764 a_n787_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A 0.02fF
C765 a_n2495_n3696# a_n2290_n2118# 0.00fF
C766 a_n2045_n5942# a_n787_n6852# 0.00fF
C767 a_n2345_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C768 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_425_n10008# 0.00fF
C769 a_n2195_n2786# a_n787_n3696# 0.00fF
C770 a_n2140_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.05fF
C771 a_n787_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C772 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_425_n5274# 0.01fF
C773 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_n787_n10008# 0.01fF
C774 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT 0.02fF
C775 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 11.92fF
C776 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_425_n7820# 0.00fF
C777 a_275_n9098# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.12fF
C778 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.42fF
C779 a_1637_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B 0.01fF
C780 a_n1990_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C781 a_n732_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C782 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 1.29fF
C783 a_n4395_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C784 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n4695_n540# 0.00fF
C785 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n2345_n6852# 0.00fF
C786 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n1990_n8430# 0.00fF
C787 a_275_n9098# a_n787_n9098# 0.00fF
C788 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C789 a_n4395_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C790 a_n732_n4664# a_n2140_n5274# 0.00fF
C791 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n787_370# 0.00fF
C792 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n1990_1038# 0.01fF
C793 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A a_n2290_n5274# 0.00fF
C794 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n1990_370# 0.00fF
C795 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_425_n4664# 0.02fF
C796 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B a_425_370# 0.00fF
C797 a_n787_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C798 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.03fF
C799 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n2495_n10008# 0.00fF
C800 a_n2290_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C801 a_n2290_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C802 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n1990_n2118# 0.00fF
C803 a_n1990_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.03fF
C804 a_n1990_n540# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A 0.00fF
C805 a_n2195_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.00fF
C806 a_n2140_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.18fF
C807 a_n1990_n4664# a_n2140_n5274# 0.03fF
C808 a_n787_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C809 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.04fF
C810 a_275_n5942# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.01fF
C811 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C812 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 12.50fF
C813 a_n4695_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C814 a_n2290_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C815 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C816 a_n4395_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C817 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n4695_n540# 0.00fF
C818 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n4395_n2118# 0.00fF
C819 a_n732_n7820# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.02fF
C820 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.00fF
C821 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n1990_370# 0.00fF
C822 a_n787_n6852# CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.10fF
C823 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.06fF
C824 a_n4695_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C825 a_n2195_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C826 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.00fF
C827 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.04fF
C828 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR 0.03fF
C829 a_n4395_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C830 a_n787_n6852# a_n732_n7820# 0.00fF
C831 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_425_n7820# 0.00fF
C832 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.44fF
C833 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.05fF
C834 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar a_n1990_n5274# 0.01fF
C835 a_n2290_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.00fF
C836 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_425_n540# 0.04fF
C837 a_n787_n6852# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.01fF
C838 a_n787_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND 0.00fF
C839 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND a_n787_n9098# 0.00fF
C840 a_n787_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C841 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C842 a_425_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C843 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_575_n3696# 0.00fF
C844 a_n2290_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.00fF
C845 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C846 a_n2140_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.15fF
C847 a_n4695_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C848 a_n2140_n5274# a_n2195_n2786# 0.00fF
C849 a_425_n1508# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.00fF
C850 a_n2195_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C851 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_n787_n540# 0.01fF
C852 a_n2345_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C853 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_n1990_n8430# 0.00fF
C854 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n2140_n8430# 0.13fF
C855 a_n787_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C856 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A a_425_370# 0.01fF
C857 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2290_n1508# 0.01fF
C858 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n2290_n5274# 0.01fF
C859 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar a_n1990_n1508# 0.01fF
C860 a_n4395_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C861 a_425_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C862 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.35fF
C863 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n2290_1038# 0.00fF
C864 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_n2290_1648# 0.02fF
C865 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.02fF
C866 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n432_n8430# 0.00fF
C867 a_n2140_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.04fF
C868 a_n432_n4664# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.03fF
C869 a_n2140_n2118# a_n2140_n540# 0.02fF
C870 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A a_n732_n5274# 0.01fF
C871 a_275_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.01fF
C872 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n432_n7820# 0.01fF
C873 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n4395_1038# 0.00fF
C874 a_n2345_n6852# a_n2290_n8430# 0.00fF
C875 a_n4695_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C876 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.74fF
C877 a_n2495_n10008# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.11fF
C878 a_n4395_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C879 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT 0.00fF
C880 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.05fF
C881 a_n2290_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C882 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_425_n1508# 0.01fF
C883 a_n2195_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C884 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_n787_1038# 0.07fF
C885 a_425_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C886 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_425_n4664# 0.00fF
C887 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B 0.00fF
C888 a_425_n540# a_425_n2118# 0.00fF
C889 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n2140_n8430# 0.06fF
C890 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n1990_1038# 0.00fF
C891 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_n432_n5274# 0.00fF
C892 a_n2290_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C893 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.04fF
C894 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n1990_n2118# 0.00fF
C895 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n787_n3696# 0.06fF
C896 a_n732_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C897 a_n2195_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C898 a_n1990_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C899 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B 0.00fF
C900 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n1990_n1508# 0.01fF
C901 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n4395_1648# 0.00fF
C902 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A a_425_n4664# 0.09fF
C903 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C904 a_425_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C905 a_n787_1648# a_n787_n540# 0.00fF
C906 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT a_n2495_n3696# 0.05fF
C907 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n732_n8430# 0.00fF
C908 a_n4695_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C909 a_n732_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C910 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 1.24fF
C911 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.90fF
C912 a_n1990_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C913 a_425_n540# a_425_1648# 0.01fF
C914 a_n787_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C915 a_n2345_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C916 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n787_370# 0.01fF
C917 a_425_n1508# a_425_370# 0.00fF
C918 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n432_n7820# 0.00fF
C919 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2495_n10008# 0.09fF
C920 a_275_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C921 a_n1990_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C922 a_n2345_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C923 a_n787_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C924 a_275_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C925 a_425_n7820# a_575_n6852# 0.00fF
C926 a_n1990_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C927 a_n2140_n2118# a_n732_n1508# 0.00fF
C928 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A a_n432_n8430# 0.01fF
C929 a_275_n2786# a_425_n3696# 0.02fF
C930 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B 0.09fF
C931 a_n2140_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.16fF
C932 a_n787_1038# a_425_1038# 0.00fF
C933 a_n2290_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C934 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n2140_n8430# 0.08fF
C935 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.00fF
C936 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C937 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.00fF
C938 a_425_n7820# a_425_n6852# 0.00fF
C939 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n1990_n5274# 0.01fF
C940 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 11.03fF
C941 a_n787_1648# a_n787_1038# 0.01fF
C942 a_n432_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C943 a_n4395_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C944 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_425_n7820# 0.01fF
C945 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT a_n2495_n10008# 0.05fF
C946 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.14fF
C947 a_n1990_n540# a_n787_n540# 0.00fF
C948 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C949 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.18fF
C950 a_n4395_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C951 a_n4395_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C952 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C953 a_n2140_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.22fF
C954 a_n4695_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C955 a_n4695_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C956 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n732_n2118# 0.01fF
C957 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.62fF
C958 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR a_n732_n8430# 0.00fF
C959 a_n2290_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C960 a_n2195_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C961 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.06fF
C962 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.01fF
C963 a_275_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.02fF
C964 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_1637_1038# 0.00fF
C965 a_425_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B 0.00fF
C966 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR a_n2290_n540# 0.00fF
C967 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT a_425_n7820# 0.00fF
C968 a_275_n9098# CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR 0.00fF
C969 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n4395_1038# 0.00fF
C970 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A 0.32fF
C971 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C972 a_n787_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.00fF
C973 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2140_n5274# 0.06fF
C974 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n2290_n5274# 0.00fF
C975 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n1990_n5274# 0.01fF
C976 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 14.38fF
C977 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C978 a_n1990_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.03fF
C979 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.03fF
C980 a_425_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C981 a_425_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C982 a_n732_n2118# a_425_n1508# 0.00fF
C983 a_425_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C984 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.24fF
C985 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.02fF
C986 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.10fF
C987 a_n2290_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C988 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n2140_n540# 0.04fF
C989 a_n4695_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C990 a_n1990_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.01fF
C991 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.02fF
C992 a_425_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C993 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n4395_n3696# 0.02fF
C994 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B 0.00fF
C995 a_275_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND 0.10fF
C996 a_n2290_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.01fF
C997 a_n732_n2118# a_n787_n3696# 0.00fF
C998 a_n787_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C999 a_n2140_n540# a_n1990_370# 0.01fF
C1000 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n2290_370# 0.01fF
C1001 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n1990_n1508# 0.00fF
C1002 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n4395_1648# 0.00fF
C1003 a_n432_n5274# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.01fF
C1004 a_n432_n7820# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C1005 a_n2195_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C1006 a_n2045_n5942# a_n2345_n6852# 0.01fF
C1007 a_425_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C1008 a_n4695_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C1009 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.00fF
C1010 a_275_n2786# a_425_n4664# 0.01fF
C1011 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n732_n1508# 0.00fF
C1012 a_425_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A 0.00fF
C1013 a_425_1038# a_1637_1038# 0.00fF
C1014 a_n787_n6852# a_n732_n5274# 0.00fF
C1015 a_n2195_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C1016 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n4395_n2118# 0.02fF
C1017 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT a_575_n10008# 0.01fF
C1018 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.12fF
C1019 a_n4695_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.01fF
C1020 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n2495_n10008# 0.04fF
C1021 a_n2140_n2118# a_n2290_n2118# 0.01fF
C1022 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.00fF
C1023 a_n1990_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C1024 a_n2140_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.25fF
C1025 a_n2195_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C1026 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_425_n1508# 0.08fF
C1027 a_n2290_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C1028 a_275_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND 0.12fF
C1029 a_425_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.00fF
C1030 a_n787_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.07fF
C1031 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR a_425_1038# 0.00fF
C1032 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C a_425_n8430# 0.00fF
C1033 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.07fF
C1034 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR 0.00fF
C1035 a_n1990_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C1036 a_n432_n1508# a_n787_n540# 0.00fF
C1037 a_n1990_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C1038 a_n2345_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C1039 a_n787_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR 0.00fF
C1040 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n1990_n7820# 0.01fF
C1041 a_n787_1038# a_n787_n540# 0.01fF
C1042 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n2290_370# 0.00fF
C1043 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_n787_n3696# 0.00fF
C1044 a_n4395_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C1045 a_n2195_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C1046 a_n732_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C1047 a_n432_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.00fF
C1048 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A a_n2290_1038# 0.01fF
C1049 a_n732_n4664# a_n787_n6852# 0.00fF
C1050 a_n4695_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C1051 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 1.22fF
C1052 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_425_n7820# 0.05fF
C1053 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n432_n7820# 0.03fF
C1054 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.15fF
C1055 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n732_n1508# 0.00fF
C1056 a_n787_1038# a_n2290_1648# 0.00fF
C1057 a_n432_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.01fF
C1058 a_n2345_n6852# a_n2290_n7820# 0.00fF
C1059 a_n2290_n8430# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C1060 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C1061 a_1637_1648# CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A 0.01fF
C1062 a_n732_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C1063 a_n4395_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C1064 a_275_n9098# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C1065 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR a_n732_n5274# 0.00fF
C1066 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2195_n9098# 0.00fF
C1067 a_n787_n6852# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.05fF
C1068 a_425_n10008# a_n787_n10008# 0.00fF
C1069 a_425_n2118# a_425_n1508# 0.01fF
C1070 a_n2345_n6852# CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.05fF
C1071 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n2140_n8430# 0.17fF
C1072 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.09fF
C1073 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A 0.04fF
C1074 a_n2345_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.01fF
C1075 a_n2290_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.02fF
C1076 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar a_n1990_n7820# 0.00fF
C1077 a_n4695_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C1078 a_n4695_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.02fF
C1079 a_n2140_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.05fF
C1080 a_n787_n5942# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C1081 a_n432_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR 0.00fF
C1082 a_425_n4664# a_n732_n5274# 0.00fF
C1083 a_1637_1648# a_425_1648# 0.00fF
C1084 a_n432_n5274# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C1085 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.00fF
C1086 a_n2045_n5942# CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C 0.00fF
C1087 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT a_n2195_n9098# 0.00fF
C1088 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B a_n732_n8430# 0.01fF
C1089 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.01fF
C1090 a_425_n7820# a_575_n10008# 0.00fF
C1091 a_n432_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.00fF
C1092 a_n732_n4664# CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR 0.01fF
C1093 a_n2290_n1508# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C1094 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.87fF
C1095 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n787_370# 0.01fF
C1096 a_425_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.00fF
C1097 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n1990_1038# 0.00fF
C1098 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT a_n2140_n8430# 0.01fF
C1099 a_n4395_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C1100 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A a_n4695_n540# 0.02fF
C1101 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.05fF
C1102 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND a_n732_n2118# 0.00fF
C1103 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C1104 a_425_1648# a_425_370# 0.00fF
C1105 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B a_n1990_n2118# 0.01fF
C1106 a_n2140_n540# a_n787_370# 0.00fF
C1107 a_n1990_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C1108 a_n787_n6852# CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND 0.07fF
C1109 a_n2495_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.08fF
C1110 a_n2140_n540# a_n1990_1038# 0.00fF
C1111 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND 0.00fF
C1112 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A a_n1990_n2118# 0.00fF
C1113 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.04fF
C1114 a_n1990_n4664# CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR 0.00fF
C1115 a_n4695_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C1116 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar a_n2290_n2118# 0.00fF
C1117 a_n4395_1038# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.02fF
C1118 a_n1990_1648# a_n2140_n540# 0.00fF
C1119 a_n2345_n6852# a_n1990_n8430# 0.00fF
C1120 a_n732_n4664# a_425_n4664# 0.00fF
C1121 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A 0.00fF
C1122 a_n4695_370# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.00fF
C1123 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar a_n1990_n5274# 0.01fF
C1124 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 1.04fF
C1125 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.01fF
C1126 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.00fF
C1127 a_425_n8430# CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND 0.01fF
C1128 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.15fF
C1129 a_n732_n7820# a_n787_n10008# 0.00fF
C1130 a_n1990_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar 0.00fF
C1131 a_275_n5942# a_575_n6852# 0.02fF
C1132 a_n2495_n3696# a_n2290_n5274# 0.00fF
C1133 a_n1990_n7820# CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR 0.00fF
C1134 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.01fF
C1135 a_n2140_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.14fF
C1136 a_n2140_n2118# a_n2495_n3696# 0.01fF
C1137 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.00fF
C1138 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND a_n787_n6852# 0.00fF
C1139 a_n4695_n2786# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar 0.00fF
C1140 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT a_275_n9098# 0.05fF
C1141 a_425_n4664# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar 0.05fF
C1142 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar 0.02fF
C1143 a_n2195_n9098# a_n2495_n10008# 0.01fF
C1144 a_n2140_n540# CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A 0.00fF
C1145 a_n787_n3696# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.03fF
C1146 a_n2140_n8430# a_n2495_n10008# 0.01fF
C1147 a_275_n5942# a_425_n6852# 0.02fF
C1148 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A a_n1990_n1508# 0.00fF
C1149 a_n4395_1648# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A 0.02fF
C1150 a_425_n2118# CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A 0.00fF
C1151 a_n2290_n540# CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B 0.01fF
C1152 a_575_n10008# GND 0.02fF
C1153 a_425_n10008# GND 0.02fF
C1154 a_n787_n9098# GND 0.03fF
C1155 a_n2195_n9098# GND 0.03fF
C1156 a_n2345_n9098# GND 0.03fF
C1157 a_275_n9098# GND 0.94fF
C1158 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT GND 0.88fF $ **FLOATING
C1159 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/AND GND 0.58fF
C1160 a_n787_n10008# GND 0.50fF
C1161 a_n2495_n10008# GND 0.71fF
C1162 a_425_n8430# GND 0.03fF
C1163 a_n432_n8430# GND 0.03fF
C1164 a_n732_n8430# GND 0.02fF
C1165 a_n1990_n8430# GND 0.02fF
C1166 a_n2290_n8430# GND 0.02fF
C1167 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/AND GND 1.99fF
C1168 a_n432_n7820# GND 0.01fF
C1169 a_n732_n7820# GND 0.01fF
C1170 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/XNOR GND 1.10fF
C1171 a_n1990_n7820# GND 0.01fF
C1172 a_n2290_n7820# GND 0.01fF
C1173 a_425_n7820# GND 0.52fF
C1174 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/A GND 1.13fF
C1175 a_n2140_n8430# GND 0.59fF
C1176 a_575_n6852# GND 0.02fF
C1177 a_425_n6852# GND 0.02fF
C1178 a_n787_n5942# GND 0.03fF
C1179 a_n2045_n5942# GND 0.03fF
C1180 a_n2195_n5942# GND 0.03fF
C1181 a_n2345_n5942# GND 0.03fF
C1182 a_275_n5942# GND 0.90fF
C1183 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C GND 1.13fF $ **FLOATING
C1184 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/AND GND 0.56fF
C1185 a_n787_n6852# GND 0.46fF
C1186 a_n2345_n6852# GND 0.47fF
C1187 a_425_n5274# GND 0.03fF
C1188 a_n432_n5274# GND 0.03fF
C1189 a_n732_n5274# GND 0.02fF
C1190 a_n1990_n5274# GND 0.02fF
C1191 a_n2290_n5274# GND 0.02fF
C1192 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/AND GND 1.98fF
C1193 a_n432_n4664# GND 0.01fF
C1194 a_n732_n4664# GND 0.01fF
C1195 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/XNOR GND 1.08fF
C1196 a_n1990_n4664# GND 0.01fF
C1197 a_n2290_n4664# GND 0.01fF
C1198 a_425_n4664# GND 0.52fF
C1199 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/A GND 1.13fF
C1200 a_n2140_n5274# GND 0.59fF
C1201 a_575_n3696# GND 0.02fF
C1202 a_425_n3696# GND 0.02fF
C1203 a_n4395_n3696# GND 0.01fF
C1204 a_n4695_n3696# GND 0.01fF
C1205 a_n787_n2786# GND 0.03fF
C1206 a_n2195_n2786# GND 0.03fF
C1207 a_n2345_n2786# GND 0.03fF
C1208 a_n4395_n2786# GND 0.02fF
C1209 a_n4695_n2786# GND 0.01fF
C1210 a_275_n2786# GND 0.90fF
C1211 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT GND 0.93fF $ **FLOATING
C1212 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/AND GND 0.56fF
C1213 a_n787_n3696# GND 0.47fF
C1214 a_n2495_n3696# GND 0.60fF
C1215 a_425_n2118# GND 0.02fF
C1216 a_n432_n2118# GND 0.03fF
C1217 a_n732_n2118# GND 0.02fF
C1218 a_n1990_n2118# GND 0.02fF
C1219 a_n2290_n2118# GND 0.02fF
C1220 a_n4395_n2118# GND 0.01fF
C1221 a_n4695_n2118# GND 0.01fF
C1222 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/AND GND 1.95fF
C1223 a_n432_n1508# GND 0.01fF
C1224 a_n732_n1508# GND 0.01fF
C1225 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/XNOR GND 1.08fF
C1226 a_n1990_n1508# GND 0.01fF
C1227 a_n2290_n1508# GND 0.01fF
C1228 a_n4395_n1508# GND 0.00fF
C1229 a_n4695_n1508# GND 0.00fF
C1230 a_425_n1508# GND 0.51fF
C1231 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/A GND 1.12fF
C1232 a_n2140_n2118# GND 0.58fF
C1233 a_n1990_n540# GND 0.00fF
C1234 a_n2290_n540# GND 0.00fF
C1235 a_n4395_n540# GND 0.00fF
C1236 a_n4695_n540# GND 0.00fF
C1237 a_425_370# GND 0.03fF
C1238 a_n787_370# GND 0.03fF
C1239 a_n1990_370# GND 0.02fF
C1240 a_n2290_370# GND 0.01fF
C1241 a_n4395_370# GND 0.01fF
C1242 a_n4695_370# GND 0.01fF
C1243 a_425_n540# GND 0.52fF
C1244 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/XNOR GND 0.87fF
C1245 a_n787_n540# GND 0.47fF
C1246 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar GND 5.75fF $ **FLOATING
C1247 a_n2140_n540# GND 0.54fF
C1248 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_1/A GND 0.95fF
C1249 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B GND 6.01fF $ **FLOATING
C1250 a_425_1038# GND 0.03fF
C1251 a_n1990_1038# GND 0.02fF
C1252 a_n2290_1038# GND 0.01fF
C1253 a_n4395_1038# GND 0.01fF
C1254 a_n4695_1038# GND 0.01fF
C1255 a_1637_1648# GND 0.02fF
C1256 a_n787_1648# GND 0.01fF
C1257 a_n1990_1648# GND 0.00fF
C1258 a_n2290_1648# GND 0.00fF
C1259 a_n4395_1648# GND 0.00fF
C1260 a_n4695_1648# GND 0.00fF
C1261 a_1637_1038# GND 0.67fF
C1262 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/B GND 1.28fF
C1263 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/A GND 0.64fF
C1264 a_425_1648# GND 0.50fF
C1265 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/A GND 1.60fF
C1266 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/OR GND 0.57fF
C1267 a_n787_1038# GND 0.61fF
C1268 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar GND 7.15fF $ **FLOATING
C1269 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A GND 8.47fF $ **FLOATING
C1270 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar GND 7.23fF $ **FLOATING
C1271 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar GND 14.03fF $ **FLOATING
C1272 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A GND 7.51fF $ **FLOATING
C1273 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B GND 4.18fF $ **FLOATING
C1274 CMOS_4in_XOR_0/XOR1_bar GND 0.53fF $ **FLOATING
C1275 CMOS_sbox_0/CMOS_s0_0/x1_bar GND 1.66fF $ **FLOATING
C1276 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t1 GND 0.67fF
C1277 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t6 GND 0.40fF
C1278 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t7 GND 0.35fF
C1279 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/A_bar GND 0.79fF $ **FLOATING
C1280 CMOS_sbox_0/CMOS_s3_0/x1_bar GND 6.20fF $ **FLOATING
C1281 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t10 GND 0.17fF
C1282 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t8 GND 0.25fF
C1283 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n0 GND 0.35fF $ **FLOATING
C1284 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_1/B GND 0.05fF $ **FLOATING
C1285 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n1 GND 0.90fF $ **FLOATING
C1286 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n2 GND 2.55fF $ **FLOATING
C1287 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t4 GND 0.40fF
C1288 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t9 GND 0.35fF
C1289 CMOS_sbox_0/CMOS_s2_0/CMOS_XOR_0/A_bar GND 0.66fF $ **FLOATING
C1290 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n3 GND 4.24fF $ **FLOATING
C1291 CMOS_sbox_0/CMOS_s2_0/x1_bar GND 2.35fF $ **FLOATING
C1292 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t11 GND 0.40fF
C1293 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t5 GND 0.35fF
C1294 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n4 GND 4.93fF $ **FLOATING
C1295 CMOS_sbox_0/CMOS_s1_0/x1_bar GND 1.42fF $ **FLOATING
C1296 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t3 GND 0.17fF
C1297 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t2 GND 0.25fF
C1298 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n5 GND 0.35fF $ **FLOATING
C1299 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_2/B GND 0.59fF $ **FLOATING
C1300 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n6 GND 3.57fF $ **FLOATING
C1301 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n7 GND 2.52fF $ **FLOATING
C1302 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.n8 GND 0.57fF $ **FLOATING
C1303 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A_bar.t0 GND 1.71fF
C1304 CMOS_4in_XOR_0/CMOS_INV_1/OUT GND 0.63fF $ **FLOATING
C1305 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t2 GND 0.10fF
C1306 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t3 GND 0.12fF
C1307 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t0 GND 0.31fF
C1308 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.t1 GND 0.29fF
C1309 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/OUT.n0 GND 0.70fF $ **FLOATING
C1310 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_OR_0/C GND 0.42fF $ **FLOATING
C1311 CMOS_4in_XOR_0/XOR2_bar GND 0.48fF $ **FLOATING
C1312 CMOS_sbox_0/CMOS_s0_0/x2_bar GND 1.15fF $ **FLOATING
C1313 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t0 GND 1.65fF
C1314 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t2 GND 0.23fF
C1315 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t5 GND 0.16fF
C1316 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n0 GND 0.32fF $ **FLOATING
C1317 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/B GND 0.04fF $ **FLOATING
C1318 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n1 GND 1.52fF $ **FLOATING
C1319 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t8 GND 0.23fF
C1320 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t11 GND 0.16fF
C1321 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n2 GND 0.32fF $ **FLOATING
C1322 CMOS_sbox_0/CMOS_s2_0/CMOS_AND_0/B GND 0.04fF $ **FLOATING
C1323 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n3 GND 1.52fF $ **FLOATING
C1324 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t4 GND 0.37fF
C1325 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t10 GND 0.33fF
C1326 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/A_bar GND 0.59fF $ **FLOATING
C1327 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t15 GND 0.26fF
C1328 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t13 GND 0.31fF
C1329 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/A GND 0.04fF $ **FLOATING
C1330 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n4 GND 0.47fF $ **FLOATING
C1331 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n5 GND 6.64fF $ **FLOATING
C1332 CMOS_sbox_0/CMOS_s3_0/x2_bar GND 2.15fF $ **FLOATING
C1333 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n6 GND 3.77fF $ **FLOATING
C1334 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t12 GND 0.27fF
C1335 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t7 GND 0.27fF
C1336 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n7 GND 0.72fF $ **FLOATING
C1337 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/B_bar GND 0.25fF $ **FLOATING
C1338 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n8 GND 1.81fF $ **FLOATING
C1339 CMOS_sbox_0/CMOS_s2_0/x2_bar GND 1.46fF $ **FLOATING
C1340 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n9 GND 3.56fF $ **FLOATING
C1341 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t3 GND 0.34fF
C1342 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t9 GND 0.28fF
C1343 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/B GND 0.56fF $ **FLOATING
C1344 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n10 GND 4.32fF $ **FLOATING
C1345 CMOS_sbox_0/CMOS_s1_0/x2_bar GND 1.79fF $ **FLOATING
C1346 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t6 GND 0.27fF
C1347 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t14 GND 0.27fF
C1348 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n11 GND 0.72fF $ **FLOATING
C1349 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n12 GND 1.24fF $ **FLOATING
C1350 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n13 GND 1.18fF $ **FLOATING
C1351 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n14 GND 0.11fF $ **FLOATING
C1352 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.t1 GND 0.63fF
C1353 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B_bar.n15 GND 0.50fF $ **FLOATING
C1354 CMOS_4in_XOR_0/CMOS_INV_3/OUT GND 0.56fF $ **FLOATING
C1355 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t3 GND 0.11fF
C1356 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t2 GND 0.14fF
C1357 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t0 GND 0.37fF
C1358 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.t1 GND 0.34fF
C1359 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/OUT GND 0.23fF $ **FLOATING
C1360 CMOS_sbox_0/CMOS_s2_0/CMOS_3in_OR_0/C.n0 GND 0.82fF $ **FLOATING
C1361 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n0 GND 0.29fF $ **FLOATING
C1362 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n1 GND 0.31fF $ **FLOATING
C1363 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n2 GND 0.08fF $ **FLOATING
C1364 CMOS_sbox_0/CMOS_s0_0/x1 GND 0.15fF $ **FLOATING
C1365 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t15 GND 0.12fF
C1366 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t16 GND 0.18fF
C1367 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n3 GND 0.25fF $ **FLOATING
C1368 CMOS_4in_XOR_0/CMOS_INV_1/A GND 0.14fF $ **FLOATING
C1369 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t19 GND 0.24fF
C1370 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t17 GND 0.09fF
C1371 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n4 GND 0.27fF $ **FLOATING
C1372 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n5 GND 1.35fF $ **FLOATING
C1373 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t10 GND 0.27fF
C1374 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t14 GND 0.22fF
C1375 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n6 GND 0.35fF $ **FLOATING
C1376 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/B GND 0.35fF $ **FLOATING
C1377 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t8 GND 0.18fF
C1378 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t11 GND 0.12fF
C1379 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n7 GND 0.25fF $ **FLOATING
C1380 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/B GND 0.03fF $ **FLOATING
C1381 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n8 GND 1.57fF $ **FLOATING
C1382 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t4 GND 0.24fF
C1383 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t7 GND 0.09fF
C1384 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n9 GND 0.27fF $ **FLOATING
C1385 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/A GND 0.35fF $ **FLOATING
C1386 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n10 GND 4.93fF $ **FLOATING
C1387 CMOS_sbox_0/CMOS_s3_0/x1 GND 1.34fF $ **FLOATING
C1388 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t9 GND 0.24fF
C1389 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t5 GND 0.09fF
C1390 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n11 GND 0.27fF $ **FLOATING
C1391 CMOS_sbox_0/CMOS_s2_0/CMOS_XOR_0/A GND 0.03fF $ **FLOATING
C1392 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n12 GND 1.29fF $ **FLOATING
C1393 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t13 GND 0.27fF
C1394 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t18 GND 0.22fF
C1395 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n13 GND 0.33fF $ **FLOATING
C1396 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/B GND 0.38fF $ **FLOATING
C1397 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n14 GND 2.30fF $ **FLOATING
C1398 CMOS_sbox_0/CMOS_s2_0/x1 GND 1.71fF $ **FLOATING
C1399 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n15 GND 2.25fF $ **FLOATING
C1400 CMOS_sbox_0/CMOS_s1_0/x1 GND 1.44fF $ **FLOATING
C1401 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t6 GND 0.18fF
C1402 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t12 GND 0.12fF
C1403 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n16 GND 0.25fF $ **FLOATING
C1404 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/A GND 0.48fF $ **FLOATING
C1405 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n17 GND 3.20fF $ **FLOATING
C1406 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n18 GND 1.86fF $ **FLOATING
C1407 CMOS_4in_XOR_0/XOR1 GND 0.30fF $ **FLOATING
C1408 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n19 GND 0.35fF $ **FLOATING
C1409 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n20 GND 0.04fF $ **FLOATING
C1410 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n21 GND 0.12fF $ **FLOATING
C1411 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n22 GND 0.05fF $ **FLOATING
C1412 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n23 GND 0.02fF $ **FLOATING
C1413 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n24 GND 0.01fF $ **FLOATING
C1414 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n25 GND 0.04fF $ **FLOATING
C1415 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n26 GND 0.04fF $ **FLOATING
C1416 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n27 GND 0.04fF $ **FLOATING
C1417 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n28 GND 0.15fF $ **FLOATING
C1418 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n29 GND 0.02fF $ **FLOATING
C1419 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t2 GND 0.12fF
C1420 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t3 GND 0.12fF
C1421 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n30 GND 0.25fF $ **FLOATING
C1422 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n31 GND 0.05fF $ **FLOATING
C1423 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n32 GND 0.01fF $ **FLOATING
C1424 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n33 GND 0.33fF $ **FLOATING
C1425 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n34 GND 0.06fF $ **FLOATING
C1426 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n35 GND 0.02fF $ **FLOATING
C1427 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n36 GND 0.01fF $ **FLOATING
C1428 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n37 GND 0.04fF $ **FLOATING
C1429 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n38 GND 0.01fF $ **FLOATING
C1430 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n39 GND 0.32fF $ **FLOATING
C1431 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n40 GND 0.08fF $ **FLOATING
C1432 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n41 GND 0.08fF $ **FLOATING
C1433 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n42 GND 0.16fF $ **FLOATING
C1434 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n43 GND 0.01fF $ **FLOATING
C1435 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n44 GND 0.04fF $ **FLOATING
C1436 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n45 GND 0.04fF $ **FLOATING
C1437 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n46 GND 0.04fF $ **FLOATING
C1438 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t0 GND 0.24fF
C1439 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.t1 GND 0.24fF
C1440 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n47 GND 0.49fF $ **FLOATING
C1441 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n48 GND 0.00fF $ **FLOATING
C1442 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n49 GND 0.04fF $ **FLOATING
C1443 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n50 GND 0.01fF $ **FLOATING
C1444 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n51 GND 0.04fF $ **FLOATING
C1445 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n52 GND 0.02fF $ **FLOATING
C1446 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n53 GND 0.01fF $ **FLOATING
C1447 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n54 GND 0.01fF $ **FLOATING
C1448 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n55 GND 0.04fF $ **FLOATING
C1449 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n56 GND 0.02fF $ **FLOATING
C1450 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n57 GND 0.01fF $ **FLOATING
C1451 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n58 GND 0.01fF $ **FLOATING
C1452 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n59 GND 0.02fF $ **FLOATING
C1453 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n60 GND 0.03fF $ **FLOATING
C1454 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/A.n61 GND 0.20fF $ **FLOATING
C1455 CMOS_4in_XOR_0/CMOS_XOR_2/XOR GND 0.12fF $ **FLOATING
C1456 CMOS_4in_XOR_0/XOR0_bar GND 0.37fF $ **FLOATING
C1457 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t0 GND 1.36fF
C1458 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t5 GND 0.31fF
C1459 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t7 GND 0.27fF
C1460 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t10 GND 0.22fF
C1461 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t4 GND 0.22fF
C1462 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n0 GND 0.59fF $ **FLOATING
C1463 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/B_bar GND 0.35fF $ **FLOATING
C1464 CMOS_sbox_0/CMOS_s3_0/x0_bar GND 5.20fF $ **FLOATING
C1465 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t9 GND 0.22fF
C1466 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t2 GND 0.20fF
C1467 CMOS_sbox_0/CMOS_s2_0/CMOS_XOR_0/B_bar GND 0.03fF $ **FLOATING
C1468 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n1 GND 1.51fF $ **FLOATING
C1469 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n2 GND 3.24fF $ **FLOATING
C1470 CMOS_sbox_0/CMOS_s2_0/x0_bar GND 1.35fF $ **FLOATING
C1471 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t8 GND 0.13fF
C1472 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t3 GND 0.20fF
C1473 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n3 GND 0.23fF $ **FLOATING
C1474 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/C GND 0.39fF $ **FLOATING
C1475 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n4 GND 1.60fF $ **FLOATING
C1476 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n5 GND 2.01fF $ **FLOATING
C1477 CMOS_sbox_0/CMOS_s1_0/x0_bar GND 1.33fF $ **FLOATING
C1478 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t13 GND 0.22fF
C1479 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t6 GND 0.22fF
C1480 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n6 GND 0.59fF $ **FLOATING
C1481 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/B_bar GND 0.34fF $ **FLOATING
C1482 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n7 GND 1.62fF $ **FLOATING
C1483 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t11 GND 0.31fF
C1484 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t12 GND 0.27fF
C1485 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/A_bar GND 0.66fF $ **FLOATING
C1486 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n8 GND 1.43fF $ **FLOATING
C1487 CMOS_sbox_0/CMOS_s0_0/x0_bar GND 0.71fF $ **FLOATING
C1488 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n9 GND 0.94fF $ **FLOATING
C1489 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.t1 GND 0.52fF
C1490 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A_bar.n10 GND 0.43fF $ **FLOATING
C1491 CMOS_4in_XOR_0/CMOS_INV_2/OUT GND 0.47fF $ **FLOATING
C1492 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n0 GND 0.29fF $ **FLOATING
C1493 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n1 GND 0.30fF $ **FLOATING
C1494 CMOS_sbox_0/CMOS_s0_0/x3 GND 0.14fF $ **FLOATING
C1495 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n2 GND 0.08fF $ **FLOATING
C1496 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t6 GND 0.12fF
C1497 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t19 GND 0.18fF
C1498 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n3 GND 0.25fF $ **FLOATING
C1499 CMOS_4in_XOR_0/CMOS_INV_0/A GND 0.14fF $ **FLOATING
C1500 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t14 GND 0.68fF
C1501 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t15 GND 0.46fF
C1502 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/B GND 0.48fF $ **FLOATING
C1503 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n4 GND 1.62fF $ **FLOATING
C1504 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t4 GND 0.09fF
C1505 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t7 GND 0.24fF
C1506 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n5 GND 0.26fF $ **FLOATING
C1507 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/A GND 0.23fF $ **FLOATING
C1508 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n6 GND 2.01fF $ **FLOATING
C1509 CMOS_sbox_0/CMOS_s1_0/x3 GND 0.65fF $ **FLOATING
C1510 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t5 GND 0.68fF
C1511 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t8 GND 0.46fF
C1512 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B GND 0.44fF $ **FLOATING
C1513 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n7 GND 2.77fF $ **FLOATING
C1514 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n8 GND 1.20fF $ **FLOATING
C1515 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t17 GND 0.12fF
C1516 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t12 GND 0.18fF
C1517 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n9 GND 0.25fF $ **FLOATING
C1518 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n10 GND 0.50fF $ **FLOATING
C1519 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t16 GND 0.12fF
C1520 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t18 GND 0.18fF
C1521 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n11 GND 0.22fF $ **FLOATING
C1522 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/C GND 0.26fF $ **FLOATING
C1523 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t10 GND 0.68fF
C1524 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t13 GND 0.46fF
C1525 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/B GND 0.44fF $ **FLOATING
C1526 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n12 GND 5.26fF $ **FLOATING
C1527 CMOS_sbox_0/CMOS_s3_0/x3 GND 1.22fF $ **FLOATING
C1528 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t9 GND 0.24fF
C1529 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t11 GND 0.09fF
C1530 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n13 GND 0.26fF $ **FLOATING
C1531 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/A GND 0.23fF $ **FLOATING
C1532 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n14 GND 2.07fF $ **FLOATING
C1533 CMOS_sbox_0/CMOS_s2_0/x3 GND 1.01fF $ **FLOATING
C1534 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n15 GND 0.50fF $ **FLOATING
C1535 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n16 GND 0.95fF $ **FLOATING
C1536 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n17 GND 0.30fF $ **FLOATING
C1537 CMOS_4in_XOR_0/XOR3 GND 0.29fF $ **FLOATING
C1538 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n18 GND 0.35fF $ **FLOATING
C1539 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n19 GND 0.04fF $ **FLOATING
C1540 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n20 GND 0.12fF $ **FLOATING
C1541 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n21 GND 0.05fF $ **FLOATING
C1542 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n22 GND 0.02fF $ **FLOATING
C1543 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n23 GND 0.01fF $ **FLOATING
C1544 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n24 GND 0.04fF $ **FLOATING
C1545 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n25 GND 0.04fF $ **FLOATING
C1546 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n26 GND 0.04fF $ **FLOATING
C1547 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n27 GND 0.15fF $ **FLOATING
C1548 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n28 GND 0.02fF $ **FLOATING
C1549 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t3 GND 0.12fF
C1550 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t2 GND 0.12fF
C1551 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n29 GND 0.24fF $ **FLOATING
C1552 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n30 GND 0.05fF $ **FLOATING
C1553 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n31 GND 0.01fF $ **FLOATING
C1554 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n32 GND 0.33fF $ **FLOATING
C1555 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n33 GND 0.05fF $ **FLOATING
C1556 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n34 GND 0.02fF $ **FLOATING
C1557 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n35 GND 0.01fF $ **FLOATING
C1558 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n36 GND 0.03fF $ **FLOATING
C1559 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n37 GND 0.01fF $ **FLOATING
C1560 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n38 GND 0.32fF $ **FLOATING
C1561 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n39 GND 0.08fF $ **FLOATING
C1562 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n40 GND 0.08fF $ **FLOATING
C1563 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n41 GND 0.15fF $ **FLOATING
C1564 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n42 GND 0.01fF $ **FLOATING
C1565 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n43 GND 0.04fF $ **FLOATING
C1566 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n44 GND 0.04fF $ **FLOATING
C1567 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n45 GND 0.04fF $ **FLOATING
C1568 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t0 GND 0.24fF
C1569 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.t1 GND 0.24fF
C1570 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n46 GND 0.48fF $ **FLOATING
C1571 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n47 GND 0.00fF $ **FLOATING
C1572 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n48 GND 0.04fF $ **FLOATING
C1573 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n49 GND 0.01fF $ **FLOATING
C1574 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n50 GND 0.04fF $ **FLOATING
C1575 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n51 GND 0.02fF $ **FLOATING
C1576 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n52 GND 0.01fF $ **FLOATING
C1577 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n53 GND 0.01fF $ **FLOATING
C1578 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n54 GND 0.03fF $ **FLOATING
C1579 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n55 GND 0.02fF $ **FLOATING
C1580 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n56 GND 0.01fF $ **FLOATING
C1581 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n57 GND 0.01fF $ **FLOATING
C1582 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n58 GND 0.02fF $ **FLOATING
C1583 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n59 GND 0.03fF $ **FLOATING
C1584 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/B.n60 GND 0.19fF $ **FLOATING
C1585 CMOS_4in_XOR_0/CMOS_XOR_1/XOR GND 0.12fF $ **FLOATING
C1586 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t3 GND 0.12fF
C1587 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t2 GND 0.14fF
C1588 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t0 GND 0.38fF
C1589 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.t1 GND 0.35fF
C1590 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/OUT.n0 GND 0.86fF $ **FLOATING
C1591 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_OR_0/C GND 0.51fF $ **FLOATING
C1592 VDD.t114 GND 0.09fF
C1593 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/VDD GND 0.01fF $ **FLOATING
C1594 VDD.n0 GND 0.16fF $ **FLOATING
C1595 VDD.n1 GND 0.02fF $ **FLOATING
C1596 VDD.t134 GND 0.09fF
C1597 VDD.t167 GND 0.09fF
C1598 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_1/VDD GND 0.01fF $ **FLOATING
C1599 VDD.t77 GND 0.09fF
C1600 VDD.t116 GND 0.09fF
C1601 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_0/VDD GND 0.01fF $ **FLOATING
C1602 VDD.t124 GND 0.09fF
C1603 VDD.t118 GND 0.09fF
C1604 CMOS_sbox_0/CMOS_s0_0/CMOS_OR_0/VDD GND 0.01fF $ **FLOATING
C1605 VDD.t66 GND 0.09fF
C1606 VDD.n2 GND 0.26fF $ **FLOATING
C1607 VDD.n3 GND 0.02fF $ **FLOATING
C1608 VDD.n4 GND 0.02fF $ **FLOATING
C1609 VDD.n5 GND 0.20fF $ **FLOATING
C1610 VDD.t65 GND 0.13fF
C1611 VDD.n6 GND 0.13fF $ **FLOATING
C1612 VDD.n7 GND 0.02fF $ **FLOATING
C1613 VDD.n8 GND 0.02fF $ **FLOATING
C1614 VDD.n9 GND 0.07fF $ **FLOATING
C1615 VDD.n10 GND 0.48fF $ **FLOATING
C1616 VDD.n11 GND 0.22fF $ **FLOATING
C1617 VDD.n12 GND 0.02fF $ **FLOATING
C1618 VDD.n13 GND 0.02fF $ **FLOATING
C1619 VDD.n14 GND 0.01fF $ **FLOATING
C1620 VDD.n15 GND 0.22fF $ **FLOATING
C1621 VDD.n16 GND 0.02fF $ **FLOATING
C1622 VDD.n17 GND 0.02fF $ **FLOATING
C1623 VDD.n18 GND 0.02fF $ **FLOATING
C1624 VDD.n19 GND 0.22fF $ **FLOATING
C1625 VDD.n20 GND 0.02fF $ **FLOATING
C1626 VDD.n21 GND 0.02fF $ **FLOATING
C1627 VDD.n22 GND 0.02fF $ **FLOATING
C1628 VDD.n23 GND 0.02fF $ **FLOATING
C1629 VDD.n24 GND 0.22fF $ **FLOATING
C1630 VDD.n25 GND 0.02fF $ **FLOATING
C1631 VDD.n26 GND 0.02fF $ **FLOATING
C1632 VDD.t55 GND 0.11fF
C1633 VDD.n27 GND 0.14fF $ **FLOATING
C1634 VDD.n28 GND 0.02fF $ **FLOATING
C1635 VDD.n29 GND 0.02fF $ **FLOATING
C1636 VDD.n30 GND 0.02fF $ **FLOATING
C1637 VDD.n31 GND 0.19fF $ **FLOATING
C1638 VDD.n32 GND 0.02fF $ **FLOATING
C1639 VDD.n33 GND 0.02fF $ **FLOATING
C1640 VDD.n34 GND 0.02fF $ **FLOATING
C1641 VDD.t117 GND 0.13fF
C1642 VDD.n35 GND 0.15fF $ **FLOATING
C1643 VDD.n36 GND 0.02fF $ **FLOATING
C1644 VDD.n37 GND 0.02fF $ **FLOATING
C1645 VDD.n38 GND 0.02fF $ **FLOATING
C1646 VDD.n39 GND 0.24fF $ **FLOATING
C1647 VDD.n40 GND 0.02fF $ **FLOATING
C1648 VDD.n41 GND 0.02fF $ **FLOATING
C1649 VDD.n42 GND 0.02fF $ **FLOATING
C1650 VDD.n43 GND 0.48fF $ **FLOATING
C1651 VDD.n44 GND 0.23fF $ **FLOATING
C1652 VDD.n45 GND 0.08fF $ **FLOATING
C1653 VDD.n46 GND 0.20fF $ **FLOATING
C1654 VDD.n47 GND 0.08fF $ **FLOATING
C1655 VDD.n48 GND 0.25fF $ **FLOATING
C1656 VDD.n49 GND 0.02fF $ **FLOATING
C1657 VDD.n50 GND 0.02fF $ **FLOATING
C1658 VDD.n51 GND 0.02fF $ **FLOATING
C1659 VDD.t123 GND 0.13fF
C1660 VDD.n52 GND 0.13fF $ **FLOATING
C1661 VDD.n53 GND 0.02fF $ **FLOATING
C1662 VDD.n54 GND 0.02fF $ **FLOATING
C1663 VDD.n55 GND 0.02fF $ **FLOATING
C1664 VDD.n56 GND 0.48fF $ **FLOATING
C1665 VDD.n57 GND 0.22fF $ **FLOATING
C1666 VDD.n58 GND 0.02fF $ **FLOATING
C1667 VDD.n59 GND 0.02fF $ **FLOATING
C1668 VDD.n60 GND 0.01fF $ **FLOATING
C1669 VDD.n61 GND 0.22fF $ **FLOATING
C1670 VDD.n62 GND 0.02fF $ **FLOATING
C1671 VDD.n63 GND 0.02fF $ **FLOATING
C1672 VDD.n64 GND 0.02fF $ **FLOATING
C1673 VDD.n65 GND 0.22fF $ **FLOATING
C1674 VDD.n66 GND 0.02fF $ **FLOATING
C1675 VDD.n67 GND 0.02fF $ **FLOATING
C1676 VDD.n68 GND 0.02fF $ **FLOATING
C1677 VDD.t60 GND 0.09fF
C1678 VDD.n69 GND 0.47fF $ **FLOATING
C1679 VDD.n70 GND 0.01fF $ **FLOATING
C1680 VDD.n71 GND 0.22fF $ **FLOATING
C1681 VDD.n72 GND 0.02fF $ **FLOATING
C1682 VDD.n73 GND 0.02fF $ **FLOATING
C1683 VDD.t59 GND 0.11fF
C1684 VDD.n74 GND 0.14fF $ **FLOATING
C1685 VDD.n75 GND 0.02fF $ **FLOATING
C1686 VDD.n76 GND 0.02fF $ **FLOATING
C1687 VDD.n77 GND 0.02fF $ **FLOATING
C1688 VDD.n78 GND 0.19fF $ **FLOATING
C1689 VDD.n79 GND 0.02fF $ **FLOATING
C1690 VDD.n80 GND 0.02fF $ **FLOATING
C1691 VDD.n81 GND 0.02fF $ **FLOATING
C1692 VDD.t115 GND 0.13fF
C1693 VDD.n82 GND 0.15fF $ **FLOATING
C1694 VDD.n83 GND 0.02fF $ **FLOATING
C1695 VDD.n84 GND 0.02fF $ **FLOATING
C1696 VDD.n85 GND 0.02fF $ **FLOATING
C1697 VDD.n86 GND 0.24fF $ **FLOATING
C1698 VDD.n87 GND 0.02fF $ **FLOATING
C1699 VDD.n88 GND 0.02fF $ **FLOATING
C1700 VDD.n89 GND 0.02fF $ **FLOATING
C1701 VDD.n90 GND 0.48fF $ **FLOATING
C1702 VDD.n91 GND 0.23fF $ **FLOATING
C1703 VDD.n92 GND 0.08fF $ **FLOATING
C1704 VDD.n93 GND 0.20fF $ **FLOATING
C1705 VDD.n94 GND 0.08fF $ **FLOATING
C1706 VDD.n95 GND 0.25fF $ **FLOATING
C1707 VDD.n96 GND 0.02fF $ **FLOATING
C1708 VDD.n97 GND 0.02fF $ **FLOATING
C1709 VDD.n98 GND 0.02fF $ **FLOATING
C1710 VDD.t76 GND 0.13fF
C1711 VDD.n99 GND 0.13fF $ **FLOATING
C1712 VDD.n100 GND 0.02fF $ **FLOATING
C1713 VDD.n101 GND 0.02fF $ **FLOATING
C1714 VDD.n102 GND 0.02fF $ **FLOATING
C1715 VDD.n103 GND 0.48fF $ **FLOATING
C1716 VDD.n104 GND 0.22fF $ **FLOATING
C1717 VDD.n105 GND 0.02fF $ **FLOATING
C1718 VDD.n106 GND 0.02fF $ **FLOATING
C1719 VDD.n107 GND 0.01fF $ **FLOATING
C1720 VDD.n108 GND 0.22fF $ **FLOATING
C1721 VDD.n109 GND 0.02fF $ **FLOATING
C1722 VDD.n110 GND 0.02fF $ **FLOATING
C1723 VDD.n111 GND 0.02fF $ **FLOATING
C1724 VDD.n112 GND 0.22fF $ **FLOATING
C1725 VDD.n113 GND 0.02fF $ **FLOATING
C1726 VDD.n114 GND 0.02fF $ **FLOATING
C1727 VDD.n115 GND 0.02fF $ **FLOATING
C1728 VDD.n116 GND 0.02fF $ **FLOATING
C1729 VDD.n117 GND 0.22fF $ **FLOATING
C1730 VDD.n118 GND 0.02fF $ **FLOATING
C1731 VDD.n119 GND 0.02fF $ **FLOATING
C1732 VDD.t69 GND 0.11fF
C1733 VDD.n120 GND 0.14fF $ **FLOATING
C1734 VDD.n121 GND 0.02fF $ **FLOATING
C1735 VDD.n122 GND 0.02fF $ **FLOATING
C1736 VDD.n123 GND 0.02fF $ **FLOATING
C1737 VDD.n124 GND 0.19fF $ **FLOATING
C1738 VDD.n125 GND 0.02fF $ **FLOATING
C1739 VDD.n126 GND 0.02fF $ **FLOATING
C1740 VDD.n127 GND 0.02fF $ **FLOATING
C1741 VDD.t166 GND 0.13fF
C1742 VDD.n128 GND 0.15fF $ **FLOATING
C1743 VDD.n129 GND 0.02fF $ **FLOATING
C1744 VDD.n130 GND 0.02fF $ **FLOATING
C1745 VDD.n131 GND 0.02fF $ **FLOATING
C1746 VDD.n132 GND 0.24fF $ **FLOATING
C1747 VDD.n133 GND 0.02fF $ **FLOATING
C1748 VDD.n134 GND 0.02fF $ **FLOATING
C1749 VDD.n135 GND 0.02fF $ **FLOATING
C1750 VDD.n136 GND 0.48fF $ **FLOATING
C1751 VDD.n137 GND 0.23fF $ **FLOATING
C1752 VDD.n138 GND 0.14fF $ **FLOATING
C1753 VDD.n139 GND 0.19fF $ **FLOATING
C1754 VDD.n140 GND 0.14fF $ **FLOATING
C1755 VDD.n141 GND 0.27fF $ **FLOATING
C1756 VDD.n142 GND 0.02fF $ **FLOATING
C1757 VDD.n143 GND 0.02fF $ **FLOATING
C1758 VDD.n144 GND 0.02fF $ **FLOATING
C1759 VDD.n145 GND 0.48fF $ **FLOATING
C1760 VDD.t133 GND 0.11fF
C1761 VDD.n146 GND 0.16fF $ **FLOATING
C1762 VDD.n147 GND 0.02fF $ **FLOATING
C1763 VDD.n148 GND 0.02fF $ **FLOATING
C1764 VDD.n149 GND 0.02fF $ **FLOATING
C1765 VDD.n150 GND 0.19fF $ **FLOATING
C1766 VDD.n151 GND 0.02fF $ **FLOATING
C1767 VDD.n152 GND 0.02fF $ **FLOATING
C1768 VDD.n153 GND 0.02fF $ **FLOATING
C1769 VDD.t159 GND 0.11fF
C1770 VDD.n154 GND 0.16fF $ **FLOATING
C1771 VDD.n155 GND 0.02fF $ **FLOATING
C1772 VDD.n156 GND 0.02fF $ **FLOATING
C1773 VDD.n157 GND 0.02fF $ **FLOATING
C1774 VDD.n158 GND 0.18fF $ **FLOATING
C1775 VDD.n159 GND 0.02fF $ **FLOATING
C1776 VDD.n160 GND 0.02fF $ **FLOATING
C1777 VDD.n161 GND 0.02fF $ **FLOATING
C1778 VDD.n162 GND 0.02fF $ **FLOATING
C1779 VDD.n163 GND 0.02fF $ **FLOATING
C1780 VDD.t182 GND 0.11fF
C1781 VDD.n164 GND 0.17fF $ **FLOATING
C1782 VDD.n165 GND 0.02fF $ **FLOATING
C1783 VDD.n166 GND 0.02fF $ **FLOATING
C1784 VDD.n167 GND 0.02fF $ **FLOATING
C1785 VDD.n168 GND 0.17fF $ **FLOATING
C1786 VDD.n169 GND 0.02fF $ **FLOATING
C1787 VDD.n170 GND 0.02fF $ **FLOATING
C1788 VDD.n171 GND 0.02fF $ **FLOATING
C1789 VDD.t113 GND 0.11fF
C1790 VDD.n172 GND 0.17fF $ **FLOATING
C1791 VDD.n173 GND 0.02fF $ **FLOATING
C1792 VDD.n174 GND 0.02fF $ **FLOATING
C1793 VDD.n175 GND 0.02fF $ **FLOATING
C1794 VDD.n176 GND 0.48fF $ **FLOATING
C1795 VDD.n177 GND 0.25fF $ **FLOATING
C1796 VDD.n178 GND 0.02fF $ **FLOATING
C1797 VDD.n179 GND 0.02fF $ **FLOATING
C1798 VDD.n180 GND 0.02fF $ **FLOATING
C1799 CMOS_sbox_0/VDD GND 0.00fF $ **FLOATING
C1800 CMOS_sbox_0/CMOS_s0_0/VDD GND 0.01fF $ **FLOATING
C1801 VDD.t181 GND 0.06fF
C1802 VDD.t132 GND 0.06fF
C1803 VDD.n181 GND 0.25fF $ **FLOATING
C1804 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/VDD GND 0.01fF $ **FLOATING
C1805 VDD.t27 GND 0.09fF
C1806 VDD.t53 GND 0.09fF
C1807 VDD.t112 GND 0.09fF
C1808 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/VDD GND 0.01fF $ **FLOATING
C1809 VDD.t120 GND 0.09fF
C1810 VDD.t100 GND 0.09fF
C1811 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_OR_0/VDD GND 0.01fF $ **FLOATING
C1812 VDD.t73 GND 0.09fF
C1813 VDD.n182 GND 0.26fF $ **FLOATING
C1814 VDD.n183 GND 0.02fF $ **FLOATING
C1815 VDD.n184 GND 0.02fF $ **FLOATING
C1816 VDD.n185 GND 0.21fF $ **FLOATING
C1817 VDD.t72 GND 0.13fF
C1818 VDD.n186 GND 0.14fF $ **FLOATING
C1819 VDD.n187 GND 0.02fF $ **FLOATING
C1820 VDD.n188 GND 0.02fF $ **FLOATING
C1821 VDD.n189 GND 0.06fF $ **FLOATING
C1822 VDD.n190 GND 0.48fF $ **FLOATING
C1823 VDD.n191 GND 0.22fF $ **FLOATING
C1824 VDD.n192 GND 0.02fF $ **FLOATING
C1825 VDD.n193 GND 0.02fF $ **FLOATING
C1826 VDD.n194 GND 0.01fF $ **FLOATING
C1827 VDD.n195 GND 0.22fF $ **FLOATING
C1828 VDD.n196 GND 0.02fF $ **FLOATING
C1829 VDD.n197 GND 0.02fF $ **FLOATING
C1830 VDD.n198 GND 0.02fF $ **FLOATING
C1831 VDD.n199 GND 0.22fF $ **FLOATING
C1832 VDD.n200 GND 0.02fF $ **FLOATING
C1833 VDD.n201 GND 0.02fF $ **FLOATING
C1834 VDD.n202 GND 0.02fF $ **FLOATING
C1835 VDD.n203 GND 0.22fF $ **FLOATING
C1836 VDD.n204 GND 0.02fF $ **FLOATING
C1837 VDD.n205 GND 0.02fF $ **FLOATING
C1838 VDD.n206 GND 0.02fF $ **FLOATING
C1839 VDD.t3 GND 0.11fF
C1840 VDD.n207 GND 0.13fF $ **FLOATING
C1841 VDD.n208 GND 0.02fF $ **FLOATING
C1842 VDD.n209 GND 0.02fF $ **FLOATING
C1843 VDD.n210 GND 0.02fF $ **FLOATING
C1844 VDD.n211 GND 0.02fF $ **FLOATING
C1845 VDD.n212 GND 0.20fF $ **FLOATING
C1846 VDD.n213 GND 0.02fF $ **FLOATING
C1847 VDD.n214 GND 0.02fF $ **FLOATING
C1848 VDD.t54 GND 0.11fF
C1849 VDD.n215 GND 0.14fF $ **FLOATING
C1850 VDD.n216 GND 0.02fF $ **FLOATING
C1851 VDD.n217 GND 0.02fF $ **FLOATING
C1852 VDD.n218 GND 0.02fF $ **FLOATING
C1853 VDD.n219 GND 0.19fF $ **FLOATING
C1854 VDD.n220 GND 0.02fF $ **FLOATING
C1855 VDD.n221 GND 0.02fF $ **FLOATING
C1856 VDD.n222 GND 0.02fF $ **FLOATING
C1857 VDD.t99 GND 0.13fF
C1858 VDD.n223 GND 0.15fF $ **FLOATING
C1859 VDD.n224 GND 0.02fF $ **FLOATING
C1860 VDD.n225 GND 0.02fF $ **FLOATING
C1861 VDD.n226 GND 0.02fF $ **FLOATING
C1862 VDD.n227 GND 0.24fF $ **FLOATING
C1863 VDD.n228 GND 0.02fF $ **FLOATING
C1864 VDD.n229 GND 0.02fF $ **FLOATING
C1865 VDD.n230 GND 0.02fF $ **FLOATING
C1866 VDD.n231 GND 0.48fF $ **FLOATING
C1867 VDD.n232 GND 0.23fF $ **FLOATING
C1868 VDD.n233 GND 0.08fF $ **FLOATING
C1869 VDD.n234 GND 0.20fF $ **FLOATING
C1870 VDD.n235 GND 0.08fF $ **FLOATING
C1871 VDD.n236 GND 0.25fF $ **FLOATING
C1872 VDD.n237 GND 0.02fF $ **FLOATING
C1873 VDD.n238 GND 0.02fF $ **FLOATING
C1874 VDD.n239 GND 0.02fF $ **FLOATING
C1875 VDD.t119 GND 0.13fF
C1876 VDD.n240 GND 0.13fF $ **FLOATING
C1877 VDD.n241 GND 0.02fF $ **FLOATING
C1878 VDD.n242 GND 0.02fF $ **FLOATING
C1879 VDD.n243 GND 0.02fF $ **FLOATING
C1880 VDD.n244 GND 0.48fF $ **FLOATING
C1881 VDD.n245 GND 0.22fF $ **FLOATING
C1882 VDD.n246 GND 0.02fF $ **FLOATING
C1883 VDD.n247 GND 0.02fF $ **FLOATING
C1884 VDD.n248 GND 0.01fF $ **FLOATING
C1885 VDD.n249 GND 0.22fF $ **FLOATING
C1886 VDD.n250 GND 0.02fF $ **FLOATING
C1887 VDD.n251 GND 0.02fF $ **FLOATING
C1888 VDD.n252 GND 0.02fF $ **FLOATING
C1889 VDD.n253 GND 0.22fF $ **FLOATING
C1890 VDD.n254 GND 0.02fF $ **FLOATING
C1891 VDD.n255 GND 0.02fF $ **FLOATING
C1892 VDD.n256 GND 0.02fF $ **FLOATING
C1893 VDD.t7 GND 0.09fF
C1894 VDD.n257 GND 0.47fF $ **FLOATING
C1895 VDD.n258 GND 0.01fF $ **FLOATING
C1896 VDD.n259 GND 0.22fF $ **FLOATING
C1897 VDD.n260 GND 0.02fF $ **FLOATING
C1898 VDD.n261 GND 0.02fF $ **FLOATING
C1899 VDD.t6 GND 0.11fF
C1900 VDD.n262 GND 0.14fF $ **FLOATING
C1901 VDD.n263 GND 0.02fF $ **FLOATING
C1902 VDD.n264 GND 0.02fF $ **FLOATING
C1903 VDD.n265 GND 0.02fF $ **FLOATING
C1904 VDD.n266 GND 0.19fF $ **FLOATING
C1905 VDD.n267 GND 0.02fF $ **FLOATING
C1906 VDD.n268 GND 0.02fF $ **FLOATING
C1907 VDD.n269 GND 0.02fF $ **FLOATING
C1908 VDD.t111 GND 0.13fF
C1909 VDD.n270 GND 0.15fF $ **FLOATING
C1910 VDD.n271 GND 0.02fF $ **FLOATING
C1911 VDD.n272 GND 0.02fF $ **FLOATING
C1912 VDD.n273 GND 0.02fF $ **FLOATING
C1913 VDD.n274 GND 0.24fF $ **FLOATING
C1914 VDD.n275 GND 0.02fF $ **FLOATING
C1915 VDD.n276 GND 0.02fF $ **FLOATING
C1916 VDD.n277 GND 0.02fF $ **FLOATING
C1917 VDD.n278 GND 0.48fF $ **FLOATING
C1918 VDD.n279 GND 0.23fF $ **FLOATING
C1919 VDD.n280 GND 0.11fF $ **FLOATING
C1920 VDD.n281 GND 0.22fF $ **FLOATING
C1921 VDD.n282 GND 0.12fF $ **FLOATING
C1922 VDD.n283 GND 0.25fF $ **FLOATING
C1923 VDD.n284 GND 0.02fF $ **FLOATING
C1924 VDD.n285 GND 0.02fF $ **FLOATING
C1925 VDD.n286 GND 0.02fF $ **FLOATING
C1926 VDD.t52 GND 0.13fF
C1927 VDD.n287 GND 0.14fF $ **FLOATING
C1928 VDD.n288 GND 0.02fF $ **FLOATING
C1929 VDD.n289 GND 0.02fF $ **FLOATING
C1930 VDD.n290 GND 0.02fF $ **FLOATING
C1931 VDD.n291 GND 0.48fF $ **FLOATING
C1932 VDD.n292 GND 0.22fF $ **FLOATING
C1933 VDD.n293 GND 0.02fF $ **FLOATING
C1934 VDD.n294 GND 0.02fF $ **FLOATING
C1935 VDD.n295 GND 0.01fF $ **FLOATING
C1936 VDD.n296 GND 0.22fF $ **FLOATING
C1937 VDD.n297 GND 0.02fF $ **FLOATING
C1938 VDD.n298 GND 0.02fF $ **FLOATING
C1939 VDD.n299 GND 0.02fF $ **FLOATING
C1940 VDD.n300 GND 0.22fF $ **FLOATING
C1941 VDD.n301 GND 0.02fF $ **FLOATING
C1942 VDD.n302 GND 0.02fF $ **FLOATING
C1943 VDD.n303 GND 0.02fF $ **FLOATING
C1944 VDD.n304 GND 0.22fF $ **FLOATING
C1945 VDD.n305 GND 0.02fF $ **FLOATING
C1946 VDD.n306 GND 0.02fF $ **FLOATING
C1947 VDD.n307 GND 0.01fF $ **FLOATING
C1948 VDD.n308 GND 0.48fF $ **FLOATING
C1949 VDD.t26 GND 0.11fF
C1950 VDD.n309 GND 0.13fF $ **FLOATING
C1951 VDD.n310 GND 0.02fF $ **FLOATING
C1952 VDD.n311 GND 0.02fF $ **FLOATING
C1953 VDD.n312 GND 0.02fF $ **FLOATING
C1954 VDD.n313 GND 0.02fF $ **FLOATING
C1955 VDD.n314 GND 0.20fF $ **FLOATING
C1956 VDD.n315 GND 0.02fF $ **FLOATING
C1957 VDD.n316 GND 0.02fF $ **FLOATING
C1958 VDD.t180 GND 0.11fF
C1959 VDD.n317 GND 0.14fF $ **FLOATING
C1960 VDD.n318 GND 0.02fF $ **FLOATING
C1961 VDD.n319 GND 0.02fF $ **FLOATING
C1962 VDD.n320 GND 0.02fF $ **FLOATING
C1963 VDD.n321 GND 0.19fF $ **FLOATING
C1964 VDD.n322 GND 0.02fF $ **FLOATING
C1965 VDD.n323 GND 0.02fF $ **FLOATING
C1966 VDD.n324 GND 0.02fF $ **FLOATING
C1967 VDD.n325 GND 0.21fF $ **FLOATING
C1968 VDD.t131 GND 0.13fF
C1969 VDD.n326 GND 0.15fF $ **FLOATING
C1970 VDD.n327 GND 0.02fF $ **FLOATING
C1971 VDD.n328 GND 0.02fF $ **FLOATING
C1972 VDD.n329 GND 0.02fF $ **FLOATING
C1973 VDD.n330 GND 0.24fF $ **FLOATING
C1974 VDD.n331 GND 0.02fF $ **FLOATING
C1975 VDD.n332 GND 0.02fF $ **FLOATING
C1976 VDD.n333 GND 0.02fF $ **FLOATING
C1977 VDD.n334 GND 0.23fF $ **FLOATING
C1978 VDD.n335 GND 0.46fF $ **FLOATING
C1979 VDD.t149 GND 0.09fF
C1980 VDD.t15 GND 0.09fF
C1981 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/VDD GND 0.01fF $ **FLOATING
C1982 VDD.t103 GND 0.09fF
C1983 VDD.t179 GND 0.09fF
C1984 VDD.t41 GND 0.09fF
C1985 VDD.t96 GND 0.09fF
C1986 VDD.t34 GND 0.09fF
C1987 VDD.t105 GND 0.09fF
C1988 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/VDD GND 0.01fF $ **FLOATING
C1989 VDD.t161 GND 0.09fF
C1990 VDD.t136 GND 0.09fF
C1991 VDD.t163 GND 0.09fF
C1992 VDD.t25 GND 0.09fF
C1993 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_0/VDD GND 0.01fF $ **FLOATING
C1994 VDD.t64 GND 0.09fF
C1995 VDD.t98 GND 0.09fF
C1996 VDD.n336 GND 0.32fF $ **FLOATING
C1997 VDD.n337 GND 0.02fF $ **FLOATING
C1998 VDD.n338 GND 0.02fF $ **FLOATING
C1999 VDD.n339 GND 0.12fF $ **FLOATING
C2000 VDD.t97 GND 0.17fF
C2001 VDD.n340 GND 0.15fF $ **FLOATING
C2002 VDD.n341 GND 0.02fF $ **FLOATING
C2003 VDD.n342 GND 0.02fF $ **FLOATING
C2004 VDD.n343 GND 0.06fF $ **FLOATING
C2005 VDD.n344 GND 0.48fF $ **FLOATING
C2006 VDD.n345 GND 0.24fF $ **FLOATING
C2007 VDD.n346 GND 0.02fF $ **FLOATING
C2008 VDD.n347 GND 0.02fF $ **FLOATING
C2009 VDD.n348 GND 0.01fF $ **FLOATING
C2010 VDD.n349 GND 0.24fF $ **FLOATING
C2011 VDD.n350 GND 0.02fF $ **FLOATING
C2012 VDD.n351 GND 0.02fF $ **FLOATING
C2013 VDD.n352 GND 0.02fF $ **FLOATING
C2014 VDD.n353 GND 0.48fF $ **FLOATING
C2015 VDD.n354 GND 0.24fF $ **FLOATING
C2016 VDD.n355 GND 0.02fF $ **FLOATING
C2017 VDD.n356 GND 0.02fF $ **FLOATING
C2018 VDD.n357 GND 0.01fF $ **FLOATING
C2019 VDD.n358 GND 0.24fF $ **FLOATING
C2020 VDD.n359 GND 0.02fF $ **FLOATING
C2021 VDD.n360 GND 0.02fF $ **FLOATING
C2022 VDD.n361 GND 0.02fF $ **FLOATING
C2023 VDD.t20 GND 0.07fF
C2024 VDD.n362 GND 0.14fF $ **FLOATING
C2025 VDD.n363 GND 0.02fF $ **FLOATING
C2026 VDD.n364 GND 0.02fF $ **FLOATING
C2027 VDD.n365 GND 0.02fF $ **FLOATING
C2028 VDD.t81 GND 0.09fF
C2029 VDD.n366 GND 0.47fF $ **FLOATING
C2030 VDD.n367 GND 0.01fF $ **FLOATING
C2031 VDD.t63 GND 0.72fF
C2032 VDD.t24 GND 0.58fF
C2033 VDD.t80 GND 0.31fF
C2034 VDD.n368 GND 0.55fF $ **FLOATING
C2035 VDD.n369 GND 0.17fF $ **FLOATING
C2036 VDD.n370 GND 0.02fF $ **FLOATING
C2037 VDD.n371 GND 0.02fF $ **FLOATING
C2038 VDD.t43 GND 0.12fF
C2039 VDD.n372 GND 0.15fF $ **FLOATING
C2040 VDD.n373 GND 0.02fF $ **FLOATING
C2041 VDD.n374 GND 0.02fF $ **FLOATING
C2042 VDD.n375 GND 0.02fF $ **FLOATING
C2043 VDD.n376 GND 0.21fF $ **FLOATING
C2044 VDD.n377 GND 0.02fF $ **FLOATING
C2045 VDD.n378 GND 0.02fF $ **FLOATING
C2046 VDD.n379 GND 0.02fF $ **FLOATING
C2047 VDD.t162 GND 0.14fF
C2048 VDD.n380 GND 0.16fF $ **FLOATING
C2049 VDD.n381 GND 0.02fF $ **FLOATING
C2050 VDD.n382 GND 0.02fF $ **FLOATING
C2051 VDD.n383 GND 0.02fF $ **FLOATING
C2052 VDD.n384 GND 0.26fF $ **FLOATING
C2053 VDD.n385 GND 0.02fF $ **FLOATING
C2054 VDD.n386 GND 0.02fF $ **FLOATING
C2055 VDD.n387 GND 0.02fF $ **FLOATING
C2056 VDD.n388 GND 0.95fF $ **FLOATING
C2057 VDD.n389 GND 0.24fF $ **FLOATING
C2058 VDD.n390 GND 0.08fF $ **FLOATING
C2059 VDD.n391 GND 0.20fF $ **FLOATING
C2060 VDD.n392 GND 0.08fF $ **FLOATING
C2061 VDD.n393 GND 0.27fF $ **FLOATING
C2062 VDD.n394 GND 0.02fF $ **FLOATING
C2063 VDD.n395 GND 0.02fF $ **FLOATING
C2064 VDD.n396 GND 0.02fF $ **FLOATING
C2065 VDD.n397 GND 0.48fF $ **FLOATING
C2066 VDD.t160 GND 0.13fF
C2067 VDD.n398 GND 0.14fF $ **FLOATING
C2068 VDD.n399 GND 0.02fF $ **FLOATING
C2069 VDD.n400 GND 0.02fF $ **FLOATING
C2070 VDD.n401 GND 0.02fF $ **FLOATING
C2071 VDD.n402 GND 0.48fF $ **FLOATING
C2072 VDD.n403 GND 0.24fF $ **FLOATING
C2073 VDD.n404 GND 0.02fF $ **FLOATING
C2074 VDD.n405 GND 0.02fF $ **FLOATING
C2075 VDD.n406 GND 0.01fF $ **FLOATING
C2076 VDD.n407 GND 0.24fF $ **FLOATING
C2077 VDD.n408 GND 0.02fF $ **FLOATING
C2078 VDD.n409 GND 0.02fF $ **FLOATING
C2079 VDD.n410 GND 0.02fF $ **FLOATING
C2080 VDD.t135 GND 0.65fF
C2081 VDD.t58 GND 0.25fF
C2082 VDD.t104 GND 0.62fF
C2083 VDD.t154 GND 0.27fF
C2084 VDD.n411 GND 0.29fF $ **FLOATING
C2085 VDD.n412 GND 0.16fF $ **FLOATING
C2086 VDD.n413 GND 0.02fF $ **FLOATING
C2087 VDD.n414 GND 0.02fF $ **FLOATING
C2088 VDD.n415 GND 0.02fF $ **FLOATING
C2089 VDD.t48 GND 0.09fF
C2090 VDD.n416 GND 0.47fF $ **FLOATING
C2091 VDD.n417 GND 0.01fF $ **FLOATING
C2092 VDD.n418 GND 0.19fF $ **FLOATING
C2093 VDD.n419 GND 0.02fF $ **FLOATING
C2094 VDD.n420 GND 0.02fF $ **FLOATING
C2095 VDD.t47 GND 0.12fF
C2096 VDD.n421 GND 0.15fF $ **FLOATING
C2097 VDD.n422 GND 0.02fF $ **FLOATING
C2098 VDD.n423 GND 0.02fF $ **FLOATING
C2099 VDD.n424 GND 0.02fF $ **FLOATING
C2100 VDD.n425 GND 0.21fF $ **FLOATING
C2101 VDD.n426 GND 0.02fF $ **FLOATING
C2102 VDD.n427 GND 0.02fF $ **FLOATING
C2103 VDD.n428 GND 0.02fF $ **FLOATING
C2104 VDD.t33 GND 0.14fF
C2105 VDD.n429 GND 0.16fF $ **FLOATING
C2106 VDD.n430 GND 0.02fF $ **FLOATING
C2107 VDD.n431 GND 0.02fF $ **FLOATING
C2108 VDD.n432 GND 0.02fF $ **FLOATING
C2109 VDD.n433 GND 0.48fF $ **FLOATING
C2110 VDD.n434 GND 0.26fF $ **FLOATING
C2111 VDD.n435 GND 0.02fF $ **FLOATING
C2112 VDD.n436 GND 0.02fF $ **FLOATING
C2113 VDD.n437 GND 0.01fF $ **FLOATING
C2114 VDD.n438 GND 0.48fF $ **FLOATING
C2115 VDD.n439 GND 0.24fF $ **FLOATING
C2116 VDD.n440 GND 0.08fF $ **FLOATING
C2117 VDD.n441 GND 0.15fF $ **FLOATING
C2118 VDD.n442 GND 0.02fF $ **FLOATING
C2119 VDD.n443 GND 0.02fF $ **FLOATING
C2120 VDD.n444 GND 0.08fF $ **FLOATING
C2121 VDD.n445 GND 0.21fF $ **FLOATING
C2122 VDD.n446 GND 0.02fF $ **FLOATING
C2123 VDD.n447 GND 0.02fF $ **FLOATING
C2124 VDD.n448 GND 0.02fF $ **FLOATING
C2125 VDD.n449 GND 0.20fF $ **FLOATING
C2126 VDD.n450 GND 0.02fF $ **FLOATING
C2127 VDD.n451 GND 0.02fF $ **FLOATING
C2128 VDD.n452 GND 0.02fF $ **FLOATING
C2129 VDD.n453 GND 0.48fF $ **FLOATING
C2130 VDD.t40 GND 0.12fF
C2131 VDD.n454 GND 0.16fF $ **FLOATING
C2132 VDD.n455 GND 0.02fF $ **FLOATING
C2133 VDD.n456 GND 0.02fF $ **FLOATING
C2134 VDD.n457 GND 0.01fF $ **FLOATING
C2135 VDD.n458 GND 0.48fF $ **FLOATING
C2136 VDD.n459 GND 0.24fF $ **FLOATING
C2137 VDD.n460 GND 0.02fF $ **FLOATING
C2138 VDD.n461 GND 0.02fF $ **FLOATING
C2139 VDD.n462 GND 0.02fF $ **FLOATING
C2140 VDD.n463 GND 0.24fF $ **FLOATING
C2141 VDD.n464 GND 0.02fF $ **FLOATING
C2142 VDD.n465 GND 0.02fF $ **FLOATING
C2143 VDD.n466 GND 0.02fF $ **FLOATING
C2144 VDD.n467 GND 0.24fF $ **FLOATING
C2145 VDD.n468 GND 0.02fF $ **FLOATING
C2146 VDD.n469 GND 0.02fF $ **FLOATING
C2147 VDD.n470 GND 0.02fF $ **FLOATING
C2148 VDD.n471 GND 0.48fF $ **FLOATING
C2149 VDD.n472 GND 0.24fF $ **FLOATING
C2150 VDD.n473 GND 0.02fF $ **FLOATING
C2151 VDD.n474 GND 0.02fF $ **FLOATING
C2152 VDD.n475 GND 0.01fF $ **FLOATING
C2153 VDD.n476 GND 0.48fF $ **FLOATING
C2154 VDD.t95 GND 0.85fF
C2155 VDD.t178 GND 0.54fF
C2156 VDD.t14 GND 0.62fF
C2157 VDD.t2 GND 0.35fF
C2158 VDD.t21 GND 0.27fF
C2159 VDD.n477 GND 0.28fF $ **FLOATING
C2160 VDD.t102 GND 0.03fF
C2161 VDD.n478 GND 0.13fF $ **FLOATING
C2162 VDD.n479 GND 0.02fF $ **FLOATING
C2163 VDD.n480 GND 0.02fF $ **FLOATING
C2164 VDD.n481 GND 0.02fF $ **FLOATING
C2165 VDD.n482 GND 0.20fF $ **FLOATING
C2166 VDD.n483 GND 0.02fF $ **FLOATING
C2167 VDD.n484 GND 0.02fF $ **FLOATING
C2168 VDD.n485 GND 0.02fF $ **FLOATING
C2169 VDD.t84 GND 0.12fF
C2170 VDD.n486 GND 0.14fF $ **FLOATING
C2171 VDD.n487 GND 0.02fF $ **FLOATING
C2172 VDD.n488 GND 0.02fF $ **FLOATING
C2173 VDD.n489 GND 0.02fF $ **FLOATING
C2174 VDD.t85 GND 0.06fF
C2175 VDD.t177 GND 0.06fF
C2176 VDD.n490 GND 0.25fF $ **FLOATING
C2177 VDD.n491 GND 0.20fF $ **FLOATING
C2178 VDD.n492 GND 0.01fF $ **FLOATING
C2179 VDD.n493 GND 0.22fF $ **FLOATING
C2180 VDD.n494 GND 0.02fF $ **FLOATING
C2181 VDD.n495 GND 0.02fF $ **FLOATING
C2182 VDD.t176 GND 0.12fF
C2183 VDD.n496 GND 0.15fF $ **FLOATING
C2184 VDD.n497 GND 0.02fF $ **FLOATING
C2185 VDD.n498 GND 0.02fF $ **FLOATING
C2186 VDD.n499 GND 0.02fF $ **FLOATING
C2187 VDD.n500 GND 0.21fF $ **FLOATING
C2188 VDD.n501 GND 0.02fF $ **FLOATING
C2189 VDD.n502 GND 0.02fF $ **FLOATING
C2190 VDD.n503 GND 0.02fF $ **FLOATING
C2191 VDD.t148 GND 0.14fF
C2192 VDD.n504 GND 0.16fF $ **FLOATING
C2193 VDD.n505 GND 0.02fF $ **FLOATING
C2194 VDD.n506 GND 0.02fF $ **FLOATING
C2195 VDD.n507 GND 0.02fF $ **FLOATING
C2196 VDD.n508 GND 0.48fF $ **FLOATING
C2197 VDD.n509 GND 0.26fF $ **FLOATING
C2198 VDD.n510 GND 0.02fF $ **FLOATING
C2199 VDD.n511 GND 0.02fF $ **FLOATING
C2200 VDD.n512 GND 0.01fF $ **FLOATING
C2201 VDD.n513 GND 0.48fF $ **FLOATING
C2202 VDD.n514 GND 0.24fF $ **FLOATING
C2203 VDD.n515 GND 0.03fF $ **FLOATING
C2204 CMOS_sbox_0/CMOS_s3_0/VDD GND 0.01fF $ **FLOATING
C2205 VDD.n516 GND 0.85fF $ **FLOATING
C2206 VDD.t29 GND 0.09fF
C2207 VDD.t1 GND 0.06fF
C2208 VDD.t39 GND 0.06fF
C2209 VDD.n517 GND 0.25fF $ **FLOATING
C2210 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/VDD GND 0.01fF $ **FLOATING
C2211 VDD.t110 GND 0.09fF
C2212 VDD.t147 GND 0.09fF
C2213 VDD.t83 GND 0.09fF
C2214 VDD.t50 GND 0.09fF
C2215 VDD.t138 GND 0.09fF
C2216 VDD.t169 GND 0.09fF
C2217 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_1/VDD GND 0.01fF $ **FLOATING
C2218 VDD.t93 GND 0.09fF
C2219 VDD.t172 GND 0.09fF
C2220 VDD.t62 GND 0.09fF
C2221 VDD.t13 GND 0.09fF
C2222 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_OR_0/VDD GND 0.01fF $ **FLOATING
C2223 VDD.t45 GND 0.09fF
C2224 VDD.t126 GND 0.09fF
C2225 VDD.n518 GND 0.32fF $ **FLOATING
C2226 VDD.n519 GND 0.02fF $ **FLOATING
C2227 VDD.n520 GND 0.02fF $ **FLOATING
C2228 VDD.n521 GND 0.12fF $ **FLOATING
C2229 VDD.t125 GND 0.17fF
C2230 VDD.n522 GND 0.15fF $ **FLOATING
C2231 VDD.n523 GND 0.02fF $ **FLOATING
C2232 VDD.n524 GND 0.02fF $ **FLOATING
C2233 VDD.n525 GND 0.06fF $ **FLOATING
C2234 VDD.n526 GND 0.48fF $ **FLOATING
C2235 VDD.n527 GND 0.24fF $ **FLOATING
C2236 VDD.n528 GND 0.02fF $ **FLOATING
C2237 VDD.n529 GND 0.02fF $ **FLOATING
C2238 VDD.n530 GND 0.01fF $ **FLOATING
C2239 VDD.n531 GND 0.24fF $ **FLOATING
C2240 VDD.n532 GND 0.02fF $ **FLOATING
C2241 VDD.n533 GND 0.02fF $ **FLOATING
C2242 VDD.n534 GND 0.02fF $ **FLOATING
C2243 VDD.n535 GND 0.48fF $ **FLOATING
C2244 VDD.n536 GND 0.24fF $ **FLOATING
C2245 VDD.n537 GND 0.02fF $ **FLOATING
C2246 VDD.n538 GND 0.02fF $ **FLOATING
C2247 VDD.n539 GND 0.01fF $ **FLOATING
C2248 VDD.n540 GND 0.24fF $ **FLOATING
C2249 VDD.n541 GND 0.02fF $ **FLOATING
C2250 VDD.n542 GND 0.02fF $ **FLOATING
C2251 VDD.n543 GND 0.02fF $ **FLOATING
C2252 VDD.t57 GND 0.07fF
C2253 VDD.n544 GND 0.14fF $ **FLOATING
C2254 VDD.n545 GND 0.02fF $ **FLOATING
C2255 VDD.n546 GND 0.02fF $ **FLOATING
C2256 VDD.n547 GND 0.02fF $ **FLOATING
C2257 VDD.t79 GND 0.09fF
C2258 VDD.n548 GND 0.47fF $ **FLOATING
C2259 VDD.n549 GND 0.01fF $ **FLOATING
C2260 VDD.t44 GND 0.72fF
C2261 VDD.t12 GND 0.58fF
C2262 VDD.t78 GND 0.31fF
C2263 VDD.n550 GND 0.55fF $ **FLOATING
C2264 VDD.n551 GND 0.17fF $ **FLOATING
C2265 VDD.n552 GND 0.02fF $ **FLOATING
C2266 VDD.n553 GND 0.02fF $ **FLOATING
C2267 VDD.t17 GND 0.12fF
C2268 VDD.n554 GND 0.15fF $ **FLOATING
C2269 VDD.n555 GND 0.02fF $ **FLOATING
C2270 VDD.n556 GND 0.02fF $ **FLOATING
C2271 VDD.n557 GND 0.02fF $ **FLOATING
C2272 VDD.n558 GND 0.21fF $ **FLOATING
C2273 VDD.n559 GND 0.02fF $ **FLOATING
C2274 VDD.n560 GND 0.02fF $ **FLOATING
C2275 VDD.n561 GND 0.02fF $ **FLOATING
C2276 VDD.t61 GND 0.14fF
C2277 VDD.n562 GND 0.16fF $ **FLOATING
C2278 VDD.n563 GND 0.02fF $ **FLOATING
C2279 VDD.n564 GND 0.02fF $ **FLOATING
C2280 VDD.n565 GND 0.02fF $ **FLOATING
C2281 VDD.n566 GND 0.26fF $ **FLOATING
C2282 VDD.n567 GND 0.02fF $ **FLOATING
C2283 VDD.n568 GND 0.02fF $ **FLOATING
C2284 VDD.n569 GND 0.02fF $ **FLOATING
C2285 VDD.n570 GND 0.95fF $ **FLOATING
C2286 VDD.n571 GND 0.24fF $ **FLOATING
C2287 VDD.n572 GND 0.08fF $ **FLOATING
C2288 VDD.n573 GND 0.20fF $ **FLOATING
C2289 VDD.n574 GND 0.08fF $ **FLOATING
C2290 VDD.n575 GND 0.27fF $ **FLOATING
C2291 VDD.n576 GND 0.02fF $ **FLOATING
C2292 VDD.n577 GND 0.02fF $ **FLOATING
C2293 VDD.n578 GND 0.02fF $ **FLOATING
C2294 VDD.n579 GND 0.48fF $ **FLOATING
C2295 VDD.t92 GND 0.13fF
C2296 VDD.n580 GND 0.14fF $ **FLOATING
C2297 VDD.n581 GND 0.02fF $ **FLOATING
C2298 VDD.n582 GND 0.02fF $ **FLOATING
C2299 VDD.n583 GND 0.02fF $ **FLOATING
C2300 VDD.n584 GND 0.48fF $ **FLOATING
C2301 VDD.n585 GND 0.24fF $ **FLOATING
C2302 VDD.n586 GND 0.02fF $ **FLOATING
C2303 VDD.n587 GND 0.02fF $ **FLOATING
C2304 VDD.n588 GND 0.01fF $ **FLOATING
C2305 VDD.n589 GND 0.24fF $ **FLOATING
C2306 VDD.n590 GND 0.02fF $ **FLOATING
C2307 VDD.n591 GND 0.02fF $ **FLOATING
C2308 VDD.n592 GND 0.02fF $ **FLOATING
C2309 VDD.t171 GND 0.65fF
C2310 VDD.t42 GND 0.25fF
C2311 VDD.t168 GND 0.62fF
C2312 VDD.t156 GND 0.27fF
C2313 VDD.n593 GND 0.29fF $ **FLOATING
C2314 VDD.n594 GND 0.16fF $ **FLOATING
C2315 VDD.n595 GND 0.02fF $ **FLOATING
C2316 VDD.n596 GND 0.02fF $ **FLOATING
C2317 VDD.n597 GND 0.02fF $ **FLOATING
C2318 VDD.t122 GND 0.09fF
C2319 VDD.n598 GND 0.47fF $ **FLOATING
C2320 VDD.n599 GND 0.01fF $ **FLOATING
C2321 VDD.n600 GND 0.19fF $ **FLOATING
C2322 VDD.n601 GND 0.02fF $ **FLOATING
C2323 VDD.n602 GND 0.02fF $ **FLOATING
C2324 VDD.t121 GND 0.12fF
C2325 VDD.n603 GND 0.15fF $ **FLOATING
C2326 VDD.n604 GND 0.02fF $ **FLOATING
C2327 VDD.n605 GND 0.02fF $ **FLOATING
C2328 VDD.n606 GND 0.02fF $ **FLOATING
C2329 VDD.n607 GND 0.21fF $ **FLOATING
C2330 VDD.n608 GND 0.02fF $ **FLOATING
C2331 VDD.n609 GND 0.02fF $ **FLOATING
C2332 VDD.n610 GND 0.02fF $ **FLOATING
C2333 VDD.t137 GND 0.14fF
C2334 VDD.n611 GND 0.16fF $ **FLOATING
C2335 VDD.n612 GND 0.02fF $ **FLOATING
C2336 VDD.n613 GND 0.02fF $ **FLOATING
C2337 VDD.n614 GND 0.02fF $ **FLOATING
C2338 VDD.n615 GND 0.48fF $ **FLOATING
C2339 VDD.n616 GND 0.26fF $ **FLOATING
C2340 VDD.n617 GND 0.02fF $ **FLOATING
C2341 VDD.n618 GND 0.02fF $ **FLOATING
C2342 VDD.n619 GND 0.01fF $ **FLOATING
C2343 VDD.n620 GND 0.48fF $ **FLOATING
C2344 VDD.n621 GND 0.24fF $ **FLOATING
C2345 VDD.n622 GND 0.08fF $ **FLOATING
C2346 VDD.n623 GND 0.03fF $ **FLOATING
C2347 VDD.n624 GND 0.08fF $ **FLOATING
C2348 VDD.t49 GND 0.26fF
C2349 VDD.n625 GND 0.21fF $ **FLOATING
C2350 VDD.n626 GND 0.16fF $ **FLOATING
C2351 VDD.n627 GND 0.01fF $ **FLOATING
C2352 VDD.n628 GND 0.02fF $ **FLOATING
C2353 VDD.n629 GND 0.02fF $ **FLOATING
C2354 VDD.n630 GND 0.02fF $ **FLOATING
C2355 VDD.n631 GND 0.02fF $ **FLOATING
C2356 VDD.n632 GND 0.02fF $ **FLOATING
C2357 VDD.n633 GND 0.02fF $ **FLOATING
C2358 VDD.n634 GND 0.48fF $ **FLOATING
C2359 VDD.n635 GND 0.30fF $ **FLOATING
C2360 VDD.n636 GND 0.02fF $ **FLOATING
C2361 VDD.n637 GND 0.02fF $ **FLOATING
C2362 VDD.n638 GND 0.01fF $ **FLOATING
C2363 VDD.n639 GND 0.21fF $ **FLOATING
C2364 VDD.n640 GND 0.02fF $ **FLOATING
C2365 VDD.n641 GND 0.02fF $ **FLOATING
C2366 VDD.n642 GND 0.02fF $ **FLOATING
C2367 VDD.t82 GND 0.12fF
C2368 VDD.n643 GND 0.15fF $ **FLOATING
C2369 VDD.n644 GND 0.02fF $ **FLOATING
C2370 VDD.n645 GND 0.02fF $ **FLOATING
C2371 VDD.n646 GND 0.02fF $ **FLOATING
C2372 VDD.n647 GND 0.48fF $ **FLOATING
C2373 VDD.n648 GND 0.24fF $ **FLOATING
C2374 VDD.n649 GND 0.02fF $ **FLOATING
C2375 VDD.n650 GND 0.02fF $ **FLOATING
C2376 VDD.n651 GND 0.01fF $ **FLOATING
C2377 VDD.n652 GND 0.48fF $ **FLOATING
C2378 VDD.n653 GND 0.24fF $ **FLOATING
C2379 VDD.n654 GND 0.02fF $ **FLOATING
C2380 VDD.n655 GND 0.02fF $ **FLOATING
C2381 VDD.n656 GND 0.02fF $ **FLOATING
C2382 VDD.n657 GND 0.24fF $ **FLOATING
C2383 VDD.n658 GND 0.02fF $ **FLOATING
C2384 VDD.n659 GND 0.02fF $ **FLOATING
C2385 VDD.n660 GND 0.02fF $ **FLOATING
C2386 VDD.t146 GND 0.99fF
C2387 VDD.t28 GND 0.62fF
C2388 VDD.t139 GND 0.35fF
C2389 VDD.t108 GND 0.18fF
C2390 VDD.n661 GND 0.29fF $ **FLOATING
C2391 VDD.n662 GND 0.15fF $ **FLOATING
C2392 VDD.n663 GND 0.02fF $ **FLOATING
C2393 VDD.n664 GND 0.02fF $ **FLOATING
C2394 VDD.n665 GND 0.01fF $ **FLOATING
C2395 VDD.n666 GND 0.48fF $ **FLOATING
C2396 VDD.t109 GND 0.12fF
C2397 VDD.n667 GND 0.10fF $ **FLOATING
C2398 VDD.n668 GND 0.02fF $ **FLOATING
C2399 VDD.n669 GND 0.02fF $ **FLOATING
C2400 VDD.n670 GND 0.02fF $ **FLOATING
C2401 VDD.n671 GND 0.02fF $ **FLOATING
C2402 VDD.n672 GND 0.22fF $ **FLOATING
C2403 VDD.n673 GND 0.02fF $ **FLOATING
C2404 VDD.n674 GND 0.02fF $ **FLOATING
C2405 VDD.t0 GND 0.12fF
C2406 VDD.n675 GND 0.15fF $ **FLOATING
C2407 VDD.n676 GND 0.02fF $ **FLOATING
C2408 VDD.n677 GND 0.02fF $ **FLOATING
C2409 VDD.n678 GND 0.02fF $ **FLOATING
C2410 VDD.n679 GND 0.21fF $ **FLOATING
C2411 VDD.n680 GND 0.02fF $ **FLOATING
C2412 VDD.n681 GND 0.02fF $ **FLOATING
C2413 VDD.n682 GND 0.02fF $ **FLOATING
C2414 VDD.n683 GND 0.21fF $ **FLOATING
C2415 VDD.t38 GND 0.14fF
C2416 VDD.n684 GND 0.16fF $ **FLOATING
C2417 VDD.n685 GND 0.02fF $ **FLOATING
C2418 VDD.n686 GND 0.02fF $ **FLOATING
C2419 VDD.n687 GND 0.02fF $ **FLOATING
C2420 VDD.n688 GND 0.48fF $ **FLOATING
C2421 VDD.n689 GND 0.26fF $ **FLOATING
C2422 VDD.n690 GND 0.02fF $ **FLOATING
C2423 VDD.n691 GND 0.02fF $ **FLOATING
C2424 VDD.n692 GND 0.02fF $ **FLOATING
C2425 VDD.n693 GND 0.40fF $ **FLOATING
C2426 VDD.n694 GND 0.03fF $ **FLOATING
C2427 CMOS_sbox_0/CMOS_s2_0/VDD GND 0.01fF $ **FLOATING
C2428 VDD.n695 GND 0.84fF $ **FLOATING
C2429 VDD.t31 GND 0.09fF
C2430 VDD.t51 GND 0.09fF
C2431 VDD.t173 GND 0.09fF
C2432 VDD.t153 GND 0.09fF
C2433 VDD.t56 GND 0.09fF
C2434 VDD.t19 GND 0.09fF
C2435 VDD.t89 GND 0.09fF
C2436 VDD.t107 GND 0.09fF
C2437 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/VDD GND 0.01fF $ **FLOATING
C2438 VDD.t128 GND 0.09fF
C2439 VDD.t141 GND 0.09fF
C2440 VDD.t9 GND 0.09fF
C2441 VDD.t46 GND 0.09fF
C2442 CMOS_sbox_0/CMOS_s1_0/CMOS_AND_0/VDD GND 0.01fF $ **FLOATING
C2443 VDD.t5 GND 0.09fF
C2444 VDD.t143 GND 0.09fF
C2445 VDD.n696 GND 0.51fF $ **FLOATING
C2446 VDD.n697 GND 0.02fF $ **FLOATING
C2447 VDD.n698 GND 0.02fF $ **FLOATING
C2448 VDD.n699 GND 0.28fF $ **FLOATING
C2449 VDD.t4 GND 0.24fF
C2450 VDD.n700 GND 0.23fF $ **FLOATING
C2451 VDD.n701 GND 0.02fF $ **FLOATING
C2452 VDD.n702 GND 0.02fF $ **FLOATING
C2453 VDD.n703 GND 0.07fF $ **FLOATING
C2454 VDD.n704 GND 0.95fF $ **FLOATING
C2455 VDD.n705 GND 0.40fF $ **FLOATING
C2456 VDD.n706 GND 0.02fF $ **FLOATING
C2457 VDD.n707 GND 0.02fF $ **FLOATING
C2458 VDD.n708 GND 0.01fF $ **FLOATING
C2459 VDD.n709 GND 0.40fF $ **FLOATING
C2460 VDD.n710 GND 0.02fF $ **FLOATING
C2461 VDD.n711 GND 0.02fF $ **FLOATING
C2462 VDD.n712 GND 0.02fF $ **FLOATING
C2463 VDD.n713 GND 0.40fF $ **FLOATING
C2464 VDD.n714 GND 0.02fF $ **FLOATING
C2465 VDD.n715 GND 0.02fF $ **FLOATING
C2466 VDD.n716 GND 0.02fF $ **FLOATING
C2467 VDD.t75 GND 0.09fF
C2468 VDD.t170 GND 0.09fF
C2469 VDD.n717 GND 0.94fF $ **FLOATING
C2470 VDD.n718 GND 0.01fF $ **FLOATING
C2471 VDD.n719 GND 0.40fF $ **FLOATING
C2472 VDD.n720 GND 0.02fF $ **FLOATING
C2473 VDD.n721 GND 0.02fF $ **FLOATING
C2474 VDD.t74 GND 0.20fF
C2475 VDD.n722 GND 0.25fF $ **FLOATING
C2476 VDD.n723 GND 0.02fF $ **FLOATING
C2477 VDD.n724 GND 0.02fF $ **FLOATING
C2478 VDD.n725 GND 0.02fF $ **FLOATING
C2479 VDD.n726 GND 0.35fF $ **FLOATING
C2480 VDD.n727 GND 0.02fF $ **FLOATING
C2481 VDD.n728 GND 0.02fF $ **FLOATING
C2482 VDD.n729 GND 0.02fF $ **FLOATING
C2483 VDD.t8 GND 0.24fF
C2484 VDD.n730 GND 0.27fF $ **FLOATING
C2485 VDD.n731 GND 0.02fF $ **FLOATING
C2486 VDD.n732 GND 0.02fF $ **FLOATING
C2487 VDD.n733 GND 0.02fF $ **FLOATING
C2488 VDD.n734 GND 0.48fF $ **FLOATING
C2489 VDD.n735 GND 0.02fF $ **FLOATING
C2490 VDD.n736 GND 0.02fF $ **FLOATING
C2491 VDD.n737 GND 0.02fF $ **FLOATING
C2492 VDD.n738 GND 0.95fF $ **FLOATING
C2493 VDD.n739 GND 0.35fF $ **FLOATING
C2494 VDD.n740 GND 0.08fF $ **FLOATING
C2495 VDD.n741 GND 0.20fF $ **FLOATING
C2496 VDD.n742 GND 0.08fF $ **FLOATING
C2497 VDD.n743 GND 0.27fF $ **FLOATING
C2498 VDD.n744 GND 0.02fF $ **FLOATING
C2499 VDD.n745 GND 0.02fF $ **FLOATING
C2500 VDD.n746 GND 0.02fF $ **FLOATING
C2501 VDD.n747 GND 0.48fF $ **FLOATING
C2502 VDD.t127 GND 0.13fF
C2503 VDD.n748 GND 0.14fF $ **FLOATING
C2504 VDD.n749 GND 0.02fF $ **FLOATING
C2505 VDD.n750 GND 0.02fF $ **FLOATING
C2506 VDD.n751 GND 0.02fF $ **FLOATING
C2507 VDD.n752 GND 0.48fF $ **FLOATING
C2508 VDD.n753 GND 0.24fF $ **FLOATING
C2509 VDD.n754 GND 0.02fF $ **FLOATING
C2510 VDD.n755 GND 0.02fF $ **FLOATING
C2511 VDD.n756 GND 0.01fF $ **FLOATING
C2512 VDD.n757 GND 0.24fF $ **FLOATING
C2513 VDD.n758 GND 0.02fF $ **FLOATING
C2514 VDD.n759 GND 0.02fF $ **FLOATING
C2515 VDD.n760 GND 0.02fF $ **FLOATING
C2516 VDD.t140 GND 0.65fF
C2517 VDD.t32 GND 0.25fF
C2518 VDD.t106 GND 0.62fF
C2519 VDD.t155 GND 0.27fF
C2520 VDD.n761 GND 0.29fF $ **FLOATING
C2521 VDD.n762 GND 0.16fF $ **FLOATING
C2522 VDD.n763 GND 0.02fF $ **FLOATING
C2523 VDD.n764 GND 0.02fF $ **FLOATING
C2524 VDD.n765 GND 0.02fF $ **FLOATING
C2525 VDD.t151 GND 0.09fF
C2526 VDD.n766 GND 0.47fF $ **FLOATING
C2527 VDD.n767 GND 0.01fF $ **FLOATING
C2528 VDD.n768 GND 0.19fF $ **FLOATING
C2529 VDD.n769 GND 0.02fF $ **FLOATING
C2530 VDD.n770 GND 0.02fF $ **FLOATING
C2531 VDD.t150 GND 0.12fF
C2532 VDD.n771 GND 0.15fF $ **FLOATING
C2533 VDD.n772 GND 0.02fF $ **FLOATING
C2534 VDD.n773 GND 0.02fF $ **FLOATING
C2535 VDD.n774 GND 0.02fF $ **FLOATING
C2536 VDD.n775 GND 0.21fF $ **FLOATING
C2537 VDD.n776 GND 0.02fF $ **FLOATING
C2538 VDD.n777 GND 0.02fF $ **FLOATING
C2539 VDD.n778 GND 0.02fF $ **FLOATING
C2540 VDD.t88 GND 0.14fF
C2541 VDD.n779 GND 0.16fF $ **FLOATING
C2542 VDD.n780 GND 0.02fF $ **FLOATING
C2543 VDD.n781 GND 0.02fF $ **FLOATING
C2544 VDD.n782 GND 0.02fF $ **FLOATING
C2545 VDD.n783 GND 0.48fF $ **FLOATING
C2546 VDD.n784 GND 0.26fF $ **FLOATING
C2547 VDD.n785 GND 0.02fF $ **FLOATING
C2548 VDD.n786 GND 0.02fF $ **FLOATING
C2549 VDD.n787 GND 0.01fF $ **FLOATING
C2550 VDD.n788 GND 0.48fF $ **FLOATING
C2551 VDD.n789 GND 0.24fF $ **FLOATING
C2552 VDD.n790 GND 0.08fF $ **FLOATING
C2553 VDD.n791 GND 0.32fF $ **FLOATING
C2554 VDD.n792 GND 0.08fF $ **FLOATING
C2555 VDD.n793 GND 0.49fF $ **FLOATING
C2556 VDD.n794 GND 0.02fF $ **FLOATING
C2557 VDD.n795 GND 0.02fF $ **FLOATING
C2558 VDD.n796 GND 0.02fF $ **FLOATING
C2559 VDD.t18 GND 0.24fF
C2560 VDD.n797 GND 0.25fF $ **FLOATING
C2561 VDD.n798 GND 0.02fF $ **FLOATING
C2562 VDD.n799 GND 0.02fF $ **FLOATING
C2563 VDD.n800 GND 0.02fF $ **FLOATING
C2564 VDD.n801 GND 0.95fF $ **FLOATING
C2565 VDD.n802 GND 0.40fF $ **FLOATING
C2566 VDD.n803 GND 0.02fF $ **FLOATING
C2567 VDD.n804 GND 0.02fF $ **FLOATING
C2568 VDD.n805 GND 0.01fF $ **FLOATING
C2569 VDD.n806 GND 0.40fF $ **FLOATING
C2570 VDD.n807 GND 0.02fF $ **FLOATING
C2571 VDD.n808 GND 0.02fF $ **FLOATING
C2572 VDD.n809 GND 0.02fF $ **FLOATING
C2573 VDD.n810 GND 0.40fF $ **FLOATING
C2574 VDD.n811 GND 0.02fF $ **FLOATING
C2575 VDD.n812 GND 0.02fF $ **FLOATING
C2576 VDD.n813 GND 0.02fF $ **FLOATING
C2577 VDD.n814 GND 0.40fF $ **FLOATING
C2578 VDD.n815 GND 0.02fF $ **FLOATING
C2579 VDD.n816 GND 0.02fF $ **FLOATING
C2580 VDD.n817 GND 0.02fF $ **FLOATING
C2581 VDD.n818 GND 0.95fF $ **FLOATING
C2582 VDD.t152 GND 0.20fF
C2583 VDD.n819 GND 0.27fF $ **FLOATING
C2584 VDD.n820 GND 0.02fF $ **FLOATING
C2585 VDD.n821 GND 0.02fF $ **FLOATING
C2586 VDD.n822 GND 0.02fF $ **FLOATING
C2587 VDD.n823 GND 0.34fF $ **FLOATING
C2588 VDD.n824 GND 0.02fF $ **FLOATING
C2589 VDD.n825 GND 0.02fF $ **FLOATING
C2590 VDD.n826 GND 0.02fF $ **FLOATING
C2591 VDD.t101 GND 0.20fF
C2592 VDD.n827 GND 0.28fF $ **FLOATING
C2593 VDD.n828 GND 0.02fF $ **FLOATING
C2594 VDD.n829 GND 0.02fF $ **FLOATING
C2595 VDD.n830 GND 0.02fF $ **FLOATING
C2596 VDD.n831 GND 0.32fF $ **FLOATING
C2597 VDD.n832 GND 0.02fF $ **FLOATING
C2598 VDD.n833 GND 0.02fF $ **FLOATING
C2599 VDD.n834 GND 0.02fF $ **FLOATING
C2600 VDD.n835 GND 0.02fF $ **FLOATING
C2601 VDD.n836 GND 0.30fF $ **FLOATING
C2602 VDD.n837 GND 0.02fF $ **FLOATING
C2603 VDD.n838 GND 0.02fF $ **FLOATING
C2604 VDD.t142 GND 0.20fF
C2605 VDD.n839 GND 0.30fF $ **FLOATING
C2606 VDD.n840 GND 0.02fF $ **FLOATING
C2607 VDD.n841 GND 0.02fF $ **FLOATING
C2608 VDD.n842 GND 0.02fF $ **FLOATING
C2609 VDD.n843 GND 0.32fF $ **FLOATING
C2610 VDD.n844 GND 0.02fF $ **FLOATING
C2611 VDD.n845 GND 0.02fF $ **FLOATING
C2612 VDD.n846 GND 0.02fF $ **FLOATING
C2613 VDD.t30 GND 0.20fF
C2614 VDD.n847 GND 0.32fF $ **FLOATING
C2615 VDD.n848 GND 0.02fF $ **FLOATING
C2616 VDD.n849 GND 0.02fF $ **FLOATING
C2617 VDD.n850 GND 0.02fF $ **FLOATING
C2618 VDD.n851 GND 0.95fF $ **FLOATING
C2619 VDD.n852 GND 0.47fF $ **FLOATING
C2620 VDD.n853 GND 0.02fF $ **FLOATING
C2621 VDD.n854 GND 0.02fF $ **FLOATING
C2622 VDD.n855 GND 0.02fF $ **FLOATING
C2623 VDD.n856 GND 0.36fF $ **FLOATING
C2624 VDD.n857 GND 0.03fF $ **FLOATING
C2625 CMOS_sbox_0/CMOS_s1_0/VDD GND 0.01fF $ **FLOATING
C2626 VDD.n858 GND 0.84fF $ **FLOATING
C2627 VDD.n859 GND 0.43fF $ **FLOATING
C2628 VDD.n860 GND 0.03fF $ **FLOATING
C2629 VDD.n861 GND 0.29fF $ **FLOATING
C2630 VDD.n862 GND 0.38fF $ **FLOATING
C2631 VDD.n863 GND 0.25fF $ **FLOATING
C2632 VDD.n864 GND 0.02fF $ **FLOATING
C2633 VDD.n865 GND 0.02fF $ **FLOATING
C2634 VDD.n866 GND 0.00fF $ **FLOATING
C2635 VDD.t174 GND 0.13fF
C2636 VDD.n867 GND 0.14fF $ **FLOATING
C2637 VDD.n868 GND 0.02fF $ **FLOATING
C2638 VDD.n869 GND 0.02fF $ **FLOATING
C2639 VDD.n870 GND 0.06fF $ **FLOATING
C2640 VDD.t175 GND 0.09fF
C2641 VDD.t158 GND 0.09fF
C2642 CMOS_4in_XOR_0/CMOS_XOR_3/VDD GND 0.01fF $ **FLOATING
C2643 VDD.t16 GND 0.11fF
C2644 VDD.n871 GND 0.16fF $ **FLOATING
C2645 VDD.n872 GND 0.02fF $ **FLOATING
C2646 VDD.t87 GND 0.09fF
C2647 VDD.t91 GND 0.09fF
C2648 CMOS_4in_XOR_0/CMOS_XOR_1/VDD GND 0.01fF $ **FLOATING
C2649 VDD.t71 GND 0.09fF
C2650 VDD.t130 GND 0.09fF
C2651 VDD.n873 GND 0.48fF $ **FLOATING
C2652 VDD.n874 GND 0.38fF $ **FLOATING
C2653 VDD.n875 GND 0.25fF $ **FLOATING
C2654 VDD.n876 GND 0.02fF $ **FLOATING
C2655 VDD.n877 GND 0.02fF $ **FLOATING
C2656 VDD.n878 GND 0.00fF $ **FLOATING
C2657 CMOS_4in_XOR_0/CMOS_INV_0/VDD GND 0.01fF $ **FLOATING
C2658 VDD.n879 GND 0.06fF $ **FLOATING
C2659 VDD.t129 GND 0.13fF
C2660 VDD.n880 GND 0.14fF $ **FLOATING
C2661 VDD.n881 GND 0.02fF $ **FLOATING
C2662 VDD.n882 GND 0.02fF $ **FLOATING
C2663 VDD.n883 GND 0.22fF $ **FLOATING
C2664 VDD.n884 GND 0.02fF $ **FLOATING
C2665 VDD.n885 GND 0.02fF $ **FLOATING
C2666 VDD.n886 GND 0.01fF $ **FLOATING
C2667 VDD.n887 GND 0.22fF $ **FLOATING
C2668 VDD.n888 GND 0.02fF $ **FLOATING
C2669 VDD.n889 GND 0.02fF $ **FLOATING
C2670 VDD.n890 GND 0.02fF $ **FLOATING
C2671 VDD.n891 GND 0.22fF $ **FLOATING
C2672 VDD.n892 GND 0.02fF $ **FLOATING
C2673 VDD.n893 GND 0.02fF $ **FLOATING
C2674 VDD.n894 GND 0.02fF $ **FLOATING
C2675 VDD.n895 GND 0.22fF $ **FLOATING
C2676 VDD.n896 GND 0.02fF $ **FLOATING
C2677 VDD.n897 GND 0.02fF $ **FLOATING
C2678 VDD.n898 GND 0.02fF $ **FLOATING
C2679 VDD.n899 GND 0.48fF $ **FLOATING
C2680 VDD.t70 GND 0.11fF
C2681 VDD.n900 GND 0.15fF $ **FLOATING
C2682 VDD.n901 GND 0.02fF $ **FLOATING
C2683 VDD.n902 GND 0.02fF $ **FLOATING
C2684 VDD.n903 GND 0.02fF $ **FLOATING
C2685 VDD.n904 GND 0.19fF $ **FLOATING
C2686 VDD.n905 GND 0.02fF $ **FLOATING
C2687 VDD.n906 GND 0.02fF $ **FLOATING
C2688 VDD.n907 GND 0.02fF $ **FLOATING
C2689 VDD.t10 GND 0.11fF
C2690 VDD.n908 GND 0.16fF $ **FLOATING
C2691 VDD.n909 GND 0.02fF $ **FLOATING
C2692 VDD.n910 GND 0.02fF $ **FLOATING
C2693 VDD.n911 GND 0.02fF $ **FLOATING
C2694 VDD.n912 GND 0.18fF $ **FLOATING
C2695 VDD.n913 GND 0.02fF $ **FLOATING
C2696 VDD.n914 GND 0.02fF $ **FLOATING
C2697 VDD.n915 GND 0.02fF $ **FLOATING
C2698 VDD.n916 GND 0.02fF $ **FLOATING
C2699 VDD.n917 GND 0.16fF $ **FLOATING
C2700 VDD.n918 GND 0.02fF $ **FLOATING
C2701 VDD.n919 GND 0.02fF $ **FLOATING
C2702 VDD.t11 GND 0.11fF
C2703 VDD.n920 GND 0.17fF $ **FLOATING
C2704 VDD.n921 GND 0.02fF $ **FLOATING
C2705 VDD.n922 GND 0.02fF $ **FLOATING
C2706 VDD.n923 GND 0.02fF $ **FLOATING
C2707 VDD.n924 GND 0.17fF $ **FLOATING
C2708 VDD.n925 GND 0.02fF $ **FLOATING
C2709 VDD.n926 GND 0.02fF $ **FLOATING
C2710 VDD.n927 GND 0.02fF $ **FLOATING
C2711 VDD.t90 GND 0.11fF
C2712 VDD.n928 GND 0.17fF $ **FLOATING
C2713 VDD.n929 GND 0.02fF $ **FLOATING
C2714 VDD.n930 GND 0.02fF $ **FLOATING
C2715 VDD.n931 GND 0.02fF $ **FLOATING
C2716 VDD.n932 GND 0.48fF $ **FLOATING
C2717 VDD.n933 GND 0.25fF $ **FLOATING
C2718 VDD.n934 GND 0.02fF $ **FLOATING
C2719 VDD.n935 GND 0.02fF $ **FLOATING
C2720 VDD.n936 GND 0.02fF $ **FLOATING
C2721 VDD.n937 GND 0.14fF $ **FLOATING
C2722 VDD.n938 GND 0.46fF $ **FLOATING
C2723 VDD.t68 GND 0.09fF
C2724 VDD.t164 GND 0.09fF
C2725 CMOS_4in_XOR_0/CMOS_XOR_0/VDD GND 0.01fF $ **FLOATING
C2726 VDD.t36 GND 0.09fF
C2727 VDD.t94 GND 0.09fF
C2728 VDD.t165 GND 0.09fF
C2729 VDD.t145 GND 0.09fF
C2730 VDD.n939 GND 0.95fF $ **FLOATING
C2731 VDD.n940 GND 0.48fF $ **FLOATING
C2732 VDD.n941 GND 0.49fF $ **FLOATING
C2733 VDD.n942 GND 0.02fF $ **FLOATING
C2734 VDD.n943 GND 0.02fF $ **FLOATING
C2735 VDD.n944 GND 0.00fF $ **FLOATING
C2736 CMOS_4in_XOR_0/CMOS_INV_1/VDD GND 0.01fF $ **FLOATING
C2737 VDD.n945 GND 0.06fF $ **FLOATING
C2738 VDD.t144 GND 0.24fF
C2739 VDD.n946 GND 0.25fF $ **FLOATING
C2740 VDD.n947 GND 0.02fF $ **FLOATING
C2741 VDD.n948 GND 0.02fF $ **FLOATING
C2742 VDD.n949 GND 0.40fF $ **FLOATING
C2743 VDD.n950 GND 0.02fF $ **FLOATING
C2744 VDD.n951 GND 0.02fF $ **FLOATING
C2745 VDD.n952 GND 0.01fF $ **FLOATING
C2746 VDD.n953 GND 0.40fF $ **FLOATING
C2747 VDD.n954 GND 0.02fF $ **FLOATING
C2748 VDD.n955 GND 0.02fF $ **FLOATING
C2749 VDD.n956 GND 0.02fF $ **FLOATING
C2750 VDD.n957 GND 0.40fF $ **FLOATING
C2751 VDD.n958 GND 0.02fF $ **FLOATING
C2752 VDD.n959 GND 0.02fF $ **FLOATING
C2753 VDD.n960 GND 0.02fF $ **FLOATING
C2754 VDD.n961 GND 0.40fF $ **FLOATING
C2755 VDD.n962 GND 0.02fF $ **FLOATING
C2756 VDD.n963 GND 0.02fF $ **FLOATING
C2757 VDD.n964 GND 0.02fF $ **FLOATING
C2758 VDD.n965 GND 0.95fF $ **FLOATING
C2759 VDD.t35 GND 0.20fF
C2760 VDD.n966 GND 0.27fF $ **FLOATING
C2761 VDD.n967 GND 0.02fF $ **FLOATING
C2762 VDD.n968 GND 0.02fF $ **FLOATING
C2763 VDD.n969 GND 0.02fF $ **FLOATING
C2764 VDD.n970 GND 0.34fF $ **FLOATING
C2765 VDD.n971 GND 0.02fF $ **FLOATING
C2766 VDD.n972 GND 0.02fF $ **FLOATING
C2767 VDD.n973 GND 0.02fF $ **FLOATING
C2768 VDD.t23 GND 0.20fF
C2769 VDD.n974 GND 0.28fF $ **FLOATING
C2770 VDD.n975 GND 0.02fF $ **FLOATING
C2771 VDD.n976 GND 0.02fF $ **FLOATING
C2772 VDD.n977 GND 0.02fF $ **FLOATING
C2773 VDD.n978 GND 0.32fF $ **FLOATING
C2774 VDD.n979 GND 0.02fF $ **FLOATING
C2775 VDD.n980 GND 0.02fF $ **FLOATING
C2776 VDD.n981 GND 0.02fF $ **FLOATING
C2777 VDD.n982 GND 0.02fF $ **FLOATING
C2778 VDD.n983 GND 0.30fF $ **FLOATING
C2779 VDD.n984 GND 0.02fF $ **FLOATING
C2780 VDD.n985 GND 0.02fF $ **FLOATING
C2781 VDD.t37 GND 0.20fF
C2782 VDD.n986 GND 0.30fF $ **FLOATING
C2783 VDD.n987 GND 0.02fF $ **FLOATING
C2784 VDD.n988 GND 0.02fF $ **FLOATING
C2785 VDD.n989 GND 0.02fF $ **FLOATING
C2786 VDD.n990 GND 0.32fF $ **FLOATING
C2787 VDD.n991 GND 0.02fF $ **FLOATING
C2788 VDD.n992 GND 0.02fF $ **FLOATING
C2789 VDD.n993 GND 0.02fF $ **FLOATING
C2790 VDD.t67 GND 0.20fF
C2791 VDD.n994 GND 0.32fF $ **FLOATING
C2792 VDD.n995 GND 0.02fF $ **FLOATING
C2793 VDD.n996 GND 0.02fF $ **FLOATING
C2794 VDD.n997 GND 0.02fF $ **FLOATING
C2795 VDD.n998 GND 0.95fF $ **FLOATING
C2796 VDD.n999 GND 0.47fF $ **FLOATING
C2797 VDD.n1000 GND 0.02fF $ **FLOATING
C2798 VDD.n1001 GND 0.02fF $ **FLOATING
C2799 VDD.n1002 GND 0.02fF $ **FLOATING
C2800 VDD.n1003 GND 0.20fF $ **FLOATING
C2801 VDD.n1004 GND 0.03fF $ **FLOATING
C2802 VDD.n1005 GND 0.86fF $ **FLOATING
C2803 CMOS_4in_XOR_0/VDD GND 0.01fF $ **FLOATING
C2804 VDD.n1006 GND 0.43fF $ **FLOATING
C2805 VDD.n1007 GND 0.14fF $ **FLOATING
C2806 VDD.n1008 GND 0.03fF $ **FLOATING
C2807 VDD.n1009 GND 0.25fF $ **FLOATING
C2808 VDD.n1010 GND 0.02fF $ **FLOATING
C2809 VDD.n1011 GND 0.02fF $ **FLOATING
C2810 VDD.n1012 GND 0.02fF $ **FLOATING
C2811 VDD.n1013 GND 0.48fF $ **FLOATING
C2812 VDD.t86 GND 0.11fF
C2813 VDD.n1014 GND 0.17fF $ **FLOATING
C2814 VDD.n1015 GND 0.02fF $ **FLOATING
C2815 VDD.n1016 GND 0.02fF $ **FLOATING
C2816 VDD.n1017 GND 0.02fF $ **FLOATING
C2817 VDD.n1018 GND 0.17fF $ **FLOATING
C2818 VDD.n1019 GND 0.02fF $ **FLOATING
C2819 VDD.n1020 GND 0.02fF $ **FLOATING
C2820 VDD.n1021 GND 0.02fF $ **FLOATING
C2821 VDD.n1022 GND 0.02fF $ **FLOATING
C2822 VDD.n1023 GND 0.17fF $ **FLOATING
C2823 VDD.n1024 GND 0.02fF $ **FLOATING
C2824 VDD.n1025 GND 0.02fF $ **FLOATING
C2825 VDD.n1026 GND 0.02fF $ **FLOATING
C2826 VDD.n1027 GND 0.02fF $ **FLOATING
C2827 VDD.n1028 GND 0.18fF $ **FLOATING
C2828 VDD.n1029 GND 0.02fF $ **FLOATING
C2829 VDD.n1030 GND 0.02fF $ **FLOATING
C2830 VDD.n1031 GND 0.02fF $ **FLOATING
C2831 VDD.t22 GND 0.11fF
C2832 VDD.n1032 GND 0.16fF $ **FLOATING
C2833 VDD.n1033 GND 0.02fF $ **FLOATING
C2834 VDD.n1034 GND 0.02fF $ **FLOATING
C2835 VDD.n1035 GND 0.02fF $ **FLOATING
C2836 VDD.n1036 GND 0.19fF $ **FLOATING
C2837 VDD.n1037 GND 0.02fF $ **FLOATING
C2838 VDD.n1038 GND 0.02fF $ **FLOATING
C2839 VDD.n1039 GND 0.02fF $ **FLOATING
C2840 VDD.t157 GND 0.11fF
C2841 VDD.n1040 GND 0.15fF $ **FLOATING
C2842 VDD.n1041 GND 0.02fF $ **FLOATING
C2843 VDD.n1042 GND 0.02fF $ **FLOATING
C2844 VDD.n1043 GND 0.02fF $ **FLOATING
C2845 VDD.n1044 GND 0.48fF $ **FLOATING
C2846 VDD.n1045 GND 0.22fF $ **FLOATING
C2847 VDD.n1046 GND 0.02fF $ **FLOATING
C2848 VDD.n1047 GND 0.02fF $ **FLOATING
C2849 VDD.n1048 GND 0.02fF $ **FLOATING
C2850 VDD.n1049 GND 0.22fF $ **FLOATING
C2851 VDD.n1050 GND 0.02fF $ **FLOATING
C2852 VDD.n1051 GND 0.02fF $ **FLOATING
C2853 VDD.n1052 GND 0.02fF $ **FLOATING
C2854 VDD.n1053 GND 0.22fF $ **FLOATING
C2855 VDD.n1054 GND 0.02fF $ **FLOATING
C2856 VDD.n1055 GND 0.02fF $ **FLOATING
C2857 VDD.n1056 GND 0.02fF $ **FLOATING
C2858 VDD.n1057 GND 0.22fF $ **FLOATING
C2859 VDD.n1058 GND 0.02fF $ **FLOATING
C2860 VDD.n1059 GND 0.02fF $ **FLOATING
C2861 VDD.n1060 GND 0.01fF $ **FLOATING
C2862 VDD.n1061 GND 0.48fF $ **FLOATING
C2863 CMOS_4in_XOR_0/CMOS_INV_2/VDD GND 0.01fF $ **FLOATING
C2864 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n0 GND 0.55fF $ **FLOATING
C2865 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n1 GND 0.32fF $ **FLOATING
C2866 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n2 GND 0.18fF $ **FLOATING
C2867 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n3 GND 0.21fF $ **FLOATING
C2868 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n4 GND 0.09fF $ **FLOATING
C2869 CMOS_sbox_0/CMOS_s0_0/x2 GND 1.13fF $ **FLOATING
C2870 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t13 GND 0.21fF
C2871 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t14 GND 0.14fF
C2872 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n5 GND 0.29fF $ **FLOATING
C2873 CMOS_4in_XOR_0/CMOS_INV_3/A GND 0.16fF $ **FLOATING
C2874 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t9 GND 0.79fF
C2875 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t12 GND 0.53fF
C2876 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/B GND 0.63fF $ **FLOATING
C2877 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t10 GND 0.23fF
C2878 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t8 GND 0.28fF
C2879 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/D GND 0.47fF $ **FLOATING
C2880 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t5 GND 0.27fF
C2881 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t4 GND 0.11fF
C2882 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n6 GND 0.30fF $ **FLOATING
C2883 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/A GND 0.04fF $ **FLOATING
C2884 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n7 GND 1.72fF $ **FLOATING
C2885 CMOS_sbox_0/CMOS_s3_0/x2 GND 4.89fF $ **FLOATING
C2886 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n8 GND 2.36fF $ **FLOATING
C2887 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n9 GND 2.50fF $ **FLOATING
C2888 CMOS_sbox_0/CMOS_s2_0/x2 GND 1.53fF $ **FLOATING
C2889 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t15 GND 0.79fF
C2890 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t6 GND 0.53fF
C2891 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t7 GND 0.30fF
C2892 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t11 GND 0.25fF
C2893 CMOS_sbox_0/CMOS_s0_0/CMOS_AND_2/A GND 0.44fF $ **FLOATING
C2894 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n10 GND 3.97fF $ **FLOATING
C2895 CMOS_sbox_0/CMOS_s1_0/x2 GND 1.01fF $ **FLOATING
C2896 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n11 GND 1.15fF $ **FLOATING
C2897 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n12 GND 2.22fF $ **FLOATING
C2898 CMOS_4in_XOR_0/XOR2 GND 0.39fF $ **FLOATING
C2899 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n13 GND 0.40fF $ **FLOATING
C2900 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n14 GND 0.10fF $ **FLOATING
C2901 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t1 GND 0.14fF
C2902 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t2 GND 0.14fF
C2903 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n15 GND 0.28fF $ **FLOATING
C2904 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n16 GND 0.06fF $ **FLOATING
C2905 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n17 GND 0.02fF $ **FLOATING
C2906 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n18 GND 0.01fF $ **FLOATING
C2907 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n19 GND 0.04fF $ **FLOATING
C2908 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n20 GND 0.04fF $ **FLOATING
C2909 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n21 GND 0.04fF $ **FLOATING
C2910 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n22 GND 0.04fF $ **FLOATING
C2911 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n23 GND 0.02fF $ **FLOATING
C2912 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n24 GND 0.06fF $ **FLOATING
C2913 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n25 GND 0.01fF $ **FLOATING
C2914 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n26 GND 0.06fF $ **FLOATING
C2915 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n27 GND 0.01fF $ **FLOATING
C2916 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n28 GND 0.04fF $ **FLOATING
C2917 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n29 GND 0.02fF $ **FLOATING
C2918 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n30 GND 0.01fF $ **FLOATING
C2919 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n31 GND 0.04fF $ **FLOATING
C2920 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n32 GND 0.02fF $ **FLOATING
C2921 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n33 GND 0.01fF $ **FLOATING
C2922 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n34 GND 0.01fF $ **FLOATING
C2923 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n35 GND 0.28fF $ **FLOATING
C2924 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n36 GND 0.04fF $ **FLOATING
C2925 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n37 GND 0.04fF $ **FLOATING
C2926 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n38 GND 0.01fF $ **FLOATING
C2927 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n39 GND 0.26fF $ **FLOATING
C2928 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t3 GND 0.28fF
C2929 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.t0 GND 0.28fF
C2930 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n40 GND 0.56fF $ **FLOATING
C2931 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n41 GND 0.00fF $ **FLOATING
C2932 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n42 GND 0.04fF $ **FLOATING
C2933 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n43 GND 0.04fF $ **FLOATING
C2934 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n44 GND 0.01fF $ **FLOATING
C2935 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n45 GND 0.18fF $ **FLOATING
C2936 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n46 GND 0.02fF $ **FLOATING
C2937 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n47 GND 0.01fF $ **FLOATING
C2938 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n48 GND 0.04fF $ **FLOATING
C2939 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n49 GND 0.01fF $ **FLOATING
C2940 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n50 GND 0.02fF $ **FLOATING
C2941 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n51 GND 0.04fF $ **FLOATING
C2942 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/B.n52 GND 0.22fF $ **FLOATING
C2943 CMOS_4in_XOR_0/CMOS_XOR_0/XOR GND 0.13fF $ **FLOATING
C2944 CMOS_sbox_0/CMOS_s0_0/x3_bar GND 0.53fF $ **FLOATING
C2945 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t17 GND 0.27fF
C2946 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t10 GND 0.24fF
C2947 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/A_bar GND 0.40fF $ **FLOATING
C2948 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t6 GND 0.20fF
C2949 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t4 GND 0.20fF
C2950 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n0 GND 0.53fF $ **FLOATING
C2951 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/B_bar GND 0.13fF $ **FLOATING
C2952 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n1 GND 1.17fF $ **FLOATING
C2953 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n2 GND 1.69fF $ **FLOATING
C2954 CMOS_sbox_0/CMOS_s1_0/x3_bar GND 1.48fF $ **FLOATING
C2955 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t3 GND 0.20fF
C2956 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t13 GND 0.18fF
C2957 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n3 GND 1.17fF $ **FLOATING
C2958 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n4 GND 2.12fF $ **FLOATING
C2959 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t11 GND 0.27fF
C2960 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t14 GND 0.24fF
C2961 CMOS_sbox_0/CMOS_s2_0/CMOS_XNOR_0/A_bar GND 0.40fF $ **FLOATING
C2962 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t2 GND 0.12fF
C2963 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t8 GND 0.17fF
C2964 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n5 GND 0.24fF $ **FLOATING
C2965 CMOS_sbox_0/CMOS_s3_0/CMOS_AND_1/B GND 0.03fF $ **FLOATING
C2966 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n6 GND 0.76fF $ **FLOATING
C2967 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t7 GND 0.20fF
C2968 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t15 GND 0.18fF
C2969 CMOS_sbox_0/CMOS_s3_0/CMOS_XOR_0/B_bar GND 0.03fF $ **FLOATING
C2970 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n7 GND 1.17fF $ **FLOATING
C2971 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n8 GND 4.21fF $ **FLOATING
C2972 CMOS_sbox_0/CMOS_s3_0/x3_bar GND 1.28fF $ **FLOATING
C2973 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t5 GND 0.09fF
C2974 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t16 GND 0.20fF
C2975 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n9 GND 0.21fF $ **FLOATING
C2976 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/A GND 0.29fF $ **FLOATING
C2977 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n10 GND 1.36fF $ **FLOATING
C2978 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n11 GND 1.52fF $ **FLOATING
C2979 CMOS_sbox_0/CMOS_s2_0/x3_bar GND 0.80fF $ **FLOATING
C2980 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t12 GND 0.19fF
C2981 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t9 GND 0.23fF
C2982 CMOS_sbox_0/CMOS_s1_0/CMOS_3in_AND_0/A GND 0.03fF $ **FLOATING
C2983 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n12 GND 0.25fF $ **FLOATING
C2984 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n13 GND 1.42fF $ **FLOATING
C2985 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n14 GND 1.25fF $ **FLOATING
C2986 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t1 GND 0.46fF
C2987 CMOS_4in_XOR_0/XOR3_bar GND 0.15fF $ **FLOATING
C2988 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.n15 GND 0.62fF $ **FLOATING
C2989 CMOS_sbox_0/CMOS_s1_0/CMOS_XOR_0/B_bar.t0 GND 1.18fF
C2990 CMOS_4in_XOR_0/CMOS_INV_0/OUT GND 0.43fF $ **FLOATING
C2991 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n0 GND 0.36fF $ **FLOATING
C2992 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n1 GND 0.21fF $ **FLOATING
C2993 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n2 GND 0.12fF $ **FLOATING
C2994 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n3 GND 0.14fF $ **FLOATING
C2995 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n4 GND 0.06fF $ **FLOATING
C2996 CMOS_sbox_0/CMOS_s0_0/x0 GND 0.38fF $ **FLOATING
C2997 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t13 GND 0.13fF
C2998 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t19 GND 0.09fF
C2999 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n5 GND 0.19fF $ **FLOATING
C3000 CMOS_4in_XOR_0/CMOS_INV_2/A GND 0.10fF $ **FLOATING
C3001 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t8 GND 0.52fF
C3002 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t14 GND 0.35fF
C3003 CMOS_sbox_0/CMOS_s0_0/CMOS_XNOR_0/B GND 0.50fF $ **FLOATING
C3004 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t6 GND 0.52fF
C3005 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t10 GND 0.35fF
C3006 CMOS_sbox_0/CMOS_s3_0/CMOS_XNOR_0/B GND 0.50fF $ **FLOATING
C3007 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t7 GND 0.20fF
C3008 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t18 GND 0.16fF
C3009 CMOS_sbox_0/CMOS_s3_0/CMOS_3in_AND_0/B GND 0.43fF $ **FLOATING
C3010 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n6 GND 3.48fF $ **FLOATING
C3011 CMOS_sbox_0/CMOS_s3_0/x0 GND 0.42fF $ **FLOATING
C3012 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t16 GND 0.09fF
C3013 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t12 GND 0.14fF
C3014 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n7 GND 0.16fF $ **FLOATING
C3015 CMOS_sbox_0/CMOS_s2_0/CMOS_4in_AND_0/C GND 0.33fF $ **FLOATING
C3016 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n8 GND 1.68fF $ **FLOATING
C3017 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t9 GND 0.52fF
C3018 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t15 GND 0.35fF
C3019 CMOS_sbox_0/CMOS_s2_0/CMOS_XOR_0/B GND 0.39fF $ **FLOATING
C3020 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n9 GND 2.32fF $ **FLOATING
C3021 CMOS_sbox_0/CMOS_s2_0/x0 GND 0.92fF $ **FLOATING
C3022 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t17 GND 0.18fF
C3023 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t4 GND 0.07fF
C3024 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n10 GND 0.20fF $ **FLOATING
C3025 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n11 GND 1.70fF $ **FLOATING
C3026 CMOS_sbox_0/CMOS_s1_0/x0 GND 0.49fF $ **FLOATING
C3027 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n12 GND 1.37fF $ **FLOATING
C3028 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t5 GND 0.18fF
C3029 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t11 GND 0.07fF
C3030 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n13 GND 0.20fF $ **FLOATING
C3031 CMOS_sbox_0/CMOS_s0_0/CMOS_XOR_0/A GND 0.31fF $ **FLOATING
C3032 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n14 GND 1.30fF $ **FLOATING
C3033 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n15 GND 0.52fF $ **FLOATING
C3034 CMOS_4in_XOR_0/XOR0 GND 0.22fF $ **FLOATING
C3035 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n16 GND 0.26fF $ **FLOATING
C3036 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n17 GND 0.07fF $ **FLOATING
C3037 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t2 GND 0.09fF
C3038 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t3 GND 0.09fF
C3039 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n18 GND 0.18fF $ **FLOATING
C3040 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n19 GND 0.04fF $ **FLOATING
C3041 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n20 GND 0.02fF $ **FLOATING
C3042 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n21 GND 0.01fF $ **FLOATING
C3043 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n22 GND 0.03fF $ **FLOATING
C3044 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n23 GND 0.03fF $ **FLOATING
C3045 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n24 GND 0.03fF $ **FLOATING
C3046 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n25 GND 0.03fF $ **FLOATING
C3047 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n26 GND 0.02fF $ **FLOATING
C3048 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n27 GND 0.04fF $ **FLOATING
C3049 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n28 GND 0.01fF $ **FLOATING
C3050 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n29 GND 0.04fF $ **FLOATING
C3051 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n30 GND 0.01fF $ **FLOATING
C3052 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n31 GND 0.03fF $ **FLOATING
C3053 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n32 GND 0.02fF $ **FLOATING
C3054 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n33 GND 0.01fF $ **FLOATING
C3055 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n34 GND 0.03fF $ **FLOATING
C3056 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n35 GND 0.02fF $ **FLOATING
C3057 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n36 GND 0.01fF $ **FLOATING
C3058 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n37 GND 0.01fF $ **FLOATING
C3059 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n38 GND 0.18fF $ **FLOATING
C3060 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n39 GND 0.03fF $ **FLOATING
C3061 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n40 GND 0.03fF $ **FLOATING
C3062 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n41 GND 0.01fF $ **FLOATING
C3063 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n42 GND 0.17fF $ **FLOATING
C3064 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t1 GND 0.18fF
C3065 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.t0 GND 0.18fF
C3066 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n43 GND 0.36fF $ **FLOATING
C3067 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n44 GND 0.00fF $ **FLOATING
C3068 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n45 GND 0.03fF $ **FLOATING
C3069 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n46 GND 0.03fF $ **FLOATING
C3070 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n47 GND 0.01fF $ **FLOATING
C3071 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n48 GND 0.12fF $ **FLOATING
C3072 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n49 GND 0.02fF $ **FLOATING
C3073 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n50 GND 0.01fF $ **FLOATING
C3074 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n51 GND 0.03fF $ **FLOATING
C3075 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n52 GND 0.01fF $ **FLOATING
C3076 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n53 GND 0.02fF $ **FLOATING
C3077 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n54 GND 0.03fF $ **FLOATING
C3078 CMOS_sbox_0/CMOS_s1_0/CMOS_XNOR_0/A.n55 GND 0.15fF $ **FLOATING
C3079 CMOS_4in_XOR_0/CMOS_XOR_3/XOR GND 0.09fF $ **FLOATING
.ends

