magic
tech sky130A
magscale 1 2
timestamp 1675192118
<< nwell >>
rect -105 1114 2255 1304
rect 2535 1114 4025 1304
rect 4285 1114 6045 1304
rect 665 724 1485 1114
rect 2875 724 3695 1114
rect 4755 724 5575 1114
rect 665 -1066 1485 -676
rect 2875 -1066 3695 -676
rect 4755 -1066 5575 -676
rect -145 -1387 2275 -1066
rect 2535 -1256 4025 -1066
rect 4285 -1256 6045 -1066
rect 665 -1777 1485 -1387
rect 2536 -1706 4026 -1516
rect 4305 -1706 6385 -1516
rect 2876 -2096 3696 -1706
rect 4935 -2096 5755 -1706
<< pwell >>
rect -91 -492 2241 540
rect 2569 -492 4001 540
rect 4299 -492 6031 540
rect -91 -2721 2241 -2281
rect -111 -2873 2261 -2721
rect 2570 -2872 4002 -2280
rect 4329 -2720 6361 -2280
rect 4319 -2872 6371 -2720
<< nmos >>
rect 55 214 85 514
rect 205 214 235 514
rect 355 214 385 514
rect 505 214 535 514
rect 835 214 865 514
rect 985 214 1015 514
rect 1135 214 1165 514
rect 1285 214 1315 514
rect 1615 214 1645 514
rect 1765 214 1795 514
rect 1915 214 1945 514
rect 2065 214 2095 514
rect 2715 214 2745 514
rect 3045 214 3075 514
rect 3195 214 3225 514
rect 3345 214 3375 514
rect 3495 214 3525 514
rect 3825 214 3855 514
rect 4445 214 4475 514
rect 4595 214 4625 514
rect 4925 214 4955 514
rect 5075 214 5105 514
rect 5225 214 5255 514
rect 5375 214 5405 514
rect 5705 214 5735 514
rect 5855 214 5885 514
rect 55 -466 85 -166
rect 205 -466 235 -166
rect 355 -466 385 -166
rect 505 -466 535 -166
rect 835 -466 865 -166
rect 985 -466 1015 -166
rect 1135 -466 1165 -166
rect 1285 -466 1315 -166
rect 1615 -466 1645 -166
rect 1765 -466 1795 -166
rect 1915 -466 1945 -166
rect 2065 -466 2095 -166
rect 2715 -466 2745 -166
rect 3045 -466 3075 -166
rect 3195 -466 3225 -166
rect 3345 -466 3375 -166
rect 3495 -466 3525 -166
rect 3825 -466 3855 -166
rect 4445 -466 4475 -166
rect 4595 -466 4625 -166
rect 4925 -466 4955 -166
rect 5075 -466 5105 -166
rect 5225 -466 5255 -166
rect 5375 -466 5405 -166
rect 5705 -466 5735 -166
rect 5855 -466 5885 -166
rect 55 -2607 85 -2307
rect 205 -2607 235 -2307
rect 355 -2607 385 -2307
rect 505 -2607 535 -2307
rect 835 -2607 865 -2307
rect 985 -2607 1015 -2307
rect 1135 -2607 1165 -2307
rect 1285 -2607 1315 -2307
rect 1615 -2607 1645 -2307
rect 1765 -2607 1795 -2307
rect 1915 -2607 1945 -2307
rect 2065 -2607 2095 -2307
rect 2716 -2606 2746 -2306
rect 3046 -2606 3076 -2306
rect 3196 -2606 3226 -2306
rect 3346 -2606 3376 -2306
rect 3496 -2606 3526 -2306
rect 3826 -2606 3856 -2306
rect 4475 -2606 4505 -2306
rect 4625 -2606 4655 -2306
rect 4775 -2606 4805 -2306
rect 5105 -2606 5135 -2306
rect 5255 -2606 5285 -2306
rect 5405 -2606 5435 -2306
rect 5555 -2606 5585 -2306
rect 5885 -2606 5915 -2306
rect 6035 -2606 6065 -2306
rect 6185 -2606 6215 -2306
<< pmos >>
rect 835 774 865 1074
rect 985 774 1015 1074
rect 1135 774 1165 1074
rect 1285 774 1315 1074
rect 3045 774 3075 1074
rect 3195 774 3225 1074
rect 3345 774 3375 1074
rect 3495 774 3525 1074
rect 4925 774 4955 1074
rect 5075 774 5105 1074
rect 5225 774 5255 1074
rect 5375 774 5405 1074
rect 835 -1026 865 -726
rect 985 -1026 1015 -726
rect 1135 -1026 1165 -726
rect 1285 -1026 1315 -726
rect 3045 -1026 3075 -726
rect 3195 -1026 3225 -726
rect 3345 -1026 3375 -726
rect 3495 -1026 3525 -726
rect 4925 -1026 4955 -726
rect 5075 -1026 5105 -726
rect 5225 -1026 5255 -726
rect 5375 -1026 5405 -726
rect 835 -1727 865 -1427
rect 985 -1727 1015 -1427
rect 1135 -1727 1165 -1427
rect 1285 -1727 1315 -1427
rect 3046 -2046 3076 -1746
rect 3196 -2046 3226 -1746
rect 3346 -2046 3376 -1746
rect 3496 -2046 3526 -1746
rect 5105 -2046 5135 -1746
rect 5255 -2046 5285 -1746
rect 5405 -2046 5435 -1746
rect 5555 -2046 5585 -1746
<< ndiff >>
rect -65 441 55 514
rect -65 407 -22 441
rect 12 407 55 441
rect -65 361 55 407
rect -65 327 -22 361
rect 12 327 55 361
rect -65 281 55 327
rect -65 247 -22 281
rect 12 247 55 281
rect -65 214 55 247
rect 85 214 205 514
rect 235 441 355 514
rect 235 407 278 441
rect 312 407 355 441
rect 235 361 355 407
rect 235 327 278 361
rect 312 327 355 361
rect 235 281 355 327
rect 235 247 278 281
rect 312 247 355 281
rect 235 214 355 247
rect 385 214 505 514
rect 535 441 655 514
rect 535 407 578 441
rect 612 407 655 441
rect 535 361 655 407
rect 535 327 578 361
rect 612 327 655 361
rect 535 281 655 327
rect 535 247 578 281
rect 612 247 655 281
rect 535 214 655 247
rect 715 441 835 514
rect 715 407 758 441
rect 792 407 835 441
rect 715 361 835 407
rect 715 327 758 361
rect 792 327 835 361
rect 715 281 835 327
rect 715 247 758 281
rect 792 247 835 281
rect 715 214 835 247
rect 865 441 985 514
rect 865 407 908 441
rect 942 407 985 441
rect 865 361 985 407
rect 865 327 908 361
rect 942 327 985 361
rect 865 281 985 327
rect 865 247 908 281
rect 942 247 985 281
rect 865 214 985 247
rect 1015 441 1135 514
rect 1015 407 1058 441
rect 1092 407 1135 441
rect 1015 361 1135 407
rect 1015 327 1058 361
rect 1092 327 1135 361
rect 1015 281 1135 327
rect 1015 247 1058 281
rect 1092 247 1135 281
rect 1015 214 1135 247
rect 1165 441 1285 514
rect 1165 407 1208 441
rect 1242 407 1285 441
rect 1165 361 1285 407
rect 1165 327 1208 361
rect 1242 327 1285 361
rect 1165 281 1285 327
rect 1165 247 1208 281
rect 1242 247 1285 281
rect 1165 214 1285 247
rect 1315 441 1435 514
rect 1315 407 1358 441
rect 1392 407 1435 441
rect 1315 361 1435 407
rect 1315 327 1358 361
rect 1392 327 1435 361
rect 1315 281 1435 327
rect 1315 247 1358 281
rect 1392 247 1435 281
rect 1315 214 1435 247
rect 1495 441 1615 514
rect 1495 407 1538 441
rect 1572 407 1615 441
rect 1495 361 1615 407
rect 1495 327 1538 361
rect 1572 327 1615 361
rect 1495 281 1615 327
rect 1495 247 1538 281
rect 1572 247 1615 281
rect 1495 214 1615 247
rect 1645 214 1765 514
rect 1795 441 1915 514
rect 1795 407 1838 441
rect 1872 407 1915 441
rect 1795 361 1915 407
rect 1795 327 1838 361
rect 1872 327 1915 361
rect 1795 281 1915 327
rect 1795 247 1838 281
rect 1872 247 1915 281
rect 1795 214 1915 247
rect 1945 214 2065 514
rect 2095 441 2215 514
rect 2095 407 2138 441
rect 2172 407 2215 441
rect 2095 361 2215 407
rect 2095 327 2138 361
rect 2172 327 2215 361
rect 2095 281 2215 327
rect 2095 247 2138 281
rect 2172 247 2215 281
rect 2095 214 2215 247
rect 2595 441 2715 514
rect 2595 407 2638 441
rect 2672 407 2715 441
rect 2595 361 2715 407
rect 2595 327 2638 361
rect 2672 327 2715 361
rect 2595 281 2715 327
rect 2595 247 2638 281
rect 2672 247 2715 281
rect 2595 214 2715 247
rect 2745 441 2865 514
rect 2745 407 2788 441
rect 2822 407 2865 441
rect 2745 361 2865 407
rect 2745 327 2788 361
rect 2822 327 2865 361
rect 2745 281 2865 327
rect 2745 247 2788 281
rect 2822 247 2865 281
rect 2745 214 2865 247
rect 2925 441 3045 514
rect 2925 407 2968 441
rect 3002 407 3045 441
rect 2925 361 3045 407
rect 2925 327 2968 361
rect 3002 327 3045 361
rect 2925 281 3045 327
rect 2925 247 2968 281
rect 3002 247 3045 281
rect 2925 214 3045 247
rect 3075 441 3195 514
rect 3075 407 3118 441
rect 3152 407 3195 441
rect 3075 361 3195 407
rect 3075 327 3118 361
rect 3152 327 3195 361
rect 3075 281 3195 327
rect 3075 247 3118 281
rect 3152 247 3195 281
rect 3075 214 3195 247
rect 3225 441 3345 514
rect 3225 407 3268 441
rect 3302 407 3345 441
rect 3225 361 3345 407
rect 3225 327 3268 361
rect 3302 327 3345 361
rect 3225 281 3345 327
rect 3225 247 3268 281
rect 3302 247 3345 281
rect 3225 214 3345 247
rect 3375 441 3495 514
rect 3375 407 3418 441
rect 3452 407 3495 441
rect 3375 361 3495 407
rect 3375 327 3418 361
rect 3452 327 3495 361
rect 3375 281 3495 327
rect 3375 247 3418 281
rect 3452 247 3495 281
rect 3375 214 3495 247
rect 3525 441 3645 514
rect 3525 407 3568 441
rect 3602 407 3645 441
rect 3525 361 3645 407
rect 3525 327 3568 361
rect 3602 327 3645 361
rect 3525 281 3645 327
rect 3525 247 3568 281
rect 3602 247 3645 281
rect 3525 214 3645 247
rect 3705 441 3825 514
rect 3705 407 3748 441
rect 3782 407 3825 441
rect 3705 361 3825 407
rect 3705 327 3748 361
rect 3782 327 3825 361
rect 3705 281 3825 327
rect 3705 247 3748 281
rect 3782 247 3825 281
rect 3705 214 3825 247
rect 3855 441 3975 514
rect 3855 407 3898 441
rect 3932 407 3975 441
rect 3855 361 3975 407
rect 3855 327 3898 361
rect 3932 327 3975 361
rect 3855 281 3975 327
rect 3855 247 3898 281
rect 3932 247 3975 281
rect 3855 214 3975 247
rect 4325 441 4445 514
rect 4325 407 4368 441
rect 4402 407 4445 441
rect 4325 361 4445 407
rect 4325 327 4368 361
rect 4402 327 4445 361
rect 4325 281 4445 327
rect 4325 247 4368 281
rect 4402 247 4445 281
rect 4325 214 4445 247
rect 4475 441 4595 514
rect 4475 407 4518 441
rect 4552 407 4595 441
rect 4475 361 4595 407
rect 4475 327 4518 361
rect 4552 327 4595 361
rect 4475 281 4595 327
rect 4475 247 4518 281
rect 4552 247 4595 281
rect 4475 214 4595 247
rect 4625 441 4745 514
rect 4625 407 4668 441
rect 4702 407 4745 441
rect 4625 361 4745 407
rect 4625 327 4668 361
rect 4702 327 4745 361
rect 4625 281 4745 327
rect 4625 247 4668 281
rect 4702 247 4745 281
rect 4625 214 4745 247
rect 4805 441 4925 514
rect 4805 407 4848 441
rect 4882 407 4925 441
rect 4805 361 4925 407
rect 4805 327 4848 361
rect 4882 327 4925 361
rect 4805 281 4925 327
rect 4805 247 4848 281
rect 4882 247 4925 281
rect 4805 214 4925 247
rect 4955 441 5075 514
rect 4955 407 4998 441
rect 5032 407 5075 441
rect 4955 361 5075 407
rect 4955 327 4998 361
rect 5032 327 5075 361
rect 4955 281 5075 327
rect 4955 247 4998 281
rect 5032 247 5075 281
rect 4955 214 5075 247
rect 5105 441 5225 514
rect 5105 407 5148 441
rect 5182 407 5225 441
rect 5105 361 5225 407
rect 5105 327 5148 361
rect 5182 327 5225 361
rect 5105 281 5225 327
rect 5105 247 5148 281
rect 5182 247 5225 281
rect 5105 214 5225 247
rect 5255 441 5375 514
rect 5255 407 5298 441
rect 5332 407 5375 441
rect 5255 361 5375 407
rect 5255 327 5298 361
rect 5332 327 5375 361
rect 5255 281 5375 327
rect 5255 247 5298 281
rect 5332 247 5375 281
rect 5255 214 5375 247
rect 5405 441 5525 514
rect 5405 407 5448 441
rect 5482 407 5525 441
rect 5405 361 5525 407
rect 5405 327 5448 361
rect 5482 327 5525 361
rect 5405 281 5525 327
rect 5405 247 5448 281
rect 5482 247 5525 281
rect 5405 214 5525 247
rect 5585 441 5705 514
rect 5585 407 5628 441
rect 5662 407 5705 441
rect 5585 361 5705 407
rect 5585 327 5628 361
rect 5662 327 5705 361
rect 5585 281 5705 327
rect 5585 247 5628 281
rect 5662 247 5705 281
rect 5585 214 5705 247
rect 5735 214 5855 514
rect 5885 441 6005 514
rect 5885 407 5928 441
rect 5962 407 6005 441
rect 5885 361 6005 407
rect 5885 327 5928 361
rect 5962 327 6005 361
rect 5885 281 6005 327
rect 5885 247 5928 281
rect 5962 247 6005 281
rect 5885 214 6005 247
rect -65 -199 55 -166
rect -65 -233 -22 -199
rect 12 -233 55 -199
rect -65 -279 55 -233
rect -65 -313 -22 -279
rect 12 -313 55 -279
rect -65 -359 55 -313
rect -65 -393 -22 -359
rect 12 -393 55 -359
rect -65 -466 55 -393
rect 85 -466 205 -166
rect 235 -199 355 -166
rect 235 -233 278 -199
rect 312 -233 355 -199
rect 235 -279 355 -233
rect 235 -313 278 -279
rect 312 -313 355 -279
rect 235 -359 355 -313
rect 235 -393 278 -359
rect 312 -393 355 -359
rect 235 -466 355 -393
rect 385 -466 505 -166
rect 535 -199 655 -166
rect 535 -233 578 -199
rect 612 -233 655 -199
rect 535 -279 655 -233
rect 535 -313 578 -279
rect 612 -313 655 -279
rect 535 -359 655 -313
rect 535 -393 578 -359
rect 612 -393 655 -359
rect 535 -466 655 -393
rect 715 -199 835 -166
rect 715 -233 758 -199
rect 792 -233 835 -199
rect 715 -279 835 -233
rect 715 -313 758 -279
rect 792 -313 835 -279
rect 715 -359 835 -313
rect 715 -393 758 -359
rect 792 -393 835 -359
rect 715 -466 835 -393
rect 865 -199 985 -166
rect 865 -233 908 -199
rect 942 -233 985 -199
rect 865 -279 985 -233
rect 865 -313 908 -279
rect 942 -313 985 -279
rect 865 -359 985 -313
rect 865 -393 908 -359
rect 942 -393 985 -359
rect 865 -466 985 -393
rect 1015 -199 1135 -166
rect 1015 -233 1058 -199
rect 1092 -233 1135 -199
rect 1015 -279 1135 -233
rect 1015 -313 1058 -279
rect 1092 -313 1135 -279
rect 1015 -359 1135 -313
rect 1015 -393 1058 -359
rect 1092 -393 1135 -359
rect 1015 -466 1135 -393
rect 1165 -199 1285 -166
rect 1165 -233 1208 -199
rect 1242 -233 1285 -199
rect 1165 -279 1285 -233
rect 1165 -313 1208 -279
rect 1242 -313 1285 -279
rect 1165 -359 1285 -313
rect 1165 -393 1208 -359
rect 1242 -393 1285 -359
rect 1165 -466 1285 -393
rect 1315 -199 1435 -166
rect 1315 -233 1358 -199
rect 1392 -233 1435 -199
rect 1315 -279 1435 -233
rect 1315 -313 1358 -279
rect 1392 -313 1435 -279
rect 1315 -359 1435 -313
rect 1315 -393 1358 -359
rect 1392 -393 1435 -359
rect 1315 -466 1435 -393
rect 1495 -199 1615 -166
rect 1495 -233 1538 -199
rect 1572 -233 1615 -199
rect 1495 -279 1615 -233
rect 1495 -313 1538 -279
rect 1572 -313 1615 -279
rect 1495 -359 1615 -313
rect 1495 -393 1538 -359
rect 1572 -393 1615 -359
rect 1495 -466 1615 -393
rect 1645 -466 1765 -166
rect 1795 -199 1915 -166
rect 1795 -233 1838 -199
rect 1872 -233 1915 -199
rect 1795 -279 1915 -233
rect 1795 -313 1838 -279
rect 1872 -313 1915 -279
rect 1795 -359 1915 -313
rect 1795 -393 1838 -359
rect 1872 -393 1915 -359
rect 1795 -466 1915 -393
rect 1945 -466 2065 -166
rect 2095 -199 2215 -166
rect 2095 -233 2138 -199
rect 2172 -233 2215 -199
rect 2095 -279 2215 -233
rect 2095 -313 2138 -279
rect 2172 -313 2215 -279
rect 2095 -359 2215 -313
rect 2095 -393 2138 -359
rect 2172 -393 2215 -359
rect 2095 -466 2215 -393
rect 2595 -199 2715 -166
rect 2595 -233 2638 -199
rect 2672 -233 2715 -199
rect 2595 -279 2715 -233
rect 2595 -313 2638 -279
rect 2672 -313 2715 -279
rect 2595 -359 2715 -313
rect 2595 -393 2638 -359
rect 2672 -393 2715 -359
rect 2595 -466 2715 -393
rect 2745 -199 2865 -166
rect 2745 -233 2788 -199
rect 2822 -233 2865 -199
rect 2745 -279 2865 -233
rect 2745 -313 2788 -279
rect 2822 -313 2865 -279
rect 2745 -359 2865 -313
rect 2745 -393 2788 -359
rect 2822 -393 2865 -359
rect 2745 -466 2865 -393
rect 2925 -199 3045 -166
rect 2925 -233 2968 -199
rect 3002 -233 3045 -199
rect 2925 -279 3045 -233
rect 2925 -313 2968 -279
rect 3002 -313 3045 -279
rect 2925 -359 3045 -313
rect 2925 -393 2968 -359
rect 3002 -393 3045 -359
rect 2925 -466 3045 -393
rect 3075 -199 3195 -166
rect 3075 -233 3118 -199
rect 3152 -233 3195 -199
rect 3075 -279 3195 -233
rect 3075 -313 3118 -279
rect 3152 -313 3195 -279
rect 3075 -359 3195 -313
rect 3075 -393 3118 -359
rect 3152 -393 3195 -359
rect 3075 -466 3195 -393
rect 3225 -199 3345 -166
rect 3225 -233 3268 -199
rect 3302 -233 3345 -199
rect 3225 -279 3345 -233
rect 3225 -313 3268 -279
rect 3302 -313 3345 -279
rect 3225 -359 3345 -313
rect 3225 -393 3268 -359
rect 3302 -393 3345 -359
rect 3225 -466 3345 -393
rect 3375 -199 3495 -166
rect 3375 -233 3418 -199
rect 3452 -233 3495 -199
rect 3375 -279 3495 -233
rect 3375 -313 3418 -279
rect 3452 -313 3495 -279
rect 3375 -359 3495 -313
rect 3375 -393 3418 -359
rect 3452 -393 3495 -359
rect 3375 -466 3495 -393
rect 3525 -199 3645 -166
rect 3525 -233 3568 -199
rect 3602 -233 3645 -199
rect 3525 -279 3645 -233
rect 3525 -313 3568 -279
rect 3602 -313 3645 -279
rect 3525 -359 3645 -313
rect 3525 -393 3568 -359
rect 3602 -393 3645 -359
rect 3525 -466 3645 -393
rect 3705 -199 3825 -166
rect 3705 -233 3748 -199
rect 3782 -233 3825 -199
rect 3705 -279 3825 -233
rect 3705 -313 3748 -279
rect 3782 -313 3825 -279
rect 3705 -359 3825 -313
rect 3705 -393 3748 -359
rect 3782 -393 3825 -359
rect 3705 -466 3825 -393
rect 3855 -199 3975 -166
rect 3855 -233 3898 -199
rect 3932 -233 3975 -199
rect 3855 -279 3975 -233
rect 3855 -313 3898 -279
rect 3932 -313 3975 -279
rect 3855 -359 3975 -313
rect 3855 -393 3898 -359
rect 3932 -393 3975 -359
rect 3855 -466 3975 -393
rect 4325 -199 4445 -166
rect 4325 -233 4368 -199
rect 4402 -233 4445 -199
rect 4325 -279 4445 -233
rect 4325 -313 4368 -279
rect 4402 -313 4445 -279
rect 4325 -359 4445 -313
rect 4325 -393 4368 -359
rect 4402 -393 4445 -359
rect 4325 -466 4445 -393
rect 4475 -199 4595 -166
rect 4475 -233 4518 -199
rect 4552 -233 4595 -199
rect 4475 -279 4595 -233
rect 4475 -313 4518 -279
rect 4552 -313 4595 -279
rect 4475 -359 4595 -313
rect 4475 -393 4518 -359
rect 4552 -393 4595 -359
rect 4475 -466 4595 -393
rect 4625 -199 4745 -166
rect 4625 -233 4668 -199
rect 4702 -233 4745 -199
rect 4625 -279 4745 -233
rect 4625 -313 4668 -279
rect 4702 -313 4745 -279
rect 4625 -359 4745 -313
rect 4625 -393 4668 -359
rect 4702 -393 4745 -359
rect 4625 -466 4745 -393
rect 4805 -199 4925 -166
rect 4805 -233 4848 -199
rect 4882 -233 4925 -199
rect 4805 -279 4925 -233
rect 4805 -313 4848 -279
rect 4882 -313 4925 -279
rect 4805 -359 4925 -313
rect 4805 -393 4848 -359
rect 4882 -393 4925 -359
rect 4805 -466 4925 -393
rect 4955 -199 5075 -166
rect 4955 -233 4998 -199
rect 5032 -233 5075 -199
rect 4955 -279 5075 -233
rect 4955 -313 4998 -279
rect 5032 -313 5075 -279
rect 4955 -359 5075 -313
rect 4955 -393 4998 -359
rect 5032 -393 5075 -359
rect 4955 -466 5075 -393
rect 5105 -199 5225 -166
rect 5105 -233 5148 -199
rect 5182 -233 5225 -199
rect 5105 -279 5225 -233
rect 5105 -313 5148 -279
rect 5182 -313 5225 -279
rect 5105 -359 5225 -313
rect 5105 -393 5148 -359
rect 5182 -393 5225 -359
rect 5105 -466 5225 -393
rect 5255 -199 5375 -166
rect 5255 -233 5298 -199
rect 5332 -233 5375 -199
rect 5255 -279 5375 -233
rect 5255 -313 5298 -279
rect 5332 -313 5375 -279
rect 5255 -359 5375 -313
rect 5255 -393 5298 -359
rect 5332 -393 5375 -359
rect 5255 -466 5375 -393
rect 5405 -199 5525 -166
rect 5405 -233 5448 -199
rect 5482 -233 5525 -199
rect 5405 -279 5525 -233
rect 5405 -313 5448 -279
rect 5482 -313 5525 -279
rect 5405 -359 5525 -313
rect 5405 -393 5448 -359
rect 5482 -393 5525 -359
rect 5405 -466 5525 -393
rect 5585 -199 5705 -166
rect 5585 -233 5628 -199
rect 5662 -233 5705 -199
rect 5585 -279 5705 -233
rect 5585 -313 5628 -279
rect 5662 -313 5705 -279
rect 5585 -359 5705 -313
rect 5585 -393 5628 -359
rect 5662 -393 5705 -359
rect 5585 -466 5705 -393
rect 5735 -466 5855 -166
rect 5885 -199 6005 -166
rect 5885 -233 5928 -199
rect 5962 -233 6005 -199
rect 5885 -279 6005 -233
rect 5885 -313 5928 -279
rect 5962 -313 6005 -279
rect 5885 -359 6005 -313
rect 5885 -393 5928 -359
rect 5962 -393 6005 -359
rect 5885 -466 6005 -393
rect -65 -2380 55 -2307
rect -65 -2414 -22 -2380
rect 12 -2414 55 -2380
rect -65 -2460 55 -2414
rect -65 -2494 -22 -2460
rect 12 -2494 55 -2460
rect -65 -2540 55 -2494
rect -65 -2574 -22 -2540
rect 12 -2574 55 -2540
rect -65 -2607 55 -2574
rect 85 -2380 205 -2307
rect 85 -2414 128 -2380
rect 162 -2414 205 -2380
rect 85 -2460 205 -2414
rect 85 -2494 128 -2460
rect 162 -2494 205 -2460
rect 85 -2540 205 -2494
rect 85 -2574 128 -2540
rect 162 -2574 205 -2540
rect 85 -2607 205 -2574
rect 235 -2380 355 -2307
rect 235 -2414 278 -2380
rect 312 -2414 355 -2380
rect 235 -2460 355 -2414
rect 235 -2494 278 -2460
rect 312 -2494 355 -2460
rect 235 -2540 355 -2494
rect 235 -2574 278 -2540
rect 312 -2574 355 -2540
rect 235 -2607 355 -2574
rect 385 -2380 505 -2307
rect 385 -2414 428 -2380
rect 462 -2414 505 -2380
rect 385 -2460 505 -2414
rect 385 -2494 428 -2460
rect 462 -2494 505 -2460
rect 385 -2540 505 -2494
rect 385 -2574 428 -2540
rect 462 -2574 505 -2540
rect 385 -2607 505 -2574
rect 535 -2380 655 -2307
rect 535 -2414 578 -2380
rect 612 -2414 655 -2380
rect 535 -2460 655 -2414
rect 535 -2494 578 -2460
rect 612 -2494 655 -2460
rect 535 -2540 655 -2494
rect 535 -2574 578 -2540
rect 612 -2574 655 -2540
rect 535 -2607 655 -2574
rect 715 -2380 835 -2307
rect 715 -2414 758 -2380
rect 792 -2414 835 -2380
rect 715 -2460 835 -2414
rect 715 -2494 758 -2460
rect 792 -2494 835 -2460
rect 715 -2540 835 -2494
rect 715 -2574 758 -2540
rect 792 -2574 835 -2540
rect 715 -2607 835 -2574
rect 865 -2380 985 -2307
rect 865 -2414 908 -2380
rect 942 -2414 985 -2380
rect 865 -2460 985 -2414
rect 865 -2494 908 -2460
rect 942 -2494 985 -2460
rect 865 -2540 985 -2494
rect 865 -2574 908 -2540
rect 942 -2574 985 -2540
rect 865 -2607 985 -2574
rect 1015 -2380 1135 -2307
rect 1015 -2414 1058 -2380
rect 1092 -2414 1135 -2380
rect 1015 -2460 1135 -2414
rect 1015 -2494 1058 -2460
rect 1092 -2494 1135 -2460
rect 1015 -2540 1135 -2494
rect 1015 -2574 1058 -2540
rect 1092 -2574 1135 -2540
rect 1015 -2607 1135 -2574
rect 1165 -2380 1285 -2307
rect 1165 -2414 1208 -2380
rect 1242 -2414 1285 -2380
rect 1165 -2460 1285 -2414
rect 1165 -2494 1208 -2460
rect 1242 -2494 1285 -2460
rect 1165 -2540 1285 -2494
rect 1165 -2574 1208 -2540
rect 1242 -2574 1285 -2540
rect 1165 -2607 1285 -2574
rect 1315 -2380 1435 -2307
rect 1315 -2414 1358 -2380
rect 1392 -2414 1435 -2380
rect 1315 -2460 1435 -2414
rect 1315 -2494 1358 -2460
rect 1392 -2494 1435 -2460
rect 1315 -2540 1435 -2494
rect 1315 -2574 1358 -2540
rect 1392 -2574 1435 -2540
rect 1315 -2607 1435 -2574
rect 1495 -2380 1615 -2307
rect 1495 -2414 1538 -2380
rect 1572 -2414 1615 -2380
rect 1495 -2460 1615 -2414
rect 1495 -2494 1538 -2460
rect 1572 -2494 1615 -2460
rect 1495 -2540 1615 -2494
rect 1495 -2574 1538 -2540
rect 1572 -2574 1615 -2540
rect 1495 -2607 1615 -2574
rect 1645 -2607 1765 -2307
rect 1795 -2607 1915 -2307
rect 1945 -2607 2065 -2307
rect 2095 -2380 2215 -2307
rect 2095 -2414 2138 -2380
rect 2172 -2414 2215 -2380
rect 2095 -2460 2215 -2414
rect 2095 -2494 2138 -2460
rect 2172 -2494 2215 -2460
rect 2095 -2540 2215 -2494
rect 2095 -2574 2138 -2540
rect 2172 -2574 2215 -2540
rect 2095 -2607 2215 -2574
rect 2596 -2379 2716 -2306
rect 2596 -2413 2639 -2379
rect 2673 -2413 2716 -2379
rect 2596 -2459 2716 -2413
rect 2596 -2493 2639 -2459
rect 2673 -2493 2716 -2459
rect 2596 -2539 2716 -2493
rect 2596 -2573 2639 -2539
rect 2673 -2573 2716 -2539
rect 2596 -2606 2716 -2573
rect 2746 -2379 2866 -2306
rect 2746 -2413 2789 -2379
rect 2823 -2413 2866 -2379
rect 2746 -2459 2866 -2413
rect 2746 -2493 2789 -2459
rect 2823 -2493 2866 -2459
rect 2746 -2539 2866 -2493
rect 2746 -2573 2789 -2539
rect 2823 -2573 2866 -2539
rect 2746 -2606 2866 -2573
rect 2926 -2379 3046 -2306
rect 2926 -2413 2969 -2379
rect 3003 -2413 3046 -2379
rect 2926 -2459 3046 -2413
rect 2926 -2493 2969 -2459
rect 3003 -2493 3046 -2459
rect 2926 -2539 3046 -2493
rect 2926 -2573 2969 -2539
rect 3003 -2573 3046 -2539
rect 2926 -2606 3046 -2573
rect 3076 -2379 3196 -2306
rect 3076 -2413 3119 -2379
rect 3153 -2413 3196 -2379
rect 3076 -2459 3196 -2413
rect 3076 -2493 3119 -2459
rect 3153 -2493 3196 -2459
rect 3076 -2539 3196 -2493
rect 3076 -2573 3119 -2539
rect 3153 -2573 3196 -2539
rect 3076 -2606 3196 -2573
rect 3226 -2379 3346 -2306
rect 3226 -2413 3269 -2379
rect 3303 -2413 3346 -2379
rect 3226 -2459 3346 -2413
rect 3226 -2493 3269 -2459
rect 3303 -2493 3346 -2459
rect 3226 -2539 3346 -2493
rect 3226 -2573 3269 -2539
rect 3303 -2573 3346 -2539
rect 3226 -2606 3346 -2573
rect 3376 -2379 3496 -2306
rect 3376 -2413 3419 -2379
rect 3453 -2413 3496 -2379
rect 3376 -2459 3496 -2413
rect 3376 -2493 3419 -2459
rect 3453 -2493 3496 -2459
rect 3376 -2539 3496 -2493
rect 3376 -2573 3419 -2539
rect 3453 -2573 3496 -2539
rect 3376 -2606 3496 -2573
rect 3526 -2379 3646 -2306
rect 3526 -2413 3569 -2379
rect 3603 -2413 3646 -2379
rect 3526 -2459 3646 -2413
rect 3526 -2493 3569 -2459
rect 3603 -2493 3646 -2459
rect 3526 -2539 3646 -2493
rect 3526 -2573 3569 -2539
rect 3603 -2573 3646 -2539
rect 3526 -2606 3646 -2573
rect 3706 -2379 3826 -2306
rect 3706 -2413 3749 -2379
rect 3783 -2413 3826 -2379
rect 3706 -2459 3826 -2413
rect 3706 -2493 3749 -2459
rect 3783 -2493 3826 -2459
rect 3706 -2539 3826 -2493
rect 3706 -2573 3749 -2539
rect 3783 -2573 3826 -2539
rect 3706 -2606 3826 -2573
rect 3856 -2379 3976 -2306
rect 3856 -2413 3899 -2379
rect 3933 -2413 3976 -2379
rect 3856 -2459 3976 -2413
rect 3856 -2493 3899 -2459
rect 3933 -2493 3976 -2459
rect 3856 -2539 3976 -2493
rect 3856 -2573 3899 -2539
rect 3933 -2573 3976 -2539
rect 3856 -2606 3976 -2573
rect 4355 -2379 4475 -2306
rect 4355 -2413 4398 -2379
rect 4432 -2413 4475 -2379
rect 4355 -2459 4475 -2413
rect 4355 -2493 4398 -2459
rect 4432 -2493 4475 -2459
rect 4355 -2539 4475 -2493
rect 4355 -2573 4398 -2539
rect 4432 -2573 4475 -2539
rect 4355 -2606 4475 -2573
rect 4505 -2379 4625 -2306
rect 4505 -2413 4548 -2379
rect 4582 -2413 4625 -2379
rect 4505 -2459 4625 -2413
rect 4505 -2493 4548 -2459
rect 4582 -2493 4625 -2459
rect 4505 -2539 4625 -2493
rect 4505 -2573 4548 -2539
rect 4582 -2573 4625 -2539
rect 4505 -2606 4625 -2573
rect 4655 -2379 4775 -2306
rect 4655 -2413 4698 -2379
rect 4732 -2413 4775 -2379
rect 4655 -2459 4775 -2413
rect 4655 -2493 4698 -2459
rect 4732 -2493 4775 -2459
rect 4655 -2539 4775 -2493
rect 4655 -2573 4698 -2539
rect 4732 -2573 4775 -2539
rect 4655 -2606 4775 -2573
rect 4805 -2379 4925 -2306
rect 4805 -2413 4848 -2379
rect 4882 -2413 4925 -2379
rect 4805 -2459 4925 -2413
rect 4805 -2493 4848 -2459
rect 4882 -2493 4925 -2459
rect 4805 -2539 4925 -2493
rect 4805 -2573 4848 -2539
rect 4882 -2573 4925 -2539
rect 4805 -2606 4925 -2573
rect 4985 -2379 5105 -2306
rect 4985 -2413 5028 -2379
rect 5062 -2413 5105 -2379
rect 4985 -2459 5105 -2413
rect 4985 -2493 5028 -2459
rect 5062 -2493 5105 -2459
rect 4985 -2539 5105 -2493
rect 4985 -2573 5028 -2539
rect 5062 -2573 5105 -2539
rect 4985 -2606 5105 -2573
rect 5135 -2379 5255 -2306
rect 5135 -2413 5178 -2379
rect 5212 -2413 5255 -2379
rect 5135 -2459 5255 -2413
rect 5135 -2493 5178 -2459
rect 5212 -2493 5255 -2459
rect 5135 -2539 5255 -2493
rect 5135 -2573 5178 -2539
rect 5212 -2573 5255 -2539
rect 5135 -2606 5255 -2573
rect 5285 -2379 5405 -2306
rect 5285 -2413 5328 -2379
rect 5362 -2413 5405 -2379
rect 5285 -2459 5405 -2413
rect 5285 -2493 5328 -2459
rect 5362 -2493 5405 -2459
rect 5285 -2539 5405 -2493
rect 5285 -2573 5328 -2539
rect 5362 -2573 5405 -2539
rect 5285 -2606 5405 -2573
rect 5435 -2379 5555 -2306
rect 5435 -2413 5478 -2379
rect 5512 -2413 5555 -2379
rect 5435 -2459 5555 -2413
rect 5435 -2493 5478 -2459
rect 5512 -2493 5555 -2459
rect 5435 -2539 5555 -2493
rect 5435 -2573 5478 -2539
rect 5512 -2573 5555 -2539
rect 5435 -2606 5555 -2573
rect 5585 -2379 5705 -2306
rect 5585 -2413 5628 -2379
rect 5662 -2413 5705 -2379
rect 5585 -2459 5705 -2413
rect 5585 -2493 5628 -2459
rect 5662 -2493 5705 -2459
rect 5585 -2539 5705 -2493
rect 5585 -2573 5628 -2539
rect 5662 -2573 5705 -2539
rect 5585 -2606 5705 -2573
rect 5765 -2379 5885 -2306
rect 5765 -2413 5808 -2379
rect 5842 -2413 5885 -2379
rect 5765 -2459 5885 -2413
rect 5765 -2493 5808 -2459
rect 5842 -2493 5885 -2459
rect 5765 -2539 5885 -2493
rect 5765 -2573 5808 -2539
rect 5842 -2573 5885 -2539
rect 5765 -2606 5885 -2573
rect 5915 -2606 6035 -2306
rect 6065 -2606 6185 -2306
rect 6215 -2379 6335 -2306
rect 6215 -2413 6258 -2379
rect 6292 -2413 6335 -2379
rect 6215 -2459 6335 -2413
rect 6215 -2493 6258 -2459
rect 6292 -2493 6335 -2459
rect 6215 -2539 6335 -2493
rect 6215 -2573 6258 -2539
rect 6292 -2573 6335 -2539
rect 6215 -2606 6335 -2573
<< pdiff >>
rect 715 1001 835 1074
rect 715 967 758 1001
rect 792 967 835 1001
rect 715 921 835 967
rect 715 887 758 921
rect 792 887 835 921
rect 715 841 835 887
rect 715 807 758 841
rect 792 807 835 841
rect 715 774 835 807
rect 865 1001 985 1074
rect 865 967 908 1001
rect 942 967 985 1001
rect 865 921 985 967
rect 865 887 908 921
rect 942 887 985 921
rect 865 841 985 887
rect 865 807 908 841
rect 942 807 985 841
rect 865 774 985 807
rect 1015 1001 1135 1074
rect 1015 967 1058 1001
rect 1092 967 1135 1001
rect 1015 921 1135 967
rect 1015 887 1058 921
rect 1092 887 1135 921
rect 1015 841 1135 887
rect 1015 807 1058 841
rect 1092 807 1135 841
rect 1015 774 1135 807
rect 1165 1001 1285 1074
rect 1165 967 1208 1001
rect 1242 967 1285 1001
rect 1165 921 1285 967
rect 1165 887 1208 921
rect 1242 887 1285 921
rect 1165 841 1285 887
rect 1165 807 1208 841
rect 1242 807 1285 841
rect 1165 774 1285 807
rect 1315 1001 1435 1074
rect 1315 967 1358 1001
rect 1392 967 1435 1001
rect 1315 921 1435 967
rect 1315 887 1358 921
rect 1392 887 1435 921
rect 1315 841 1435 887
rect 1315 807 1358 841
rect 1392 807 1435 841
rect 1315 774 1435 807
rect 2925 1001 3045 1074
rect 2925 967 2968 1001
rect 3002 967 3045 1001
rect 2925 921 3045 967
rect 2925 887 2968 921
rect 3002 887 3045 921
rect 2925 841 3045 887
rect 2925 807 2968 841
rect 3002 807 3045 841
rect 2925 774 3045 807
rect 3075 1001 3195 1074
rect 3075 967 3118 1001
rect 3152 967 3195 1001
rect 3075 921 3195 967
rect 3075 887 3118 921
rect 3152 887 3195 921
rect 3075 841 3195 887
rect 3075 807 3118 841
rect 3152 807 3195 841
rect 3075 774 3195 807
rect 3225 1001 3345 1074
rect 3225 967 3268 1001
rect 3302 967 3345 1001
rect 3225 921 3345 967
rect 3225 887 3268 921
rect 3302 887 3345 921
rect 3225 841 3345 887
rect 3225 807 3268 841
rect 3302 807 3345 841
rect 3225 774 3345 807
rect 3375 1001 3495 1074
rect 3375 967 3418 1001
rect 3452 967 3495 1001
rect 3375 921 3495 967
rect 3375 887 3418 921
rect 3452 887 3495 921
rect 3375 841 3495 887
rect 3375 807 3418 841
rect 3452 807 3495 841
rect 3375 774 3495 807
rect 3525 1001 3645 1074
rect 3525 967 3568 1001
rect 3602 967 3645 1001
rect 3525 921 3645 967
rect 3525 887 3568 921
rect 3602 887 3645 921
rect 3525 841 3645 887
rect 4805 1001 4925 1074
rect 4805 967 4848 1001
rect 4882 967 4925 1001
rect 4805 921 4925 967
rect 4805 887 4848 921
rect 4882 887 4925 921
rect 3525 807 3568 841
rect 3602 807 3645 841
rect 3525 774 3645 807
rect 4805 841 4925 887
rect 4805 807 4848 841
rect 4882 807 4925 841
rect 4805 774 4925 807
rect 4955 1001 5075 1074
rect 4955 967 4998 1001
rect 5032 967 5075 1001
rect 4955 921 5075 967
rect 4955 887 4998 921
rect 5032 887 5075 921
rect 4955 841 5075 887
rect 4955 807 4998 841
rect 5032 807 5075 841
rect 4955 774 5075 807
rect 5105 1001 5225 1074
rect 5105 967 5148 1001
rect 5182 967 5225 1001
rect 5105 921 5225 967
rect 5105 887 5148 921
rect 5182 887 5225 921
rect 5105 841 5225 887
rect 5105 807 5148 841
rect 5182 807 5225 841
rect 5105 774 5225 807
rect 5255 1001 5375 1074
rect 5255 967 5298 1001
rect 5332 967 5375 1001
rect 5255 921 5375 967
rect 5255 887 5298 921
rect 5332 887 5375 921
rect 5255 841 5375 887
rect 5255 807 5298 841
rect 5332 807 5375 841
rect 5255 774 5375 807
rect 5405 1001 5525 1074
rect 5405 967 5448 1001
rect 5482 967 5525 1001
rect 5405 921 5525 967
rect 5405 887 5448 921
rect 5482 887 5525 921
rect 5405 841 5525 887
rect 5405 807 5448 841
rect 5482 807 5525 841
rect 5405 774 5525 807
rect 715 -759 835 -726
rect 715 -793 758 -759
rect 792 -793 835 -759
rect 715 -839 835 -793
rect 715 -873 758 -839
rect 792 -873 835 -839
rect 715 -919 835 -873
rect 715 -953 758 -919
rect 792 -953 835 -919
rect 715 -1026 835 -953
rect 865 -759 985 -726
rect 865 -793 908 -759
rect 942 -793 985 -759
rect 865 -839 985 -793
rect 865 -873 908 -839
rect 942 -873 985 -839
rect 865 -919 985 -873
rect 865 -953 908 -919
rect 942 -953 985 -919
rect 865 -1026 985 -953
rect 1015 -759 1135 -726
rect 1015 -793 1058 -759
rect 1092 -793 1135 -759
rect 1015 -839 1135 -793
rect 1015 -873 1058 -839
rect 1092 -873 1135 -839
rect 1015 -919 1135 -873
rect 1015 -953 1058 -919
rect 1092 -953 1135 -919
rect 1015 -1026 1135 -953
rect 1165 -759 1285 -726
rect 1165 -793 1208 -759
rect 1242 -793 1285 -759
rect 1165 -839 1285 -793
rect 1165 -873 1208 -839
rect 1242 -873 1285 -839
rect 1165 -919 1285 -873
rect 1165 -953 1208 -919
rect 1242 -953 1285 -919
rect 1165 -1026 1285 -953
rect 1315 -759 1435 -726
rect 1315 -793 1358 -759
rect 1392 -793 1435 -759
rect 1315 -839 1435 -793
rect 1315 -873 1358 -839
rect 1392 -873 1435 -839
rect 1315 -919 1435 -873
rect 1315 -953 1358 -919
rect 1392 -953 1435 -919
rect 1315 -1026 1435 -953
rect 2925 -759 3045 -726
rect 2925 -793 2968 -759
rect 3002 -793 3045 -759
rect 2925 -839 3045 -793
rect 2925 -873 2968 -839
rect 3002 -873 3045 -839
rect 2925 -919 3045 -873
rect 2925 -953 2968 -919
rect 3002 -953 3045 -919
rect 2925 -1026 3045 -953
rect 3075 -759 3195 -726
rect 3075 -793 3118 -759
rect 3152 -793 3195 -759
rect 3075 -839 3195 -793
rect 3075 -873 3118 -839
rect 3152 -873 3195 -839
rect 3075 -919 3195 -873
rect 3075 -953 3118 -919
rect 3152 -953 3195 -919
rect 3075 -1026 3195 -953
rect 3225 -759 3345 -726
rect 3225 -793 3268 -759
rect 3302 -793 3345 -759
rect 3225 -839 3345 -793
rect 3225 -873 3268 -839
rect 3302 -873 3345 -839
rect 3225 -919 3345 -873
rect 3225 -953 3268 -919
rect 3302 -953 3345 -919
rect 3225 -1026 3345 -953
rect 3375 -759 3495 -726
rect 3375 -793 3418 -759
rect 3452 -793 3495 -759
rect 3375 -839 3495 -793
rect 3375 -873 3418 -839
rect 3452 -873 3495 -839
rect 3375 -919 3495 -873
rect 3375 -953 3418 -919
rect 3452 -953 3495 -919
rect 3375 -1026 3495 -953
rect 3525 -759 3645 -726
rect 3525 -793 3568 -759
rect 3602 -793 3645 -759
rect 3525 -839 3645 -793
rect 4805 -759 4925 -726
rect 4805 -793 4848 -759
rect 4882 -793 4925 -759
rect 3525 -873 3568 -839
rect 3602 -873 3645 -839
rect 3525 -919 3645 -873
rect 3525 -953 3568 -919
rect 3602 -953 3645 -919
rect 3525 -1026 3645 -953
rect 4805 -839 4925 -793
rect 4805 -873 4848 -839
rect 4882 -873 4925 -839
rect 4805 -919 4925 -873
rect 4805 -953 4848 -919
rect 4882 -953 4925 -919
rect 4805 -1026 4925 -953
rect 4955 -759 5075 -726
rect 4955 -793 4998 -759
rect 5032 -793 5075 -759
rect 4955 -839 5075 -793
rect 4955 -873 4998 -839
rect 5032 -873 5075 -839
rect 4955 -919 5075 -873
rect 4955 -953 4998 -919
rect 5032 -953 5075 -919
rect 4955 -1026 5075 -953
rect 5105 -759 5225 -726
rect 5105 -793 5148 -759
rect 5182 -793 5225 -759
rect 5105 -839 5225 -793
rect 5105 -873 5148 -839
rect 5182 -873 5225 -839
rect 5105 -919 5225 -873
rect 5105 -953 5148 -919
rect 5182 -953 5225 -919
rect 5105 -1026 5225 -953
rect 5255 -759 5375 -726
rect 5255 -793 5298 -759
rect 5332 -793 5375 -759
rect 5255 -839 5375 -793
rect 5255 -873 5298 -839
rect 5332 -873 5375 -839
rect 5255 -919 5375 -873
rect 5255 -953 5298 -919
rect 5332 -953 5375 -919
rect 5255 -1026 5375 -953
rect 5405 -759 5525 -726
rect 5405 -793 5448 -759
rect 5482 -793 5525 -759
rect 5405 -839 5525 -793
rect 5405 -873 5448 -839
rect 5482 -873 5525 -839
rect 5405 -919 5525 -873
rect 5405 -953 5448 -919
rect 5482 -953 5525 -919
rect 5405 -1026 5525 -953
rect 715 -1500 835 -1427
rect 715 -1534 758 -1500
rect 792 -1534 835 -1500
rect 715 -1580 835 -1534
rect 715 -1614 758 -1580
rect 792 -1614 835 -1580
rect 715 -1660 835 -1614
rect 715 -1694 758 -1660
rect 792 -1694 835 -1660
rect 715 -1727 835 -1694
rect 865 -1500 985 -1427
rect 865 -1534 908 -1500
rect 942 -1534 985 -1500
rect 865 -1580 985 -1534
rect 865 -1614 908 -1580
rect 942 -1614 985 -1580
rect 865 -1660 985 -1614
rect 865 -1694 908 -1660
rect 942 -1694 985 -1660
rect 865 -1727 985 -1694
rect 1015 -1500 1135 -1427
rect 1015 -1534 1058 -1500
rect 1092 -1534 1135 -1500
rect 1015 -1580 1135 -1534
rect 1015 -1614 1058 -1580
rect 1092 -1614 1135 -1580
rect 1015 -1660 1135 -1614
rect 1015 -1694 1058 -1660
rect 1092 -1694 1135 -1660
rect 1015 -1727 1135 -1694
rect 1165 -1500 1285 -1427
rect 1165 -1534 1208 -1500
rect 1242 -1534 1285 -1500
rect 1165 -1580 1285 -1534
rect 1165 -1614 1208 -1580
rect 1242 -1614 1285 -1580
rect 1165 -1660 1285 -1614
rect 1165 -1694 1208 -1660
rect 1242 -1694 1285 -1660
rect 1165 -1727 1285 -1694
rect 1315 -1500 1435 -1427
rect 1315 -1534 1358 -1500
rect 1392 -1534 1435 -1500
rect 1315 -1580 1435 -1534
rect 1315 -1614 1358 -1580
rect 1392 -1614 1435 -1580
rect 1315 -1660 1435 -1614
rect 1315 -1694 1358 -1660
rect 1392 -1694 1435 -1660
rect 1315 -1727 1435 -1694
rect 2926 -1819 3046 -1746
rect 2926 -1853 2969 -1819
rect 3003 -1853 3046 -1819
rect 2926 -1899 3046 -1853
rect 2926 -1933 2969 -1899
rect 3003 -1933 3046 -1899
rect 2926 -1979 3046 -1933
rect 2926 -2013 2969 -1979
rect 3003 -2013 3046 -1979
rect 2926 -2046 3046 -2013
rect 3076 -1819 3196 -1746
rect 3076 -1853 3119 -1819
rect 3153 -1853 3196 -1819
rect 3076 -1899 3196 -1853
rect 3076 -1933 3119 -1899
rect 3153 -1933 3196 -1899
rect 3076 -1979 3196 -1933
rect 3076 -2013 3119 -1979
rect 3153 -2013 3196 -1979
rect 3076 -2046 3196 -2013
rect 3226 -1819 3346 -1746
rect 3226 -1853 3269 -1819
rect 3303 -1853 3346 -1819
rect 3226 -1899 3346 -1853
rect 3226 -1933 3269 -1899
rect 3303 -1933 3346 -1899
rect 3226 -1979 3346 -1933
rect 3226 -2013 3269 -1979
rect 3303 -2013 3346 -1979
rect 3226 -2046 3346 -2013
rect 3376 -1819 3496 -1746
rect 3376 -1853 3419 -1819
rect 3453 -1853 3496 -1819
rect 3376 -1899 3496 -1853
rect 3376 -1933 3419 -1899
rect 3453 -1933 3496 -1899
rect 3376 -1979 3496 -1933
rect 3376 -2013 3419 -1979
rect 3453 -2013 3496 -1979
rect 3376 -2046 3496 -2013
rect 3526 -1819 3646 -1746
rect 3526 -1853 3569 -1819
rect 3603 -1853 3646 -1819
rect 3526 -1899 3646 -1853
rect 3526 -1933 3569 -1899
rect 3603 -1933 3646 -1899
rect 3526 -1979 3646 -1933
rect 3526 -2013 3569 -1979
rect 3603 -2013 3646 -1979
rect 3526 -2046 3646 -2013
rect 4985 -1819 5105 -1746
rect 4985 -1853 5028 -1819
rect 5062 -1853 5105 -1819
rect 4985 -1899 5105 -1853
rect 4985 -1933 5028 -1899
rect 5062 -1933 5105 -1899
rect 4985 -1979 5105 -1933
rect 4985 -2013 5028 -1979
rect 5062 -2013 5105 -1979
rect 4985 -2046 5105 -2013
rect 5135 -1819 5255 -1746
rect 5135 -1853 5178 -1819
rect 5212 -1853 5255 -1819
rect 5135 -1899 5255 -1853
rect 5135 -1933 5178 -1899
rect 5212 -1933 5255 -1899
rect 5135 -1979 5255 -1933
rect 5135 -2013 5178 -1979
rect 5212 -2013 5255 -1979
rect 5135 -2046 5255 -2013
rect 5285 -1819 5405 -1746
rect 5285 -1853 5328 -1819
rect 5362 -1853 5405 -1819
rect 5285 -1899 5405 -1853
rect 5285 -1933 5328 -1899
rect 5362 -1933 5405 -1899
rect 5285 -1979 5405 -1933
rect 5285 -2013 5328 -1979
rect 5362 -2013 5405 -1979
rect 5285 -2046 5405 -2013
rect 5435 -1819 5555 -1746
rect 5435 -1853 5478 -1819
rect 5512 -1853 5555 -1819
rect 5435 -1899 5555 -1853
rect 5435 -1933 5478 -1899
rect 5512 -1933 5555 -1899
rect 5435 -1979 5555 -1933
rect 5435 -2013 5478 -1979
rect 5512 -2013 5555 -1979
rect 5435 -2046 5555 -2013
rect 5585 -1819 5705 -1746
rect 5585 -1853 5628 -1819
rect 5662 -1853 5705 -1819
rect 5585 -1899 5705 -1853
rect 5585 -1933 5628 -1899
rect 5662 -1933 5705 -1899
rect 5585 -1979 5705 -1933
rect 5585 -2013 5628 -1979
rect 5662 -2013 5705 -1979
rect 5585 -2046 5705 -2013
<< ndiffc >>
rect -22 407 12 441
rect -22 327 12 361
rect -22 247 12 281
rect 278 407 312 441
rect 278 327 312 361
rect 278 247 312 281
rect 578 407 612 441
rect 578 327 612 361
rect 578 247 612 281
rect 758 407 792 441
rect 758 327 792 361
rect 758 247 792 281
rect 908 407 942 441
rect 908 327 942 361
rect 908 247 942 281
rect 1058 407 1092 441
rect 1058 327 1092 361
rect 1058 247 1092 281
rect 1208 407 1242 441
rect 1208 327 1242 361
rect 1208 247 1242 281
rect 1358 407 1392 441
rect 1358 327 1392 361
rect 1358 247 1392 281
rect 1538 407 1572 441
rect 1538 327 1572 361
rect 1538 247 1572 281
rect 1838 407 1872 441
rect 1838 327 1872 361
rect 1838 247 1872 281
rect 2138 407 2172 441
rect 2138 327 2172 361
rect 2138 247 2172 281
rect 2638 407 2672 441
rect 2638 327 2672 361
rect 2638 247 2672 281
rect 2788 407 2822 441
rect 2788 327 2822 361
rect 2788 247 2822 281
rect 2968 407 3002 441
rect 2968 327 3002 361
rect 2968 247 3002 281
rect 3118 407 3152 441
rect 3118 327 3152 361
rect 3118 247 3152 281
rect 3268 407 3302 441
rect 3268 327 3302 361
rect 3268 247 3302 281
rect 3418 407 3452 441
rect 3418 327 3452 361
rect 3418 247 3452 281
rect 3568 407 3602 441
rect 3568 327 3602 361
rect 3568 247 3602 281
rect 3748 407 3782 441
rect 3748 327 3782 361
rect 3748 247 3782 281
rect 3898 407 3932 441
rect 3898 327 3932 361
rect 3898 247 3932 281
rect 4368 407 4402 441
rect 4368 327 4402 361
rect 4368 247 4402 281
rect 4518 407 4552 441
rect 4518 327 4552 361
rect 4518 247 4552 281
rect 4668 407 4702 441
rect 4668 327 4702 361
rect 4668 247 4702 281
rect 4848 407 4882 441
rect 4848 327 4882 361
rect 4848 247 4882 281
rect 4998 407 5032 441
rect 4998 327 5032 361
rect 4998 247 5032 281
rect 5148 407 5182 441
rect 5148 327 5182 361
rect 5148 247 5182 281
rect 5298 407 5332 441
rect 5298 327 5332 361
rect 5298 247 5332 281
rect 5448 407 5482 441
rect 5448 327 5482 361
rect 5448 247 5482 281
rect 5628 407 5662 441
rect 5628 327 5662 361
rect 5628 247 5662 281
rect 5928 407 5962 441
rect 5928 327 5962 361
rect 5928 247 5962 281
rect -22 -233 12 -199
rect -22 -313 12 -279
rect -22 -393 12 -359
rect 278 -233 312 -199
rect 278 -313 312 -279
rect 278 -393 312 -359
rect 578 -233 612 -199
rect 578 -313 612 -279
rect 578 -393 612 -359
rect 758 -233 792 -199
rect 758 -313 792 -279
rect 758 -393 792 -359
rect 908 -233 942 -199
rect 908 -313 942 -279
rect 908 -393 942 -359
rect 1058 -233 1092 -199
rect 1058 -313 1092 -279
rect 1058 -393 1092 -359
rect 1208 -233 1242 -199
rect 1208 -313 1242 -279
rect 1208 -393 1242 -359
rect 1358 -233 1392 -199
rect 1358 -313 1392 -279
rect 1358 -393 1392 -359
rect 1538 -233 1572 -199
rect 1538 -313 1572 -279
rect 1538 -393 1572 -359
rect 1838 -233 1872 -199
rect 1838 -313 1872 -279
rect 1838 -393 1872 -359
rect 2138 -233 2172 -199
rect 2138 -313 2172 -279
rect 2138 -393 2172 -359
rect 2638 -233 2672 -199
rect 2638 -313 2672 -279
rect 2638 -393 2672 -359
rect 2788 -233 2822 -199
rect 2788 -313 2822 -279
rect 2788 -393 2822 -359
rect 2968 -233 3002 -199
rect 2968 -313 3002 -279
rect 2968 -393 3002 -359
rect 3118 -233 3152 -199
rect 3118 -313 3152 -279
rect 3118 -393 3152 -359
rect 3268 -233 3302 -199
rect 3268 -313 3302 -279
rect 3268 -393 3302 -359
rect 3418 -233 3452 -199
rect 3418 -313 3452 -279
rect 3418 -393 3452 -359
rect 3568 -233 3602 -199
rect 3568 -313 3602 -279
rect 3568 -393 3602 -359
rect 3748 -233 3782 -199
rect 3748 -313 3782 -279
rect 3748 -393 3782 -359
rect 3898 -233 3932 -199
rect 3898 -313 3932 -279
rect 3898 -393 3932 -359
rect 4368 -233 4402 -199
rect 4368 -313 4402 -279
rect 4368 -393 4402 -359
rect 4518 -233 4552 -199
rect 4518 -313 4552 -279
rect 4518 -393 4552 -359
rect 4668 -233 4702 -199
rect 4668 -313 4702 -279
rect 4668 -393 4702 -359
rect 4848 -233 4882 -199
rect 4848 -313 4882 -279
rect 4848 -393 4882 -359
rect 4998 -233 5032 -199
rect 4998 -313 5032 -279
rect 4998 -393 5032 -359
rect 5148 -233 5182 -199
rect 5148 -313 5182 -279
rect 5148 -393 5182 -359
rect 5298 -233 5332 -199
rect 5298 -313 5332 -279
rect 5298 -393 5332 -359
rect 5448 -233 5482 -199
rect 5448 -313 5482 -279
rect 5448 -393 5482 -359
rect 5628 -233 5662 -199
rect 5628 -313 5662 -279
rect 5628 -393 5662 -359
rect 5928 -233 5962 -199
rect 5928 -313 5962 -279
rect 5928 -393 5962 -359
rect -22 -2414 12 -2380
rect -22 -2494 12 -2460
rect -22 -2574 12 -2540
rect 128 -2414 162 -2380
rect 128 -2494 162 -2460
rect 128 -2574 162 -2540
rect 278 -2414 312 -2380
rect 278 -2494 312 -2460
rect 278 -2574 312 -2540
rect 428 -2414 462 -2380
rect 428 -2494 462 -2460
rect 428 -2574 462 -2540
rect 578 -2414 612 -2380
rect 578 -2494 612 -2460
rect 578 -2574 612 -2540
rect 758 -2414 792 -2380
rect 758 -2494 792 -2460
rect 758 -2574 792 -2540
rect 908 -2414 942 -2380
rect 908 -2494 942 -2460
rect 908 -2574 942 -2540
rect 1058 -2414 1092 -2380
rect 1058 -2494 1092 -2460
rect 1058 -2574 1092 -2540
rect 1208 -2414 1242 -2380
rect 1208 -2494 1242 -2460
rect 1208 -2574 1242 -2540
rect 1358 -2414 1392 -2380
rect 1358 -2494 1392 -2460
rect 1358 -2574 1392 -2540
rect 1538 -2414 1572 -2380
rect 1538 -2494 1572 -2460
rect 1538 -2574 1572 -2540
rect 2138 -2414 2172 -2380
rect 2138 -2494 2172 -2460
rect 2138 -2574 2172 -2540
rect 2639 -2413 2673 -2379
rect 2639 -2493 2673 -2459
rect 2639 -2573 2673 -2539
rect 2789 -2413 2823 -2379
rect 2789 -2493 2823 -2459
rect 2789 -2573 2823 -2539
rect 2969 -2413 3003 -2379
rect 2969 -2493 3003 -2459
rect 2969 -2573 3003 -2539
rect 3119 -2413 3153 -2379
rect 3119 -2493 3153 -2459
rect 3119 -2573 3153 -2539
rect 3269 -2413 3303 -2379
rect 3269 -2493 3303 -2459
rect 3269 -2573 3303 -2539
rect 3419 -2413 3453 -2379
rect 3419 -2493 3453 -2459
rect 3419 -2573 3453 -2539
rect 3569 -2413 3603 -2379
rect 3569 -2493 3603 -2459
rect 3569 -2573 3603 -2539
rect 3749 -2413 3783 -2379
rect 3749 -2493 3783 -2459
rect 3749 -2573 3783 -2539
rect 3899 -2413 3933 -2379
rect 3899 -2493 3933 -2459
rect 3899 -2573 3933 -2539
rect 4398 -2413 4432 -2379
rect 4398 -2493 4432 -2459
rect 4398 -2573 4432 -2539
rect 4548 -2413 4582 -2379
rect 4548 -2493 4582 -2459
rect 4548 -2573 4582 -2539
rect 4698 -2413 4732 -2379
rect 4698 -2493 4732 -2459
rect 4698 -2573 4732 -2539
rect 4848 -2413 4882 -2379
rect 4848 -2493 4882 -2459
rect 4848 -2573 4882 -2539
rect 5028 -2413 5062 -2379
rect 5028 -2493 5062 -2459
rect 5028 -2573 5062 -2539
rect 5178 -2413 5212 -2379
rect 5178 -2493 5212 -2459
rect 5178 -2573 5212 -2539
rect 5328 -2413 5362 -2379
rect 5328 -2493 5362 -2459
rect 5328 -2573 5362 -2539
rect 5478 -2413 5512 -2379
rect 5478 -2493 5512 -2459
rect 5478 -2573 5512 -2539
rect 5628 -2413 5662 -2379
rect 5628 -2493 5662 -2459
rect 5628 -2573 5662 -2539
rect 5808 -2413 5842 -2379
rect 5808 -2493 5842 -2459
rect 5808 -2573 5842 -2539
rect 6258 -2413 6292 -2379
rect 6258 -2493 6292 -2459
rect 6258 -2573 6292 -2539
<< pdiffc >>
rect 758 967 792 1001
rect 758 887 792 921
rect 758 807 792 841
rect 908 967 942 1001
rect 908 887 942 921
rect 908 807 942 841
rect 1058 967 1092 1001
rect 1058 887 1092 921
rect 1058 807 1092 841
rect 1208 967 1242 1001
rect 1208 887 1242 921
rect 1208 807 1242 841
rect 1358 967 1392 1001
rect 1358 887 1392 921
rect 1358 807 1392 841
rect 2968 967 3002 1001
rect 2968 887 3002 921
rect 2968 807 3002 841
rect 3118 967 3152 1001
rect 3118 887 3152 921
rect 3118 807 3152 841
rect 3268 967 3302 1001
rect 3268 887 3302 921
rect 3268 807 3302 841
rect 3418 967 3452 1001
rect 3418 887 3452 921
rect 3418 807 3452 841
rect 3568 967 3602 1001
rect 3568 887 3602 921
rect 4848 967 4882 1001
rect 4848 887 4882 921
rect 3568 807 3602 841
rect 4848 807 4882 841
rect 4998 967 5032 1001
rect 4998 887 5032 921
rect 4998 807 5032 841
rect 5148 967 5182 1001
rect 5148 887 5182 921
rect 5148 807 5182 841
rect 5298 967 5332 1001
rect 5298 887 5332 921
rect 5298 807 5332 841
rect 5448 967 5482 1001
rect 5448 887 5482 921
rect 5448 807 5482 841
rect 758 -793 792 -759
rect 758 -873 792 -839
rect 758 -953 792 -919
rect 908 -793 942 -759
rect 908 -873 942 -839
rect 908 -953 942 -919
rect 1058 -793 1092 -759
rect 1058 -873 1092 -839
rect 1058 -953 1092 -919
rect 1208 -793 1242 -759
rect 1208 -873 1242 -839
rect 1208 -953 1242 -919
rect 1358 -793 1392 -759
rect 1358 -873 1392 -839
rect 1358 -953 1392 -919
rect 2968 -793 3002 -759
rect 2968 -873 3002 -839
rect 2968 -953 3002 -919
rect 3118 -793 3152 -759
rect 3118 -873 3152 -839
rect 3118 -953 3152 -919
rect 3268 -793 3302 -759
rect 3268 -873 3302 -839
rect 3268 -953 3302 -919
rect 3418 -793 3452 -759
rect 3418 -873 3452 -839
rect 3418 -953 3452 -919
rect 3568 -793 3602 -759
rect 4848 -793 4882 -759
rect 3568 -873 3602 -839
rect 3568 -953 3602 -919
rect 4848 -873 4882 -839
rect 4848 -953 4882 -919
rect 4998 -793 5032 -759
rect 4998 -873 5032 -839
rect 4998 -953 5032 -919
rect 5148 -793 5182 -759
rect 5148 -873 5182 -839
rect 5148 -953 5182 -919
rect 5298 -793 5332 -759
rect 5298 -873 5332 -839
rect 5298 -953 5332 -919
rect 5448 -793 5482 -759
rect 5448 -873 5482 -839
rect 5448 -953 5482 -919
rect 758 -1534 792 -1500
rect 758 -1614 792 -1580
rect 758 -1694 792 -1660
rect 908 -1534 942 -1500
rect 908 -1614 942 -1580
rect 908 -1694 942 -1660
rect 1058 -1534 1092 -1500
rect 1058 -1614 1092 -1580
rect 1058 -1694 1092 -1660
rect 1208 -1534 1242 -1500
rect 1208 -1614 1242 -1580
rect 1208 -1694 1242 -1660
rect 1358 -1534 1392 -1500
rect 1358 -1614 1392 -1580
rect 1358 -1694 1392 -1660
rect 2969 -1853 3003 -1819
rect 2969 -1933 3003 -1899
rect 2969 -2013 3003 -1979
rect 3119 -1853 3153 -1819
rect 3119 -1933 3153 -1899
rect 3119 -2013 3153 -1979
rect 3269 -1853 3303 -1819
rect 3269 -1933 3303 -1899
rect 3269 -2013 3303 -1979
rect 3419 -1853 3453 -1819
rect 3419 -1933 3453 -1899
rect 3419 -2013 3453 -1979
rect 3569 -1853 3603 -1819
rect 3569 -1933 3603 -1899
rect 3569 -2013 3603 -1979
rect 5028 -1853 5062 -1819
rect 5028 -1933 5062 -1899
rect 5028 -2013 5062 -1979
rect 5178 -1853 5212 -1819
rect 5178 -1933 5212 -1899
rect 5178 -2013 5212 -1979
rect 5328 -1853 5362 -1819
rect 5328 -1933 5362 -1899
rect 5328 -2013 5362 -1979
rect 5478 -1853 5512 -1819
rect 5478 -1933 5512 -1899
rect 5478 -2013 5512 -1979
rect 5628 -1853 5662 -1819
rect 5628 -1933 5662 -1899
rect 5628 -2013 5662 -1979
<< psubdiff >>
rect -65 41 2215 74
rect -65 7 18 41
rect 52 7 98 41
rect 132 7 178 41
rect 212 7 258 41
rect 292 7 338 41
rect 372 7 418 41
rect 452 7 498 41
rect 532 7 578 41
rect 612 7 658 41
rect 692 7 738 41
rect 772 7 818 41
rect 852 7 898 41
rect 932 7 978 41
rect 1012 7 1058 41
rect 1092 7 1138 41
rect 1172 7 1218 41
rect 1252 7 1298 41
rect 1332 7 1378 41
rect 1412 7 1458 41
rect 1492 7 1538 41
rect 1572 7 1618 41
rect 1652 7 1698 41
rect 1732 7 1778 41
rect 1812 7 1858 41
rect 1892 7 1938 41
rect 1972 7 2018 41
rect 2052 7 2098 41
rect 2132 7 2215 41
rect -65 -26 2215 7
rect 2595 41 3975 74
rect 2595 7 2628 41
rect 2662 7 2708 41
rect 2742 7 2788 41
rect 2822 7 2868 41
rect 2902 7 2948 41
rect 2982 7 3028 41
rect 3062 7 3108 41
rect 3142 7 3188 41
rect 3222 7 3268 41
rect 3302 7 3348 41
rect 3382 7 3428 41
rect 3462 7 3508 41
rect 3542 7 3588 41
rect 3622 7 3668 41
rect 3702 7 3748 41
rect 3782 7 3828 41
rect 3862 7 3908 41
rect 3942 7 3975 41
rect 2595 -26 3975 7
rect 4325 41 6005 74
rect 4325 7 4348 41
rect 4382 7 4428 41
rect 4462 7 4508 41
rect 4542 7 4588 41
rect 4622 7 4668 41
rect 4702 7 4748 41
rect 4782 7 4828 41
rect 4862 7 4908 41
rect 4942 7 4988 41
rect 5022 7 5068 41
rect 5102 7 5148 41
rect 5182 7 5228 41
rect 5262 7 5308 41
rect 5342 7 5388 41
rect 5422 7 5468 41
rect 5502 7 5548 41
rect 5582 7 5628 41
rect 5662 7 5708 41
rect 5742 7 5788 41
rect 5822 7 5868 41
rect 5902 7 5948 41
rect 5982 7 6005 41
rect 4325 -26 6005 7
rect -85 -2780 2235 -2747
rect -85 -2814 -62 -2780
rect -28 -2814 18 -2780
rect 52 -2814 98 -2780
rect 132 -2814 178 -2780
rect 212 -2814 258 -2780
rect 292 -2814 338 -2780
rect 372 -2814 418 -2780
rect 452 -2814 498 -2780
rect 532 -2814 578 -2780
rect 612 -2814 658 -2780
rect 692 -2814 738 -2780
rect 772 -2814 818 -2780
rect 852 -2814 898 -2780
rect 932 -2814 978 -2780
rect 1012 -2814 1058 -2780
rect 1092 -2814 1138 -2780
rect 1172 -2814 1218 -2780
rect 1252 -2814 1298 -2780
rect 1332 -2814 1378 -2780
rect 1412 -2814 1458 -2780
rect 1492 -2814 1538 -2780
rect 1572 -2814 1618 -2780
rect 1652 -2814 1698 -2780
rect 1732 -2814 1778 -2780
rect 1812 -2814 1858 -2780
rect 1892 -2814 1938 -2780
rect 1972 -2814 2018 -2780
rect 2052 -2814 2098 -2780
rect 2132 -2814 2178 -2780
rect 2212 -2814 2235 -2780
rect -85 -2847 2235 -2814
rect 2596 -2779 3976 -2746
rect 2596 -2813 2629 -2779
rect 2663 -2813 2709 -2779
rect 2743 -2813 2789 -2779
rect 2823 -2813 2869 -2779
rect 2903 -2813 2949 -2779
rect 2983 -2813 3029 -2779
rect 3063 -2813 3109 -2779
rect 3143 -2813 3189 -2779
rect 3223 -2813 3269 -2779
rect 3303 -2813 3349 -2779
rect 3383 -2813 3429 -2779
rect 3463 -2813 3509 -2779
rect 3543 -2813 3589 -2779
rect 3623 -2813 3669 -2779
rect 3703 -2813 3749 -2779
rect 3783 -2813 3829 -2779
rect 3863 -2813 3909 -2779
rect 3943 -2813 3976 -2779
rect 2596 -2846 3976 -2813
rect 4345 -2779 6345 -2746
rect 4345 -2813 4368 -2779
rect 4402 -2813 4448 -2779
rect 4482 -2813 4528 -2779
rect 4562 -2813 4608 -2779
rect 4642 -2813 4688 -2779
rect 4722 -2813 4768 -2779
rect 4802 -2813 4848 -2779
rect 4882 -2813 4928 -2779
rect 4962 -2813 5008 -2779
rect 5042 -2813 5088 -2779
rect 5122 -2813 5168 -2779
rect 5202 -2813 5248 -2779
rect 5282 -2813 5328 -2779
rect 5362 -2813 5408 -2779
rect 5442 -2813 5488 -2779
rect 5522 -2813 5568 -2779
rect 5602 -2813 5648 -2779
rect 5682 -2813 5728 -2779
rect 5762 -2813 5808 -2779
rect 5842 -2813 5888 -2779
rect 5922 -2813 5968 -2779
rect 6002 -2813 6048 -2779
rect 6082 -2813 6128 -2779
rect 6162 -2813 6208 -2779
rect 6242 -2813 6288 -2779
rect 6322 -2813 6345 -2779
rect 4345 -2846 6345 -2813
<< nsubdiff >>
rect -65 1221 2215 1254
rect -65 1187 18 1221
rect 52 1187 98 1221
rect 132 1187 178 1221
rect 212 1187 258 1221
rect 292 1187 338 1221
rect 372 1187 418 1221
rect 452 1187 498 1221
rect 532 1187 578 1221
rect 612 1187 658 1221
rect 692 1187 738 1221
rect 772 1187 818 1221
rect 852 1187 898 1221
rect 932 1187 978 1221
rect 1012 1187 1058 1221
rect 1092 1187 1138 1221
rect 1172 1187 1218 1221
rect 1252 1187 1298 1221
rect 1332 1187 1378 1221
rect 1412 1187 1458 1221
rect 1492 1187 1538 1221
rect 1572 1187 1618 1221
rect 1652 1187 1698 1221
rect 1732 1187 1778 1221
rect 1812 1187 1858 1221
rect 1892 1187 1938 1221
rect 1972 1187 2018 1221
rect 2052 1187 2098 1221
rect 2132 1187 2215 1221
rect -65 1154 2215 1187
rect 2595 1221 3975 1254
rect 2595 1187 2628 1221
rect 2662 1187 2708 1221
rect 2742 1187 2788 1221
rect 2822 1187 2868 1221
rect 2902 1187 2948 1221
rect 2982 1187 3028 1221
rect 3062 1187 3108 1221
rect 3142 1187 3188 1221
rect 3222 1187 3268 1221
rect 3302 1187 3348 1221
rect 3382 1187 3428 1221
rect 3462 1187 3508 1221
rect 3542 1187 3588 1221
rect 3622 1187 3668 1221
rect 3702 1187 3748 1221
rect 3782 1187 3828 1221
rect 3862 1187 3908 1221
rect 3942 1187 3975 1221
rect 2595 1154 3975 1187
rect 4325 1221 6005 1254
rect 4325 1187 4348 1221
rect 4382 1187 4428 1221
rect 4462 1187 4508 1221
rect 4542 1187 4588 1221
rect 4622 1187 4668 1221
rect 4702 1187 4748 1221
rect 4782 1187 4828 1221
rect 4862 1187 4908 1221
rect 4942 1187 4988 1221
rect 5022 1187 5068 1221
rect 5102 1187 5148 1221
rect 5182 1187 5228 1221
rect 5262 1187 5308 1221
rect 5342 1187 5388 1221
rect 5422 1187 5468 1221
rect 5502 1187 5548 1221
rect 5582 1187 5628 1221
rect 5662 1187 5708 1221
rect 5742 1187 5788 1221
rect 5822 1187 5868 1221
rect 5902 1187 5948 1221
rect 5982 1187 6005 1221
rect 4325 1154 6005 1187
rect -85 -1139 2235 -1106
rect -85 -1173 -62 -1139
rect -28 -1173 18 -1139
rect 52 -1173 98 -1139
rect 132 -1173 178 -1139
rect 212 -1173 258 -1139
rect 292 -1173 338 -1139
rect 372 -1173 418 -1139
rect 452 -1173 498 -1139
rect 532 -1173 578 -1139
rect 612 -1173 658 -1139
rect 692 -1173 738 -1139
rect 772 -1173 818 -1139
rect 852 -1173 898 -1139
rect 932 -1173 978 -1139
rect 1012 -1173 1058 -1139
rect 1092 -1173 1138 -1139
rect 1172 -1173 1218 -1139
rect 1252 -1173 1298 -1139
rect 1332 -1173 1378 -1139
rect 1412 -1173 1458 -1139
rect 1492 -1173 1538 -1139
rect 1572 -1173 1618 -1139
rect 1652 -1173 1698 -1139
rect 1732 -1173 1778 -1139
rect 1812 -1173 1858 -1139
rect 1892 -1173 1938 -1139
rect 1972 -1173 2018 -1139
rect 2052 -1173 2098 -1139
rect 2132 -1173 2178 -1139
rect 2212 -1173 2235 -1139
rect -85 -1280 2235 -1173
rect 2595 -1139 3975 -1106
rect 2595 -1173 2628 -1139
rect 2662 -1173 2708 -1139
rect 2742 -1173 2788 -1139
rect 2822 -1173 2868 -1139
rect 2902 -1173 2948 -1139
rect 2982 -1173 3028 -1139
rect 3062 -1173 3108 -1139
rect 3142 -1173 3188 -1139
rect 3222 -1173 3268 -1139
rect 3302 -1173 3348 -1139
rect 3382 -1173 3428 -1139
rect 3462 -1173 3508 -1139
rect 3542 -1173 3588 -1139
rect 3622 -1173 3668 -1139
rect 3702 -1173 3748 -1139
rect 3782 -1173 3828 -1139
rect 3862 -1173 3908 -1139
rect 3942 -1173 3975 -1139
rect 2595 -1206 3975 -1173
rect 4325 -1139 6005 -1106
rect 4325 -1173 4348 -1139
rect 4382 -1173 4428 -1139
rect 4462 -1173 4508 -1139
rect 4542 -1173 4588 -1139
rect 4622 -1173 4668 -1139
rect 4702 -1173 4748 -1139
rect 4782 -1173 4828 -1139
rect 4862 -1173 4908 -1139
rect 4942 -1173 4988 -1139
rect 5022 -1173 5068 -1139
rect 5102 -1173 5148 -1139
rect 5182 -1173 5228 -1139
rect 5262 -1173 5308 -1139
rect 5342 -1173 5388 -1139
rect 5422 -1173 5468 -1139
rect 5502 -1173 5548 -1139
rect 5582 -1173 5628 -1139
rect 5662 -1173 5708 -1139
rect 5742 -1173 5788 -1139
rect 5822 -1173 5868 -1139
rect 5902 -1173 5948 -1139
rect 5982 -1173 6005 -1139
rect 4325 -1206 6005 -1173
rect -85 -1314 -62 -1280
rect -28 -1314 18 -1280
rect 52 -1314 98 -1280
rect 132 -1314 178 -1280
rect 212 -1314 258 -1280
rect 292 -1314 338 -1280
rect 372 -1314 418 -1280
rect 452 -1314 498 -1280
rect 532 -1314 578 -1280
rect 612 -1314 658 -1280
rect 692 -1314 738 -1280
rect 772 -1314 818 -1280
rect 852 -1314 898 -1280
rect 932 -1314 978 -1280
rect 1012 -1314 1058 -1280
rect 1092 -1314 1138 -1280
rect 1172 -1314 1218 -1280
rect 1252 -1314 1298 -1280
rect 1332 -1314 1378 -1280
rect 1412 -1314 1458 -1280
rect 1492 -1314 1538 -1280
rect 1572 -1314 1618 -1280
rect 1652 -1314 1698 -1280
rect 1732 -1314 1778 -1280
rect 1812 -1314 1858 -1280
rect 1892 -1314 1938 -1280
rect 1972 -1314 2018 -1280
rect 2052 -1314 2098 -1280
rect 2132 -1314 2178 -1280
rect 2212 -1314 2235 -1280
rect -85 -1347 2235 -1314
rect 2596 -1599 3976 -1566
rect 2596 -1633 2629 -1599
rect 2663 -1633 2709 -1599
rect 2743 -1633 2789 -1599
rect 2823 -1633 2869 -1599
rect 2903 -1633 2949 -1599
rect 2983 -1633 3029 -1599
rect 3063 -1633 3109 -1599
rect 3143 -1633 3189 -1599
rect 3223 -1633 3269 -1599
rect 3303 -1633 3349 -1599
rect 3383 -1633 3429 -1599
rect 3463 -1633 3509 -1599
rect 3543 -1633 3589 -1599
rect 3623 -1633 3669 -1599
rect 3703 -1633 3749 -1599
rect 3783 -1633 3829 -1599
rect 3863 -1633 3909 -1599
rect 3943 -1633 3976 -1599
rect 2596 -1666 3976 -1633
rect 4345 -1599 6345 -1566
rect 4345 -1633 4368 -1599
rect 4402 -1633 4448 -1599
rect 4482 -1633 4528 -1599
rect 4562 -1633 4608 -1599
rect 4642 -1633 4688 -1599
rect 4722 -1633 4768 -1599
rect 4802 -1633 4848 -1599
rect 4882 -1633 4928 -1599
rect 4962 -1633 5008 -1599
rect 5042 -1633 5088 -1599
rect 5122 -1633 5168 -1599
rect 5202 -1633 5248 -1599
rect 5282 -1633 5328 -1599
rect 5362 -1633 5408 -1599
rect 5442 -1633 5488 -1599
rect 5522 -1633 5568 -1599
rect 5602 -1633 5648 -1599
rect 5682 -1633 5728 -1599
rect 5762 -1633 5808 -1599
rect 5842 -1633 5888 -1599
rect 5922 -1633 5968 -1599
rect 6002 -1633 6048 -1599
rect 6082 -1633 6128 -1599
rect 6162 -1633 6208 -1599
rect 6242 -1633 6288 -1599
rect 6322 -1633 6345 -1599
rect 4345 -1666 6345 -1633
<< psubdiffcont >>
rect 18 7 52 41
rect 98 7 132 41
rect 178 7 212 41
rect 258 7 292 41
rect 338 7 372 41
rect 418 7 452 41
rect 498 7 532 41
rect 578 7 612 41
rect 658 7 692 41
rect 738 7 772 41
rect 818 7 852 41
rect 898 7 932 41
rect 978 7 1012 41
rect 1058 7 1092 41
rect 1138 7 1172 41
rect 1218 7 1252 41
rect 1298 7 1332 41
rect 1378 7 1412 41
rect 1458 7 1492 41
rect 1538 7 1572 41
rect 1618 7 1652 41
rect 1698 7 1732 41
rect 1778 7 1812 41
rect 1858 7 1892 41
rect 1938 7 1972 41
rect 2018 7 2052 41
rect 2098 7 2132 41
rect 2628 7 2662 41
rect 2708 7 2742 41
rect 2788 7 2822 41
rect 2868 7 2902 41
rect 2948 7 2982 41
rect 3028 7 3062 41
rect 3108 7 3142 41
rect 3188 7 3222 41
rect 3268 7 3302 41
rect 3348 7 3382 41
rect 3428 7 3462 41
rect 3508 7 3542 41
rect 3588 7 3622 41
rect 3668 7 3702 41
rect 3748 7 3782 41
rect 3828 7 3862 41
rect 3908 7 3942 41
rect 4348 7 4382 41
rect 4428 7 4462 41
rect 4508 7 4542 41
rect 4588 7 4622 41
rect 4668 7 4702 41
rect 4748 7 4782 41
rect 4828 7 4862 41
rect 4908 7 4942 41
rect 4988 7 5022 41
rect 5068 7 5102 41
rect 5148 7 5182 41
rect 5228 7 5262 41
rect 5308 7 5342 41
rect 5388 7 5422 41
rect 5468 7 5502 41
rect 5548 7 5582 41
rect 5628 7 5662 41
rect 5708 7 5742 41
rect 5788 7 5822 41
rect 5868 7 5902 41
rect 5948 7 5982 41
rect -62 -2814 -28 -2780
rect 18 -2814 52 -2780
rect 98 -2814 132 -2780
rect 178 -2814 212 -2780
rect 258 -2814 292 -2780
rect 338 -2814 372 -2780
rect 418 -2814 452 -2780
rect 498 -2814 532 -2780
rect 578 -2814 612 -2780
rect 658 -2814 692 -2780
rect 738 -2814 772 -2780
rect 818 -2814 852 -2780
rect 898 -2814 932 -2780
rect 978 -2814 1012 -2780
rect 1058 -2814 1092 -2780
rect 1138 -2814 1172 -2780
rect 1218 -2814 1252 -2780
rect 1298 -2814 1332 -2780
rect 1378 -2814 1412 -2780
rect 1458 -2814 1492 -2780
rect 1538 -2814 1572 -2780
rect 1618 -2814 1652 -2780
rect 1698 -2814 1732 -2780
rect 1778 -2814 1812 -2780
rect 1858 -2814 1892 -2780
rect 1938 -2814 1972 -2780
rect 2018 -2814 2052 -2780
rect 2098 -2814 2132 -2780
rect 2178 -2814 2212 -2780
rect 2629 -2813 2663 -2779
rect 2709 -2813 2743 -2779
rect 2789 -2813 2823 -2779
rect 2869 -2813 2903 -2779
rect 2949 -2813 2983 -2779
rect 3029 -2813 3063 -2779
rect 3109 -2813 3143 -2779
rect 3189 -2813 3223 -2779
rect 3269 -2813 3303 -2779
rect 3349 -2813 3383 -2779
rect 3429 -2813 3463 -2779
rect 3509 -2813 3543 -2779
rect 3589 -2813 3623 -2779
rect 3669 -2813 3703 -2779
rect 3749 -2813 3783 -2779
rect 3829 -2813 3863 -2779
rect 3909 -2813 3943 -2779
rect 4368 -2813 4402 -2779
rect 4448 -2813 4482 -2779
rect 4528 -2813 4562 -2779
rect 4608 -2813 4642 -2779
rect 4688 -2813 4722 -2779
rect 4768 -2813 4802 -2779
rect 4848 -2813 4882 -2779
rect 4928 -2813 4962 -2779
rect 5008 -2813 5042 -2779
rect 5088 -2813 5122 -2779
rect 5168 -2813 5202 -2779
rect 5248 -2813 5282 -2779
rect 5328 -2813 5362 -2779
rect 5408 -2813 5442 -2779
rect 5488 -2813 5522 -2779
rect 5568 -2813 5602 -2779
rect 5648 -2813 5682 -2779
rect 5728 -2813 5762 -2779
rect 5808 -2813 5842 -2779
rect 5888 -2813 5922 -2779
rect 5968 -2813 6002 -2779
rect 6048 -2813 6082 -2779
rect 6128 -2813 6162 -2779
rect 6208 -2813 6242 -2779
rect 6288 -2813 6322 -2779
<< nsubdiffcont >>
rect 18 1187 52 1221
rect 98 1187 132 1221
rect 178 1187 212 1221
rect 258 1187 292 1221
rect 338 1187 372 1221
rect 418 1187 452 1221
rect 498 1187 532 1221
rect 578 1187 612 1221
rect 658 1187 692 1221
rect 738 1187 772 1221
rect 818 1187 852 1221
rect 898 1187 932 1221
rect 978 1187 1012 1221
rect 1058 1187 1092 1221
rect 1138 1187 1172 1221
rect 1218 1187 1252 1221
rect 1298 1187 1332 1221
rect 1378 1187 1412 1221
rect 1458 1187 1492 1221
rect 1538 1187 1572 1221
rect 1618 1187 1652 1221
rect 1698 1187 1732 1221
rect 1778 1187 1812 1221
rect 1858 1187 1892 1221
rect 1938 1187 1972 1221
rect 2018 1187 2052 1221
rect 2098 1187 2132 1221
rect 2628 1187 2662 1221
rect 2708 1187 2742 1221
rect 2788 1187 2822 1221
rect 2868 1187 2902 1221
rect 2948 1187 2982 1221
rect 3028 1187 3062 1221
rect 3108 1187 3142 1221
rect 3188 1187 3222 1221
rect 3268 1187 3302 1221
rect 3348 1187 3382 1221
rect 3428 1187 3462 1221
rect 3508 1187 3542 1221
rect 3588 1187 3622 1221
rect 3668 1187 3702 1221
rect 3748 1187 3782 1221
rect 3828 1187 3862 1221
rect 3908 1187 3942 1221
rect 4348 1187 4382 1221
rect 4428 1187 4462 1221
rect 4508 1187 4542 1221
rect 4588 1187 4622 1221
rect 4668 1187 4702 1221
rect 4748 1187 4782 1221
rect 4828 1187 4862 1221
rect 4908 1187 4942 1221
rect 4988 1187 5022 1221
rect 5068 1187 5102 1221
rect 5148 1187 5182 1221
rect 5228 1187 5262 1221
rect 5308 1187 5342 1221
rect 5388 1187 5422 1221
rect 5468 1187 5502 1221
rect 5548 1187 5582 1221
rect 5628 1187 5662 1221
rect 5708 1187 5742 1221
rect 5788 1187 5822 1221
rect 5868 1187 5902 1221
rect 5948 1187 5982 1221
rect -62 -1173 -28 -1139
rect 18 -1173 52 -1139
rect 98 -1173 132 -1139
rect 178 -1173 212 -1139
rect 258 -1173 292 -1139
rect 338 -1173 372 -1139
rect 418 -1173 452 -1139
rect 498 -1173 532 -1139
rect 578 -1173 612 -1139
rect 658 -1173 692 -1139
rect 738 -1173 772 -1139
rect 818 -1173 852 -1139
rect 898 -1173 932 -1139
rect 978 -1173 1012 -1139
rect 1058 -1173 1092 -1139
rect 1138 -1173 1172 -1139
rect 1218 -1173 1252 -1139
rect 1298 -1173 1332 -1139
rect 1378 -1173 1412 -1139
rect 1458 -1173 1492 -1139
rect 1538 -1173 1572 -1139
rect 1618 -1173 1652 -1139
rect 1698 -1173 1732 -1139
rect 1778 -1173 1812 -1139
rect 1858 -1173 1892 -1139
rect 1938 -1173 1972 -1139
rect 2018 -1173 2052 -1139
rect 2098 -1173 2132 -1139
rect 2178 -1173 2212 -1139
rect 2628 -1173 2662 -1139
rect 2708 -1173 2742 -1139
rect 2788 -1173 2822 -1139
rect 2868 -1173 2902 -1139
rect 2948 -1173 2982 -1139
rect 3028 -1173 3062 -1139
rect 3108 -1173 3142 -1139
rect 3188 -1173 3222 -1139
rect 3268 -1173 3302 -1139
rect 3348 -1173 3382 -1139
rect 3428 -1173 3462 -1139
rect 3508 -1173 3542 -1139
rect 3588 -1173 3622 -1139
rect 3668 -1173 3702 -1139
rect 3748 -1173 3782 -1139
rect 3828 -1173 3862 -1139
rect 3908 -1173 3942 -1139
rect 4348 -1173 4382 -1139
rect 4428 -1173 4462 -1139
rect 4508 -1173 4542 -1139
rect 4588 -1173 4622 -1139
rect 4668 -1173 4702 -1139
rect 4748 -1173 4782 -1139
rect 4828 -1173 4862 -1139
rect 4908 -1173 4942 -1139
rect 4988 -1173 5022 -1139
rect 5068 -1173 5102 -1139
rect 5148 -1173 5182 -1139
rect 5228 -1173 5262 -1139
rect 5308 -1173 5342 -1139
rect 5388 -1173 5422 -1139
rect 5468 -1173 5502 -1139
rect 5548 -1173 5582 -1139
rect 5628 -1173 5662 -1139
rect 5708 -1173 5742 -1139
rect 5788 -1173 5822 -1139
rect 5868 -1173 5902 -1139
rect 5948 -1173 5982 -1139
rect -62 -1314 -28 -1280
rect 18 -1314 52 -1280
rect 98 -1314 132 -1280
rect 178 -1314 212 -1280
rect 258 -1314 292 -1280
rect 338 -1314 372 -1280
rect 418 -1314 452 -1280
rect 498 -1314 532 -1280
rect 578 -1314 612 -1280
rect 658 -1314 692 -1280
rect 738 -1314 772 -1280
rect 818 -1314 852 -1280
rect 898 -1314 932 -1280
rect 978 -1314 1012 -1280
rect 1058 -1314 1092 -1280
rect 1138 -1314 1172 -1280
rect 1218 -1314 1252 -1280
rect 1298 -1314 1332 -1280
rect 1378 -1314 1412 -1280
rect 1458 -1314 1492 -1280
rect 1538 -1314 1572 -1280
rect 1618 -1314 1652 -1280
rect 1698 -1314 1732 -1280
rect 1778 -1314 1812 -1280
rect 1858 -1314 1892 -1280
rect 1938 -1314 1972 -1280
rect 2018 -1314 2052 -1280
rect 2098 -1314 2132 -1280
rect 2178 -1314 2212 -1280
rect 2629 -1633 2663 -1599
rect 2709 -1633 2743 -1599
rect 2789 -1633 2823 -1599
rect 2869 -1633 2903 -1599
rect 2949 -1633 2983 -1599
rect 3029 -1633 3063 -1599
rect 3109 -1633 3143 -1599
rect 3189 -1633 3223 -1599
rect 3269 -1633 3303 -1599
rect 3349 -1633 3383 -1599
rect 3429 -1633 3463 -1599
rect 3509 -1633 3543 -1599
rect 3589 -1633 3623 -1599
rect 3669 -1633 3703 -1599
rect 3749 -1633 3783 -1599
rect 3829 -1633 3863 -1599
rect 3909 -1633 3943 -1599
rect 4368 -1633 4402 -1599
rect 4448 -1633 4482 -1599
rect 4528 -1633 4562 -1599
rect 4608 -1633 4642 -1599
rect 4688 -1633 4722 -1599
rect 4768 -1633 4802 -1599
rect 4848 -1633 4882 -1599
rect 4928 -1633 4962 -1599
rect 5008 -1633 5042 -1599
rect 5088 -1633 5122 -1599
rect 5168 -1633 5202 -1599
rect 5248 -1633 5282 -1599
rect 5328 -1633 5362 -1599
rect 5408 -1633 5442 -1599
rect 5488 -1633 5522 -1599
rect 5568 -1633 5602 -1599
rect 5648 -1633 5682 -1599
rect 5728 -1633 5762 -1599
rect 5808 -1633 5842 -1599
rect 5888 -1633 5922 -1599
rect 5968 -1633 6002 -1599
rect 6048 -1633 6082 -1599
rect 6128 -1633 6162 -1599
rect 6208 -1633 6242 -1599
rect 6288 -1633 6322 -1599
<< poly >>
rect 325 1091 405 1114
rect 325 1057 348 1091
rect 382 1057 405 1091
rect 835 1104 1015 1134
rect 835 1074 865 1104
rect 985 1074 1015 1104
rect 1135 1104 1315 1134
rect 1135 1074 1165 1104
rect 1285 1074 1315 1104
rect 1715 1091 1795 1114
rect 325 1034 405 1057
rect 205 991 285 1014
rect 205 957 228 991
rect 262 957 285 991
rect 205 934 285 957
rect 5 791 85 814
rect 5 757 28 791
rect 62 757 85 791
rect 5 734 85 757
rect 55 514 85 734
rect 205 514 235 934
rect 355 514 385 1034
rect 455 891 535 914
rect 455 857 478 891
rect 512 857 535 891
rect 455 834 535 857
rect 505 514 535 834
rect 1715 1057 1738 1091
rect 1772 1057 1795 1091
rect 3045 1104 3225 1134
rect 3045 1074 3075 1104
rect 3195 1074 3225 1104
rect 3345 1104 3525 1134
rect 3345 1074 3375 1104
rect 3495 1074 3525 1104
rect 4925 1104 5105 1134
rect 4925 1074 4955 1104
rect 5075 1074 5105 1104
rect 5225 1104 5405 1134
rect 5225 1074 5255 1104
rect 5375 1074 5405 1104
rect 1715 1034 1795 1057
rect 1615 791 1695 814
rect 835 744 865 774
rect 985 619 1015 774
rect 1135 744 1165 774
rect 1285 744 1315 774
rect 1615 757 1638 791
rect 1672 757 1695 791
rect 1085 721 1165 744
rect 1085 687 1108 721
rect 1142 687 1165 721
rect 1085 664 1165 687
rect 985 596 1065 619
rect 985 562 1008 596
rect 1042 562 1065 596
rect 835 514 865 544
rect 985 539 1065 562
rect 985 514 1015 539
rect 1135 514 1165 664
rect 1615 734 1695 757
rect 1285 514 1315 544
rect 1615 514 1645 734
rect 1765 514 1795 1034
rect 1915 991 1995 1014
rect 1915 957 1938 991
rect 1972 957 1995 991
rect 1915 934 1995 957
rect 1915 514 1945 934
rect 2065 891 2145 914
rect 2065 857 2088 891
rect 2122 857 2145 891
rect 2065 834 2145 857
rect 2065 514 2095 834
rect 3825 841 3905 864
rect 3825 807 3848 841
rect 3882 807 3905 841
rect 3825 784 3905 807
rect 3045 744 3075 774
rect 2665 601 2745 624
rect 2665 567 2688 601
rect 2722 567 2745 601
rect 2665 544 2745 567
rect 3195 619 3225 774
rect 3345 744 3375 774
rect 3495 744 3525 774
rect 3295 721 3375 744
rect 3295 687 3318 721
rect 3352 687 3375 721
rect 3295 664 3375 687
rect 3195 596 3275 619
rect 3195 562 3218 596
rect 3252 562 3275 596
rect 2715 514 2745 544
rect 3045 514 3075 544
rect 3195 539 3275 562
rect 3195 514 3225 539
rect 3345 514 3375 664
rect 3495 514 3525 544
rect 3825 514 3855 784
rect 4545 771 4625 794
rect 5805 991 5885 1014
rect 5805 957 5828 991
rect 5862 957 5885 991
rect 5805 934 5885 957
rect 5655 871 5735 894
rect 5655 837 5678 871
rect 5712 837 5735 871
rect 5655 814 5735 837
rect 4545 737 4568 771
rect 4602 737 4625 771
rect 4925 744 4955 774
rect 4545 714 4625 737
rect 4395 671 4475 694
rect 4395 637 4418 671
rect 4452 637 4475 671
rect 4395 614 4475 637
rect 4445 514 4475 614
rect 4595 514 4625 714
rect 5075 619 5105 774
rect 5225 744 5255 774
rect 5375 744 5405 774
rect 5175 721 5255 744
rect 5175 687 5198 721
rect 5232 687 5255 721
rect 5175 664 5255 687
rect 5075 596 5155 619
rect 5075 562 5098 596
rect 5132 562 5155 596
rect 4925 514 4955 544
rect 5075 539 5155 562
rect 5075 514 5105 539
rect 5225 514 5255 664
rect 5375 514 5405 544
rect 5705 514 5735 814
rect 5855 514 5885 934
rect 55 184 85 214
rect 205 184 235 214
rect 355 184 385 214
rect 505 184 535 214
rect 835 184 865 214
rect 985 184 1015 214
rect 1135 184 1165 214
rect 1285 184 1315 214
rect 1615 184 1645 214
rect 835 161 915 184
rect 835 127 858 161
rect 892 127 915 161
rect 835 104 915 127
rect 1235 161 1315 184
rect 1765 174 1795 214
rect 1915 174 1945 214
rect 2065 174 2095 214
rect 2715 184 2745 214
rect 3045 184 3075 214
rect 3195 184 3225 214
rect 3345 184 3375 214
rect 3495 184 3525 214
rect 3825 184 3855 214
rect 4445 184 4475 214
rect 4595 184 4625 214
rect 4925 184 4955 214
rect 5075 184 5105 214
rect 5225 184 5255 214
rect 5375 184 5405 214
rect 5705 184 5735 214
rect 5855 184 5885 214
rect 1235 127 1258 161
rect 1292 127 1315 161
rect 1235 104 1315 127
rect 3045 161 3125 184
rect 3045 127 3068 161
rect 3102 127 3125 161
rect 3045 104 3125 127
rect 3445 161 3525 184
rect 3445 127 3468 161
rect 3502 127 3525 161
rect 3445 104 3525 127
rect 4925 161 5005 184
rect 4925 127 4948 161
rect 4982 127 5005 161
rect 4925 104 5005 127
rect 5325 161 5405 184
rect 5325 127 5348 161
rect 5382 127 5405 161
rect 5325 104 5405 127
rect 835 -79 915 -56
rect 835 -113 858 -79
rect 892 -113 915 -79
rect 835 -136 915 -113
rect 1235 -79 1315 -56
rect 1235 -113 1258 -79
rect 1292 -113 1315 -79
rect 1235 -136 1315 -113
rect 3045 -79 3125 -56
rect 3045 -113 3068 -79
rect 3102 -113 3125 -79
rect 55 -166 85 -136
rect 205 -166 235 -136
rect 355 -166 385 -136
rect 505 -166 535 -136
rect 835 -166 865 -136
rect 985 -166 1015 -136
rect 1135 -166 1165 -136
rect 1285 -166 1315 -136
rect 1615 -166 1645 -136
rect 1765 -166 1795 -126
rect 1915 -166 1945 -126
rect 2065 -166 2095 -126
rect 3045 -136 3125 -113
rect 3445 -79 3525 -56
rect 3445 -113 3468 -79
rect 3502 -113 3525 -79
rect 3445 -136 3525 -113
rect 4925 -79 5005 -56
rect 4925 -113 4948 -79
rect 4982 -113 5005 -79
rect 4925 -136 5005 -113
rect 5325 -79 5405 -56
rect 5325 -113 5348 -79
rect 5382 -113 5405 -79
rect 5325 -136 5405 -113
rect 2715 -166 2745 -136
rect 3045 -166 3075 -136
rect 3195 -166 3225 -136
rect 3345 -166 3375 -136
rect 3495 -166 3525 -136
rect 3825 -166 3855 -136
rect 4445 -166 4475 -136
rect 4595 -166 4625 -136
rect 4925 -166 4955 -136
rect 5075 -166 5105 -136
rect 5225 -166 5255 -136
rect 5375 -166 5405 -136
rect 5705 -166 5735 -136
rect 5855 -166 5885 -136
rect 55 -686 85 -466
rect 5 -709 85 -686
rect 5 -743 28 -709
rect 62 -743 85 -709
rect 5 -766 85 -743
rect 205 -886 235 -466
rect 205 -909 285 -886
rect 205 -943 228 -909
rect 262 -943 285 -909
rect 205 -966 285 -943
rect 355 -986 385 -466
rect 505 -786 535 -466
rect 835 -496 865 -466
rect 985 -491 1015 -466
rect 985 -514 1065 -491
rect 985 -548 1008 -514
rect 1042 -548 1065 -514
rect 985 -571 1065 -548
rect 835 -726 865 -696
rect 985 -726 1015 -571
rect 1135 -616 1165 -466
rect 1285 -496 1315 -466
rect 1085 -639 1165 -616
rect 1085 -673 1108 -639
rect 1142 -673 1165 -639
rect 1085 -696 1165 -673
rect 1615 -686 1645 -466
rect 1135 -726 1165 -696
rect 1285 -726 1315 -696
rect 1615 -709 1695 -686
rect 455 -809 535 -786
rect 455 -843 478 -809
rect 512 -843 535 -809
rect 455 -866 535 -843
rect 325 -1009 405 -986
rect 325 -1043 348 -1009
rect 382 -1043 405 -1009
rect 1615 -743 1638 -709
rect 1672 -743 1695 -709
rect 1615 -766 1695 -743
rect 1765 -986 1795 -466
rect 1915 -886 1945 -466
rect 2065 -786 2095 -466
rect 2715 -496 2745 -466
rect 3045 -496 3075 -466
rect 3195 -491 3225 -466
rect 2665 -519 2745 -496
rect 2665 -553 2688 -519
rect 2722 -553 2745 -519
rect 2665 -576 2745 -553
rect 3195 -514 3275 -491
rect 3195 -548 3218 -514
rect 3252 -548 3275 -514
rect 3195 -571 3275 -548
rect 3045 -726 3075 -696
rect 3195 -726 3225 -571
rect 3345 -616 3375 -466
rect 3495 -496 3525 -466
rect 3295 -639 3375 -616
rect 3295 -673 3318 -639
rect 3352 -673 3375 -639
rect 3295 -696 3375 -673
rect 3345 -726 3375 -696
rect 3495 -726 3525 -696
rect 2065 -809 2145 -786
rect 2065 -843 2088 -809
rect 2122 -843 2145 -809
rect 2065 -866 2145 -843
rect 1915 -909 1995 -886
rect 1915 -943 1938 -909
rect 1972 -943 1995 -909
rect 1915 -966 1995 -943
rect 1715 -1009 1795 -986
rect 325 -1066 405 -1043
rect 835 -1056 865 -1026
rect 985 -1056 1015 -1026
rect 835 -1086 1015 -1056
rect 1135 -1056 1165 -1026
rect 1285 -1056 1315 -1026
rect 1135 -1086 1315 -1056
rect 1715 -1043 1738 -1009
rect 1772 -1043 1795 -1009
rect 3825 -736 3855 -466
rect 4445 -566 4475 -466
rect 4395 -589 4475 -566
rect 4395 -623 4418 -589
rect 4452 -623 4475 -589
rect 4395 -646 4475 -623
rect 4595 -666 4625 -466
rect 4925 -496 4955 -466
rect 5075 -491 5105 -466
rect 4545 -689 4625 -666
rect 4545 -723 4568 -689
rect 4602 -723 4625 -689
rect 5075 -514 5155 -491
rect 5075 -548 5098 -514
rect 5132 -548 5155 -514
rect 5075 -571 5155 -548
rect 3825 -759 3905 -736
rect 4545 -746 4625 -723
rect 4925 -726 4955 -696
rect 5075 -726 5105 -571
rect 5225 -616 5255 -466
rect 5375 -496 5405 -466
rect 5175 -639 5255 -616
rect 5175 -673 5198 -639
rect 5232 -673 5255 -639
rect 5175 -696 5255 -673
rect 5225 -726 5255 -696
rect 5375 -726 5405 -696
rect 3825 -793 3848 -759
rect 3882 -793 3905 -759
rect 3825 -816 3905 -793
rect 5705 -766 5735 -466
rect 5655 -789 5735 -766
rect 5655 -823 5678 -789
rect 5712 -823 5735 -789
rect 5655 -846 5735 -823
rect 5855 -886 5885 -466
rect 5805 -909 5885 -886
rect 5805 -943 5828 -909
rect 5862 -943 5885 -909
rect 5805 -966 5885 -943
rect 1715 -1066 1795 -1043
rect 3045 -1056 3075 -1026
rect 3195 -1056 3225 -1026
rect 3045 -1086 3225 -1056
rect 3345 -1056 3375 -1026
rect 3495 -1056 3525 -1026
rect 3345 -1086 3525 -1056
rect 4925 -1056 4955 -1026
rect 5075 -1056 5105 -1026
rect 4925 -1086 5105 -1056
rect 5225 -1056 5255 -1026
rect 5375 -1056 5405 -1026
rect 5225 -1086 5405 -1056
rect 835 -1397 1015 -1367
rect 835 -1427 865 -1397
rect 985 -1427 1015 -1397
rect 1135 -1397 1315 -1367
rect 1135 -1427 1165 -1397
rect 1285 -1427 1315 -1397
rect 3046 -1716 3226 -1686
rect 835 -1757 865 -1727
rect 455 -1870 535 -1847
rect 455 -1904 478 -1870
rect 512 -1904 535 -1870
rect 455 -1927 535 -1904
rect 305 -1970 385 -1947
rect 305 -2004 328 -1970
rect 362 -2004 385 -1970
rect 305 -2027 385 -2004
rect 155 -2070 235 -2047
rect 155 -2104 178 -2070
rect 212 -2104 235 -2070
rect 155 -2127 235 -2104
rect 5 -2170 85 -2147
rect 5 -2204 28 -2170
rect 62 -2204 85 -2170
rect 5 -2227 85 -2204
rect 55 -2307 85 -2227
rect 205 -2307 235 -2127
rect 355 -2307 385 -2027
rect 505 -2307 535 -1927
rect 985 -1987 1015 -1727
rect 1135 -1847 1165 -1727
rect 1285 -1757 1315 -1727
rect 3046 -1746 3076 -1716
rect 3196 -1746 3226 -1716
rect 3346 -1716 3526 -1686
rect 3346 -1746 3376 -1716
rect 3496 -1746 3526 -1716
rect 4475 -1729 4555 -1706
rect 1085 -1870 1165 -1847
rect 1085 -1904 1108 -1870
rect 1142 -1904 1165 -1870
rect 1085 -1927 1165 -1904
rect 985 -2010 1065 -1987
rect 985 -2044 1008 -2010
rect 1042 -2044 1065 -2010
rect 985 -2067 1065 -2044
rect 835 -2307 865 -2277
rect 985 -2307 1015 -2067
rect 1135 -2307 1165 -1927
rect 4475 -1763 4498 -1729
rect 4532 -1763 4555 -1729
rect 5105 -1716 5285 -1686
rect 5105 -1746 5135 -1716
rect 5255 -1746 5285 -1716
rect 5405 -1716 5585 -1686
rect 5405 -1746 5435 -1716
rect 5555 -1746 5585 -1716
rect 4475 -1786 4555 -1763
rect 3826 -1979 3906 -1956
rect 3826 -2013 3849 -1979
rect 3883 -2013 3906 -1979
rect 3826 -2036 3906 -2013
rect 3046 -2076 3076 -2046
rect 1565 -2170 1645 -2147
rect 1565 -2204 1588 -2170
rect 1622 -2204 1645 -2170
rect 1565 -2227 1645 -2204
rect 1715 -2170 1795 -2147
rect 1715 -2204 1738 -2170
rect 1772 -2204 1795 -2170
rect 1715 -2227 1795 -2204
rect 1865 -2170 1945 -2147
rect 1865 -2204 1888 -2170
rect 1922 -2204 1945 -2170
rect 1865 -2227 1945 -2204
rect 2015 -2170 2095 -2147
rect 2015 -2204 2038 -2170
rect 2072 -2204 2095 -2170
rect 2015 -2227 2095 -2204
rect 1285 -2307 1315 -2277
rect 1615 -2307 1645 -2227
rect 1765 -2307 1795 -2227
rect 1915 -2307 1945 -2227
rect 2065 -2307 2095 -2227
rect 2666 -2219 2746 -2196
rect 2666 -2253 2689 -2219
rect 2723 -2253 2746 -2219
rect 2666 -2276 2746 -2253
rect 3196 -2201 3226 -2046
rect 3346 -2076 3376 -2046
rect 3496 -2076 3526 -2046
rect 3296 -2099 3376 -2076
rect 3296 -2133 3319 -2099
rect 3353 -2133 3376 -2099
rect 3296 -2156 3376 -2133
rect 3196 -2224 3276 -2201
rect 3196 -2258 3219 -2224
rect 3253 -2258 3276 -2224
rect 2716 -2306 2746 -2276
rect 3046 -2306 3076 -2276
rect 3196 -2281 3276 -2258
rect 3196 -2306 3226 -2281
rect 3346 -2306 3376 -2156
rect 3496 -2306 3526 -2276
rect 3826 -2306 3856 -2036
rect 4475 -2306 4505 -1786
rect 4587 -1849 4667 -1826
rect 4587 -1883 4610 -1849
rect 4644 -1883 4667 -1849
rect 4587 -1906 4667 -1883
rect 4625 -2306 4655 -1906
rect 4775 -1939 4855 -1916
rect 4775 -1973 4798 -1939
rect 4832 -1973 4855 -1939
rect 4775 -1996 4855 -1973
rect 4775 -2306 4805 -1996
rect 5105 -2076 5135 -2046
rect 5255 -2076 5285 -2046
rect 5255 -2099 5335 -2076
rect 5255 -2133 5278 -2099
rect 5312 -2133 5335 -2099
rect 5255 -2156 5335 -2133
rect 5105 -2306 5135 -2276
rect 5255 -2306 5285 -2156
rect 5405 -2201 5435 -2046
rect 5555 -2076 5585 -2046
rect 6175 -2049 6255 -2026
rect 6175 -2083 6198 -2049
rect 6232 -2083 6255 -2049
rect 6175 -2106 6255 -2083
rect 5355 -2224 5435 -2201
rect 6035 -2149 6115 -2126
rect 6035 -2183 6058 -2149
rect 6092 -2183 6115 -2149
rect 6035 -2206 6115 -2183
rect 5355 -2258 5378 -2224
rect 5412 -2258 5435 -2224
rect 5355 -2281 5435 -2258
rect 5885 -2229 5965 -2206
rect 5885 -2263 5908 -2229
rect 5942 -2263 5965 -2229
rect 5405 -2306 5435 -2281
rect 5555 -2306 5585 -2276
rect 5885 -2286 5965 -2263
rect 5885 -2306 5915 -2286
rect 6035 -2306 6065 -2206
rect 6185 -2306 6215 -2106
rect 55 -2637 85 -2607
rect 205 -2637 235 -2607
rect 355 -2637 385 -2607
rect 505 -2637 535 -2607
rect 835 -2637 865 -2607
rect 985 -2637 1015 -2607
rect 1135 -2637 1165 -2607
rect 1285 -2637 1315 -2607
rect 1615 -2637 1645 -2607
rect 1765 -2637 1795 -2607
rect 1915 -2637 1945 -2607
rect 2065 -2637 2095 -2607
rect 2716 -2636 2746 -2606
rect 3046 -2636 3076 -2606
rect 3196 -2636 3226 -2606
rect 3346 -2636 3376 -2606
rect 3496 -2636 3526 -2606
rect 3826 -2636 3856 -2606
rect 4475 -2636 4505 -2606
rect 4625 -2636 4655 -2606
rect 4775 -2636 4805 -2606
rect 5105 -2636 5135 -2606
rect 5255 -2636 5285 -2606
rect 5405 -2636 5435 -2606
rect 5555 -2636 5585 -2606
rect 5885 -2636 5915 -2606
rect 6035 -2636 6065 -2606
rect 6185 -2636 6215 -2606
rect 835 -2660 915 -2637
rect 835 -2694 858 -2660
rect 892 -2694 915 -2660
rect 835 -2717 915 -2694
rect 1235 -2660 1315 -2637
rect 1235 -2694 1258 -2660
rect 1292 -2694 1315 -2660
rect 1235 -2717 1315 -2694
rect 3046 -2659 3126 -2636
rect 3046 -2693 3069 -2659
rect 3103 -2693 3126 -2659
rect 3046 -2716 3126 -2693
rect 3446 -2659 3526 -2636
rect 3446 -2693 3469 -2659
rect 3503 -2693 3526 -2659
rect 3446 -2716 3526 -2693
rect 5105 -2659 5185 -2636
rect 5105 -2693 5128 -2659
rect 5162 -2693 5185 -2659
rect 5105 -2716 5185 -2693
rect 5505 -2659 5585 -2636
rect 5505 -2693 5528 -2659
rect 5562 -2693 5585 -2659
rect 5505 -2716 5585 -2693
<< polycont >>
rect 348 1057 382 1091
rect 228 957 262 991
rect 28 757 62 791
rect 478 857 512 891
rect 1738 1057 1772 1091
rect 1638 757 1672 791
rect 1108 687 1142 721
rect 1008 562 1042 596
rect 1938 957 1972 991
rect 2088 857 2122 891
rect 3848 807 3882 841
rect 2688 567 2722 601
rect 3318 687 3352 721
rect 3218 562 3252 596
rect 5828 957 5862 991
rect 5678 837 5712 871
rect 4568 737 4602 771
rect 4418 637 4452 671
rect 5198 687 5232 721
rect 5098 562 5132 596
rect 858 127 892 161
rect 1258 127 1292 161
rect 3068 127 3102 161
rect 3468 127 3502 161
rect 4948 127 4982 161
rect 5348 127 5382 161
rect 858 -113 892 -79
rect 1258 -113 1292 -79
rect 3068 -113 3102 -79
rect 3468 -113 3502 -79
rect 4948 -113 4982 -79
rect 5348 -113 5382 -79
rect 28 -743 62 -709
rect 228 -943 262 -909
rect 1008 -548 1042 -514
rect 1108 -673 1142 -639
rect 478 -843 512 -809
rect 348 -1043 382 -1009
rect 1638 -743 1672 -709
rect 2688 -553 2722 -519
rect 3218 -548 3252 -514
rect 3318 -673 3352 -639
rect 2088 -843 2122 -809
rect 1938 -943 1972 -909
rect 1738 -1043 1772 -1009
rect 4418 -623 4452 -589
rect 4568 -723 4602 -689
rect 5098 -548 5132 -514
rect 5198 -673 5232 -639
rect 3848 -793 3882 -759
rect 5678 -823 5712 -789
rect 5828 -943 5862 -909
rect 478 -1904 512 -1870
rect 328 -2004 362 -1970
rect 178 -2104 212 -2070
rect 28 -2204 62 -2170
rect 1108 -1904 1142 -1870
rect 1008 -2044 1042 -2010
rect 4498 -1763 4532 -1729
rect 3849 -2013 3883 -1979
rect 1588 -2204 1622 -2170
rect 1738 -2204 1772 -2170
rect 1888 -2204 1922 -2170
rect 2038 -2204 2072 -2170
rect 2689 -2253 2723 -2219
rect 3319 -2133 3353 -2099
rect 3219 -2258 3253 -2224
rect 4610 -1883 4644 -1849
rect 4798 -1973 4832 -1939
rect 5278 -2133 5312 -2099
rect 6198 -2083 6232 -2049
rect 6058 -2183 6092 -2149
rect 5378 -2258 5412 -2224
rect 5908 -2263 5942 -2229
rect 858 -2694 892 -2660
rect 1258 -2694 1292 -2660
rect 3069 -2693 3103 -2659
rect 3469 -2693 3503 -2659
rect 5128 -2693 5162 -2659
rect 5528 -2693 5562 -2659
<< locali >>
rect -65 1221 2215 1244
rect -65 1187 18 1221
rect 52 1187 98 1221
rect 132 1187 178 1221
rect 212 1187 258 1221
rect 292 1187 338 1221
rect 372 1187 418 1221
rect 452 1187 498 1221
rect 532 1187 578 1221
rect 612 1187 658 1221
rect 692 1187 738 1221
rect 772 1187 818 1221
rect 852 1187 898 1221
rect 932 1187 978 1221
rect 1012 1187 1058 1221
rect 1092 1187 1138 1221
rect 1172 1187 1218 1221
rect 1252 1187 1298 1221
rect 1332 1187 1378 1221
rect 1412 1187 1458 1221
rect 1492 1187 1538 1221
rect 1572 1187 1618 1221
rect 1652 1187 1698 1221
rect 1732 1187 1778 1221
rect 1812 1187 1858 1221
rect 1892 1187 1938 1221
rect 1972 1187 2018 1221
rect 2052 1187 2098 1221
rect 2132 1187 2215 1221
rect -65 1164 2215 1187
rect 2595 1221 3975 1244
rect 2595 1187 2628 1221
rect 2662 1187 2708 1221
rect 2742 1187 2788 1221
rect 2822 1187 2868 1221
rect 2902 1187 2948 1221
rect 2982 1187 3028 1221
rect 3062 1187 3108 1221
rect 3142 1187 3188 1221
rect 3222 1187 3268 1221
rect 3302 1187 3348 1221
rect 3382 1187 3428 1221
rect 3462 1187 3508 1221
rect 3542 1187 3588 1221
rect 3622 1187 3668 1221
rect 3702 1187 3748 1221
rect 3782 1187 3828 1221
rect 3862 1187 3908 1221
rect 3942 1187 3975 1221
rect 2595 1164 3975 1187
rect 4325 1221 6005 1244
rect 4325 1187 4348 1221
rect 4382 1187 4428 1221
rect 4462 1187 4508 1221
rect 4542 1187 4588 1221
rect 4622 1187 4668 1221
rect 4702 1187 4748 1221
rect 4782 1187 4828 1221
rect 4862 1187 4908 1221
rect 4942 1187 4988 1221
rect 5022 1187 5068 1221
rect 5102 1187 5148 1221
rect 5182 1187 5228 1221
rect 5262 1187 5308 1221
rect 5342 1187 5388 1221
rect 5422 1187 5468 1221
rect 5502 1187 5548 1221
rect 5582 1187 5628 1221
rect 5662 1187 5708 1221
rect 5742 1187 5788 1221
rect 5822 1187 5868 1221
rect 5902 1187 5948 1221
rect 5982 1187 6005 1221
rect 4325 1164 6005 1187
rect 325 1094 405 1114
rect 455 1094 535 1114
rect -441 1091 535 1094
rect -441 1071 348 1091
rect -441 1037 -418 1071
rect -384 1057 348 1071
rect 382 1057 478 1091
rect 512 1057 535 1091
rect -384 1054 535 1057
rect -384 1037 -361 1054
rect -441 1014 -361 1037
rect 325 1034 405 1054
rect 455 1034 535 1054
rect 1715 1091 1795 1114
rect 1715 1057 1738 1091
rect 1772 1057 1795 1091
rect 1715 1034 1795 1057
rect -327 994 -247 1012
rect 205 994 285 1014
rect 585 994 665 1014
rect -327 991 665 994
rect -327 989 228 991
rect -327 955 -304 989
rect -270 957 228 989
rect 262 957 608 991
rect 642 957 665 991
rect -270 955 665 957
rect -327 954 665 955
rect -327 932 -247 954
rect 205 934 285 954
rect 585 934 665 954
rect 735 1001 815 1034
rect 735 967 758 1001
rect 792 967 815 1001
rect 735 921 815 967
rect 455 894 535 914
rect -669 891 535 894
rect -669 871 478 891
rect -669 837 -646 871
rect -612 857 478 871
rect 512 857 535 891
rect -612 854 535 857
rect -612 837 -589 854
rect -669 814 -589 837
rect 455 834 535 854
rect 735 887 758 921
rect 792 887 815 921
rect 735 841 815 887
rect 5 794 85 814
rect 585 794 665 814
rect -555 791 665 794
rect -555 771 28 791
rect -555 737 -532 771
rect -498 757 28 771
rect 62 757 608 791
rect 642 757 665 791
rect 735 807 758 841
rect 792 807 815 841
rect 735 784 815 807
rect 885 1001 965 1034
rect 885 967 908 1001
rect 942 967 965 1001
rect 885 921 965 967
rect 885 887 908 921
rect 942 887 965 921
rect 885 841 965 887
rect 885 807 908 841
rect 942 807 965 841
rect 885 774 965 807
rect 1035 1001 1115 1034
rect 1035 967 1058 1001
rect 1092 967 1115 1001
rect 1035 921 1115 967
rect 1035 887 1058 921
rect 1092 887 1115 921
rect 1035 841 1115 887
rect 1035 807 1058 841
rect 1092 807 1115 841
rect 1035 784 1115 807
rect 1185 1001 1265 1034
rect 1185 967 1208 1001
rect 1242 967 1265 1001
rect 1185 921 1265 967
rect 1185 887 1208 921
rect 1242 887 1265 921
rect 1185 841 1265 887
rect 1185 807 1208 841
rect 1242 807 1265 841
rect 1185 774 1265 807
rect 1335 1001 1415 1034
rect 2507 1028 2587 1048
rect 2179 1025 2587 1028
rect 1335 967 1358 1001
rect 1392 967 1415 1001
rect 1335 921 1415 967
rect 1915 991 1995 1014
rect 1915 957 1938 991
rect 1972 957 1995 991
rect 1915 934 1995 957
rect 2179 991 2530 1025
rect 2564 991 2587 1025
rect 2179 988 2587 991
rect 1335 887 1358 921
rect 1392 887 1415 921
rect 1335 841 1415 887
rect 1335 807 1358 841
rect 1392 807 1415 841
rect 2065 891 2145 914
rect 2065 857 2088 891
rect 2122 857 2145 891
rect 2065 834 2145 857
rect 1335 784 1415 807
rect 1615 791 1695 814
rect -498 754 665 757
rect -498 737 -475 754
rect -555 714 -475 737
rect 5 734 85 754
rect 585 734 665 754
rect 905 724 945 774
rect 1085 724 1165 744
rect 905 721 1165 724
rect 905 687 1108 721
rect 1142 687 1165 721
rect 905 684 1165 687
rect 905 554 945 684
rect 1085 664 1165 684
rect -25 514 945 554
rect 985 604 1065 619
rect 1205 604 1245 774
rect 1615 757 1638 791
rect 1672 757 1695 791
rect 1615 734 1695 757
rect 1455 711 1535 734
rect 1455 677 1478 711
rect 1512 694 1535 711
rect 2179 694 2219 988
rect 2507 968 2587 988
rect 2945 1001 3025 1034
rect 2945 967 2968 1001
rect 3002 967 3025 1001
rect 2945 921 3025 967
rect 2945 887 2968 921
rect 3002 887 3025 921
rect 2795 844 2875 864
rect 2595 841 2875 844
rect 2595 807 2818 841
rect 2852 807 2875 841
rect 2595 804 2875 807
rect 2795 784 2875 804
rect 2945 841 3025 887
rect 2945 807 2968 841
rect 3002 807 3025 841
rect 2945 784 3025 807
rect 3095 1001 3175 1034
rect 3095 967 3118 1001
rect 3152 967 3175 1001
rect 3095 921 3175 967
rect 3095 887 3118 921
rect 3152 887 3175 921
rect 3095 841 3175 887
rect 3095 807 3118 841
rect 3152 807 3175 841
rect 3095 774 3175 807
rect 3245 1001 3325 1034
rect 3245 967 3268 1001
rect 3302 967 3325 1001
rect 3245 921 3325 967
rect 3245 887 3268 921
rect 3302 887 3325 921
rect 3245 841 3325 887
rect 3245 807 3268 841
rect 3302 807 3325 841
rect 3245 784 3325 807
rect 3395 1001 3475 1034
rect 3395 967 3418 1001
rect 3452 967 3475 1001
rect 3395 921 3475 967
rect 3395 887 3418 921
rect 3452 887 3475 921
rect 3395 841 3475 887
rect 3395 807 3418 841
rect 3452 807 3475 841
rect 3395 774 3475 807
rect 3545 1001 3625 1034
rect 3545 967 3568 1001
rect 3602 967 3625 1001
rect 3983 1025 4063 1048
rect 3983 991 4006 1025
rect 4040 1008 4063 1025
rect 4040 994 4345 1008
rect 4675 994 4755 1014
rect 4040 991 4755 994
rect 3983 968 4698 991
rect 3545 921 3625 967
rect 4305 957 4698 968
rect 4732 957 4755 991
rect 4305 954 4755 957
rect 4675 934 4755 954
rect 4825 1001 4905 1034
rect 4825 967 4848 1001
rect 4882 967 4905 1001
rect 3545 887 3568 921
rect 3602 887 3625 921
rect 3545 841 3625 887
rect 3983 910 4063 933
rect 4825 921 4905 967
rect 3983 876 4006 910
rect 4040 876 4063 910
rect 3545 807 3568 841
rect 3602 807 3625 841
rect 3545 784 3625 807
rect 3695 844 3775 864
rect 3825 844 3905 864
rect 3983 853 4063 876
rect 4245 891 4325 914
rect 4245 857 4268 891
rect 4302 874 4325 891
rect 4675 874 4755 894
rect 4302 871 4755 874
rect 4302 857 4698 871
rect 3695 841 3905 844
rect 3695 807 3718 841
rect 3752 807 3848 841
rect 3882 807 3905 841
rect 3695 804 3905 807
rect 3695 784 3775 804
rect 3825 784 3905 804
rect 4004 798 4044 853
rect 4245 837 4698 857
rect 4732 837 4755 871
rect 4245 834 4755 837
rect 4675 814 4755 834
rect 4825 887 4848 921
rect 4882 887 4905 921
rect 4825 841 4905 887
rect 4825 807 4848 841
rect 4882 807 4905 841
rect 4004 774 4231 798
rect 4545 774 4625 794
rect 4825 784 4905 807
rect 4975 1001 5055 1034
rect 4975 967 4998 1001
rect 5032 967 5055 1001
rect 4975 921 5055 967
rect 4975 887 4998 921
rect 5032 887 5055 921
rect 4975 841 5055 887
rect 4975 807 4998 841
rect 5032 807 5055 841
rect 4975 774 5055 807
rect 5125 1001 5205 1034
rect 5125 967 5148 1001
rect 5182 967 5205 1001
rect 5125 921 5205 967
rect 5125 887 5148 921
rect 5182 887 5205 921
rect 5125 841 5205 887
rect 5125 807 5148 841
rect 5182 807 5205 841
rect 5125 784 5205 807
rect 5275 1001 5355 1034
rect 5275 967 5298 1001
rect 5332 967 5355 1001
rect 5275 921 5355 967
rect 5275 887 5298 921
rect 5332 887 5355 921
rect 5275 841 5355 887
rect 5275 807 5298 841
rect 5332 807 5355 841
rect 5275 774 5355 807
rect 5425 1001 5505 1034
rect 5425 967 5448 1001
rect 5482 967 5505 1001
rect 5425 921 5505 967
rect 5805 991 5885 1014
rect 5805 957 5828 991
rect 5862 957 5885 991
rect 5805 934 5885 957
rect 5425 887 5448 921
rect 5482 887 5505 921
rect 5425 841 5505 887
rect 5425 807 5448 841
rect 5482 807 5505 841
rect 5655 871 5735 894
rect 5655 837 5678 871
rect 5712 837 5735 871
rect 5655 814 5735 837
rect 5425 784 5505 807
rect 1512 677 2219 694
rect 1455 654 2219 677
rect 3115 724 3155 774
rect 3295 724 3375 744
rect 3115 721 3375 724
rect 3115 687 3318 721
rect 3352 687 3375 721
rect 3115 684 3375 687
rect 2215 604 2295 620
rect 2665 604 2745 624
rect 985 597 2295 604
rect 985 596 2238 597
rect 985 562 1008 596
rect 1042 564 2238 596
rect 1042 562 1065 564
rect 985 539 1065 562
rect -25 474 15 514
rect 575 474 615 514
rect 905 474 945 514
rect 1205 474 1245 564
rect 1535 474 1575 564
rect 2135 474 2175 564
rect 2215 563 2238 564
rect 2272 563 2295 597
rect 2215 540 2295 563
rect 2541 601 2745 604
rect 2541 567 2688 601
rect 2722 567 2745 601
rect 2541 564 2745 567
rect -45 441 35 474
rect -45 407 -22 441
rect 12 407 35 441
rect -45 361 35 407
rect -45 327 -22 361
rect 12 327 35 361
rect -45 281 35 327
rect -45 247 -22 281
rect 12 247 35 281
rect -45 224 35 247
rect 255 441 335 474
rect 255 407 278 441
rect 312 407 335 441
rect 255 361 335 407
rect 255 327 278 361
rect 312 327 335 361
rect 255 281 335 327
rect 255 247 278 281
rect 312 247 335 281
rect 255 224 335 247
rect 555 441 635 474
rect 555 407 578 441
rect 612 407 635 441
rect 555 361 635 407
rect 555 327 578 361
rect 612 327 635 361
rect 555 281 635 327
rect 555 247 578 281
rect 612 247 635 281
rect 555 224 635 247
rect 735 441 815 474
rect 735 407 758 441
rect 792 407 815 441
rect 735 361 815 407
rect 735 327 758 361
rect 792 327 815 361
rect 735 281 815 327
rect 735 247 758 281
rect 792 247 815 281
rect 735 224 815 247
rect 885 441 965 474
rect 885 407 908 441
rect 942 407 965 441
rect 885 361 965 407
rect 885 327 908 361
rect 942 327 965 361
rect 885 281 965 327
rect 885 247 908 281
rect 942 247 965 281
rect 885 224 965 247
rect 1035 441 1115 474
rect 1035 407 1058 441
rect 1092 407 1115 441
rect 1035 361 1115 407
rect 1035 327 1058 361
rect 1092 327 1115 361
rect 1035 281 1115 327
rect 1035 247 1058 281
rect 1092 247 1115 281
rect 1035 224 1115 247
rect 1185 441 1265 474
rect 1185 407 1208 441
rect 1242 407 1265 441
rect 1185 361 1265 407
rect 1185 327 1208 361
rect 1242 327 1265 361
rect 1185 281 1265 327
rect 1185 247 1208 281
rect 1242 247 1265 281
rect 1185 224 1265 247
rect 1335 441 1415 474
rect 1335 407 1358 441
rect 1392 407 1415 441
rect 1335 361 1415 407
rect 1335 327 1358 361
rect 1392 327 1415 361
rect 1335 281 1415 327
rect 1335 247 1358 281
rect 1392 247 1415 281
rect 1335 224 1415 247
rect 1515 441 1595 474
rect 1515 407 1538 441
rect 1572 407 1595 441
rect 1515 361 1595 407
rect 1515 327 1538 361
rect 1572 327 1595 361
rect 1515 281 1595 327
rect 1515 247 1538 281
rect 1572 247 1595 281
rect 1515 224 1595 247
rect 1815 441 1895 474
rect 1815 407 1838 441
rect 1872 407 1895 441
rect 1815 361 1895 407
rect 1815 327 1838 361
rect 1872 327 1895 361
rect 1815 281 1895 327
rect 1815 247 1838 281
rect 1872 247 1895 281
rect 1815 224 1895 247
rect 2115 441 2195 474
rect 2115 407 2138 441
rect 2172 407 2195 441
rect 2115 361 2195 407
rect 2115 327 2138 361
rect 2172 327 2195 361
rect 2115 281 2195 327
rect 2229 361 2309 381
rect 2541 361 2581 564
rect 2665 544 2745 564
rect 3115 554 3155 684
rect 3295 664 3375 684
rect 2785 514 3155 554
rect 3195 604 3275 619
rect 3415 604 3455 774
rect 4004 771 4625 774
rect 4004 758 4568 771
rect 3695 724 3775 744
rect 4191 737 4568 758
rect 4602 737 4625 771
rect 4191 734 4625 737
rect 3695 721 4157 724
rect 3695 687 3718 721
rect 3752 687 4157 721
rect 4545 714 4625 734
rect 4995 724 5035 774
rect 5175 724 5255 744
rect 4995 721 5255 724
rect 3695 684 4157 687
rect 3695 664 3775 684
rect 4117 674 4157 684
rect 4395 674 4475 694
rect 4117 671 4475 674
rect 4117 637 4418 671
rect 4452 637 4475 671
rect 4117 634 4475 637
rect 4395 614 4475 634
rect 4995 687 5198 721
rect 5232 687 5255 721
rect 4995 684 5255 687
rect 3195 596 3455 604
rect 3195 562 3218 596
rect 3252 564 3455 596
rect 3252 562 3275 564
rect 3195 539 3275 562
rect 3415 554 3455 564
rect 3983 571 4063 594
rect 3983 554 4006 571
rect 3415 537 4006 554
rect 4040 537 4063 571
rect 4995 554 5035 684
rect 5175 664 5255 684
rect 3415 514 4063 537
rect 4365 514 5035 554
rect 5075 604 5155 619
rect 5295 604 5335 774
rect 5575 724 5655 744
rect 5575 721 6197 724
rect 5575 687 5598 721
rect 5632 687 6197 721
rect 5575 684 6197 687
rect 5575 664 5655 684
rect 6008 604 6088 623
rect 5075 600 6088 604
rect 5075 596 6031 600
rect 5075 562 5098 596
rect 5132 566 6031 596
rect 6065 566 6088 600
rect 5132 564 6088 566
rect 5132 562 5155 564
rect 5075 539 5155 562
rect 2785 474 2825 514
rect 3115 474 3155 514
rect 2229 359 2581 361
rect 2229 325 2252 359
rect 2286 325 2581 359
rect 2229 321 2581 325
rect 2615 441 2695 474
rect 2615 407 2638 441
rect 2672 407 2695 441
rect 2615 361 2695 407
rect 2615 327 2638 361
rect 2672 327 2695 361
rect 2229 301 2309 321
rect 2115 247 2138 281
rect 2172 247 2195 281
rect 2115 224 2195 247
rect 2615 281 2695 327
rect 2615 247 2638 281
rect 2672 247 2695 281
rect 2615 224 2695 247
rect 2765 441 2845 474
rect 2765 407 2788 441
rect 2822 407 2845 441
rect 2765 361 2845 407
rect 2765 327 2788 361
rect 2822 327 2845 361
rect 2765 281 2845 327
rect 2765 247 2788 281
rect 2822 247 2845 281
rect 2765 224 2845 247
rect 2945 441 3025 474
rect 2945 407 2968 441
rect 3002 407 3025 441
rect 2945 361 3025 407
rect 2945 327 2968 361
rect 3002 327 3025 361
rect 2945 281 3025 327
rect 2945 247 2968 281
rect 3002 247 3025 281
rect 2945 224 3025 247
rect 3095 441 3175 474
rect 3095 407 3118 441
rect 3152 407 3175 441
rect 3095 361 3175 407
rect 3095 327 3118 361
rect 3152 327 3175 361
rect 3095 281 3175 327
rect 3095 247 3118 281
rect 3152 247 3175 281
rect 3095 224 3175 247
rect 3245 441 3325 474
rect 3245 407 3268 441
rect 3302 407 3325 441
rect 3245 361 3325 407
rect 3245 327 3268 361
rect 3302 327 3325 361
rect 3245 281 3325 327
rect 3245 247 3268 281
rect 3302 247 3325 281
rect 3245 224 3325 247
rect 3395 441 3475 514
rect 3745 474 3785 514
rect 4365 474 4405 514
rect 4665 474 4705 514
rect 4996 474 5035 514
rect 5295 474 5335 564
rect 5625 474 5665 564
rect 6008 543 6088 564
rect 3395 407 3418 441
rect 3452 407 3475 441
rect 3395 361 3475 407
rect 3395 327 3418 361
rect 3452 327 3475 361
rect 3395 281 3475 327
rect 3395 247 3418 281
rect 3452 247 3475 281
rect 3395 224 3475 247
rect 3545 441 3625 474
rect 3545 407 3568 441
rect 3602 407 3625 441
rect 3545 361 3625 407
rect 3545 327 3568 361
rect 3602 327 3625 361
rect 3545 281 3625 327
rect 3545 247 3568 281
rect 3602 247 3625 281
rect 3545 224 3625 247
rect 3725 441 3805 474
rect 3725 407 3748 441
rect 3782 407 3805 441
rect 3725 361 3805 407
rect 3725 327 3748 361
rect 3782 327 3805 361
rect 3725 281 3805 327
rect 3725 247 3748 281
rect 3782 247 3805 281
rect 3725 224 3805 247
rect 3875 441 3955 474
rect 3875 407 3898 441
rect 3932 407 3955 441
rect 3875 361 3955 407
rect 3875 327 3898 361
rect 3932 327 3955 361
rect 3875 281 3955 327
rect 3875 247 3898 281
rect 3932 247 3955 281
rect 3875 224 3955 247
rect 4345 441 4425 474
rect 4345 407 4368 441
rect 4402 407 4425 441
rect 4345 361 4425 407
rect 4345 327 4368 361
rect 4402 327 4425 361
rect 4345 281 4425 327
rect 4345 247 4368 281
rect 4402 247 4425 281
rect 4345 224 4425 247
rect 4495 441 4575 474
rect 4495 407 4518 441
rect 4552 407 4575 441
rect 4495 361 4575 407
rect 4495 327 4518 361
rect 4552 327 4575 361
rect 4495 281 4575 327
rect 4495 247 4518 281
rect 4552 247 4575 281
rect 4495 224 4575 247
rect 4645 441 4725 474
rect 4645 407 4668 441
rect 4702 407 4725 441
rect 4645 361 4725 407
rect 4645 327 4668 361
rect 4702 327 4725 361
rect 4645 281 4725 327
rect 4645 247 4668 281
rect 4702 247 4725 281
rect 4645 224 4725 247
rect 4825 441 4905 474
rect 4825 407 4848 441
rect 4882 407 4905 441
rect 4825 361 4905 407
rect 4825 327 4848 361
rect 4882 327 4905 361
rect 4825 281 4905 327
rect 4825 247 4848 281
rect 4882 247 4905 281
rect 4825 224 4905 247
rect 4975 441 5055 474
rect 4975 407 4998 441
rect 5032 407 5055 441
rect 4975 361 5055 407
rect 4975 327 4998 361
rect 5032 327 5055 361
rect 4975 281 5055 327
rect 4975 247 4998 281
rect 5032 247 5055 281
rect 4975 224 5055 247
rect 5125 441 5205 474
rect 5125 407 5148 441
rect 5182 407 5205 441
rect 5125 361 5205 407
rect 5125 327 5148 361
rect 5182 327 5205 361
rect 5125 281 5205 327
rect 5125 247 5148 281
rect 5182 247 5205 281
rect 5125 224 5205 247
rect 5275 441 5355 474
rect 5275 407 5298 441
rect 5332 407 5355 441
rect 5275 361 5355 407
rect 5275 327 5298 361
rect 5332 327 5355 361
rect 5275 281 5355 327
rect 5275 247 5298 281
rect 5332 247 5355 281
rect 5275 224 5355 247
rect 5425 441 5505 474
rect 5425 407 5448 441
rect 5482 407 5505 441
rect 5425 361 5505 407
rect 5425 327 5448 361
rect 5482 327 5505 361
rect 5425 281 5505 327
rect 5425 247 5448 281
rect 5482 247 5505 281
rect 5425 224 5505 247
rect 5605 441 5685 474
rect 5605 407 5628 441
rect 5662 407 5685 441
rect 5605 361 5685 407
rect 5605 327 5628 361
rect 5662 327 5685 361
rect 5605 281 5685 327
rect 5605 247 5628 281
rect 5662 247 5685 281
rect 5605 224 5685 247
rect 5905 441 5985 474
rect 5905 407 5928 441
rect 5962 407 5985 441
rect 5905 361 5985 407
rect 5905 327 5928 361
rect 5962 327 5985 361
rect 5905 281 5985 327
rect 5905 247 5928 281
rect 5962 247 5985 281
rect 5905 224 5985 247
rect 367 164 447 184
rect 835 164 915 184
rect 1235 164 1315 184
rect 3045 164 3125 184
rect 3445 164 3525 184
rect 4333 164 4413 184
rect 4925 164 5005 184
rect 5325 164 5405 184
rect -65 161 3525 164
rect -65 127 390 161
rect 424 127 858 161
rect 892 127 1258 161
rect 1292 127 3068 161
rect 3102 127 3468 161
rect 3502 127 3525 161
rect -65 124 3525 127
rect 4325 161 5405 164
rect 4325 127 4356 161
rect 4390 127 4948 161
rect 4982 127 5348 161
rect 5382 127 5405 161
rect 4325 124 5405 127
rect 367 104 447 124
rect 835 104 915 124
rect 1235 104 1315 124
rect 3045 104 3125 124
rect 3445 104 3525 124
rect 4333 104 4413 124
rect 4925 104 5005 124
rect 5325 104 5405 124
rect -213 41 2215 64
rect -213 7 -190 41
rect -156 7 18 41
rect 52 7 98 41
rect 132 7 178 41
rect 212 7 258 41
rect 292 7 338 41
rect 372 7 418 41
rect 452 7 498 41
rect 532 7 578 41
rect 612 7 658 41
rect 692 7 738 41
rect 772 7 818 41
rect 852 7 898 41
rect 932 7 978 41
rect 1012 7 1058 41
rect 1092 7 1138 41
rect 1172 7 1218 41
rect 1252 7 1298 41
rect 1332 7 1378 41
rect 1412 7 1458 41
rect 1492 7 1538 41
rect 1572 7 1618 41
rect 1652 7 1698 41
rect 1732 7 1778 41
rect 1812 7 1858 41
rect 1892 7 1938 41
rect 1972 7 2018 41
rect 2052 7 2098 41
rect 2132 7 2215 41
rect -213 -16 2215 7
rect 2595 41 3975 64
rect 2595 7 2628 41
rect 2662 7 2708 41
rect 2742 7 2788 41
rect 2822 7 2868 41
rect 2902 7 2948 41
rect 2982 7 3028 41
rect 3062 7 3108 41
rect 3142 7 3188 41
rect 3222 7 3268 41
rect 3302 7 3348 41
rect 3382 7 3428 41
rect 3462 7 3508 41
rect 3542 7 3588 41
rect 3622 7 3668 41
rect 3702 7 3748 41
rect 3782 7 3828 41
rect 3862 7 3908 41
rect 3942 7 3975 41
rect 2595 -16 3975 7
rect 4325 41 6005 64
rect 4325 7 4348 41
rect 4382 7 4428 41
rect 4462 7 4508 41
rect 4542 7 4588 41
rect 4622 7 4668 41
rect 4702 7 4748 41
rect 4782 7 4828 41
rect 4862 7 4908 41
rect 4942 7 4988 41
rect 5022 7 5068 41
rect 5102 7 5148 41
rect 5182 7 5228 41
rect 5262 7 5308 41
rect 5342 7 5388 41
rect 5422 7 5468 41
rect 5502 7 5548 41
rect 5582 7 5628 41
rect 5662 7 5708 41
rect 5742 7 5788 41
rect 5822 7 5868 41
rect 5902 7 5948 41
rect 5982 7 6005 41
rect 4325 -16 6005 7
rect 367 -76 447 -56
rect 835 -76 915 -56
rect 1235 -76 1315 -56
rect 3045 -76 3125 -56
rect 3445 -76 3525 -56
rect 4333 -76 4413 -56
rect 4925 -76 5005 -56
rect 5325 -76 5405 -56
rect -65 -79 3525 -76
rect -65 -113 390 -79
rect 424 -113 858 -79
rect 892 -113 1258 -79
rect 1292 -113 3068 -79
rect 3102 -113 3468 -79
rect 3502 -113 3525 -79
rect -65 -116 3525 -113
rect 4325 -79 5405 -76
rect 4325 -113 4356 -79
rect 4390 -113 4948 -79
rect 4982 -113 5348 -79
rect 5382 -113 5405 -79
rect 4325 -116 5405 -113
rect 367 -136 447 -116
rect 835 -136 915 -116
rect 1235 -136 1315 -116
rect 3045 -136 3125 -116
rect 3445 -136 3525 -116
rect 4333 -136 4413 -116
rect 4925 -136 5005 -116
rect 5325 -136 5405 -116
rect -45 -199 35 -176
rect -45 -233 -22 -199
rect 12 -233 35 -199
rect -45 -279 35 -233
rect -45 -313 -22 -279
rect 12 -313 35 -279
rect -45 -359 35 -313
rect -45 -393 -22 -359
rect 12 -393 35 -359
rect -45 -426 35 -393
rect 255 -199 335 -176
rect 255 -233 278 -199
rect 312 -233 335 -199
rect 255 -279 335 -233
rect 255 -313 278 -279
rect 312 -313 335 -279
rect 255 -359 335 -313
rect 255 -393 278 -359
rect 312 -393 335 -359
rect 255 -426 335 -393
rect 555 -199 635 -176
rect 555 -233 578 -199
rect 612 -233 635 -199
rect 555 -279 635 -233
rect 555 -313 578 -279
rect 612 -313 635 -279
rect 555 -359 635 -313
rect 555 -393 578 -359
rect 612 -393 635 -359
rect 555 -426 635 -393
rect 735 -199 815 -176
rect 735 -233 758 -199
rect 792 -233 815 -199
rect 735 -279 815 -233
rect 735 -313 758 -279
rect 792 -313 815 -279
rect 735 -359 815 -313
rect 735 -393 758 -359
rect 792 -393 815 -359
rect 735 -426 815 -393
rect 885 -199 965 -176
rect 885 -233 908 -199
rect 942 -233 965 -199
rect 885 -279 965 -233
rect 885 -313 908 -279
rect 942 -313 965 -279
rect 885 -359 965 -313
rect 885 -393 908 -359
rect 942 -393 965 -359
rect 885 -426 965 -393
rect 1035 -199 1115 -176
rect 1035 -233 1058 -199
rect 1092 -233 1115 -199
rect 1035 -279 1115 -233
rect 1035 -313 1058 -279
rect 1092 -313 1115 -279
rect 1035 -359 1115 -313
rect 1035 -393 1058 -359
rect 1092 -393 1115 -359
rect 1035 -426 1115 -393
rect 1185 -199 1265 -176
rect 1185 -233 1208 -199
rect 1242 -233 1265 -199
rect 1185 -279 1265 -233
rect 1185 -313 1208 -279
rect 1242 -313 1265 -279
rect 1185 -359 1265 -313
rect 1185 -393 1208 -359
rect 1242 -393 1265 -359
rect 1185 -426 1265 -393
rect 1335 -199 1415 -176
rect 1335 -233 1358 -199
rect 1392 -233 1415 -199
rect 1335 -279 1415 -233
rect 1335 -313 1358 -279
rect 1392 -313 1415 -279
rect 1335 -359 1415 -313
rect 1335 -393 1358 -359
rect 1392 -393 1415 -359
rect 1335 -426 1415 -393
rect 1515 -199 1595 -176
rect 1515 -233 1538 -199
rect 1572 -233 1595 -199
rect 1515 -279 1595 -233
rect 1515 -313 1538 -279
rect 1572 -313 1595 -279
rect 1515 -359 1595 -313
rect 1515 -393 1538 -359
rect 1572 -393 1595 -359
rect 1515 -426 1595 -393
rect 1815 -199 1895 -176
rect 1815 -233 1838 -199
rect 1872 -233 1895 -199
rect 1815 -279 1895 -233
rect 1815 -313 1838 -279
rect 1872 -313 1895 -279
rect 1815 -359 1895 -313
rect 1815 -393 1838 -359
rect 1872 -393 1895 -359
rect 1815 -426 1895 -393
rect 2115 -199 2195 -176
rect 2115 -233 2138 -199
rect 2172 -233 2195 -199
rect 2115 -279 2195 -233
rect 2615 -199 2695 -176
rect 2615 -233 2638 -199
rect 2672 -233 2695 -199
rect 2115 -313 2138 -279
rect 2172 -313 2195 -279
rect 2115 -359 2195 -313
rect 2229 -276 2309 -257
rect 2229 -279 2581 -276
rect 2229 -313 2252 -279
rect 2286 -313 2581 -279
rect 2229 -316 2581 -313
rect 2229 -337 2309 -316
rect 2115 -393 2138 -359
rect 2172 -393 2195 -359
rect 2115 -426 2195 -393
rect -25 -466 15 -426
rect 575 -466 615 -426
rect 905 -466 945 -426
rect -25 -506 945 -466
rect 905 -636 945 -506
rect 985 -514 1065 -491
rect 985 -548 1008 -514
rect 1042 -516 1065 -514
rect 1205 -516 1245 -426
rect 1535 -516 1575 -426
rect 2135 -516 2175 -426
rect 2541 -516 2581 -316
rect 2615 -279 2695 -233
rect 2615 -313 2638 -279
rect 2672 -313 2695 -279
rect 2615 -359 2695 -313
rect 2615 -393 2638 -359
rect 2672 -393 2695 -359
rect 2615 -426 2695 -393
rect 2765 -199 2845 -176
rect 2765 -233 2788 -199
rect 2822 -233 2845 -199
rect 2765 -279 2845 -233
rect 2765 -313 2788 -279
rect 2822 -313 2845 -279
rect 2765 -359 2845 -313
rect 2765 -393 2788 -359
rect 2822 -393 2845 -359
rect 2765 -426 2845 -393
rect 2945 -199 3025 -176
rect 2945 -233 2968 -199
rect 3002 -233 3025 -199
rect 2945 -279 3025 -233
rect 2945 -313 2968 -279
rect 3002 -313 3025 -279
rect 2945 -359 3025 -313
rect 2945 -393 2968 -359
rect 3002 -393 3025 -359
rect 2945 -426 3025 -393
rect 3095 -199 3175 -176
rect 3095 -233 3118 -199
rect 3152 -233 3175 -199
rect 3095 -279 3175 -233
rect 3095 -313 3118 -279
rect 3152 -313 3175 -279
rect 3095 -359 3175 -313
rect 3095 -393 3118 -359
rect 3152 -393 3175 -359
rect 3095 -426 3175 -393
rect 3245 -199 3325 -176
rect 3245 -233 3268 -199
rect 3302 -233 3325 -199
rect 3245 -279 3325 -233
rect 3245 -313 3268 -279
rect 3302 -313 3325 -279
rect 3245 -359 3325 -313
rect 3245 -393 3268 -359
rect 3302 -393 3325 -359
rect 3245 -426 3325 -393
rect 3395 -199 3475 -176
rect 3395 -233 3418 -199
rect 3452 -233 3475 -199
rect 3395 -279 3475 -233
rect 3395 -313 3418 -279
rect 3452 -313 3475 -279
rect 3395 -359 3475 -313
rect 3395 -393 3418 -359
rect 3452 -393 3475 -359
rect 2785 -466 2825 -426
rect 3115 -466 3155 -426
rect 3395 -466 3475 -393
rect 3545 -199 3625 -176
rect 3545 -233 3568 -199
rect 3602 -233 3625 -199
rect 3545 -279 3625 -233
rect 3545 -313 3568 -279
rect 3602 -313 3625 -279
rect 3545 -359 3625 -313
rect 3545 -393 3568 -359
rect 3602 -393 3625 -359
rect 3545 -426 3625 -393
rect 3725 -199 3805 -176
rect 3725 -233 3748 -199
rect 3782 -233 3805 -199
rect 3725 -279 3805 -233
rect 3725 -313 3748 -279
rect 3782 -313 3805 -279
rect 3725 -359 3805 -313
rect 3725 -393 3748 -359
rect 3782 -393 3805 -359
rect 3725 -426 3805 -393
rect 3875 -199 3955 -176
rect 3875 -233 3898 -199
rect 3932 -233 3955 -199
rect 3875 -279 3955 -233
rect 3875 -313 3898 -279
rect 3932 -313 3955 -279
rect 3875 -359 3955 -313
rect 3875 -393 3898 -359
rect 3932 -393 3955 -359
rect 3875 -426 3955 -393
rect 4345 -199 4425 -176
rect 4345 -233 4368 -199
rect 4402 -233 4425 -199
rect 4345 -279 4425 -233
rect 4345 -313 4368 -279
rect 4402 -313 4425 -279
rect 4345 -359 4425 -313
rect 4345 -393 4368 -359
rect 4402 -393 4425 -359
rect 4345 -426 4425 -393
rect 4495 -199 4575 -176
rect 4495 -233 4518 -199
rect 4552 -233 4575 -199
rect 4495 -279 4575 -233
rect 4495 -313 4518 -279
rect 4552 -313 4575 -279
rect 4495 -359 4575 -313
rect 4495 -393 4518 -359
rect 4552 -393 4575 -359
rect 4495 -426 4575 -393
rect 4645 -199 4725 -176
rect 4645 -233 4668 -199
rect 4702 -233 4725 -199
rect 4645 -279 4725 -233
rect 4645 -313 4668 -279
rect 4702 -313 4725 -279
rect 4645 -359 4725 -313
rect 4645 -393 4668 -359
rect 4702 -393 4725 -359
rect 4645 -426 4725 -393
rect 4825 -199 4905 -176
rect 4825 -233 4848 -199
rect 4882 -233 4905 -199
rect 4825 -279 4905 -233
rect 4825 -313 4848 -279
rect 4882 -313 4905 -279
rect 4825 -359 4905 -313
rect 4825 -393 4848 -359
rect 4882 -393 4905 -359
rect 4825 -426 4905 -393
rect 4975 -199 5055 -176
rect 4975 -233 4998 -199
rect 5032 -233 5055 -199
rect 4975 -279 5055 -233
rect 4975 -313 4998 -279
rect 5032 -313 5055 -279
rect 4975 -359 5055 -313
rect 4975 -393 4998 -359
rect 5032 -393 5055 -359
rect 4975 -426 5055 -393
rect 5125 -199 5205 -176
rect 5125 -233 5148 -199
rect 5182 -233 5205 -199
rect 5125 -279 5205 -233
rect 5125 -313 5148 -279
rect 5182 -313 5205 -279
rect 5125 -359 5205 -313
rect 5125 -393 5148 -359
rect 5182 -393 5205 -359
rect 5125 -426 5205 -393
rect 5275 -199 5355 -176
rect 5275 -233 5298 -199
rect 5332 -233 5355 -199
rect 5275 -279 5355 -233
rect 5275 -313 5298 -279
rect 5332 -313 5355 -279
rect 5275 -359 5355 -313
rect 5275 -393 5298 -359
rect 5332 -393 5355 -359
rect 5275 -426 5355 -393
rect 5425 -199 5505 -176
rect 5425 -233 5448 -199
rect 5482 -233 5505 -199
rect 5425 -279 5505 -233
rect 5425 -313 5448 -279
rect 5482 -313 5505 -279
rect 5425 -359 5505 -313
rect 5425 -393 5448 -359
rect 5482 -393 5505 -359
rect 5425 -426 5505 -393
rect 5605 -199 5685 -176
rect 5605 -233 5628 -199
rect 5662 -233 5685 -199
rect 5605 -279 5685 -233
rect 5605 -313 5628 -279
rect 5662 -313 5685 -279
rect 5605 -359 5685 -313
rect 5605 -393 5628 -359
rect 5662 -393 5685 -359
rect 5605 -426 5685 -393
rect 5905 -199 5985 -176
rect 5905 -233 5928 -199
rect 5962 -233 5985 -199
rect 5905 -279 5985 -233
rect 5905 -313 5928 -279
rect 5962 -313 5985 -279
rect 5905 -359 5985 -313
rect 5905 -393 5928 -359
rect 5962 -393 5985 -359
rect 5905 -426 5985 -393
rect 3745 -466 3785 -426
rect 3983 -466 4063 -446
rect 2665 -516 2745 -496
rect 2785 -506 3155 -466
rect 3415 -469 4063 -466
rect 1042 -548 2394 -516
rect 985 -556 2394 -548
rect 2541 -519 2745 -516
rect 2541 -553 2688 -519
rect 2722 -553 2745 -519
rect 2541 -556 2745 -553
rect 985 -571 1065 -556
rect 1085 -636 1165 -616
rect 905 -639 1165 -636
rect -1011 -689 -931 -666
rect 905 -673 1108 -639
rect 1142 -673 1165 -639
rect 905 -676 1165 -673
rect -1011 -723 -988 -689
rect -954 -706 -931 -689
rect 5 -706 85 -686
rect 585 -706 665 -686
rect -954 -709 665 -706
rect -954 -723 28 -709
rect -1011 -743 28 -723
rect 62 -743 608 -709
rect 642 -743 665 -709
rect 905 -726 945 -676
rect 1085 -696 1165 -676
rect 1205 -726 1245 -556
rect 1455 -629 2295 -606
rect 1455 -663 1478 -629
rect 1512 -646 2238 -629
rect 1512 -663 1535 -646
rect 1455 -686 1535 -663
rect 2215 -663 2238 -646
rect 2272 -663 2295 -629
rect 2215 -686 2295 -663
rect 1615 -709 1695 -686
rect -1011 -746 665 -743
rect 5 -766 85 -746
rect 585 -766 665 -746
rect 735 -759 815 -736
rect -1125 -806 -1045 -785
rect 455 -806 535 -786
rect -1125 -808 535 -806
rect -1125 -842 -1102 -808
rect -1068 -809 535 -808
rect -1068 -842 478 -809
rect -1125 -843 478 -842
rect 512 -843 535 -809
rect -1125 -846 535 -843
rect -1125 -865 -1045 -846
rect 455 -866 535 -846
rect 735 -793 758 -759
rect 792 -793 815 -759
rect 735 -839 815 -793
rect 735 -873 758 -839
rect 792 -873 815 -839
rect -783 -906 -703 -892
rect 205 -906 285 -886
rect 585 -906 665 -886
rect -783 -909 665 -906
rect -783 -915 228 -909
rect -783 -949 -760 -915
rect -726 -943 228 -915
rect 262 -943 608 -909
rect 642 -943 665 -909
rect -726 -946 665 -943
rect -726 -949 -703 -946
rect -783 -972 -703 -949
rect 205 -966 285 -946
rect 585 -966 665 -946
rect 735 -919 815 -873
rect 735 -953 758 -919
rect 792 -953 815 -919
rect 735 -986 815 -953
rect 885 -759 965 -726
rect 885 -793 908 -759
rect 942 -793 965 -759
rect 885 -839 965 -793
rect 885 -873 908 -839
rect 942 -873 965 -839
rect 885 -919 965 -873
rect 885 -953 908 -919
rect 942 -953 965 -919
rect 885 -986 965 -953
rect 1035 -759 1115 -736
rect 1035 -793 1058 -759
rect 1092 -793 1115 -759
rect 1035 -839 1115 -793
rect 1035 -873 1058 -839
rect 1092 -873 1115 -839
rect 1035 -919 1115 -873
rect 1035 -953 1058 -919
rect 1092 -953 1115 -919
rect 1035 -986 1115 -953
rect 1185 -759 1265 -726
rect 1185 -793 1208 -759
rect 1242 -793 1265 -759
rect 1185 -839 1265 -793
rect 1185 -873 1208 -839
rect 1242 -873 1265 -839
rect 1185 -919 1265 -873
rect 1185 -953 1208 -919
rect 1242 -953 1265 -919
rect 1185 -986 1265 -953
rect 1335 -759 1415 -736
rect 1335 -793 1358 -759
rect 1392 -793 1415 -759
rect 1615 -743 1638 -709
rect 1672 -743 1695 -709
rect 1615 -766 1695 -743
rect 1335 -839 1415 -793
rect 1335 -873 1358 -839
rect 1392 -873 1415 -839
rect 2065 -809 2145 -786
rect 2065 -843 2088 -809
rect 2122 -843 2145 -809
rect 2065 -866 2145 -843
rect 1335 -919 1415 -873
rect 1335 -953 1358 -919
rect 1392 -953 1415 -919
rect 1335 -986 1415 -953
rect 1915 -909 1995 -886
rect 1915 -943 1938 -909
rect 1972 -943 1995 -909
rect 1915 -966 1995 -943
rect 2354 -906 2394 -556
rect 2665 -576 2745 -556
rect 3115 -636 3155 -506
rect 3195 -514 3275 -491
rect 3195 -548 3218 -514
rect 3252 -516 3275 -514
rect 3415 -503 4006 -469
rect 4040 -503 4063 -469
rect 3415 -506 4063 -503
rect 4365 -466 4405 -426
rect 4665 -466 4705 -426
rect 4996 -466 5035 -426
rect 4365 -506 5035 -466
rect 3415 -516 3455 -506
rect 3252 -548 3455 -516
rect 3983 -526 4063 -506
rect 3195 -556 3455 -548
rect 3195 -571 3275 -556
rect 3295 -636 3375 -616
rect 3115 -639 3375 -636
rect 3115 -673 3318 -639
rect 3352 -673 3375 -639
rect 3115 -676 3375 -673
rect 3115 -726 3155 -676
rect 3295 -696 3375 -676
rect 3415 -726 3455 -556
rect 4395 -586 4475 -566
rect 4104 -589 4475 -586
rect 3695 -636 3775 -616
rect 4104 -623 4418 -589
rect 4452 -623 4475 -589
rect 4104 -626 4475 -623
rect 4104 -636 4144 -626
rect 3695 -639 4144 -636
rect 3695 -673 3718 -639
rect 3752 -673 4144 -639
rect 4395 -646 4475 -626
rect 4995 -636 5035 -506
rect 5075 -514 5155 -491
rect 5075 -548 5098 -514
rect 5132 -516 5155 -514
rect 5295 -516 5335 -426
rect 5625 -516 5665 -426
rect 6008 -516 6088 -496
rect 5132 -519 6088 -516
rect 5132 -548 6031 -519
rect 5075 -553 6031 -548
rect 6065 -553 6088 -519
rect 5075 -556 6088 -553
rect 5075 -571 5155 -556
rect 5175 -636 5255 -616
rect 4995 -639 5255 -636
rect 3695 -676 4144 -673
rect 3695 -696 3775 -676
rect 4245 -686 4325 -666
rect 4545 -686 4625 -666
rect 4245 -689 4625 -686
rect 4245 -723 4268 -689
rect 4302 -723 4568 -689
rect 4602 -723 4625 -689
rect 4245 -726 4625 -723
rect 4995 -673 5198 -639
rect 5232 -673 5255 -639
rect 4995 -676 5255 -673
rect 4995 -726 5035 -676
rect 5175 -696 5255 -676
rect 5295 -726 5335 -556
rect 6008 -576 6088 -556
rect 5575 -636 5655 -616
rect 5575 -639 6079 -636
rect 5575 -673 5598 -639
rect 5632 -673 6079 -639
rect 5575 -676 6079 -673
rect 5575 -696 5655 -676
rect 2795 -756 2875 -736
rect 2595 -759 2875 -756
rect 2595 -793 2818 -759
rect 2852 -793 2875 -759
rect 2595 -796 2875 -793
rect 2795 -816 2875 -796
rect 2945 -759 3025 -736
rect 2945 -793 2968 -759
rect 3002 -793 3025 -759
rect 2945 -839 3025 -793
rect 2945 -873 2968 -839
rect 3002 -873 3025 -839
rect 2507 -906 2587 -886
rect 2354 -909 2587 -906
rect 2354 -943 2530 -909
rect 2564 -943 2587 -909
rect 2354 -946 2587 -943
rect 2507 -966 2587 -946
rect 2945 -919 3025 -873
rect 2945 -953 2968 -919
rect 3002 -953 3025 -919
rect 2945 -986 3025 -953
rect 3095 -759 3175 -726
rect 3095 -793 3118 -759
rect 3152 -793 3175 -759
rect 3095 -839 3175 -793
rect 3095 -873 3118 -839
rect 3152 -873 3175 -839
rect 3095 -919 3175 -873
rect 3095 -953 3118 -919
rect 3152 -953 3175 -919
rect 3095 -986 3175 -953
rect 3245 -759 3325 -736
rect 3245 -793 3268 -759
rect 3302 -793 3325 -759
rect 3245 -839 3325 -793
rect 3245 -873 3268 -839
rect 3302 -873 3325 -839
rect 3245 -919 3325 -873
rect 3245 -953 3268 -919
rect 3302 -953 3325 -919
rect 3245 -986 3325 -953
rect 3395 -759 3475 -726
rect 3395 -793 3418 -759
rect 3452 -793 3475 -759
rect 3395 -839 3475 -793
rect 3395 -873 3418 -839
rect 3452 -873 3475 -839
rect 3395 -919 3475 -873
rect 3395 -953 3418 -919
rect 3452 -953 3475 -919
rect 3395 -986 3475 -953
rect 3545 -759 3625 -736
rect 3545 -793 3568 -759
rect 3602 -793 3625 -759
rect 3545 -839 3625 -793
rect 3695 -756 3775 -736
rect 3825 -756 3905 -736
rect 4245 -746 4325 -726
rect 4545 -746 4625 -726
rect 3695 -759 3905 -756
rect 3695 -793 3718 -759
rect 3752 -793 3848 -759
rect 3882 -793 3905 -759
rect 4825 -759 4905 -736
rect 4675 -786 4755 -766
rect 3695 -796 3905 -793
rect 3695 -816 3775 -796
rect 3825 -816 3905 -796
rect 4245 -789 4755 -786
rect 4245 -809 4698 -789
rect 3545 -873 3568 -839
rect 3602 -873 3625 -839
rect 4245 -843 4268 -809
rect 4302 -823 4698 -809
rect 4732 -823 4755 -789
rect 4302 -826 4755 -823
rect 4302 -843 4325 -826
rect 4245 -866 4325 -843
rect 4675 -846 4755 -826
rect 4825 -793 4848 -759
rect 4882 -793 4905 -759
rect 4825 -839 4905 -793
rect 3545 -919 3625 -873
rect 4825 -873 4848 -839
rect 4882 -873 4905 -839
rect 3545 -953 3568 -919
rect 3602 -953 3625 -919
rect 3545 -986 3625 -953
rect 3695 -906 3775 -886
rect 4675 -906 4755 -886
rect 3695 -909 4755 -906
rect 3695 -943 3718 -909
rect 3752 -943 4698 -909
rect 4732 -943 4755 -909
rect 3695 -946 4755 -943
rect 3695 -966 3775 -946
rect 4675 -966 4755 -946
rect 4825 -919 4905 -873
rect 4825 -953 4848 -919
rect 4882 -953 4905 -919
rect 4825 -986 4905 -953
rect 4975 -759 5055 -726
rect 4975 -793 4998 -759
rect 5032 -793 5055 -759
rect 4975 -839 5055 -793
rect 4975 -873 4998 -839
rect 5032 -873 5055 -839
rect 4975 -919 5055 -873
rect 4975 -953 4998 -919
rect 5032 -953 5055 -919
rect 4975 -986 5055 -953
rect 5125 -759 5205 -736
rect 5125 -793 5148 -759
rect 5182 -793 5205 -759
rect 5125 -839 5205 -793
rect 5125 -873 5148 -839
rect 5182 -873 5205 -839
rect 5125 -919 5205 -873
rect 5125 -953 5148 -919
rect 5182 -953 5205 -919
rect 5125 -986 5205 -953
rect 5275 -759 5355 -726
rect 5275 -793 5298 -759
rect 5332 -793 5355 -759
rect 5275 -839 5355 -793
rect 5275 -873 5298 -839
rect 5332 -873 5355 -839
rect 5275 -919 5355 -873
rect 5275 -953 5298 -919
rect 5332 -953 5355 -919
rect 5275 -986 5355 -953
rect 5425 -759 5505 -736
rect 5425 -793 5448 -759
rect 5482 -793 5505 -759
rect 5425 -839 5505 -793
rect 5425 -873 5448 -839
rect 5482 -873 5505 -839
rect 5655 -789 5735 -766
rect 5655 -823 5678 -789
rect 5712 -823 5735 -789
rect 5655 -846 5735 -823
rect 5425 -919 5505 -873
rect 5425 -953 5448 -919
rect 5482 -953 5505 -919
rect 5425 -986 5505 -953
rect 5805 -909 5885 -886
rect 5805 -943 5828 -909
rect 5862 -943 5885 -909
rect 5805 -966 5885 -943
rect 325 -1006 405 -986
rect 455 -1006 535 -986
rect -897 -1009 535 -1006
rect -897 -1029 348 -1009
rect -897 -1063 -874 -1029
rect -840 -1043 348 -1029
rect 382 -1043 478 -1009
rect 512 -1043 535 -1009
rect -840 -1046 535 -1043
rect -840 -1063 -817 -1046
rect -897 -1086 -817 -1063
rect 325 -1066 405 -1046
rect 455 -1066 535 -1046
rect 1715 -1009 1795 -986
rect 1715 -1043 1738 -1009
rect 1772 -1043 1795 -1009
rect 1715 -1066 1795 -1043
rect -85 -1139 2235 -1116
rect -85 -1173 -62 -1139
rect -28 -1173 18 -1139
rect 52 -1173 98 -1139
rect 132 -1173 178 -1139
rect 212 -1173 258 -1139
rect 292 -1173 338 -1139
rect 372 -1173 418 -1139
rect 452 -1173 498 -1139
rect 532 -1173 578 -1139
rect 612 -1173 658 -1139
rect 692 -1173 738 -1139
rect 772 -1173 818 -1139
rect 852 -1173 898 -1139
rect 932 -1173 978 -1139
rect 1012 -1173 1058 -1139
rect 1092 -1173 1138 -1139
rect 1172 -1173 1218 -1139
rect 1252 -1173 1298 -1139
rect 1332 -1173 1378 -1139
rect 1412 -1173 1458 -1139
rect 1492 -1173 1538 -1139
rect 1572 -1173 1618 -1139
rect 1652 -1173 1698 -1139
rect 1732 -1173 1778 -1139
rect 1812 -1173 1858 -1139
rect 1892 -1173 1938 -1139
rect 1972 -1173 2018 -1139
rect 2052 -1173 2098 -1139
rect 2132 -1173 2178 -1139
rect 2212 -1173 2235 -1139
rect -85 -1280 2235 -1173
rect 2595 -1139 3975 -1116
rect 2595 -1173 2628 -1139
rect 2662 -1173 2708 -1139
rect 2742 -1173 2788 -1139
rect 2822 -1173 2868 -1139
rect 2902 -1173 2948 -1139
rect 2982 -1173 3028 -1139
rect 3062 -1173 3108 -1139
rect 3142 -1173 3188 -1139
rect 3222 -1173 3268 -1139
rect 3302 -1173 3348 -1139
rect 3382 -1173 3428 -1139
rect 3462 -1173 3508 -1139
rect 3542 -1173 3588 -1139
rect 3622 -1173 3668 -1139
rect 3702 -1173 3748 -1139
rect 3782 -1173 3828 -1139
rect 3862 -1173 3908 -1139
rect 3942 -1173 3975 -1139
rect 2595 -1196 3975 -1173
rect 4325 -1139 6005 -1116
rect 4325 -1173 4348 -1139
rect 4382 -1173 4428 -1139
rect 4462 -1173 4508 -1139
rect 4542 -1173 4588 -1139
rect 4622 -1173 4668 -1139
rect 4702 -1173 4748 -1139
rect 4782 -1173 4828 -1139
rect 4862 -1173 4908 -1139
rect 4942 -1173 4988 -1139
rect 5022 -1173 5068 -1139
rect 5102 -1173 5148 -1139
rect 5182 -1173 5228 -1139
rect 5262 -1173 5308 -1139
rect 5342 -1173 5388 -1139
rect 5422 -1173 5468 -1139
rect 5502 -1173 5548 -1139
rect 5582 -1173 5628 -1139
rect 5662 -1173 5708 -1139
rect 5742 -1173 5788 -1139
rect 5822 -1173 5868 -1139
rect 5902 -1173 5948 -1139
rect 5982 -1173 6005 -1139
rect 4325 -1196 6005 -1173
rect -85 -1314 -62 -1280
rect -28 -1314 18 -1280
rect 52 -1314 98 -1280
rect 132 -1314 178 -1280
rect 212 -1314 258 -1280
rect 292 -1314 338 -1280
rect 372 -1314 418 -1280
rect 452 -1314 498 -1280
rect 532 -1314 578 -1280
rect 612 -1314 658 -1280
rect 692 -1314 738 -1280
rect 772 -1314 818 -1280
rect 852 -1314 898 -1280
rect 932 -1314 978 -1280
rect 1012 -1314 1058 -1280
rect 1092 -1314 1138 -1280
rect 1172 -1314 1218 -1280
rect 1252 -1314 1298 -1280
rect 1332 -1314 1378 -1280
rect 1412 -1314 1458 -1280
rect 1492 -1314 1538 -1280
rect 1572 -1314 1618 -1280
rect 1652 -1314 1698 -1280
rect 1732 -1314 1778 -1280
rect 1812 -1314 1858 -1280
rect 1892 -1314 1938 -1280
rect 1972 -1314 2018 -1280
rect 2052 -1314 2098 -1280
rect 2132 -1314 2178 -1280
rect 2212 -1314 2235 -1280
rect -85 -1337 2235 -1314
rect -327 -1390 -247 -1367
rect 4333 -1370 4413 -1350
rect 4010 -1373 4413 -1370
rect -327 -1424 -304 -1390
rect -270 -1407 -247 -1390
rect 5 -1407 85 -1387
rect -270 -1410 85 -1407
rect -270 -1424 28 -1410
rect -327 -1444 28 -1424
rect 62 -1444 85 -1410
rect -327 -1447 85 -1444
rect 5 -1467 85 -1447
rect 4010 -1407 4356 -1373
rect 4390 -1407 4413 -1373
rect 4010 -1410 4413 -1407
rect 735 -1500 815 -1467
rect 5 -1527 85 -1507
rect -897 -1530 85 -1527
rect -897 -1550 28 -1530
rect -897 -1584 -874 -1550
rect -840 -1564 28 -1550
rect 62 -1564 85 -1530
rect -840 -1567 85 -1564
rect -840 -1584 -817 -1567
rect -897 -1607 -817 -1584
rect 5 -1587 85 -1567
rect 735 -1534 758 -1500
rect 792 -1534 815 -1500
rect 735 -1580 815 -1534
rect 735 -1614 758 -1580
rect 792 -1614 815 -1580
rect 5 -1647 85 -1627
rect -1125 -1650 85 -1647
rect -1125 -1670 28 -1650
rect -1125 -1704 -1102 -1670
rect -1068 -1684 28 -1670
rect 62 -1684 85 -1650
rect -1068 -1687 85 -1684
rect -1068 -1704 -1045 -1687
rect -1125 -1727 -1045 -1704
rect 5 -1707 85 -1687
rect 735 -1660 815 -1614
rect 735 -1694 758 -1660
rect 792 -1694 815 -1660
rect 735 -1717 815 -1694
rect 885 -1500 965 -1467
rect 885 -1534 908 -1500
rect 942 -1534 965 -1500
rect 885 -1580 965 -1534
rect 885 -1614 908 -1580
rect 942 -1614 965 -1580
rect 885 -1660 965 -1614
rect 885 -1694 908 -1660
rect 942 -1694 965 -1660
rect 885 -1727 965 -1694
rect 1035 -1500 1115 -1467
rect 1035 -1534 1058 -1500
rect 1092 -1534 1115 -1500
rect 1035 -1580 1115 -1534
rect 1035 -1614 1058 -1580
rect 1092 -1614 1115 -1580
rect 1035 -1660 1115 -1614
rect 1035 -1694 1058 -1660
rect 1092 -1694 1115 -1660
rect 1035 -1717 1115 -1694
rect 1185 -1500 1265 -1467
rect 1185 -1534 1208 -1500
rect 1242 -1534 1265 -1500
rect 1185 -1580 1265 -1534
rect 1185 -1614 1208 -1580
rect 1242 -1614 1265 -1580
rect 1185 -1660 1265 -1614
rect 1185 -1694 1208 -1660
rect 1242 -1694 1265 -1660
rect 1185 -1727 1265 -1694
rect 1335 -1500 1415 -1467
rect 1335 -1534 1358 -1500
rect 1392 -1534 1415 -1500
rect 1335 -1580 1415 -1534
rect 1335 -1614 1358 -1580
rect 1392 -1614 1415 -1580
rect 1335 -1660 1415 -1614
rect 2596 -1599 3976 -1576
rect 2596 -1633 2629 -1599
rect 2663 -1633 2709 -1599
rect 2743 -1633 2789 -1599
rect 2823 -1633 2869 -1599
rect 2903 -1633 2949 -1599
rect 2983 -1633 3029 -1599
rect 3063 -1633 3109 -1599
rect 3143 -1633 3189 -1599
rect 3223 -1633 3269 -1599
rect 3303 -1633 3349 -1599
rect 3383 -1633 3429 -1599
rect 3463 -1633 3509 -1599
rect 3543 -1633 3589 -1599
rect 3623 -1633 3669 -1599
rect 3703 -1633 3749 -1599
rect 3783 -1633 3829 -1599
rect 3863 -1633 3909 -1599
rect 3943 -1633 3976 -1599
rect 2596 -1656 3976 -1633
rect 1335 -1694 1358 -1660
rect 1392 -1694 1415 -1660
rect 1335 -1717 1415 -1694
rect 5 -1767 85 -1747
rect -669 -1770 85 -1767
rect -669 -1790 28 -1770
rect -669 -1824 -646 -1790
rect -612 -1804 28 -1790
rect 62 -1804 85 -1770
rect -612 -1807 85 -1804
rect -612 -1824 -589 -1807
rect -669 -1847 -589 -1824
rect 5 -1827 85 -1807
rect -441 -1867 -361 -1847
rect 455 -1867 535 -1847
rect -441 -1870 535 -1867
rect -441 -1904 -418 -1870
rect -384 -1904 478 -1870
rect 512 -1904 535 -1870
rect -441 -1907 535 -1904
rect -441 -1927 -361 -1907
rect 455 -1927 535 -1907
rect 905 -1867 945 -1727
rect 1085 -1867 1165 -1847
rect 905 -1870 1165 -1867
rect 905 -1904 1108 -1870
rect 1142 -1904 1165 -1870
rect 905 -1907 1165 -1904
rect -783 -1950 -703 -1927
rect -783 -1984 -760 -1950
rect -726 -1967 -703 -1950
rect 305 -1967 385 -1947
rect -726 -1970 385 -1967
rect -726 -1984 328 -1970
rect -783 -2004 328 -1984
rect 362 -2004 385 -1970
rect -783 -2007 385 -2004
rect 305 -2027 385 -2007
rect -1011 -2050 -931 -2027
rect -1011 -2084 -988 -2050
rect -954 -2067 -931 -2050
rect 155 -2067 235 -2047
rect -954 -2070 235 -2067
rect -954 -2084 178 -2070
rect -1011 -2104 178 -2084
rect 212 -2104 235 -2070
rect -1011 -2107 235 -2104
rect 155 -2127 235 -2107
rect 5 -2167 85 -2147
rect -555 -2170 85 -2167
rect -555 -2190 28 -2170
rect -555 -2224 -532 -2190
rect -498 -2204 28 -2190
rect 62 -2204 85 -2170
rect -498 -2207 85 -2204
rect -498 -2224 -475 -2207
rect -555 -2247 -475 -2224
rect 5 -2227 85 -2207
rect 905 -2267 945 -1907
rect 1085 -1927 1165 -1907
rect 1205 -1987 1245 -1727
rect 4010 -1783 4050 -1410
rect 4333 -1430 4413 -1410
rect 6039 -1497 6079 -676
rect 6157 -1402 6197 684
rect 6369 -1402 6449 -1382
rect 6157 -1405 6449 -1402
rect 6157 -1439 6392 -1405
rect 6426 -1439 6449 -1405
rect 6157 -1442 6449 -1439
rect 6369 -1462 6449 -1442
rect 6039 -1537 6429 -1497
rect 4345 -1599 6345 -1576
rect 4345 -1633 4368 -1599
rect 4402 -1633 4448 -1599
rect 4482 -1633 4528 -1599
rect 4562 -1633 4608 -1599
rect 4642 -1633 4688 -1599
rect 4722 -1633 4768 -1599
rect 4802 -1633 4848 -1599
rect 4882 -1633 4928 -1599
rect 4962 -1633 5008 -1599
rect 5042 -1633 5088 -1599
rect 5122 -1633 5168 -1599
rect 5202 -1633 5248 -1599
rect 5282 -1633 5328 -1599
rect 5362 -1633 5408 -1599
rect 5442 -1633 5488 -1599
rect 5522 -1633 5568 -1599
rect 5602 -1633 5648 -1599
rect 5682 -1633 5728 -1599
rect 5762 -1633 5808 -1599
rect 5842 -1633 5888 -1599
rect 5922 -1633 5968 -1599
rect 6002 -1633 6048 -1599
rect 6082 -1633 6128 -1599
rect 6162 -1633 6208 -1599
rect 6242 -1633 6288 -1599
rect 6322 -1633 6345 -1599
rect 4345 -1656 6345 -1633
rect 4475 -1729 4555 -1706
rect 4475 -1763 4498 -1729
rect 4532 -1763 4555 -1729
rect 2946 -1819 3026 -1786
rect 1285 -1867 1365 -1847
rect 2215 -1867 2295 -1846
rect 1285 -1869 2295 -1867
rect 1285 -1870 2238 -1869
rect 1285 -1904 1308 -1870
rect 1342 -1903 2238 -1870
rect 2272 -1903 2295 -1869
rect 1342 -1904 2295 -1903
rect 1285 -1907 2295 -1904
rect 1285 -1927 1365 -1907
rect 2215 -1926 2295 -1907
rect 2946 -1853 2969 -1819
rect 3003 -1853 3026 -1819
rect 2946 -1899 3026 -1853
rect 2946 -1933 2969 -1899
rect 3003 -1933 3026 -1899
rect 2796 -1976 2876 -1956
rect 2388 -1979 2876 -1976
rect 2388 -1987 2819 -1979
rect 985 -2010 2819 -1987
rect 985 -2044 1008 -2010
rect 1042 -2013 2819 -2010
rect 2853 -2013 2876 -1979
rect 1042 -2016 2876 -2013
rect 1042 -2027 2428 -2016
rect 1042 -2044 1065 -2027
rect 985 -2067 1065 -2044
rect -25 -2307 945 -2267
rect -25 -2347 15 -2307
rect 275 -2347 315 -2307
rect 575 -2347 615 -2307
rect 905 -2347 945 -2307
rect 1205 -2267 1245 -2027
rect 2796 -2036 2876 -2016
rect 2946 -1979 3026 -1933
rect 2946 -2013 2969 -1979
rect 3003 -2013 3026 -1979
rect 2946 -2036 3026 -2013
rect 3096 -1819 3176 -1786
rect 3096 -1853 3119 -1819
rect 3153 -1853 3176 -1819
rect 3096 -1899 3176 -1853
rect 3096 -1933 3119 -1899
rect 3153 -1933 3176 -1899
rect 3096 -1979 3176 -1933
rect 3096 -2013 3119 -1979
rect 3153 -2013 3176 -1979
rect 3096 -2046 3176 -2013
rect 3246 -1819 3326 -1786
rect 3246 -1853 3269 -1819
rect 3303 -1853 3326 -1819
rect 3246 -1899 3326 -1853
rect 3246 -1933 3269 -1899
rect 3303 -1933 3326 -1899
rect 3246 -1979 3326 -1933
rect 3246 -2013 3269 -1979
rect 3303 -2013 3326 -1979
rect 3246 -2036 3326 -2013
rect 3396 -1819 3476 -1786
rect 3396 -1853 3419 -1819
rect 3453 -1853 3476 -1819
rect 3396 -1899 3476 -1853
rect 3396 -1933 3419 -1899
rect 3453 -1933 3476 -1899
rect 3396 -1979 3476 -1933
rect 3396 -2013 3419 -1979
rect 3453 -2013 3476 -1979
rect 3396 -2046 3476 -2013
rect 3546 -1819 3626 -1786
rect 3546 -1853 3569 -1819
rect 3603 -1853 3626 -1819
rect 3546 -1899 3626 -1853
rect 3990 -1806 4070 -1783
rect 4475 -1786 4555 -1763
rect 5755 -1726 5835 -1706
rect 6147 -1726 6227 -1706
rect 5755 -1729 6335 -1726
rect 5755 -1763 5778 -1729
rect 5812 -1763 6170 -1729
rect 6204 -1763 6335 -1729
rect 5755 -1766 6335 -1763
rect 5755 -1786 5835 -1766
rect 6147 -1786 6227 -1766
rect 3990 -1840 4013 -1806
rect 4047 -1840 4070 -1806
rect 5005 -1819 5085 -1786
rect 3990 -1863 4070 -1840
rect 4587 -1849 4667 -1826
rect 3546 -1933 3569 -1899
rect 3603 -1933 3626 -1899
rect 4587 -1883 4610 -1849
rect 4644 -1883 4667 -1849
rect 4587 -1906 4667 -1883
rect 5005 -1853 5028 -1819
rect 5062 -1853 5085 -1819
rect 5005 -1899 5085 -1853
rect 3546 -1979 3626 -1933
rect 4775 -1939 4855 -1916
rect 3546 -2013 3569 -1979
rect 3603 -2013 3626 -1979
rect 3546 -2036 3626 -2013
rect 3696 -1976 3776 -1956
rect 3826 -1976 3906 -1956
rect 3696 -1979 3906 -1976
rect 3696 -2013 3719 -1979
rect 3753 -2013 3849 -1979
rect 3883 -2013 3906 -1979
rect 4275 -1991 4355 -1968
rect 4275 -2004 4298 -1991
rect 3696 -2016 3906 -2013
rect 3696 -2036 3776 -2016
rect 3826 -2036 3906 -2016
rect 4090 -2025 4298 -2004
rect 4332 -2025 4355 -1991
rect 4775 -1973 4798 -1939
rect 4832 -1973 4855 -1939
rect 4775 -1996 4855 -1973
rect 5005 -1933 5028 -1899
rect 5062 -1933 5085 -1899
rect 5005 -1979 5085 -1933
rect 4090 -2044 4355 -2025
rect 5005 -2013 5028 -1979
rect 5062 -2013 5085 -1979
rect 5005 -2036 5085 -2013
rect 5155 -1819 5235 -1786
rect 5155 -1853 5178 -1819
rect 5212 -1853 5235 -1819
rect 5155 -1899 5235 -1853
rect 5155 -1933 5178 -1899
rect 5212 -1933 5235 -1899
rect 5155 -1979 5235 -1933
rect 5155 -2013 5178 -1979
rect 5212 -2013 5235 -1979
rect 3116 -2096 3156 -2046
rect 3296 -2096 3376 -2076
rect 3116 -2099 3376 -2096
rect 3116 -2133 3319 -2099
rect 3353 -2133 3376 -2099
rect 3116 -2136 3376 -2133
rect 1565 -2170 1645 -2147
rect 1565 -2204 1588 -2170
rect 1622 -2204 1645 -2170
rect 1565 -2227 1645 -2204
rect 1715 -2170 1795 -2147
rect 1715 -2204 1738 -2170
rect 1772 -2204 1795 -2170
rect 1715 -2227 1795 -2204
rect 1865 -2170 1945 -2147
rect 1865 -2204 1888 -2170
rect 1922 -2204 1945 -2170
rect 1865 -2227 1945 -2204
rect 2015 -2170 2095 -2147
rect 2015 -2204 2038 -2170
rect 2072 -2204 2095 -2170
rect 2015 -2227 2095 -2204
rect 2508 -2216 2588 -2196
rect 2666 -2216 2746 -2196
rect 2508 -2219 2746 -2216
rect 2508 -2253 2531 -2219
rect 2565 -2253 2689 -2219
rect 2723 -2253 2746 -2219
rect 2508 -2256 2746 -2253
rect 1205 -2307 1555 -2267
rect 2508 -2276 2588 -2256
rect 2666 -2276 2746 -2256
rect 3116 -2266 3156 -2136
rect 3296 -2156 3376 -2136
rect 1205 -2347 1245 -2307
rect 1515 -2347 1555 -2307
rect 2786 -2306 3156 -2266
rect 3196 -2216 3276 -2201
rect 3416 -2216 3456 -2046
rect 3696 -2096 3776 -2076
rect 4090 -2096 4130 -2044
rect 4275 -2048 4355 -2044
rect 5155 -2046 5235 -2013
rect 5305 -1819 5385 -1786
rect 5305 -1853 5328 -1819
rect 5362 -1853 5385 -1819
rect 5305 -1899 5385 -1853
rect 5305 -1933 5328 -1899
rect 5362 -1933 5385 -1899
rect 5305 -1979 5385 -1933
rect 5305 -2013 5328 -1979
rect 5362 -2013 5385 -1979
rect 5305 -2036 5385 -2013
rect 5455 -1819 5535 -1786
rect 5455 -1853 5478 -1819
rect 5512 -1853 5535 -1819
rect 5455 -1899 5535 -1853
rect 5455 -1933 5478 -1899
rect 5512 -1933 5535 -1899
rect 5455 -1979 5535 -1933
rect 5455 -2013 5478 -1979
rect 5512 -2013 5535 -1979
rect 5455 -2046 5535 -2013
rect 5605 -1819 5685 -1786
rect 5605 -1853 5628 -1819
rect 5662 -1853 5685 -1819
rect 5605 -1899 5685 -1853
rect 5875 -1836 5955 -1816
rect 6007 -1836 6087 -1817
rect 5875 -1839 6335 -1836
rect 5875 -1873 5898 -1839
rect 5932 -1840 6335 -1839
rect 5932 -1873 6030 -1840
rect 5875 -1874 6030 -1873
rect 6064 -1874 6335 -1840
rect 5875 -1876 6335 -1874
rect 5875 -1896 5955 -1876
rect 6007 -1897 6087 -1876
rect 5605 -1933 5628 -1899
rect 5662 -1933 5685 -1899
rect 5605 -1979 5685 -1933
rect 5605 -2013 5628 -1979
rect 5662 -2013 5685 -1979
rect 5755 -1936 5835 -1916
rect 6389 -1929 6429 -1537
rect 5755 -1939 6335 -1936
rect 5755 -1973 5778 -1939
rect 5812 -1973 6335 -1939
rect 6389 -1969 6523 -1929
rect 5755 -1976 6335 -1973
rect 5755 -1996 5835 -1976
rect 5605 -2036 5685 -2013
rect 6369 -2026 6449 -2003
rect 4855 -2096 4935 -2076
rect 3696 -2099 4130 -2096
rect 3696 -2133 3719 -2099
rect 3753 -2133 4130 -2099
rect 3696 -2136 4130 -2133
rect 4275 -2099 4935 -2096
rect 4275 -2119 4878 -2099
rect 3696 -2156 3776 -2136
rect 4275 -2153 4298 -2119
rect 4332 -2133 4878 -2119
rect 4912 -2133 4935 -2099
rect 4332 -2136 4935 -2133
rect 4332 -2153 4355 -2136
rect 4275 -2176 4355 -2153
rect 4855 -2156 4935 -2136
rect 5175 -2216 5215 -2046
rect 5255 -2096 5335 -2076
rect 5475 -2096 5515 -2046
rect 5255 -2099 5515 -2096
rect 5255 -2133 5278 -2099
rect 5312 -2133 5515 -2099
rect 6175 -2049 6392 -2026
rect 6175 -2083 6198 -2049
rect 6232 -2060 6392 -2049
rect 6426 -2060 6449 -2026
rect 6232 -2066 6449 -2060
rect 6232 -2083 6255 -2066
rect 6369 -2083 6449 -2066
rect 6175 -2106 6255 -2083
rect 5255 -2136 5515 -2133
rect 5255 -2156 5335 -2136
rect 5355 -2216 5435 -2201
rect 3196 -2224 3456 -2216
rect 3196 -2258 3219 -2224
rect 3253 -2256 3456 -2224
rect 4275 -2224 5435 -2216
rect 4275 -2239 5378 -2224
rect 3253 -2258 3276 -2256
rect 3196 -2281 3276 -2258
rect 3416 -2266 3456 -2256
rect 3990 -2266 4070 -2246
rect 3416 -2269 4070 -2266
rect 3416 -2303 4013 -2269
rect 4047 -2303 4070 -2269
rect 4275 -2273 4298 -2239
rect 4332 -2256 5378 -2239
rect 4332 -2273 4355 -2256
rect 4275 -2296 4355 -2273
rect 3416 -2306 4070 -2303
rect 2786 -2346 2826 -2306
rect 3116 -2346 3156 -2306
rect -45 -2380 35 -2347
rect -45 -2414 -22 -2380
rect 12 -2414 35 -2380
rect -45 -2460 35 -2414
rect -45 -2494 -22 -2460
rect 12 -2494 35 -2460
rect -45 -2540 35 -2494
rect -45 -2574 -22 -2540
rect 12 -2574 35 -2540
rect -45 -2597 35 -2574
rect 105 -2380 185 -2347
rect 105 -2414 128 -2380
rect 162 -2414 185 -2380
rect 105 -2460 185 -2414
rect 105 -2494 128 -2460
rect 162 -2494 185 -2460
rect 105 -2540 185 -2494
rect 105 -2574 128 -2540
rect 162 -2574 185 -2540
rect 105 -2597 185 -2574
rect 255 -2380 335 -2347
rect 255 -2414 278 -2380
rect 312 -2414 335 -2380
rect 255 -2460 335 -2414
rect 255 -2494 278 -2460
rect 312 -2494 335 -2460
rect 255 -2540 335 -2494
rect 255 -2574 278 -2540
rect 312 -2574 335 -2540
rect 255 -2597 335 -2574
rect 405 -2380 485 -2347
rect 405 -2414 428 -2380
rect 462 -2414 485 -2380
rect 405 -2460 485 -2414
rect 405 -2494 428 -2460
rect 462 -2494 485 -2460
rect 405 -2540 485 -2494
rect 405 -2574 428 -2540
rect 462 -2574 485 -2540
rect 405 -2597 485 -2574
rect 555 -2380 635 -2347
rect 555 -2414 578 -2380
rect 612 -2414 635 -2380
rect 555 -2460 635 -2414
rect 555 -2494 578 -2460
rect 612 -2494 635 -2460
rect 555 -2540 635 -2494
rect 555 -2574 578 -2540
rect 612 -2574 635 -2540
rect 555 -2597 635 -2574
rect 735 -2380 815 -2347
rect 735 -2414 758 -2380
rect 792 -2414 815 -2380
rect 735 -2460 815 -2414
rect 735 -2494 758 -2460
rect 792 -2494 815 -2460
rect 735 -2540 815 -2494
rect 735 -2574 758 -2540
rect 792 -2574 815 -2540
rect 735 -2597 815 -2574
rect 885 -2380 965 -2347
rect 885 -2414 908 -2380
rect 942 -2414 965 -2380
rect 885 -2460 965 -2414
rect 885 -2494 908 -2460
rect 942 -2494 965 -2460
rect 885 -2540 965 -2494
rect 885 -2574 908 -2540
rect 942 -2574 965 -2540
rect 885 -2597 965 -2574
rect 1035 -2380 1115 -2347
rect 1035 -2414 1058 -2380
rect 1092 -2414 1115 -2380
rect 1035 -2460 1115 -2414
rect 1035 -2494 1058 -2460
rect 1092 -2494 1115 -2460
rect 1035 -2540 1115 -2494
rect 1035 -2574 1058 -2540
rect 1092 -2574 1115 -2540
rect 1035 -2597 1115 -2574
rect 1185 -2380 1265 -2347
rect 1185 -2414 1208 -2380
rect 1242 -2414 1265 -2380
rect 1185 -2460 1265 -2414
rect 1185 -2494 1208 -2460
rect 1242 -2494 1265 -2460
rect 1185 -2540 1265 -2494
rect 1185 -2574 1208 -2540
rect 1242 -2574 1265 -2540
rect 1185 -2597 1265 -2574
rect 1335 -2380 1415 -2347
rect 1335 -2414 1358 -2380
rect 1392 -2414 1415 -2380
rect 1335 -2460 1415 -2414
rect 1335 -2494 1358 -2460
rect 1392 -2494 1415 -2460
rect 1335 -2540 1415 -2494
rect 1335 -2574 1358 -2540
rect 1392 -2574 1415 -2540
rect 1335 -2597 1415 -2574
rect 1515 -2380 1595 -2347
rect 1515 -2414 1538 -2380
rect 1572 -2414 1595 -2380
rect 1515 -2460 1595 -2414
rect 1515 -2494 1538 -2460
rect 1572 -2494 1595 -2460
rect 1515 -2540 1595 -2494
rect 1515 -2574 1538 -2540
rect 1572 -2574 1595 -2540
rect 1515 -2597 1595 -2574
rect 2115 -2380 2195 -2347
rect 2115 -2414 2138 -2380
rect 2172 -2414 2195 -2380
rect 2115 -2460 2195 -2414
rect 2115 -2494 2138 -2460
rect 2172 -2494 2195 -2460
rect 2115 -2540 2195 -2494
rect 2115 -2574 2138 -2540
rect 2172 -2574 2195 -2540
rect 2115 -2597 2195 -2574
rect 2616 -2379 2696 -2346
rect 2616 -2413 2639 -2379
rect 2673 -2413 2696 -2379
rect 2616 -2459 2696 -2413
rect 2616 -2493 2639 -2459
rect 2673 -2493 2696 -2459
rect 2616 -2539 2696 -2493
rect 2616 -2573 2639 -2539
rect 2673 -2573 2696 -2539
rect 2616 -2596 2696 -2573
rect 2766 -2379 2846 -2346
rect 2766 -2413 2789 -2379
rect 2823 -2413 2846 -2379
rect 2766 -2459 2846 -2413
rect 2766 -2493 2789 -2459
rect 2823 -2493 2846 -2459
rect 2766 -2539 2846 -2493
rect 2766 -2573 2789 -2539
rect 2823 -2573 2846 -2539
rect 2766 -2596 2846 -2573
rect 2946 -2379 3026 -2346
rect 2946 -2413 2969 -2379
rect 3003 -2413 3026 -2379
rect 2946 -2459 3026 -2413
rect 2946 -2493 2969 -2459
rect 3003 -2493 3026 -2459
rect 2946 -2539 3026 -2493
rect 2946 -2573 2969 -2539
rect 3003 -2573 3026 -2539
rect 2946 -2596 3026 -2573
rect 3096 -2379 3176 -2346
rect 3096 -2413 3119 -2379
rect 3153 -2413 3176 -2379
rect 3096 -2459 3176 -2413
rect 3096 -2493 3119 -2459
rect 3153 -2493 3176 -2459
rect 3096 -2539 3176 -2493
rect 3096 -2573 3119 -2539
rect 3153 -2573 3176 -2539
rect 3096 -2596 3176 -2573
rect 3246 -2379 3326 -2346
rect 3246 -2413 3269 -2379
rect 3303 -2413 3326 -2379
rect 3246 -2459 3326 -2413
rect 3246 -2493 3269 -2459
rect 3303 -2493 3326 -2459
rect 3246 -2539 3326 -2493
rect 3246 -2573 3269 -2539
rect 3303 -2573 3326 -2539
rect 3246 -2596 3326 -2573
rect 3396 -2379 3476 -2306
rect 3746 -2346 3786 -2306
rect 3990 -2326 4070 -2306
rect 4545 -2346 4585 -2256
rect 4845 -2346 4885 -2256
rect 5175 -2346 5215 -2256
rect 5355 -2258 5378 -2256
rect 5412 -2258 5435 -2224
rect 5355 -2281 5435 -2258
rect 5475 -2266 5515 -2136
rect 6035 -2146 6115 -2126
rect 6483 -2146 6523 -1969
rect 6035 -2149 6523 -2146
rect 6035 -2183 6058 -2149
rect 6092 -2183 6523 -2149
rect 6035 -2186 6523 -2183
rect 6035 -2206 6115 -2186
rect 5885 -2229 5965 -2206
rect 5885 -2263 5908 -2229
rect 5942 -2246 5965 -2229
rect 5942 -2263 6335 -2246
rect 5475 -2306 5825 -2266
rect 5885 -2286 6335 -2263
rect 5475 -2346 5515 -2306
rect 5785 -2346 5825 -2306
rect 3396 -2413 3419 -2379
rect 3453 -2413 3476 -2379
rect 3396 -2459 3476 -2413
rect 3396 -2493 3419 -2459
rect 3453 -2493 3476 -2459
rect 3396 -2539 3476 -2493
rect 3396 -2573 3419 -2539
rect 3453 -2573 3476 -2539
rect 3396 -2596 3476 -2573
rect 3546 -2379 3626 -2346
rect 3546 -2413 3569 -2379
rect 3603 -2413 3626 -2379
rect 3546 -2459 3626 -2413
rect 3546 -2493 3569 -2459
rect 3603 -2493 3626 -2459
rect 3546 -2539 3626 -2493
rect 3546 -2573 3569 -2539
rect 3603 -2573 3626 -2539
rect 3546 -2596 3626 -2573
rect 3726 -2379 3806 -2346
rect 3726 -2413 3749 -2379
rect 3783 -2413 3806 -2379
rect 3726 -2459 3806 -2413
rect 3726 -2493 3749 -2459
rect 3783 -2493 3806 -2459
rect 3726 -2539 3806 -2493
rect 3726 -2573 3749 -2539
rect 3783 -2573 3806 -2539
rect 3726 -2596 3806 -2573
rect 3876 -2379 3956 -2346
rect 3876 -2413 3899 -2379
rect 3933 -2413 3956 -2379
rect 3876 -2459 3956 -2413
rect 3876 -2493 3899 -2459
rect 3933 -2493 3956 -2459
rect 3876 -2539 3956 -2493
rect 3876 -2573 3899 -2539
rect 3933 -2573 3956 -2539
rect 3876 -2596 3956 -2573
rect 4375 -2379 4455 -2346
rect 4375 -2413 4398 -2379
rect 4432 -2413 4455 -2379
rect 4375 -2459 4455 -2413
rect 4375 -2493 4398 -2459
rect 4432 -2493 4455 -2459
rect 4375 -2539 4455 -2493
rect 4375 -2573 4398 -2539
rect 4432 -2573 4455 -2539
rect 4375 -2596 4455 -2573
rect 4525 -2379 4605 -2346
rect 4525 -2413 4548 -2379
rect 4582 -2413 4605 -2379
rect 4525 -2459 4605 -2413
rect 4525 -2493 4548 -2459
rect 4582 -2493 4605 -2459
rect 4525 -2539 4605 -2493
rect 4525 -2573 4548 -2539
rect 4582 -2573 4605 -2539
rect 4525 -2596 4605 -2573
rect 4675 -2379 4755 -2346
rect 4675 -2413 4698 -2379
rect 4732 -2413 4755 -2379
rect 4675 -2459 4755 -2413
rect 4675 -2493 4698 -2459
rect 4732 -2493 4755 -2459
rect 4675 -2539 4755 -2493
rect 4675 -2573 4698 -2539
rect 4732 -2573 4755 -2539
rect 4675 -2596 4755 -2573
rect 4825 -2379 4905 -2346
rect 4825 -2413 4848 -2379
rect 4882 -2413 4905 -2379
rect 4825 -2459 4905 -2413
rect 4825 -2493 4848 -2459
rect 4882 -2493 4905 -2459
rect 4825 -2539 4905 -2493
rect 4825 -2573 4848 -2539
rect 4882 -2573 4905 -2539
rect 4825 -2596 4905 -2573
rect 5005 -2379 5085 -2346
rect 5005 -2413 5028 -2379
rect 5062 -2413 5085 -2379
rect 5005 -2459 5085 -2413
rect 5005 -2493 5028 -2459
rect 5062 -2493 5085 -2459
rect 5005 -2539 5085 -2493
rect 5005 -2573 5028 -2539
rect 5062 -2573 5085 -2539
rect 5005 -2596 5085 -2573
rect 5155 -2379 5235 -2346
rect 5155 -2413 5178 -2379
rect 5212 -2413 5235 -2379
rect 5155 -2459 5235 -2413
rect 5155 -2493 5178 -2459
rect 5212 -2493 5235 -2459
rect 5155 -2539 5235 -2493
rect 5155 -2573 5178 -2539
rect 5212 -2573 5235 -2539
rect 5155 -2596 5235 -2573
rect 5305 -2379 5385 -2346
rect 5305 -2413 5328 -2379
rect 5362 -2413 5385 -2379
rect 5305 -2459 5385 -2413
rect 5305 -2493 5328 -2459
rect 5362 -2493 5385 -2459
rect 5305 -2539 5385 -2493
rect 5305 -2573 5328 -2539
rect 5362 -2573 5385 -2539
rect 5305 -2596 5385 -2573
rect 5455 -2379 5535 -2346
rect 5455 -2413 5478 -2379
rect 5512 -2413 5535 -2379
rect 5455 -2459 5535 -2413
rect 5455 -2493 5478 -2459
rect 5512 -2493 5535 -2459
rect 5455 -2539 5535 -2493
rect 5455 -2573 5478 -2539
rect 5512 -2573 5535 -2539
rect 5455 -2596 5535 -2573
rect 5605 -2379 5685 -2346
rect 5605 -2413 5628 -2379
rect 5662 -2413 5685 -2379
rect 5605 -2459 5685 -2413
rect 5605 -2493 5628 -2459
rect 5662 -2493 5685 -2459
rect 5605 -2539 5685 -2493
rect 5605 -2573 5628 -2539
rect 5662 -2573 5685 -2539
rect 5605 -2596 5685 -2573
rect 5785 -2379 5865 -2346
rect 5785 -2413 5808 -2379
rect 5842 -2413 5865 -2379
rect 5785 -2459 5865 -2413
rect 5785 -2493 5808 -2459
rect 5842 -2493 5865 -2459
rect 5785 -2539 5865 -2493
rect 5785 -2573 5808 -2539
rect 5842 -2573 5865 -2539
rect 5785 -2596 5865 -2573
rect 6235 -2379 6315 -2346
rect 6235 -2413 6258 -2379
rect 6292 -2413 6315 -2379
rect 6235 -2459 6315 -2413
rect 6235 -2493 6258 -2459
rect 6292 -2493 6315 -2459
rect 6235 -2539 6315 -2493
rect 6235 -2573 6258 -2539
rect 6292 -2573 6315 -2539
rect 6235 -2596 6315 -2573
rect -83 -2657 -3 -2636
rect 835 -2657 915 -2637
rect 1235 -2657 1315 -2637
rect 3046 -2656 3126 -2636
rect 3446 -2656 3526 -2636
rect 3990 -2656 4070 -2636
rect -83 -2659 1315 -2657
rect -83 -2693 -60 -2659
rect -26 -2660 1315 -2659
rect -26 -2693 858 -2660
rect -83 -2694 858 -2693
rect 892 -2694 1258 -2660
rect 1292 -2694 1315 -2660
rect -83 -2697 1315 -2694
rect 2596 -2659 4070 -2656
rect 2596 -2693 3069 -2659
rect 3103 -2693 3469 -2659
rect 3503 -2693 4013 -2659
rect 4047 -2693 4070 -2659
rect 2596 -2696 4070 -2693
rect -83 -2716 -3 -2697
rect 835 -2717 915 -2697
rect 1235 -2717 1315 -2697
rect 3046 -2716 3126 -2696
rect 3446 -2716 3526 -2696
rect 3990 -2716 4070 -2696
rect 4187 -2656 4267 -2636
rect 5105 -2656 5185 -2636
rect 5505 -2656 5585 -2636
rect 4187 -2659 6335 -2656
rect 4187 -2693 4210 -2659
rect 4244 -2693 5128 -2659
rect 5162 -2693 5528 -2659
rect 5562 -2693 6335 -2659
rect 4187 -2696 6335 -2693
rect 4187 -2716 4267 -2696
rect 5105 -2716 5185 -2696
rect 5505 -2716 5585 -2696
rect -213 -2780 2235 -2757
rect -213 -2814 -190 -2780
rect -156 -2814 -62 -2780
rect -28 -2814 18 -2780
rect 52 -2814 98 -2780
rect 132 -2814 178 -2780
rect 212 -2814 258 -2780
rect 292 -2814 338 -2780
rect 372 -2814 418 -2780
rect 452 -2814 498 -2780
rect 532 -2814 578 -2780
rect 612 -2814 658 -2780
rect 692 -2814 738 -2780
rect 772 -2814 818 -2780
rect 852 -2814 898 -2780
rect 932 -2814 978 -2780
rect 1012 -2814 1058 -2780
rect 1092 -2814 1138 -2780
rect 1172 -2814 1218 -2780
rect 1252 -2814 1298 -2780
rect 1332 -2814 1378 -2780
rect 1412 -2814 1458 -2780
rect 1492 -2814 1538 -2780
rect 1572 -2814 1618 -2780
rect 1652 -2814 1698 -2780
rect 1732 -2814 1778 -2780
rect 1812 -2814 1858 -2780
rect 1892 -2814 1938 -2780
rect 1972 -2814 2018 -2780
rect 2052 -2814 2098 -2780
rect 2132 -2814 2178 -2780
rect 2212 -2814 2235 -2780
rect -213 -2837 2235 -2814
rect 2596 -2779 3976 -2756
rect 2596 -2813 2629 -2779
rect 2663 -2813 2709 -2779
rect 2743 -2813 2789 -2779
rect 2823 -2813 2869 -2779
rect 2903 -2813 2949 -2779
rect 2983 -2813 3029 -2779
rect 3063 -2813 3109 -2779
rect 3143 -2813 3189 -2779
rect 3223 -2813 3269 -2779
rect 3303 -2813 3349 -2779
rect 3383 -2813 3429 -2779
rect 3463 -2813 3509 -2779
rect 3543 -2813 3589 -2779
rect 3623 -2813 3669 -2779
rect 3703 -2813 3749 -2779
rect 3783 -2813 3829 -2779
rect 3863 -2813 3909 -2779
rect 3943 -2813 3976 -2779
rect 2596 -2836 3976 -2813
rect 4345 -2779 6345 -2756
rect 4345 -2813 4368 -2779
rect 4402 -2813 4448 -2779
rect 4482 -2813 4528 -2779
rect 4562 -2813 4608 -2779
rect 4642 -2813 4688 -2779
rect 4722 -2813 4768 -2779
rect 4802 -2813 4848 -2779
rect 4882 -2813 4928 -2779
rect 4962 -2813 5008 -2779
rect 5042 -2813 5088 -2779
rect 5122 -2813 5168 -2779
rect 5202 -2813 5248 -2779
rect 5282 -2813 5328 -2779
rect 5362 -2813 5408 -2779
rect 5442 -2813 5488 -2779
rect 5522 -2813 5568 -2779
rect 5602 -2813 5648 -2779
rect 5682 -2813 5728 -2779
rect 5762 -2813 5808 -2779
rect 5842 -2813 5888 -2779
rect 5922 -2813 5968 -2779
rect 6002 -2813 6048 -2779
rect 6082 -2813 6128 -2779
rect 6162 -2813 6208 -2779
rect 6242 -2813 6288 -2779
rect 6322 -2813 6345 -2779
rect 4345 -2836 6345 -2813
<< viali >>
rect 18 1187 52 1221
rect 98 1187 132 1221
rect 178 1187 212 1221
rect 258 1187 292 1221
rect 338 1187 372 1221
rect 418 1187 452 1221
rect 498 1187 532 1221
rect 578 1187 612 1221
rect 658 1187 692 1221
rect 738 1187 772 1221
rect 818 1187 852 1221
rect 898 1187 932 1221
rect 978 1187 1012 1221
rect 1058 1187 1092 1221
rect 1138 1187 1172 1221
rect 1218 1187 1252 1221
rect 1298 1187 1332 1221
rect 1378 1187 1412 1221
rect 1458 1187 1492 1221
rect 1538 1187 1572 1221
rect 1618 1187 1652 1221
rect 1698 1187 1732 1221
rect 1778 1187 1812 1221
rect 1858 1187 1892 1221
rect 1938 1187 1972 1221
rect 2018 1187 2052 1221
rect 2098 1187 2132 1221
rect 2628 1187 2662 1221
rect 2708 1187 2742 1221
rect 2788 1187 2822 1221
rect 2868 1187 2902 1221
rect 2948 1187 2982 1221
rect 3028 1187 3062 1221
rect 3108 1187 3142 1221
rect 3188 1187 3222 1221
rect 3268 1187 3302 1221
rect 3348 1187 3382 1221
rect 3428 1187 3462 1221
rect 3508 1187 3542 1221
rect 3588 1187 3622 1221
rect 3668 1187 3702 1221
rect 3748 1187 3782 1221
rect 3828 1187 3862 1221
rect 3908 1187 3942 1221
rect 4348 1187 4382 1221
rect 4428 1187 4462 1221
rect 4508 1187 4542 1221
rect 4588 1187 4622 1221
rect 4668 1187 4702 1221
rect 4748 1187 4782 1221
rect 4828 1187 4862 1221
rect 4908 1187 4942 1221
rect 4988 1187 5022 1221
rect 5068 1187 5102 1221
rect 5148 1187 5182 1221
rect 5228 1187 5262 1221
rect 5308 1187 5342 1221
rect 5388 1187 5422 1221
rect 5468 1187 5502 1221
rect 5548 1187 5582 1221
rect 5628 1187 5662 1221
rect 5708 1187 5742 1221
rect 5788 1187 5822 1221
rect 5868 1187 5902 1221
rect 5948 1187 5982 1221
rect -418 1037 -384 1071
rect 478 1057 512 1091
rect 1738 1057 1772 1091
rect -304 955 -270 989
rect 608 957 642 991
rect 758 967 792 1001
rect -646 837 -612 871
rect 478 857 512 891
rect 758 887 792 921
rect -532 737 -498 771
rect 608 757 642 791
rect 758 807 792 841
rect 1058 967 1092 1001
rect 1058 887 1092 921
rect 1058 807 1092 841
rect 1358 967 1392 1001
rect 1938 957 1972 991
rect 2530 991 2564 1025
rect 1358 887 1392 921
rect 1358 807 1392 841
rect 2088 857 2122 891
rect 1108 687 1142 721
rect 1638 757 1672 791
rect 1478 677 1512 711
rect 2968 967 3002 1001
rect 2968 887 3002 921
rect 2818 807 2852 841
rect 2968 807 3002 841
rect 3268 967 3302 1001
rect 3268 887 3302 921
rect 3268 807 3302 841
rect 3568 967 3602 1001
rect 4006 991 4040 1025
rect 4698 957 4732 991
rect 4848 967 4882 1001
rect 3568 887 3602 921
rect 4006 876 4040 910
rect 3568 807 3602 841
rect 4268 857 4302 891
rect 3718 807 3752 841
rect 4698 837 4732 871
rect 4848 887 4882 921
rect 4848 807 4882 841
rect 5148 967 5182 1001
rect 5148 887 5182 921
rect 5148 807 5182 841
rect 5448 967 5482 1001
rect 5828 957 5862 991
rect 5448 887 5482 921
rect 5448 807 5482 841
rect 5678 837 5712 871
rect 3318 687 3352 721
rect 2238 563 2272 597
rect 278 407 312 441
rect 278 327 312 361
rect 278 247 312 281
rect 758 407 792 441
rect 758 327 792 361
rect 758 247 792 281
rect 1058 407 1092 441
rect 1058 327 1092 361
rect 1058 247 1092 281
rect 1358 407 1392 441
rect 1358 327 1392 361
rect 1358 247 1392 281
rect 1838 407 1872 441
rect 1838 327 1872 361
rect 1838 247 1872 281
rect 3718 687 3752 721
rect 5198 687 5232 721
rect 4006 537 4040 571
rect 5598 687 5632 721
rect 6031 566 6065 600
rect 2252 325 2286 359
rect 2638 407 2672 441
rect 2638 327 2672 361
rect 2638 247 2672 281
rect 2968 407 3002 441
rect 2968 327 3002 361
rect 2968 247 3002 281
rect 3268 407 3302 441
rect 3268 327 3302 361
rect 3268 247 3302 281
rect 3568 407 3602 441
rect 3568 327 3602 361
rect 3568 247 3602 281
rect 3898 407 3932 441
rect 3898 327 3932 361
rect 3898 247 3932 281
rect 4518 407 4552 441
rect 4518 327 4552 361
rect 4518 247 4552 281
rect 4848 407 4882 441
rect 4848 327 4882 361
rect 4848 247 4882 281
rect 5148 407 5182 441
rect 5148 327 5182 361
rect 5148 247 5182 281
rect 5448 407 5482 441
rect 5448 327 5482 361
rect 5448 247 5482 281
rect 5928 407 5962 441
rect 5928 327 5962 361
rect 5928 247 5962 281
rect 390 127 424 161
rect 4356 127 4390 161
rect -190 7 -156 41
rect 18 7 52 41
rect 98 7 132 41
rect 178 7 212 41
rect 258 7 292 41
rect 338 7 372 41
rect 418 7 452 41
rect 498 7 532 41
rect 578 7 612 41
rect 658 7 692 41
rect 738 7 772 41
rect 818 7 852 41
rect 898 7 932 41
rect 978 7 1012 41
rect 1058 7 1092 41
rect 1138 7 1172 41
rect 1218 7 1252 41
rect 1298 7 1332 41
rect 1378 7 1412 41
rect 1458 7 1492 41
rect 1538 7 1572 41
rect 1618 7 1652 41
rect 1698 7 1732 41
rect 1778 7 1812 41
rect 1858 7 1892 41
rect 1938 7 1972 41
rect 2018 7 2052 41
rect 2098 7 2132 41
rect 2628 7 2662 41
rect 2708 7 2742 41
rect 2788 7 2822 41
rect 2868 7 2902 41
rect 2948 7 2982 41
rect 3028 7 3062 41
rect 3108 7 3142 41
rect 3188 7 3222 41
rect 3268 7 3302 41
rect 3348 7 3382 41
rect 3428 7 3462 41
rect 3508 7 3542 41
rect 3588 7 3622 41
rect 3668 7 3702 41
rect 3748 7 3782 41
rect 3828 7 3862 41
rect 3908 7 3942 41
rect 4348 7 4382 41
rect 4428 7 4462 41
rect 4508 7 4542 41
rect 4588 7 4622 41
rect 4668 7 4702 41
rect 4748 7 4782 41
rect 4828 7 4862 41
rect 4908 7 4942 41
rect 4988 7 5022 41
rect 5068 7 5102 41
rect 5148 7 5182 41
rect 5228 7 5262 41
rect 5308 7 5342 41
rect 5388 7 5422 41
rect 5468 7 5502 41
rect 5548 7 5582 41
rect 5628 7 5662 41
rect 5708 7 5742 41
rect 5788 7 5822 41
rect 5868 7 5902 41
rect 5948 7 5982 41
rect 390 -113 424 -79
rect 4356 -113 4390 -79
rect 278 -233 312 -199
rect 278 -313 312 -279
rect 278 -393 312 -359
rect 758 -233 792 -199
rect 758 -313 792 -279
rect 758 -393 792 -359
rect 1058 -233 1092 -199
rect 1058 -313 1092 -279
rect 1058 -393 1092 -359
rect 1358 -233 1392 -199
rect 1358 -313 1392 -279
rect 1358 -393 1392 -359
rect 1838 -233 1872 -199
rect 1838 -313 1872 -279
rect 1838 -393 1872 -359
rect 2638 -233 2672 -199
rect 2252 -313 2286 -279
rect 2638 -313 2672 -279
rect 2638 -393 2672 -359
rect 2968 -233 3002 -199
rect 2968 -313 3002 -279
rect 2968 -393 3002 -359
rect 3268 -233 3302 -199
rect 3268 -313 3302 -279
rect 3268 -393 3302 -359
rect 3568 -233 3602 -199
rect 3568 -313 3602 -279
rect 3568 -393 3602 -359
rect 3898 -233 3932 -199
rect 3898 -313 3932 -279
rect 3898 -393 3932 -359
rect 4518 -233 4552 -199
rect 4518 -313 4552 -279
rect 4518 -393 4552 -359
rect 4848 -233 4882 -199
rect 4848 -313 4882 -279
rect 4848 -393 4882 -359
rect 5148 -233 5182 -199
rect 5148 -313 5182 -279
rect 5148 -393 5182 -359
rect 5448 -233 5482 -199
rect 5448 -313 5482 -279
rect 5448 -393 5482 -359
rect 5928 -233 5962 -199
rect 5928 -313 5962 -279
rect 5928 -393 5962 -359
rect 1108 -673 1142 -639
rect -988 -723 -954 -689
rect 608 -743 642 -709
rect 1478 -663 1512 -629
rect 2238 -663 2272 -629
rect -1102 -842 -1068 -808
rect 478 -843 512 -809
rect 758 -793 792 -759
rect 758 -873 792 -839
rect -760 -949 -726 -915
rect 608 -943 642 -909
rect 758 -953 792 -919
rect 1058 -793 1092 -759
rect 1058 -873 1092 -839
rect 1058 -953 1092 -919
rect 1358 -793 1392 -759
rect 1638 -743 1672 -709
rect 1358 -873 1392 -839
rect 2088 -843 2122 -809
rect 1358 -953 1392 -919
rect 1938 -943 1972 -909
rect 4006 -503 4040 -469
rect 3318 -673 3352 -639
rect 3718 -673 3752 -639
rect 6031 -553 6065 -519
rect 4268 -723 4302 -689
rect 5198 -673 5232 -639
rect 5598 -673 5632 -639
rect 2818 -793 2852 -759
rect 2968 -793 3002 -759
rect 2968 -873 3002 -839
rect 2530 -943 2564 -909
rect 2968 -953 3002 -919
rect 3268 -793 3302 -759
rect 3268 -873 3302 -839
rect 3268 -953 3302 -919
rect 3568 -793 3602 -759
rect 3718 -793 3752 -759
rect 3568 -873 3602 -839
rect 4268 -843 4302 -809
rect 4698 -823 4732 -789
rect 4848 -793 4882 -759
rect 4848 -873 4882 -839
rect 3568 -953 3602 -919
rect 3718 -943 3752 -909
rect 4698 -943 4732 -909
rect 4848 -953 4882 -919
rect 5148 -793 5182 -759
rect 5148 -873 5182 -839
rect 5148 -953 5182 -919
rect 5448 -793 5482 -759
rect 5448 -873 5482 -839
rect 5678 -823 5712 -789
rect 5448 -953 5482 -919
rect 5828 -943 5862 -909
rect -874 -1063 -840 -1029
rect 478 -1043 512 -1009
rect 1738 -1043 1772 -1009
rect -62 -1173 -28 -1139
rect 18 -1173 52 -1139
rect 98 -1173 132 -1139
rect 178 -1173 212 -1139
rect 258 -1173 292 -1139
rect 338 -1173 372 -1139
rect 418 -1173 452 -1139
rect 498 -1173 532 -1139
rect 578 -1173 612 -1139
rect 658 -1173 692 -1139
rect 738 -1173 772 -1139
rect 818 -1173 852 -1139
rect 898 -1173 932 -1139
rect 978 -1173 1012 -1139
rect 1058 -1173 1092 -1139
rect 1138 -1173 1172 -1139
rect 1218 -1173 1252 -1139
rect 1298 -1173 1332 -1139
rect 1378 -1173 1412 -1139
rect 1458 -1173 1492 -1139
rect 1538 -1173 1572 -1139
rect 1618 -1173 1652 -1139
rect 1698 -1173 1732 -1139
rect 1778 -1173 1812 -1139
rect 1858 -1173 1892 -1139
rect 1938 -1173 1972 -1139
rect 2018 -1173 2052 -1139
rect 2098 -1173 2132 -1139
rect 2178 -1173 2212 -1139
rect 2628 -1173 2662 -1139
rect 2708 -1173 2742 -1139
rect 2788 -1173 2822 -1139
rect 2868 -1173 2902 -1139
rect 2948 -1173 2982 -1139
rect 3028 -1173 3062 -1139
rect 3108 -1173 3142 -1139
rect 3188 -1173 3222 -1139
rect 3268 -1173 3302 -1139
rect 3348 -1173 3382 -1139
rect 3428 -1173 3462 -1139
rect 3508 -1173 3542 -1139
rect 3588 -1173 3622 -1139
rect 3668 -1173 3702 -1139
rect 3748 -1173 3782 -1139
rect 3828 -1173 3862 -1139
rect 3908 -1173 3942 -1139
rect 4348 -1173 4382 -1139
rect 4428 -1173 4462 -1139
rect 4508 -1173 4542 -1139
rect 4588 -1173 4622 -1139
rect 4668 -1173 4702 -1139
rect 4748 -1173 4782 -1139
rect 4828 -1173 4862 -1139
rect 4908 -1173 4942 -1139
rect 4988 -1173 5022 -1139
rect 5068 -1173 5102 -1139
rect 5148 -1173 5182 -1139
rect 5228 -1173 5262 -1139
rect 5308 -1173 5342 -1139
rect 5388 -1173 5422 -1139
rect 5468 -1173 5502 -1139
rect 5548 -1173 5582 -1139
rect 5628 -1173 5662 -1139
rect 5708 -1173 5742 -1139
rect 5788 -1173 5822 -1139
rect 5868 -1173 5902 -1139
rect 5948 -1173 5982 -1139
rect -62 -1314 -28 -1280
rect 18 -1314 52 -1280
rect 98 -1314 132 -1280
rect 178 -1314 212 -1280
rect 258 -1314 292 -1280
rect 338 -1314 372 -1280
rect 418 -1314 452 -1280
rect 498 -1314 532 -1280
rect 578 -1314 612 -1280
rect 658 -1314 692 -1280
rect 738 -1314 772 -1280
rect 818 -1314 852 -1280
rect 898 -1314 932 -1280
rect 978 -1314 1012 -1280
rect 1058 -1314 1092 -1280
rect 1138 -1314 1172 -1280
rect 1218 -1314 1252 -1280
rect 1298 -1314 1332 -1280
rect 1378 -1314 1412 -1280
rect 1458 -1314 1492 -1280
rect 1538 -1314 1572 -1280
rect 1618 -1314 1652 -1280
rect 1698 -1314 1732 -1280
rect 1778 -1314 1812 -1280
rect 1858 -1314 1892 -1280
rect 1938 -1314 1972 -1280
rect 2018 -1314 2052 -1280
rect 2098 -1314 2132 -1280
rect 2178 -1314 2212 -1280
rect -304 -1424 -270 -1390
rect 28 -1444 62 -1410
rect 4356 -1407 4390 -1373
rect -874 -1584 -840 -1550
rect 28 -1564 62 -1530
rect 758 -1534 792 -1500
rect 758 -1614 792 -1580
rect -1102 -1704 -1068 -1670
rect 28 -1684 62 -1650
rect 758 -1694 792 -1660
rect 1058 -1534 1092 -1500
rect 1058 -1614 1092 -1580
rect 1058 -1694 1092 -1660
rect 1358 -1534 1392 -1500
rect 1358 -1614 1392 -1580
rect 2629 -1633 2663 -1599
rect 2709 -1633 2743 -1599
rect 2789 -1633 2823 -1599
rect 2869 -1633 2903 -1599
rect 2949 -1633 2983 -1599
rect 3029 -1633 3063 -1599
rect 3109 -1633 3143 -1599
rect 3189 -1633 3223 -1599
rect 3269 -1633 3303 -1599
rect 3349 -1633 3383 -1599
rect 3429 -1633 3463 -1599
rect 3509 -1633 3543 -1599
rect 3589 -1633 3623 -1599
rect 3669 -1633 3703 -1599
rect 3749 -1633 3783 -1599
rect 3829 -1633 3863 -1599
rect 3909 -1633 3943 -1599
rect 1358 -1694 1392 -1660
rect -646 -1824 -612 -1790
rect 28 -1804 62 -1770
rect -418 -1904 -384 -1870
rect 1108 -1904 1142 -1870
rect -760 -1984 -726 -1950
rect -988 -2084 -954 -2050
rect -532 -2224 -498 -2190
rect 6392 -1439 6426 -1405
rect 4368 -1633 4402 -1599
rect 4448 -1633 4482 -1599
rect 4528 -1633 4562 -1599
rect 4608 -1633 4642 -1599
rect 4688 -1633 4722 -1599
rect 4768 -1633 4802 -1599
rect 4848 -1633 4882 -1599
rect 4928 -1633 4962 -1599
rect 5008 -1633 5042 -1599
rect 5088 -1633 5122 -1599
rect 5168 -1633 5202 -1599
rect 5248 -1633 5282 -1599
rect 5328 -1633 5362 -1599
rect 5408 -1633 5442 -1599
rect 5488 -1633 5522 -1599
rect 5568 -1633 5602 -1599
rect 5648 -1633 5682 -1599
rect 5728 -1633 5762 -1599
rect 5808 -1633 5842 -1599
rect 5888 -1633 5922 -1599
rect 5968 -1633 6002 -1599
rect 6048 -1633 6082 -1599
rect 6128 -1633 6162 -1599
rect 6208 -1633 6242 -1599
rect 6288 -1633 6322 -1599
rect 4498 -1763 4532 -1729
rect 1308 -1904 1342 -1870
rect 2238 -1903 2272 -1869
rect 2969 -1853 3003 -1819
rect 2969 -1933 3003 -1899
rect 2819 -2013 2853 -1979
rect 2969 -2013 3003 -1979
rect 3269 -1853 3303 -1819
rect 3269 -1933 3303 -1899
rect 3269 -2013 3303 -1979
rect 3569 -1853 3603 -1819
rect 5778 -1763 5812 -1729
rect 6170 -1763 6204 -1729
rect 4013 -1840 4047 -1806
rect 3569 -1933 3603 -1899
rect 4610 -1883 4644 -1849
rect 5028 -1853 5062 -1819
rect 3569 -2013 3603 -1979
rect 3719 -2013 3753 -1979
rect 4298 -2025 4332 -1991
rect 4798 -1973 4832 -1939
rect 5028 -1933 5062 -1899
rect 5028 -2013 5062 -1979
rect 3319 -2133 3353 -2099
rect 1588 -2204 1622 -2170
rect 1738 -2204 1772 -2170
rect 1888 -2204 1922 -2170
rect 2038 -2204 2072 -2170
rect 2531 -2253 2565 -2219
rect 5328 -1853 5362 -1819
rect 5328 -1933 5362 -1899
rect 5328 -2013 5362 -1979
rect 5628 -1853 5662 -1819
rect 5898 -1873 5932 -1839
rect 6030 -1874 6064 -1840
rect 5628 -1933 5662 -1899
rect 5628 -2013 5662 -1979
rect 5778 -1973 5812 -1939
rect 3719 -2133 3753 -2099
rect 4298 -2153 4332 -2119
rect 4878 -2133 4912 -2099
rect 5278 -2133 5312 -2099
rect 6392 -2060 6426 -2026
rect 4013 -2303 4047 -2269
rect 4298 -2273 4332 -2239
rect 128 -2414 162 -2380
rect 128 -2494 162 -2460
rect 128 -2574 162 -2540
rect 428 -2414 462 -2380
rect 428 -2494 462 -2460
rect 428 -2574 462 -2540
rect 758 -2414 792 -2380
rect 758 -2494 792 -2460
rect 758 -2574 792 -2540
rect 1058 -2414 1092 -2380
rect 1058 -2494 1092 -2460
rect 1058 -2574 1092 -2540
rect 1358 -2414 1392 -2380
rect 1358 -2494 1392 -2460
rect 1358 -2574 1392 -2540
rect 2138 -2414 2172 -2380
rect 2138 -2494 2172 -2460
rect 2138 -2574 2172 -2540
rect 2639 -2413 2673 -2379
rect 2639 -2493 2673 -2459
rect 2639 -2573 2673 -2539
rect 2969 -2413 3003 -2379
rect 2969 -2493 3003 -2459
rect 2969 -2573 3003 -2539
rect 3269 -2413 3303 -2379
rect 3269 -2493 3303 -2459
rect 3269 -2573 3303 -2539
rect 5908 -2263 5942 -2229
rect 3569 -2413 3603 -2379
rect 3569 -2493 3603 -2459
rect 3569 -2573 3603 -2539
rect 3899 -2413 3933 -2379
rect 3899 -2493 3933 -2459
rect 3899 -2573 3933 -2539
rect 4398 -2413 4432 -2379
rect 4398 -2493 4432 -2459
rect 4398 -2573 4432 -2539
rect 4698 -2413 4732 -2379
rect 4698 -2493 4732 -2459
rect 4698 -2573 4732 -2539
rect 5028 -2413 5062 -2379
rect 5028 -2493 5062 -2459
rect 5028 -2573 5062 -2539
rect 5328 -2413 5362 -2379
rect 5328 -2493 5362 -2459
rect 5328 -2573 5362 -2539
rect 5628 -2413 5662 -2379
rect 5628 -2493 5662 -2459
rect 5628 -2573 5662 -2539
rect 6258 -2413 6292 -2379
rect 6258 -2493 6292 -2459
rect 6258 -2573 6292 -2539
rect -60 -2693 -26 -2659
rect 4013 -2693 4047 -2659
rect 4210 -2693 4244 -2659
rect -190 -2814 -156 -2780
rect -62 -2814 -28 -2780
rect 18 -2814 52 -2780
rect 98 -2814 132 -2780
rect 178 -2814 212 -2780
rect 258 -2814 292 -2780
rect 338 -2814 372 -2780
rect 418 -2814 452 -2780
rect 498 -2814 532 -2780
rect 578 -2814 612 -2780
rect 658 -2814 692 -2780
rect 738 -2814 772 -2780
rect 818 -2814 852 -2780
rect 898 -2814 932 -2780
rect 978 -2814 1012 -2780
rect 1058 -2814 1092 -2780
rect 1138 -2814 1172 -2780
rect 1218 -2814 1252 -2780
rect 1298 -2814 1332 -2780
rect 1378 -2814 1412 -2780
rect 1458 -2814 1492 -2780
rect 1538 -2814 1572 -2780
rect 1618 -2814 1652 -2780
rect 1698 -2814 1732 -2780
rect 1778 -2814 1812 -2780
rect 1858 -2814 1892 -2780
rect 1938 -2814 1972 -2780
rect 2018 -2814 2052 -2780
rect 2098 -2814 2132 -2780
rect 2178 -2814 2212 -2780
rect 2629 -2813 2663 -2779
rect 2709 -2813 2743 -2779
rect 2789 -2813 2823 -2779
rect 2869 -2813 2903 -2779
rect 2949 -2813 2983 -2779
rect 3029 -2813 3063 -2779
rect 3109 -2813 3143 -2779
rect 3189 -2813 3223 -2779
rect 3269 -2813 3303 -2779
rect 3349 -2813 3383 -2779
rect 3429 -2813 3463 -2779
rect 3509 -2813 3543 -2779
rect 3589 -2813 3623 -2779
rect 3669 -2813 3703 -2779
rect 3749 -2813 3783 -2779
rect 3829 -2813 3863 -2779
rect 3909 -2813 3943 -2779
rect 4368 -2813 4402 -2779
rect 4448 -2813 4482 -2779
rect 4528 -2813 4562 -2779
rect 4608 -2813 4642 -2779
rect 4688 -2813 4722 -2779
rect 4768 -2813 4802 -2779
rect 4848 -2813 4882 -2779
rect 4928 -2813 4962 -2779
rect 5008 -2813 5042 -2779
rect 5088 -2813 5122 -2779
rect 5168 -2813 5202 -2779
rect 5248 -2813 5282 -2779
rect 5328 -2813 5362 -2779
rect 5408 -2813 5442 -2779
rect 5488 -2813 5522 -2779
rect 5568 -2813 5602 -2779
rect 5648 -2813 5682 -2779
rect 5728 -2813 5762 -2779
rect 5808 -2813 5842 -2779
rect 5888 -2813 5922 -2779
rect 5968 -2813 6002 -2779
rect 6048 -2813 6082 -2779
rect 6128 -2813 6162 -2779
rect 6208 -2813 6242 -2779
rect 6288 -2813 6322 -2779
<< metal1 >>
rect -65 1230 3975 1254
rect -65 1178 9 1230
rect 61 1221 3975 1230
rect 61 1187 98 1221
rect 132 1187 178 1221
rect 212 1187 258 1221
rect 292 1187 338 1221
rect 372 1187 418 1221
rect 452 1187 498 1221
rect 532 1187 578 1221
rect 612 1187 658 1221
rect 692 1187 738 1221
rect 772 1187 818 1221
rect 852 1187 898 1221
rect 932 1187 978 1221
rect 1012 1187 1058 1221
rect 1092 1187 1138 1221
rect 1172 1187 1218 1221
rect 1252 1187 1298 1221
rect 1332 1187 1378 1221
rect 1412 1187 1458 1221
rect 1492 1187 1538 1221
rect 1572 1187 1618 1221
rect 1652 1187 1698 1221
rect 1732 1187 1778 1221
rect 1812 1187 1858 1221
rect 1892 1187 1938 1221
rect 1972 1187 2018 1221
rect 2052 1187 2098 1221
rect 2132 1187 2628 1221
rect 2662 1187 2708 1221
rect 2742 1187 2788 1221
rect 2822 1187 2868 1221
rect 2902 1187 2948 1221
rect 2982 1187 3028 1221
rect 3062 1187 3108 1221
rect 3142 1187 3188 1221
rect 3222 1187 3268 1221
rect 3302 1187 3348 1221
rect 3382 1187 3428 1221
rect 3462 1187 3508 1221
rect 3542 1187 3588 1221
rect 3622 1187 3668 1221
rect 3702 1187 3748 1221
rect 3782 1187 3828 1221
rect 3862 1187 3908 1221
rect 3942 1187 3975 1221
rect 61 1178 3975 1187
rect -65 1154 3975 1178
rect 4325 1230 6005 1254
rect 4325 1221 4579 1230
rect 4631 1221 6005 1230
rect 4325 1187 4348 1221
rect 4382 1187 4428 1221
rect 4462 1187 4508 1221
rect 4542 1187 4579 1221
rect 4631 1187 4668 1221
rect 4702 1187 4748 1221
rect 4782 1187 4828 1221
rect 4862 1187 4908 1221
rect 4942 1187 4988 1221
rect 5022 1187 5068 1221
rect 5102 1187 5148 1221
rect 5182 1187 5228 1221
rect 5262 1187 5308 1221
rect 5342 1187 5388 1221
rect 5422 1187 5468 1221
rect 5502 1187 5548 1221
rect 5582 1187 5628 1221
rect 5662 1187 5708 1221
rect 5742 1187 5788 1221
rect 5822 1187 5868 1221
rect 5902 1187 5948 1221
rect 5982 1187 6005 1221
rect 4325 1178 4579 1187
rect 4631 1178 6005 1187
rect 4325 1154 6005 1178
rect -783 1103 -703 1116
rect -1125 -808 -1045 1094
rect -1125 -842 -1102 -808
rect -1068 -842 -1045 -808
rect -1125 -1670 -1045 -842
rect -1125 -1704 -1102 -1670
rect -1068 -1704 -1045 -1670
rect -1125 -2836 -1045 -1704
rect -1011 -689 -931 1094
rect -1011 -723 -988 -689
rect -954 -723 -931 -689
rect -1011 -2050 -931 -723
rect -1011 -2084 -988 -2050
rect -954 -2084 -931 -2050
rect -1011 -2836 -931 -2084
rect -897 368 -817 1094
rect -897 316 -883 368
rect -831 316 -817 368
rect -897 -1029 -817 316
rect -897 -1063 -874 -1029
rect -840 -1063 -817 -1029
rect -897 -1550 -817 -1063
rect -897 -1584 -874 -1550
rect -840 -1584 -817 -1550
rect -897 -2837 -817 -1584
rect -783 1051 -769 1103
rect -717 1051 -703 1103
rect -783 -915 -703 1051
rect -783 -949 -760 -915
rect -726 -949 -703 -915
rect -783 -1950 -703 -949
rect -783 -1984 -760 -1950
rect -726 -1984 -703 -1950
rect -783 -2837 -703 -1984
rect -669 871 -589 1094
rect -669 837 -646 871
rect -612 837 -589 871
rect -669 -270 -589 837
rect -669 -322 -655 -270
rect -603 -322 -589 -270
rect -669 -1790 -589 -322
rect -669 -1824 -646 -1790
rect -612 -1824 -589 -1790
rect -669 -2837 -589 -1824
rect -555 771 -475 1094
rect -555 737 -532 771
rect -498 737 -475 771
rect -555 -1001 -475 737
rect -555 -1053 -541 -1001
rect -489 -1053 -475 -1001
rect -555 -2190 -475 -1053
rect -555 -2224 -532 -2190
rect -498 -2224 -475 -2190
rect -555 -2837 -475 -2224
rect -441 1071 -361 1094
rect -441 1037 -418 1071
rect -384 1037 -361 1071
rect -441 -1870 -361 1037
rect -441 -1904 -418 -1870
rect -384 -1904 -361 -1870
rect -441 -2837 -361 -1904
rect -327 989 -247 1094
rect -327 955 -304 989
rect -270 955 -247 989
rect -327 -1390 -247 955
rect -327 -1424 -304 -1390
rect -270 -1424 -247 -1390
rect -327 -2837 -247 -1424
rect -213 41 -133 1094
rect 275 474 315 1154
rect 455 1100 535 1114
rect 455 1048 469 1100
rect 521 1048 535 1100
rect 455 1034 535 1048
rect 585 1000 665 1014
rect 585 948 599 1000
rect 651 948 665 1000
rect 585 934 665 948
rect 735 1001 815 1154
rect 735 967 758 1001
rect 792 967 815 1001
rect 735 921 815 967
rect 455 900 535 914
rect 455 848 469 900
rect 521 848 535 900
rect 455 834 535 848
rect 735 887 758 921
rect 792 887 815 921
rect 735 841 815 887
rect 585 800 665 814
rect 585 748 599 800
rect 651 748 665 800
rect 735 807 758 841
rect 792 807 815 841
rect 735 784 815 807
rect 1035 1001 1115 1154
rect 1035 967 1058 1001
rect 1092 967 1115 1001
rect 1035 921 1115 967
rect 1035 887 1058 921
rect 1092 887 1115 921
rect 1035 841 1115 887
rect 1035 807 1058 841
rect 1092 807 1115 841
rect 1035 784 1115 807
rect 1335 1001 1415 1154
rect 1715 1100 1795 1114
rect 1715 1048 1729 1100
rect 1781 1048 1795 1100
rect 1715 1034 1795 1048
rect 1335 967 1358 1001
rect 1392 967 1415 1001
rect 1335 921 1415 967
rect 1335 887 1358 921
rect 1392 887 1415 921
rect 1335 841 1415 887
rect 1335 807 1358 841
rect 1392 807 1415 841
rect 1335 784 1415 807
rect 1615 800 1695 814
rect 585 734 665 748
rect 1615 748 1629 800
rect 1681 748 1695 800
rect 1085 721 1165 744
rect 1615 734 1695 748
rect 1085 687 1108 721
rect 1142 704 1165 721
rect 1455 711 1535 734
rect 1455 704 1478 711
rect 1142 687 1478 704
rect 1085 677 1478 687
rect 1512 677 1535 711
rect 1085 664 1535 677
rect 1455 654 1535 664
rect 1835 474 1875 1154
rect 2507 1034 2587 1048
rect 1915 1000 1995 1014
rect 1915 948 1929 1000
rect 1981 948 1995 1000
rect 2507 982 2521 1034
rect 2573 982 2587 1034
rect 2507 968 2587 982
rect 1915 934 1995 948
rect 2507 926 2587 940
rect 2065 900 2145 914
rect 2065 848 2079 900
rect 2131 848 2145 900
rect 2507 874 2521 926
rect 2573 874 2587 926
rect 2507 860 2587 874
rect 2065 834 2145 848
rect 2215 599 2295 620
rect 2527 599 2567 860
rect 2215 597 2567 599
rect 2215 563 2238 597
rect 2272 563 2567 597
rect 2215 559 2567 563
rect 2215 540 2295 559
rect 255 441 335 474
rect 255 407 278 441
rect 312 407 335 441
rect 255 361 335 407
rect 255 327 278 361
rect 312 327 335 361
rect 255 281 335 327
rect 255 247 278 281
rect 312 247 335 281
rect 255 224 335 247
rect 735 441 815 474
rect 735 407 758 441
rect 792 407 815 441
rect 735 361 815 407
rect 735 327 758 361
rect 792 327 815 361
rect 735 281 815 327
rect 735 247 758 281
rect 792 247 815 281
rect 735 224 815 247
rect 1035 441 1115 474
rect 1035 407 1058 441
rect 1092 407 1115 441
rect 1035 361 1115 407
rect 1035 327 1058 361
rect 1092 327 1115 361
rect 1035 281 1115 327
rect 1035 247 1058 281
rect 1092 247 1115 281
rect 1035 224 1115 247
rect 1335 441 1415 474
rect 1335 407 1358 441
rect 1392 407 1415 441
rect 1335 361 1415 407
rect 1335 327 1358 361
rect 1392 327 1415 361
rect 1335 281 1415 327
rect 1335 247 1358 281
rect 1392 247 1415 281
rect 1335 224 1415 247
rect 1815 441 1895 474
rect 1815 407 1838 441
rect 1872 407 1895 441
rect 1815 361 1895 407
rect 2615 441 2695 1154
rect 2795 1103 2875 1116
rect 2795 1051 2809 1103
rect 2861 1051 2875 1103
rect 2795 1036 2875 1051
rect 2815 864 2855 1036
rect 2945 1001 3025 1154
rect 2945 967 2968 1001
rect 3002 967 3025 1001
rect 2945 921 3025 967
rect 2945 887 2968 921
rect 3002 887 3025 921
rect 2795 850 2875 864
rect 2795 798 2809 850
rect 2861 798 2875 850
rect 2795 784 2875 798
rect 2945 841 3025 887
rect 2945 807 2968 841
rect 3002 807 3025 841
rect 2945 784 3025 807
rect 3245 1001 3325 1154
rect 3245 967 3268 1001
rect 3302 967 3325 1001
rect 3245 921 3325 967
rect 3245 887 3268 921
rect 3302 887 3325 921
rect 3245 841 3325 887
rect 3245 807 3268 841
rect 3302 807 3325 841
rect 3245 784 3325 807
rect 3545 1001 3625 1154
rect 3545 967 3568 1001
rect 3602 967 3625 1001
rect 3545 921 3625 967
rect 3545 887 3568 921
rect 3602 887 3625 921
rect 3545 841 3625 887
rect 3545 807 3568 841
rect 3602 807 3625 841
rect 3545 784 3625 807
rect 3695 850 3775 864
rect 3695 798 3709 850
rect 3761 798 3775 850
rect 3695 784 3775 798
rect 3295 724 3375 744
rect 3695 724 3775 744
rect 3295 721 3775 724
rect 3295 687 3318 721
rect 3352 687 3718 721
rect 3752 687 3775 721
rect 3295 684 3775 687
rect 3295 664 3375 684
rect 3695 664 3775 684
rect 2615 407 2638 441
rect 2672 407 2695 441
rect 1815 327 1838 361
rect 1872 327 1895 361
rect 1815 290 1895 327
rect 2229 368 2309 381
rect 2229 316 2243 368
rect 2295 316 2309 368
rect 2229 301 2309 316
rect 2615 361 2695 407
rect 2615 327 2638 361
rect 2672 327 2695 361
rect 1815 238 1829 290
rect 1881 238 1895 290
rect 1815 224 1895 238
rect 2615 281 2695 327
rect 2615 247 2638 281
rect 2672 247 2695 281
rect 2615 224 2695 247
rect 2945 441 3025 474
rect 2945 407 2968 441
rect 3002 407 3025 441
rect 2945 361 3025 407
rect 2945 327 2968 361
rect 3002 327 3025 361
rect 2945 281 3025 327
rect 2945 247 2968 281
rect 3002 247 3025 281
rect 2945 224 3025 247
rect 3245 441 3325 474
rect 3245 407 3268 441
rect 3302 407 3325 441
rect 3245 361 3325 407
rect 3245 327 3268 361
rect 3302 327 3325 361
rect 3245 281 3325 327
rect 3245 247 3268 281
rect 3302 247 3325 281
rect 3245 224 3325 247
rect 3545 441 3625 474
rect 3545 407 3568 441
rect 3602 407 3625 441
rect 3545 361 3625 407
rect 3545 327 3568 361
rect 3602 327 3625 361
rect 3545 281 3625 327
rect 3545 247 3568 281
rect 3602 247 3625 281
rect 3545 224 3625 247
rect 3875 441 3955 1154
rect 3983 1034 4063 1048
rect 3983 982 3997 1034
rect 4049 982 4063 1034
rect 3983 968 4063 982
rect 3983 919 4063 933
rect 3983 867 3997 919
rect 4049 867 4063 919
rect 3983 853 4063 867
rect 4245 891 4325 914
rect 4245 857 4268 891
rect 4302 857 4325 891
rect 4245 834 4325 857
rect 3983 574 4063 594
rect 4265 574 4305 834
rect 3983 571 4305 574
rect 3983 537 4006 571
rect 4040 537 4305 571
rect 3983 534 4305 537
rect 3983 514 4063 534
rect 4515 474 4555 1154
rect 4675 1000 4755 1014
rect 4675 948 4689 1000
rect 4741 948 4755 1000
rect 4675 934 4755 948
rect 4825 1001 4905 1154
rect 4825 967 4848 1001
rect 4882 967 4905 1001
rect 4825 921 4905 967
rect 4675 880 4755 894
rect 4675 828 4689 880
rect 4741 828 4755 880
rect 4675 814 4755 828
rect 4825 887 4848 921
rect 4882 887 4905 921
rect 4825 841 4905 887
rect 4825 807 4848 841
rect 4882 807 4905 841
rect 4825 784 4905 807
rect 5125 1001 5205 1154
rect 5125 967 5148 1001
rect 5182 967 5205 1001
rect 5125 921 5205 967
rect 5125 887 5148 921
rect 5182 887 5205 921
rect 5125 841 5205 887
rect 5125 807 5148 841
rect 5182 807 5205 841
rect 5125 784 5205 807
rect 5425 1001 5505 1154
rect 5425 967 5448 1001
rect 5482 967 5505 1001
rect 5425 921 5505 967
rect 5805 1000 5885 1014
rect 5805 948 5819 1000
rect 5871 948 5885 1000
rect 5805 934 5885 948
rect 5425 887 5448 921
rect 5482 887 5505 921
rect 5425 841 5505 887
rect 5425 807 5448 841
rect 5482 807 5505 841
rect 5655 880 5735 894
rect 5655 828 5669 880
rect 5721 828 5735 880
rect 5655 814 5735 828
rect 5425 784 5505 807
rect 5175 724 5255 744
rect 5575 724 5655 744
rect 5175 721 5655 724
rect 5175 687 5198 721
rect 5232 687 5598 721
rect 5632 687 5655 721
rect 5175 684 5655 687
rect 5175 664 5255 684
rect 5575 664 5655 684
rect 5925 474 5965 1154
rect 6008 609 6088 623
rect 6008 557 6022 609
rect 6074 557 6088 609
rect 6008 543 6088 557
rect 3875 407 3898 441
rect 3932 407 3955 441
rect 3875 361 3955 407
rect 3875 327 3898 361
rect 3932 327 3955 361
rect 3875 281 3955 327
rect 3875 247 3898 281
rect 3932 247 3955 281
rect 3875 224 3955 247
rect 4495 441 4575 474
rect 4495 407 4518 441
rect 4552 407 4575 441
rect 4495 361 4575 407
rect 4495 327 4518 361
rect 4552 327 4575 361
rect 4495 281 4575 327
rect 4495 247 4518 281
rect 4552 247 4575 281
rect 4495 224 4575 247
rect 4825 441 4905 474
rect 4825 407 4848 441
rect 4882 407 4905 441
rect 4825 361 4905 407
rect 4825 327 4848 361
rect 4882 327 4905 361
rect 4825 281 4905 327
rect 4825 247 4848 281
rect 4882 247 4905 281
rect 4825 224 4905 247
rect 5125 441 5205 474
rect 5125 407 5148 441
rect 5182 407 5205 441
rect 5125 361 5205 407
rect 5125 327 5148 361
rect 5182 327 5205 361
rect 5125 281 5205 327
rect 5125 247 5148 281
rect 5182 247 5205 281
rect 5125 224 5205 247
rect 5425 441 5505 474
rect 5425 407 5448 441
rect 5482 407 5505 441
rect 5425 361 5505 407
rect 5425 327 5448 361
rect 5482 327 5505 361
rect 5425 281 5505 327
rect 5425 247 5448 281
rect 5482 247 5505 281
rect 5425 224 5505 247
rect 5905 441 5985 474
rect 5905 407 5928 441
rect 5962 407 5985 441
rect 5905 361 5985 407
rect 5905 327 5928 361
rect 5962 327 5985 361
rect 5905 290 5985 327
rect 5905 238 5919 290
rect 5971 238 5985 290
rect 5905 224 5985 238
rect 367 170 447 184
rect 367 118 381 170
rect 433 118 447 170
rect 367 104 447 118
rect 755 74 795 224
rect 1055 74 1095 224
rect 1355 74 1395 224
rect 2965 74 3005 224
rect 3265 74 3305 224
rect 3565 74 3605 224
rect 4333 170 4413 184
rect 4333 118 4347 170
rect 4399 118 4413 170
rect 4333 104 4413 118
rect 4845 74 4885 224
rect 5145 74 5185 224
rect 5445 74 5485 224
rect -213 7 -190 41
rect -156 7 -133 41
rect -213 -2780 -133 7
rect -65 41 6005 74
rect -65 7 18 41
rect 52 7 98 41
rect 132 7 178 41
rect 212 7 258 41
rect 292 7 338 41
rect 372 7 418 41
rect 452 7 498 41
rect 532 7 578 41
rect 612 7 658 41
rect 692 7 738 41
rect 772 7 818 41
rect 852 7 898 41
rect 932 7 978 41
rect 1012 7 1058 41
rect 1092 7 1138 41
rect 1172 7 1218 41
rect 1252 7 1298 41
rect 1332 7 1378 41
rect 1412 7 1458 41
rect 1492 7 1538 41
rect 1572 7 1618 41
rect 1652 7 1698 41
rect 1732 7 1778 41
rect 1812 7 1858 41
rect 1892 7 1938 41
rect 1972 7 2018 41
rect 2052 7 2098 41
rect 2132 7 2628 41
rect 2662 7 2708 41
rect 2742 7 2788 41
rect 2822 7 2868 41
rect 2902 7 2948 41
rect 2982 7 3028 41
rect 3062 7 3108 41
rect 3142 7 3188 41
rect 3222 7 3268 41
rect 3302 7 3348 41
rect 3382 7 3428 41
rect 3462 7 3508 41
rect 3542 7 3588 41
rect 3622 7 3668 41
rect 3702 7 3748 41
rect 3782 7 3828 41
rect 3862 7 3908 41
rect 3942 7 4348 41
rect 4382 7 4428 41
rect 4462 7 4508 41
rect 4542 7 4588 41
rect 4622 7 4668 41
rect 4702 7 4748 41
rect 4782 7 4828 41
rect 4862 7 4908 41
rect 4942 7 4988 41
rect 5022 7 5068 41
rect 5102 7 5148 41
rect 5182 7 5228 41
rect 5262 7 5308 41
rect 5342 7 5388 41
rect 5422 7 5468 41
rect 5502 7 5548 41
rect 5582 7 5628 41
rect 5662 7 5708 41
rect 5742 7 5788 41
rect 5822 7 5868 41
rect 5902 7 5948 41
rect 5982 7 6005 41
rect -65 -26 6005 7
rect 367 -70 447 -56
rect 367 -122 381 -70
rect 433 -122 447 -70
rect 367 -136 447 -122
rect 755 -176 795 -26
rect 1055 -176 1095 -26
rect 1355 -176 1395 -26
rect 2965 -176 3005 -26
rect 3265 -176 3305 -26
rect 3565 -176 3605 -26
rect 4333 -70 4413 -56
rect 4333 -122 4347 -70
rect 4399 -122 4413 -70
rect 4333 -136 4413 -122
rect 4845 -176 4885 -26
rect 5145 -176 5185 -26
rect 5445 -176 5485 -26
rect 255 -199 335 -176
rect 255 -233 278 -199
rect 312 -233 335 -199
rect 255 -279 335 -233
rect 255 -313 278 -279
rect 312 -313 335 -279
rect 255 -359 335 -313
rect 255 -393 278 -359
rect 312 -393 335 -359
rect 255 -426 335 -393
rect 735 -199 815 -176
rect 735 -233 758 -199
rect 792 -233 815 -199
rect 735 -279 815 -233
rect 735 -313 758 -279
rect 792 -313 815 -279
rect 735 -359 815 -313
rect 735 -393 758 -359
rect 792 -393 815 -359
rect 735 -426 815 -393
rect 1035 -199 1115 -176
rect 1035 -233 1058 -199
rect 1092 -233 1115 -199
rect 1035 -279 1115 -233
rect 1035 -313 1058 -279
rect 1092 -313 1115 -279
rect 1035 -359 1115 -313
rect 1035 -393 1058 -359
rect 1092 -393 1115 -359
rect 1035 -426 1115 -393
rect 1335 -199 1415 -176
rect 1335 -233 1358 -199
rect 1392 -233 1415 -199
rect 1335 -279 1415 -233
rect 1335 -313 1358 -279
rect 1392 -313 1415 -279
rect 1335 -359 1415 -313
rect 1335 -393 1358 -359
rect 1392 -393 1415 -359
rect 1335 -426 1415 -393
rect 1815 -190 1895 -176
rect 1815 -242 1829 -190
rect 1881 -242 1895 -190
rect 1815 -279 1895 -242
rect 2615 -199 2695 -176
rect 2615 -233 2638 -199
rect 2672 -233 2695 -199
rect 1815 -313 1838 -279
rect 1872 -313 1895 -279
rect 1815 -359 1895 -313
rect 2229 -270 2309 -257
rect 2229 -322 2243 -270
rect 2295 -322 2309 -270
rect 2229 -337 2309 -322
rect 2615 -279 2695 -233
rect 2615 -313 2638 -279
rect 2672 -313 2695 -279
rect 1815 -393 1838 -359
rect 1872 -393 1895 -359
rect 1815 -426 1895 -393
rect 2506 -341 2586 -327
rect 2506 -393 2520 -341
rect 2572 -393 2586 -341
rect 2506 -407 2586 -393
rect 2615 -359 2695 -313
rect 2615 -393 2638 -359
rect 2672 -393 2695 -359
rect 275 -1106 315 -426
rect 1455 -616 1535 -606
rect 1085 -629 1535 -616
rect 1085 -639 1478 -629
rect 1085 -673 1108 -639
rect 1142 -656 1478 -639
rect 1142 -673 1165 -656
rect 585 -700 665 -686
rect 1085 -696 1165 -673
rect 1455 -663 1478 -656
rect 1512 -663 1535 -629
rect 1455 -686 1535 -663
rect 585 -752 599 -700
rect 651 -752 665 -700
rect 1615 -700 1695 -686
rect 585 -766 665 -752
rect 735 -759 815 -736
rect 455 -800 535 -786
rect 455 -852 469 -800
rect 521 -852 535 -800
rect 455 -866 535 -852
rect 735 -793 758 -759
rect 792 -793 815 -759
rect 735 -839 815 -793
rect 735 -873 758 -839
rect 792 -873 815 -839
rect 585 -900 665 -886
rect 585 -952 599 -900
rect 651 -952 665 -900
rect 585 -966 665 -952
rect 735 -919 815 -873
rect 735 -953 758 -919
rect 792 -953 815 -919
rect 455 -1000 535 -986
rect 455 -1052 469 -1000
rect 521 -1052 535 -1000
rect 455 -1066 535 -1052
rect 735 -1106 815 -953
rect 1035 -759 1115 -736
rect 1035 -793 1058 -759
rect 1092 -793 1115 -759
rect 1035 -839 1115 -793
rect 1035 -873 1058 -839
rect 1092 -873 1115 -839
rect 1035 -919 1115 -873
rect 1035 -953 1058 -919
rect 1092 -953 1115 -919
rect 1035 -1106 1115 -953
rect 1335 -759 1415 -736
rect 1335 -793 1358 -759
rect 1392 -793 1415 -759
rect 1615 -752 1629 -700
rect 1681 -752 1695 -700
rect 1615 -766 1695 -752
rect 1335 -839 1415 -793
rect 1335 -873 1358 -839
rect 1392 -873 1415 -839
rect 1335 -919 1415 -873
rect 1335 -953 1358 -919
rect 1392 -953 1415 -919
rect 1335 -1106 1415 -953
rect 1715 -1000 1795 -986
rect 1715 -1052 1729 -1000
rect 1781 -1052 1795 -1000
rect 1715 -1066 1795 -1052
rect 1835 -1106 1875 -426
rect 2215 -629 2295 -606
rect 2215 -663 2238 -629
rect 2272 -646 2295 -629
rect 2527 -646 2567 -407
rect 2272 -663 2567 -646
rect 2215 -686 2567 -663
rect 2065 -800 2145 -786
rect 2065 -852 2079 -800
rect 2131 -852 2145 -800
rect 2065 -866 2145 -852
rect 1915 -900 1995 -886
rect 1915 -952 1929 -900
rect 1981 -952 1995 -900
rect 1915 -966 1995 -952
rect 2507 -900 2587 -886
rect 2507 -952 2521 -900
rect 2573 -952 2587 -900
rect 2507 -966 2587 -952
rect 2615 -1106 2695 -393
rect 2945 -199 3025 -176
rect 2945 -233 2968 -199
rect 3002 -233 3025 -199
rect 2945 -279 3025 -233
rect 2945 -313 2968 -279
rect 3002 -313 3025 -279
rect 2945 -359 3025 -313
rect 2945 -393 2968 -359
rect 3002 -393 3025 -359
rect 2945 -426 3025 -393
rect 3245 -199 3325 -176
rect 3245 -233 3268 -199
rect 3302 -233 3325 -199
rect 3245 -279 3325 -233
rect 3245 -313 3268 -279
rect 3302 -313 3325 -279
rect 3245 -359 3325 -313
rect 3245 -393 3268 -359
rect 3302 -393 3325 -359
rect 3245 -426 3325 -393
rect 3545 -199 3625 -176
rect 3545 -233 3568 -199
rect 3602 -233 3625 -199
rect 3545 -279 3625 -233
rect 3545 -313 3568 -279
rect 3602 -313 3625 -279
rect 3545 -359 3625 -313
rect 3545 -393 3568 -359
rect 3602 -393 3625 -359
rect 3545 -426 3625 -393
rect 3875 -199 3955 -176
rect 3875 -233 3898 -199
rect 3932 -233 3955 -199
rect 3875 -279 3955 -233
rect 3875 -313 3898 -279
rect 3932 -313 3955 -279
rect 3875 -359 3955 -313
rect 4495 -199 4575 -176
rect 4495 -233 4518 -199
rect 4552 -233 4575 -199
rect 4495 -279 4575 -233
rect 4495 -313 4518 -279
rect 4552 -313 4575 -279
rect 3875 -393 3898 -359
rect 3932 -393 3955 -359
rect 3295 -636 3375 -616
rect 3695 -636 3775 -616
rect 3295 -639 3775 -636
rect 3295 -673 3318 -639
rect 3352 -673 3718 -639
rect 3752 -673 3775 -639
rect 3295 -676 3775 -673
rect 3295 -696 3375 -676
rect 3695 -696 3775 -676
rect 2795 -750 2875 -736
rect 2795 -802 2809 -750
rect 2861 -802 2875 -750
rect 2795 -816 2875 -802
rect 2945 -759 3025 -736
rect 2945 -793 2968 -759
rect 3002 -793 3025 -759
rect 2815 -988 2855 -816
rect 2945 -839 3025 -793
rect 2945 -873 2968 -839
rect 3002 -873 3025 -839
rect 2945 -919 3025 -873
rect 2945 -953 2968 -919
rect 3002 -953 3025 -919
rect 2795 -1001 2875 -988
rect 2795 -1053 2809 -1001
rect 2861 -1053 2875 -1001
rect 2795 -1068 2875 -1053
rect 2945 -1106 3025 -953
rect 3245 -759 3325 -736
rect 3245 -793 3268 -759
rect 3302 -793 3325 -759
rect 3245 -839 3325 -793
rect 3245 -873 3268 -839
rect 3302 -873 3325 -839
rect 3245 -919 3325 -873
rect 3245 -953 3268 -919
rect 3302 -953 3325 -919
rect 3245 -1106 3325 -953
rect 3545 -759 3625 -736
rect 3545 -793 3568 -759
rect 3602 -793 3625 -759
rect 3545 -839 3625 -793
rect 3695 -750 3775 -736
rect 3695 -802 3709 -750
rect 3761 -802 3775 -750
rect 3695 -816 3775 -802
rect 3545 -873 3568 -839
rect 3602 -873 3625 -839
rect 3545 -919 3625 -873
rect 3545 -953 3568 -919
rect 3602 -953 3625 -919
rect 3545 -1106 3625 -953
rect 3695 -900 3775 -886
rect 3695 -952 3709 -900
rect 3761 -952 3775 -900
rect 3695 -966 3775 -952
rect 3875 -1106 3955 -393
rect 3983 -340 4063 -326
rect 3983 -392 3997 -340
rect 4049 -346 4063 -340
rect 4049 -386 4131 -346
rect 4049 -392 4063 -386
rect 3983 -406 4063 -392
rect 3983 -469 4063 -446
rect 3983 -503 4006 -469
rect 4040 -503 4063 -469
rect 3983 -526 4063 -503
rect 4003 -806 4043 -526
rect 4091 -686 4131 -386
rect 4495 -359 4575 -313
rect 4495 -393 4518 -359
rect 4552 -393 4575 -359
rect 4495 -426 4575 -393
rect 4825 -199 4905 -176
rect 4825 -233 4848 -199
rect 4882 -233 4905 -199
rect 4825 -279 4905 -233
rect 4825 -313 4848 -279
rect 4882 -313 4905 -279
rect 4825 -359 4905 -313
rect 4825 -393 4848 -359
rect 4882 -393 4905 -359
rect 4825 -426 4905 -393
rect 5125 -199 5205 -176
rect 5125 -233 5148 -199
rect 5182 -233 5205 -199
rect 5125 -279 5205 -233
rect 5125 -313 5148 -279
rect 5182 -313 5205 -279
rect 5125 -359 5205 -313
rect 5125 -393 5148 -359
rect 5182 -393 5205 -359
rect 5125 -426 5205 -393
rect 5425 -199 5505 -176
rect 5425 -233 5448 -199
rect 5482 -233 5505 -199
rect 5425 -279 5505 -233
rect 5425 -313 5448 -279
rect 5482 -313 5505 -279
rect 5425 -359 5505 -313
rect 5425 -393 5448 -359
rect 5482 -393 5505 -359
rect 5425 -426 5505 -393
rect 5905 -190 5985 -176
rect 5905 -242 5919 -190
rect 5971 -242 5985 -190
rect 5905 -279 5985 -242
rect 5905 -313 5928 -279
rect 5962 -313 5985 -279
rect 5905 -359 5985 -313
rect 5905 -393 5928 -359
rect 5962 -393 5985 -359
rect 5905 -426 5985 -393
rect 4245 -686 4325 -666
rect 4091 -689 4325 -686
rect 4091 -723 4268 -689
rect 4302 -723 4325 -689
rect 4091 -726 4325 -723
rect 4245 -746 4325 -726
rect 4245 -806 4325 -786
rect 4003 -809 4325 -806
rect 4003 -843 4268 -809
rect 4302 -843 4325 -809
rect 4003 -846 4325 -843
rect 4245 -866 4325 -846
rect 4515 -1106 4555 -426
rect 5175 -636 5255 -616
rect 5575 -636 5655 -616
rect 5175 -639 5655 -636
rect 5175 -673 5198 -639
rect 5232 -673 5598 -639
rect 5632 -673 5655 -639
rect 5175 -676 5655 -673
rect 5175 -696 5255 -676
rect 5575 -696 5655 -676
rect 4825 -759 4905 -736
rect 4675 -780 4755 -766
rect 4675 -832 4689 -780
rect 4741 -832 4755 -780
rect 4675 -846 4755 -832
rect 4825 -793 4848 -759
rect 4882 -793 4905 -759
rect 4825 -839 4905 -793
rect 4825 -873 4848 -839
rect 4882 -873 4905 -839
rect 4675 -900 4755 -886
rect 4675 -952 4689 -900
rect 4741 -952 4755 -900
rect 4675 -966 4755 -952
rect 4825 -919 4905 -873
rect 4825 -953 4848 -919
rect 4882 -953 4905 -919
rect 4825 -1106 4905 -953
rect 5125 -759 5205 -736
rect 5125 -793 5148 -759
rect 5182 -793 5205 -759
rect 5125 -839 5205 -793
rect 5125 -873 5148 -839
rect 5182 -873 5205 -839
rect 5125 -919 5205 -873
rect 5125 -953 5148 -919
rect 5182 -953 5205 -919
rect 5125 -1106 5205 -953
rect 5425 -759 5505 -736
rect 5425 -793 5448 -759
rect 5482 -793 5505 -759
rect 5425 -839 5505 -793
rect 5425 -873 5448 -839
rect 5482 -873 5505 -839
rect 5655 -780 5735 -766
rect 5655 -832 5669 -780
rect 5721 -832 5735 -780
rect 5655 -846 5735 -832
rect 5425 -919 5505 -873
rect 5425 -953 5448 -919
rect 5482 -953 5505 -919
rect 5425 -1106 5505 -953
rect 5805 -900 5885 -886
rect 5805 -952 5819 -900
rect 5871 -952 5885 -900
rect 5805 -966 5885 -952
rect 5925 -1106 5965 -426
rect 6008 -510 6088 -496
rect 6008 -562 6022 -510
rect 6074 -562 6088 -510
rect 6008 -576 6088 -562
rect -85 -1139 3975 -1106
rect -85 -1173 -62 -1139
rect -28 -1173 18 -1139
rect 52 -1173 98 -1139
rect 132 -1173 178 -1139
rect 212 -1173 258 -1139
rect 292 -1173 338 -1139
rect 372 -1173 418 -1139
rect 452 -1173 498 -1139
rect 532 -1173 578 -1139
rect 612 -1173 658 -1139
rect 692 -1173 738 -1139
rect 772 -1173 818 -1139
rect 852 -1173 898 -1139
rect 932 -1173 978 -1139
rect 1012 -1173 1058 -1139
rect 1092 -1173 1138 -1139
rect 1172 -1173 1218 -1139
rect 1252 -1173 1298 -1139
rect 1332 -1173 1378 -1139
rect 1412 -1173 1458 -1139
rect 1492 -1173 1538 -1139
rect 1572 -1173 1618 -1139
rect 1652 -1173 1698 -1139
rect 1732 -1173 1778 -1139
rect 1812 -1173 1858 -1139
rect 1892 -1173 1938 -1139
rect 1972 -1173 2018 -1139
rect 2052 -1173 2098 -1139
rect 2132 -1173 2178 -1139
rect 2212 -1173 2628 -1139
rect 2662 -1173 2708 -1139
rect 2742 -1173 2788 -1139
rect 2822 -1173 2868 -1139
rect 2902 -1173 2948 -1139
rect 2982 -1173 3028 -1139
rect 3062 -1173 3108 -1139
rect 3142 -1173 3188 -1139
rect 3222 -1173 3268 -1139
rect 3302 -1173 3348 -1139
rect 3382 -1173 3428 -1139
rect 3462 -1173 3508 -1139
rect 3542 -1173 3588 -1139
rect 3622 -1173 3668 -1139
rect 3702 -1173 3748 -1139
rect 3782 -1173 3828 -1139
rect 3862 -1173 3908 -1139
rect 3942 -1173 3975 -1139
rect -85 -1206 3975 -1173
rect 4105 -1139 6005 -1106
rect 4105 -1173 4348 -1139
rect 4382 -1173 4428 -1139
rect 4462 -1173 4508 -1139
rect 4542 -1173 4588 -1139
rect 4622 -1173 4668 -1139
rect 4702 -1173 4748 -1139
rect 4782 -1173 4828 -1139
rect 4862 -1173 4908 -1139
rect 4942 -1173 4988 -1139
rect 5022 -1173 5068 -1139
rect 5102 -1173 5148 -1139
rect 5182 -1173 5228 -1139
rect 5262 -1173 5308 -1139
rect 5342 -1173 5388 -1139
rect 5422 -1173 5468 -1139
rect 5502 -1173 5548 -1139
rect 5582 -1173 5628 -1139
rect 5662 -1173 5708 -1139
rect 5742 -1173 5788 -1139
rect 5822 -1173 5868 -1139
rect 5902 -1173 5948 -1139
rect 5982 -1173 6005 -1139
rect 4105 -1206 6005 -1173
rect -85 -1280 2235 -1206
rect -85 -1314 -62 -1280
rect -28 -1314 18 -1280
rect 52 -1314 98 -1280
rect 132 -1314 178 -1280
rect 212 -1314 258 -1280
rect 292 -1314 338 -1280
rect 372 -1314 418 -1280
rect 452 -1314 498 -1280
rect 532 -1314 578 -1280
rect 612 -1314 658 -1280
rect 692 -1314 738 -1280
rect 772 -1314 818 -1280
rect 852 -1314 898 -1280
rect 932 -1314 978 -1280
rect 1012 -1314 1058 -1280
rect 1092 -1314 1138 -1280
rect 1172 -1314 1218 -1280
rect 1252 -1314 1298 -1280
rect 1332 -1314 1378 -1280
rect 1412 -1314 1458 -1280
rect 1492 -1314 1538 -1280
rect 1572 -1314 1618 -1280
rect 1652 -1314 1698 -1280
rect 1732 -1314 1778 -1280
rect 1812 -1314 1858 -1280
rect 1892 -1314 1938 -1280
rect 1972 -1314 2018 -1280
rect 2052 -1314 2098 -1280
rect 2132 -1314 2178 -1280
rect 2212 -1314 2235 -1280
rect -85 -1347 2235 -1314
rect 4105 -1336 4205 -1206
rect 5 -1401 85 -1387
rect 5 -1453 19 -1401
rect 71 -1453 85 -1401
rect 5 -1467 85 -1453
rect 5 -1521 85 -1507
rect 5 -1573 19 -1521
rect 71 -1573 85 -1521
rect 5 -1587 85 -1573
rect 5 -1641 85 -1627
rect 5 -1693 19 -1641
rect 71 -1693 85 -1641
rect 5 -1707 85 -1693
rect 5 -1761 85 -1747
rect 5 -1813 19 -1761
rect 71 -1813 85 -1761
rect 5 -1827 85 -1813
rect 125 -2347 165 -1347
rect 425 -2347 465 -1347
rect 735 -1500 815 -1347
rect 735 -1534 758 -1500
rect 792 -1534 815 -1500
rect 735 -1580 815 -1534
rect 735 -1614 758 -1580
rect 792 -1614 815 -1580
rect 735 -1660 815 -1614
rect 735 -1694 758 -1660
rect 792 -1694 815 -1660
rect 735 -1717 815 -1694
rect 1035 -1500 1115 -1347
rect 1035 -1534 1058 -1500
rect 1092 -1534 1115 -1500
rect 1035 -1580 1115 -1534
rect 1035 -1614 1058 -1580
rect 1092 -1614 1115 -1580
rect 1035 -1660 1115 -1614
rect 1035 -1694 1058 -1660
rect 1092 -1694 1115 -1660
rect 1035 -1717 1115 -1694
rect 1335 -1500 1415 -1347
rect 2015 -1401 2095 -1387
rect 2015 -1453 2029 -1401
rect 2081 -1453 2095 -1401
rect 2015 -1467 2095 -1453
rect 1335 -1534 1358 -1500
rect 1392 -1534 1415 -1500
rect 1335 -1580 1415 -1534
rect 1335 -1614 1358 -1580
rect 1392 -1614 1415 -1580
rect 1865 -1521 1945 -1507
rect 1865 -1573 1879 -1521
rect 1931 -1573 1945 -1521
rect 1865 -1587 1945 -1573
rect 1335 -1660 1415 -1614
rect 1335 -1694 1358 -1660
rect 1392 -1694 1415 -1660
rect 1335 -1717 1415 -1694
rect 1715 -1641 1795 -1627
rect 1715 -1693 1729 -1641
rect 1781 -1693 1795 -1641
rect 1715 -1707 1795 -1693
rect 1565 -1761 1645 -1747
rect 1565 -1813 1579 -1761
rect 1631 -1813 1645 -1761
rect 1565 -1827 1645 -1813
rect 1085 -1867 1165 -1847
rect 1285 -1867 1365 -1847
rect 1085 -1870 1365 -1867
rect 1085 -1904 1108 -1870
rect 1142 -1904 1308 -1870
rect 1342 -1904 1365 -1870
rect 1085 -1907 1365 -1904
rect 1085 -1927 1165 -1907
rect 1285 -1927 1365 -1907
rect 1585 -2147 1625 -1827
rect 1735 -2147 1775 -1707
rect 1885 -2147 1925 -1587
rect 2035 -2147 2075 -1467
rect 1565 -2170 1645 -2147
rect 1565 -2204 1588 -2170
rect 1622 -2204 1645 -2170
rect 1565 -2227 1645 -2204
rect 1715 -2170 1795 -2147
rect 1715 -2204 1738 -2170
rect 1772 -2204 1795 -2170
rect 1715 -2227 1795 -2204
rect 1865 -2170 1945 -2147
rect 1865 -2204 1888 -2170
rect 1922 -2204 1945 -2170
rect 1865 -2227 1945 -2204
rect 2015 -2170 2095 -2147
rect 2015 -2204 2038 -2170
rect 2072 -2204 2095 -2170
rect 2015 -2227 2095 -2204
rect 2135 -2347 2175 -1347
rect 3736 -1436 4205 -1336
rect 4333 -1364 4413 -1350
rect 4333 -1416 4347 -1364
rect 4399 -1416 4413 -1364
rect 4333 -1430 4413 -1416
rect 6369 -1396 6449 -1382
rect 3736 -1566 3836 -1436
rect 6369 -1448 6383 -1396
rect 6435 -1448 6449 -1396
rect 6369 -1462 6449 -1448
rect 2596 -1599 3976 -1566
rect 2596 -1633 2629 -1599
rect 2663 -1633 2709 -1599
rect 2743 -1633 2789 -1599
rect 2823 -1633 2869 -1599
rect 2903 -1633 2949 -1599
rect 2983 -1633 3029 -1599
rect 3063 -1633 3109 -1599
rect 3143 -1633 3189 -1599
rect 3223 -1633 3269 -1599
rect 3303 -1633 3349 -1599
rect 3383 -1633 3429 -1599
rect 3463 -1633 3509 -1599
rect 3543 -1633 3589 -1599
rect 3623 -1633 3669 -1599
rect 3703 -1633 3749 -1599
rect 3783 -1633 3829 -1599
rect 3863 -1633 3909 -1599
rect 3943 -1633 3976 -1599
rect 2596 -1666 3976 -1633
rect 4345 -1590 6345 -1566
rect 4345 -1599 4435 -1590
rect 4487 -1599 6345 -1590
rect 4345 -1633 4368 -1599
rect 4402 -1633 4435 -1599
rect 4487 -1633 4528 -1599
rect 4562 -1633 4608 -1599
rect 4642 -1633 4688 -1599
rect 4722 -1633 4768 -1599
rect 4802 -1633 4848 -1599
rect 4882 -1633 4928 -1599
rect 4962 -1633 5008 -1599
rect 5042 -1633 5088 -1599
rect 5122 -1633 5168 -1599
rect 5202 -1633 5248 -1599
rect 5282 -1633 5328 -1599
rect 5362 -1633 5408 -1599
rect 5442 -1633 5488 -1599
rect 5522 -1633 5568 -1599
rect 5602 -1633 5648 -1599
rect 5682 -1633 5728 -1599
rect 5762 -1633 5808 -1599
rect 5842 -1633 5888 -1599
rect 5922 -1633 5968 -1599
rect 6002 -1633 6048 -1599
rect 6082 -1633 6128 -1599
rect 6162 -1633 6208 -1599
rect 6242 -1633 6288 -1599
rect 6322 -1633 6345 -1599
rect 4345 -1642 4435 -1633
rect 4487 -1642 6345 -1633
rect 4345 -1666 6345 -1642
rect 2215 -1869 2295 -1846
rect 2215 -1903 2238 -1869
rect 2272 -1903 2295 -1869
rect 2215 -1926 2295 -1903
rect 2235 -2216 2275 -1926
rect 2508 -2216 2588 -2196
rect 2235 -2219 2588 -2216
rect 2235 -2253 2531 -2219
rect 2565 -2253 2588 -2219
rect 2235 -2256 2588 -2253
rect 2508 -2276 2588 -2256
rect 105 -2380 185 -2347
rect 105 -2414 128 -2380
rect 162 -2414 185 -2380
rect 105 -2460 185 -2414
rect 105 -2494 128 -2460
rect 162 -2494 185 -2460
rect 105 -2540 185 -2494
rect 105 -2574 128 -2540
rect 162 -2574 185 -2540
rect 105 -2597 185 -2574
rect 405 -2380 485 -2347
rect 405 -2414 428 -2380
rect 462 -2414 485 -2380
rect 405 -2460 485 -2414
rect 405 -2494 428 -2460
rect 462 -2494 485 -2460
rect 405 -2540 485 -2494
rect 405 -2574 428 -2540
rect 462 -2574 485 -2540
rect 405 -2597 485 -2574
rect 735 -2380 815 -2347
rect 735 -2414 758 -2380
rect 792 -2414 815 -2380
rect 735 -2460 815 -2414
rect 735 -2494 758 -2460
rect 792 -2494 815 -2460
rect 735 -2540 815 -2494
rect 735 -2574 758 -2540
rect 792 -2574 815 -2540
rect 735 -2597 815 -2574
rect 1035 -2380 1115 -2347
rect 1035 -2414 1058 -2380
rect 1092 -2414 1115 -2380
rect 1035 -2460 1115 -2414
rect 1035 -2494 1058 -2460
rect 1092 -2494 1115 -2460
rect 1035 -2540 1115 -2494
rect 1035 -2574 1058 -2540
rect 1092 -2574 1115 -2540
rect 1035 -2597 1115 -2574
rect 1335 -2380 1415 -2347
rect 1335 -2414 1358 -2380
rect 1392 -2414 1415 -2380
rect 1335 -2460 1415 -2414
rect 1335 -2494 1358 -2460
rect 1392 -2494 1415 -2460
rect 1335 -2540 1415 -2494
rect 1335 -2574 1358 -2540
rect 1392 -2574 1415 -2540
rect 1335 -2597 1415 -2574
rect 2115 -2380 2195 -2347
rect 2115 -2414 2138 -2380
rect 2172 -2414 2195 -2380
rect 2115 -2460 2195 -2414
rect 2115 -2494 2138 -2460
rect 2172 -2494 2195 -2460
rect 2115 -2540 2195 -2494
rect 2115 -2574 2138 -2540
rect 2172 -2574 2195 -2540
rect 2115 -2597 2195 -2574
rect 2616 -2379 2696 -1666
rect 2946 -1819 3026 -1666
rect 2946 -1853 2969 -1819
rect 3003 -1853 3026 -1819
rect 2946 -1899 3026 -1853
rect 2946 -1933 2969 -1899
rect 3003 -1933 3026 -1899
rect 2796 -1970 2876 -1956
rect 2796 -2022 2810 -1970
rect 2862 -2022 2876 -1970
rect 2796 -2036 2876 -2022
rect 2946 -1979 3026 -1933
rect 2946 -2013 2969 -1979
rect 3003 -2013 3026 -1979
rect 2946 -2036 3026 -2013
rect 3246 -1819 3326 -1666
rect 3246 -1853 3269 -1819
rect 3303 -1853 3326 -1819
rect 3246 -1899 3326 -1853
rect 3246 -1933 3269 -1899
rect 3303 -1933 3326 -1899
rect 3246 -1979 3326 -1933
rect 3246 -2013 3269 -1979
rect 3303 -2013 3326 -1979
rect 3246 -2036 3326 -2013
rect 3546 -1819 3626 -1666
rect 3546 -1853 3569 -1819
rect 3603 -1853 3626 -1819
rect 3546 -1899 3626 -1853
rect 3546 -1933 3569 -1899
rect 3603 -1933 3626 -1899
rect 3546 -1979 3626 -1933
rect 3546 -2013 3569 -1979
rect 3603 -2013 3626 -1979
rect 3546 -2036 3626 -2013
rect 3696 -1970 3776 -1956
rect 3696 -2022 3710 -1970
rect 3762 -2022 3776 -1970
rect 3696 -2036 3776 -2022
rect 3296 -2096 3376 -2076
rect 3696 -2096 3776 -2076
rect 3296 -2099 3776 -2096
rect 3296 -2133 3319 -2099
rect 3353 -2133 3719 -2099
rect 3753 -2133 3776 -2099
rect 3296 -2136 3776 -2133
rect 3296 -2156 3376 -2136
rect 3696 -2156 3776 -2136
rect 2616 -2413 2639 -2379
rect 2673 -2413 2696 -2379
rect 2616 -2459 2696 -2413
rect 2616 -2493 2639 -2459
rect 2673 -2493 2696 -2459
rect 2616 -2539 2696 -2493
rect 2616 -2573 2639 -2539
rect 2673 -2573 2696 -2539
rect 2616 -2596 2696 -2573
rect 2946 -2379 3026 -2346
rect 2946 -2413 2969 -2379
rect 3003 -2413 3026 -2379
rect 2946 -2459 3026 -2413
rect 2946 -2493 2969 -2459
rect 3003 -2493 3026 -2459
rect 2946 -2539 3026 -2493
rect 2946 -2573 2969 -2539
rect 3003 -2573 3026 -2539
rect 2946 -2596 3026 -2573
rect 3246 -2379 3326 -2346
rect 3246 -2413 3269 -2379
rect 3303 -2413 3326 -2379
rect 3246 -2459 3326 -2413
rect 3246 -2493 3269 -2459
rect 3303 -2493 3326 -2459
rect 3246 -2539 3326 -2493
rect 3246 -2573 3269 -2539
rect 3303 -2573 3326 -2539
rect 3246 -2596 3326 -2573
rect 3546 -2379 3626 -2346
rect 3546 -2413 3569 -2379
rect 3603 -2413 3626 -2379
rect 3546 -2459 3626 -2413
rect 3546 -2493 3569 -2459
rect 3603 -2493 3626 -2459
rect 3546 -2539 3626 -2493
rect 3546 -2573 3569 -2539
rect 3603 -2573 3626 -2539
rect 3546 -2596 3626 -2573
rect 3876 -2379 3956 -1666
rect 3990 -1797 4070 -1783
rect 3990 -1849 4004 -1797
rect 4056 -1849 4070 -1797
rect 3990 -1863 4070 -1849
rect 4275 -1867 4355 -1853
rect 4275 -1893 4289 -1867
rect 4010 -1919 4289 -1893
rect 4341 -1919 4355 -1867
rect 4010 -1933 4355 -1919
rect 4010 -2246 4050 -1933
rect 4275 -1982 4355 -1968
rect 4275 -2034 4289 -1982
rect 4341 -2034 4355 -1982
rect 4275 -2048 4355 -2034
rect 4275 -2110 4355 -2096
rect 4275 -2162 4289 -2110
rect 4341 -2162 4355 -2110
rect 4275 -2176 4355 -2162
rect 4275 -2230 4355 -2216
rect 3990 -2269 4070 -2246
rect 3990 -2303 4013 -2269
rect 4047 -2303 4070 -2269
rect 4275 -2282 4289 -2230
rect 4341 -2282 4355 -2230
rect 4275 -2296 4355 -2282
rect 3990 -2326 4070 -2303
rect 4395 -2346 4435 -1666
rect 4475 -1720 4555 -1706
rect 4475 -1772 4489 -1720
rect 4541 -1772 4555 -1720
rect 4475 -1786 4555 -1772
rect 4587 -1840 4667 -1826
rect 4587 -1892 4601 -1840
rect 4653 -1892 4667 -1840
rect 4587 -1906 4667 -1892
rect 4695 -2346 4735 -1666
rect 5005 -1819 5085 -1666
rect 5005 -1853 5028 -1819
rect 5062 -1853 5085 -1819
rect 5005 -1899 5085 -1853
rect 4775 -1930 4855 -1916
rect 4775 -1982 4789 -1930
rect 4841 -1982 4855 -1930
rect 4775 -1996 4855 -1982
rect 5005 -1933 5028 -1899
rect 5062 -1933 5085 -1899
rect 5005 -1979 5085 -1933
rect 5005 -2013 5028 -1979
rect 5062 -2013 5085 -1979
rect 5005 -2036 5085 -2013
rect 5305 -1819 5385 -1666
rect 5305 -1853 5328 -1819
rect 5362 -1853 5385 -1819
rect 5305 -1899 5385 -1853
rect 5305 -1933 5328 -1899
rect 5362 -1933 5385 -1899
rect 5305 -1979 5385 -1933
rect 5305 -2013 5328 -1979
rect 5362 -2013 5385 -1979
rect 5305 -2036 5385 -2013
rect 5605 -1819 5685 -1666
rect 5755 -1720 5835 -1706
rect 5755 -1772 5769 -1720
rect 5821 -1772 5835 -1720
rect 5755 -1786 5835 -1772
rect 6147 -1720 6227 -1706
rect 6147 -1772 6161 -1720
rect 6213 -1772 6227 -1720
rect 6147 -1786 6227 -1772
rect 5605 -1853 5628 -1819
rect 5662 -1853 5685 -1819
rect 5605 -1899 5685 -1853
rect 5875 -1830 5955 -1816
rect 5875 -1882 5889 -1830
rect 5941 -1882 5955 -1830
rect 5875 -1896 5955 -1882
rect 6007 -1831 6087 -1817
rect 6007 -1883 6021 -1831
rect 6073 -1883 6087 -1831
rect 6007 -1897 6087 -1883
rect 5605 -1933 5628 -1899
rect 5662 -1933 5685 -1899
rect 5605 -1979 5685 -1933
rect 5605 -2013 5628 -1979
rect 5662 -2013 5685 -1979
rect 5755 -1930 5835 -1916
rect 5755 -1982 5769 -1930
rect 5821 -1982 5835 -1930
rect 5755 -1996 5835 -1982
rect 5605 -2036 5685 -2013
rect 5885 -2017 5965 -2003
rect 5885 -2069 5899 -2017
rect 5951 -2069 5965 -2017
rect 4855 -2096 4935 -2076
rect 5255 -2096 5335 -2076
rect 5885 -2083 5965 -2069
rect 4855 -2099 5335 -2096
rect 4855 -2133 4878 -2099
rect 4912 -2133 5278 -2099
rect 5312 -2133 5335 -2099
rect 4855 -2136 5335 -2133
rect 4855 -2156 4935 -2136
rect 5255 -2156 5335 -2136
rect 5905 -2206 5945 -2083
rect 5885 -2229 5965 -2206
rect 5885 -2263 5908 -2229
rect 5942 -2263 5965 -2229
rect 5885 -2286 5965 -2263
rect 6255 -2346 6295 -1666
rect 6369 -2017 6449 -2003
rect 6369 -2069 6383 -2017
rect 6435 -2069 6449 -2017
rect 6369 -2083 6449 -2069
rect 3876 -2413 3899 -2379
rect 3933 -2413 3956 -2379
rect 3876 -2459 3956 -2413
rect 3876 -2493 3899 -2459
rect 3933 -2493 3956 -2459
rect 3876 -2539 3956 -2493
rect 3876 -2573 3899 -2539
rect 3933 -2573 3956 -2539
rect 3876 -2596 3956 -2573
rect 4375 -2379 4455 -2346
rect 4375 -2413 4398 -2379
rect 4432 -2413 4455 -2379
rect 4375 -2459 4455 -2413
rect 4375 -2493 4398 -2459
rect 4432 -2493 4455 -2459
rect 4375 -2539 4455 -2493
rect 4375 -2573 4398 -2539
rect 4432 -2573 4455 -2539
rect 4375 -2596 4455 -2573
rect 4675 -2379 4755 -2346
rect 4675 -2413 4698 -2379
rect 4732 -2413 4755 -2379
rect 4675 -2459 4755 -2413
rect 4675 -2493 4698 -2459
rect 4732 -2493 4755 -2459
rect 4675 -2539 4755 -2493
rect 4675 -2573 4698 -2539
rect 4732 -2573 4755 -2539
rect 4675 -2596 4755 -2573
rect 5005 -2379 5085 -2346
rect 5005 -2413 5028 -2379
rect 5062 -2413 5085 -2379
rect 5005 -2459 5085 -2413
rect 5005 -2493 5028 -2459
rect 5062 -2493 5085 -2459
rect 5005 -2539 5085 -2493
rect 5005 -2573 5028 -2539
rect 5062 -2573 5085 -2539
rect 5005 -2596 5085 -2573
rect 5305 -2379 5385 -2346
rect 5305 -2413 5328 -2379
rect 5362 -2413 5385 -2379
rect 5305 -2459 5385 -2413
rect 5305 -2493 5328 -2459
rect 5362 -2493 5385 -2459
rect 5305 -2539 5385 -2493
rect 5305 -2573 5328 -2539
rect 5362 -2573 5385 -2539
rect 5305 -2596 5385 -2573
rect 5605 -2379 5685 -2346
rect 5605 -2413 5628 -2379
rect 5662 -2413 5685 -2379
rect 5605 -2459 5685 -2413
rect 5605 -2493 5628 -2459
rect 5662 -2493 5685 -2459
rect 5605 -2539 5685 -2493
rect 5605 -2573 5628 -2539
rect 5662 -2573 5685 -2539
rect 5605 -2596 5685 -2573
rect 6235 -2379 6315 -2346
rect 6235 -2413 6258 -2379
rect 6292 -2413 6315 -2379
rect 6235 -2459 6315 -2413
rect 6235 -2493 6258 -2459
rect 6292 -2493 6315 -2459
rect 6235 -2539 6315 -2493
rect 6235 -2573 6258 -2539
rect 6292 -2573 6315 -2539
rect 6235 -2596 6315 -2573
rect -83 -2650 -3 -2636
rect -83 -2702 -69 -2650
rect -17 -2702 -3 -2650
rect -83 -2716 -3 -2702
rect 755 -2747 795 -2597
rect 1055 -2747 1095 -2597
rect 1355 -2747 1395 -2597
rect 2966 -2746 3006 -2596
rect 3266 -2746 3306 -2596
rect 3566 -2746 3606 -2596
rect 3990 -2650 4070 -2636
rect 3990 -2702 4004 -2650
rect 4056 -2702 4070 -2650
rect 3990 -2716 4070 -2702
rect 4187 -2650 4267 -2636
rect 4187 -2702 4201 -2650
rect 4253 -2702 4267 -2650
rect 4187 -2716 4267 -2702
rect 5025 -2746 5065 -2596
rect 5325 -2746 5365 -2596
rect 5625 -2746 5665 -2596
rect 2235 -2747 6345 -2746
rect -213 -2814 -190 -2780
rect -156 -2814 -133 -2780
rect -213 -2837 -133 -2814
rect -85 -2779 6345 -2747
rect -85 -2780 2629 -2779
rect -85 -2814 -62 -2780
rect -28 -2814 18 -2780
rect 52 -2814 98 -2780
rect 132 -2814 178 -2780
rect 212 -2814 258 -2780
rect 292 -2814 338 -2780
rect 372 -2814 418 -2780
rect 452 -2814 498 -2780
rect 532 -2814 578 -2780
rect 612 -2814 658 -2780
rect 692 -2814 738 -2780
rect 772 -2814 818 -2780
rect 852 -2814 898 -2780
rect 932 -2814 978 -2780
rect 1012 -2814 1058 -2780
rect 1092 -2814 1138 -2780
rect 1172 -2814 1218 -2780
rect 1252 -2814 1298 -2780
rect 1332 -2814 1378 -2780
rect 1412 -2814 1458 -2780
rect 1492 -2814 1538 -2780
rect 1572 -2814 1618 -2780
rect 1652 -2814 1698 -2780
rect 1732 -2814 1778 -2780
rect 1812 -2814 1858 -2780
rect 1892 -2814 1938 -2780
rect 1972 -2814 2018 -2780
rect 2052 -2814 2098 -2780
rect 2132 -2814 2178 -2780
rect 2212 -2813 2629 -2780
rect 2663 -2813 2709 -2779
rect 2743 -2813 2789 -2779
rect 2823 -2813 2869 -2779
rect 2903 -2813 2949 -2779
rect 2983 -2813 3029 -2779
rect 3063 -2813 3109 -2779
rect 3143 -2813 3189 -2779
rect 3223 -2813 3269 -2779
rect 3303 -2813 3349 -2779
rect 3383 -2813 3429 -2779
rect 3463 -2813 3509 -2779
rect 3543 -2813 3589 -2779
rect 3623 -2813 3669 -2779
rect 3703 -2813 3749 -2779
rect 3783 -2813 3829 -2779
rect 3863 -2813 3909 -2779
rect 3943 -2813 4368 -2779
rect 4402 -2813 4448 -2779
rect 4482 -2813 4528 -2779
rect 4562 -2813 4608 -2779
rect 4642 -2813 4688 -2779
rect 4722 -2813 4768 -2779
rect 4802 -2813 4848 -2779
rect 4882 -2813 4928 -2779
rect 4962 -2813 5008 -2779
rect 5042 -2813 5088 -2779
rect 5122 -2813 5168 -2779
rect 5202 -2813 5248 -2779
rect 5282 -2813 5328 -2779
rect 5362 -2813 5408 -2779
rect 5442 -2813 5488 -2779
rect 5522 -2813 5568 -2779
rect 5602 -2813 5648 -2779
rect 5682 -2813 5728 -2779
rect 5762 -2813 5808 -2779
rect 5842 -2813 5888 -2779
rect 5922 -2813 5968 -2779
rect 6002 -2813 6048 -2779
rect 6082 -2813 6128 -2779
rect 6162 -2813 6208 -2779
rect 6242 -2813 6288 -2779
rect 6322 -2813 6345 -2779
rect 2212 -2814 6345 -2813
rect -85 -2846 6345 -2814
rect -85 -2847 2235 -2846
<< via1 >>
rect 9 1221 61 1230
rect 9 1187 18 1221
rect 18 1187 52 1221
rect 52 1187 61 1221
rect 9 1178 61 1187
rect 4579 1221 4631 1230
rect 4579 1187 4588 1221
rect 4588 1187 4622 1221
rect 4622 1187 4631 1221
rect 4579 1178 4631 1187
rect -883 316 -831 368
rect -769 1051 -717 1103
rect -655 -322 -603 -270
rect -541 -1053 -489 -1001
rect 469 1091 521 1100
rect 469 1057 478 1091
rect 478 1057 512 1091
rect 512 1057 521 1091
rect 469 1048 521 1057
rect 599 991 651 1000
rect 599 957 608 991
rect 608 957 642 991
rect 642 957 651 991
rect 599 948 651 957
rect 469 891 521 900
rect 469 857 478 891
rect 478 857 512 891
rect 512 857 521 891
rect 469 848 521 857
rect 599 791 651 800
rect 599 757 608 791
rect 608 757 642 791
rect 642 757 651 791
rect 599 748 651 757
rect 1729 1091 1781 1100
rect 1729 1057 1738 1091
rect 1738 1057 1772 1091
rect 1772 1057 1781 1091
rect 1729 1048 1781 1057
rect 1629 791 1681 800
rect 1629 757 1638 791
rect 1638 757 1672 791
rect 1672 757 1681 791
rect 1629 748 1681 757
rect 1929 991 1981 1000
rect 1929 957 1938 991
rect 1938 957 1972 991
rect 1972 957 1981 991
rect 1929 948 1981 957
rect 2521 1025 2573 1034
rect 2521 991 2530 1025
rect 2530 991 2564 1025
rect 2564 991 2573 1025
rect 2521 982 2573 991
rect 2079 891 2131 900
rect 2079 857 2088 891
rect 2088 857 2122 891
rect 2122 857 2131 891
rect 2079 848 2131 857
rect 2521 874 2573 926
rect 2809 1051 2861 1103
rect 2809 841 2861 850
rect 2809 807 2818 841
rect 2818 807 2852 841
rect 2852 807 2861 841
rect 2809 798 2861 807
rect 3709 841 3761 850
rect 3709 807 3718 841
rect 3718 807 3752 841
rect 3752 807 3761 841
rect 3709 798 3761 807
rect 2243 359 2295 368
rect 2243 325 2252 359
rect 2252 325 2286 359
rect 2286 325 2295 359
rect 2243 316 2295 325
rect 1829 281 1881 290
rect 1829 247 1838 281
rect 1838 247 1872 281
rect 1872 247 1881 281
rect 1829 238 1881 247
rect 3997 1025 4049 1034
rect 3997 991 4006 1025
rect 4006 991 4040 1025
rect 4040 991 4049 1025
rect 3997 982 4049 991
rect 3997 910 4049 919
rect 3997 876 4006 910
rect 4006 876 4040 910
rect 4040 876 4049 910
rect 3997 867 4049 876
rect 4689 991 4741 1000
rect 4689 957 4698 991
rect 4698 957 4732 991
rect 4732 957 4741 991
rect 4689 948 4741 957
rect 4689 871 4741 880
rect 4689 837 4698 871
rect 4698 837 4732 871
rect 4732 837 4741 871
rect 4689 828 4741 837
rect 5819 991 5871 1000
rect 5819 957 5828 991
rect 5828 957 5862 991
rect 5862 957 5871 991
rect 5819 948 5871 957
rect 5669 871 5721 880
rect 5669 837 5678 871
rect 5678 837 5712 871
rect 5712 837 5721 871
rect 5669 828 5721 837
rect 6022 600 6074 609
rect 6022 566 6031 600
rect 6031 566 6065 600
rect 6065 566 6074 600
rect 6022 557 6074 566
rect 5919 281 5971 290
rect 5919 247 5928 281
rect 5928 247 5962 281
rect 5962 247 5971 281
rect 5919 238 5971 247
rect 381 161 433 170
rect 381 127 390 161
rect 390 127 424 161
rect 424 127 433 161
rect 381 118 433 127
rect 4347 161 4399 170
rect 4347 127 4356 161
rect 4356 127 4390 161
rect 4390 127 4399 161
rect 4347 118 4399 127
rect 381 -79 433 -70
rect 381 -113 390 -79
rect 390 -113 424 -79
rect 424 -113 433 -79
rect 381 -122 433 -113
rect 4347 -79 4399 -70
rect 4347 -113 4356 -79
rect 4356 -113 4390 -79
rect 4390 -113 4399 -79
rect 4347 -122 4399 -113
rect 1829 -199 1881 -190
rect 1829 -233 1838 -199
rect 1838 -233 1872 -199
rect 1872 -233 1881 -199
rect 1829 -242 1881 -233
rect 2243 -279 2295 -270
rect 2243 -313 2252 -279
rect 2252 -313 2286 -279
rect 2286 -313 2295 -279
rect 2243 -322 2295 -313
rect 2520 -393 2572 -341
rect 599 -709 651 -700
rect 599 -743 608 -709
rect 608 -743 642 -709
rect 642 -743 651 -709
rect 599 -752 651 -743
rect 469 -809 521 -800
rect 469 -843 478 -809
rect 478 -843 512 -809
rect 512 -843 521 -809
rect 469 -852 521 -843
rect 599 -909 651 -900
rect 599 -943 608 -909
rect 608 -943 642 -909
rect 642 -943 651 -909
rect 599 -952 651 -943
rect 469 -1009 521 -1000
rect 469 -1043 478 -1009
rect 478 -1043 512 -1009
rect 512 -1043 521 -1009
rect 469 -1052 521 -1043
rect 1629 -709 1681 -700
rect 1629 -743 1638 -709
rect 1638 -743 1672 -709
rect 1672 -743 1681 -709
rect 1629 -752 1681 -743
rect 1729 -1009 1781 -1000
rect 1729 -1043 1738 -1009
rect 1738 -1043 1772 -1009
rect 1772 -1043 1781 -1009
rect 1729 -1052 1781 -1043
rect 2079 -809 2131 -800
rect 2079 -843 2088 -809
rect 2088 -843 2122 -809
rect 2122 -843 2131 -809
rect 2079 -852 2131 -843
rect 1929 -909 1981 -900
rect 1929 -943 1938 -909
rect 1938 -943 1972 -909
rect 1972 -943 1981 -909
rect 1929 -952 1981 -943
rect 2521 -909 2573 -900
rect 2521 -943 2530 -909
rect 2530 -943 2564 -909
rect 2564 -943 2573 -909
rect 2521 -952 2573 -943
rect 2809 -759 2861 -750
rect 2809 -793 2818 -759
rect 2818 -793 2852 -759
rect 2852 -793 2861 -759
rect 2809 -802 2861 -793
rect 2809 -1053 2861 -1001
rect 3709 -759 3761 -750
rect 3709 -793 3718 -759
rect 3718 -793 3752 -759
rect 3752 -793 3761 -759
rect 3709 -802 3761 -793
rect 3709 -909 3761 -900
rect 3709 -943 3718 -909
rect 3718 -943 3752 -909
rect 3752 -943 3761 -909
rect 3709 -952 3761 -943
rect 3997 -392 4049 -340
rect 5919 -199 5971 -190
rect 5919 -233 5928 -199
rect 5928 -233 5962 -199
rect 5962 -233 5971 -199
rect 5919 -242 5971 -233
rect 4689 -789 4741 -780
rect 4689 -823 4698 -789
rect 4698 -823 4732 -789
rect 4732 -823 4741 -789
rect 4689 -832 4741 -823
rect 4689 -909 4741 -900
rect 4689 -943 4698 -909
rect 4698 -943 4732 -909
rect 4732 -943 4741 -909
rect 4689 -952 4741 -943
rect 5669 -789 5721 -780
rect 5669 -823 5678 -789
rect 5678 -823 5712 -789
rect 5712 -823 5721 -789
rect 5669 -832 5721 -823
rect 5819 -909 5871 -900
rect 5819 -943 5828 -909
rect 5828 -943 5862 -909
rect 5862 -943 5871 -909
rect 5819 -952 5871 -943
rect 6022 -519 6074 -510
rect 6022 -553 6031 -519
rect 6031 -553 6065 -519
rect 6065 -553 6074 -519
rect 6022 -562 6074 -553
rect 19 -1410 71 -1401
rect 19 -1444 28 -1410
rect 28 -1444 62 -1410
rect 62 -1444 71 -1410
rect 19 -1453 71 -1444
rect 19 -1530 71 -1521
rect 19 -1564 28 -1530
rect 28 -1564 62 -1530
rect 62 -1564 71 -1530
rect 19 -1573 71 -1564
rect 19 -1650 71 -1641
rect 19 -1684 28 -1650
rect 28 -1684 62 -1650
rect 62 -1684 71 -1650
rect 19 -1693 71 -1684
rect 19 -1770 71 -1761
rect 19 -1804 28 -1770
rect 28 -1804 62 -1770
rect 62 -1804 71 -1770
rect 19 -1813 71 -1804
rect 2029 -1453 2081 -1401
rect 1879 -1573 1931 -1521
rect 1729 -1693 1781 -1641
rect 1579 -1813 1631 -1761
rect 4347 -1373 4399 -1364
rect 4347 -1407 4356 -1373
rect 4356 -1407 4390 -1373
rect 4390 -1407 4399 -1373
rect 4347 -1416 4399 -1407
rect 6383 -1405 6435 -1396
rect 6383 -1439 6392 -1405
rect 6392 -1439 6426 -1405
rect 6426 -1439 6435 -1405
rect 6383 -1448 6435 -1439
rect 4435 -1599 4487 -1590
rect 4435 -1633 4448 -1599
rect 4448 -1633 4482 -1599
rect 4482 -1633 4487 -1599
rect 4435 -1642 4487 -1633
rect 2810 -1979 2862 -1970
rect 2810 -2013 2819 -1979
rect 2819 -2013 2853 -1979
rect 2853 -2013 2862 -1979
rect 2810 -2022 2862 -2013
rect 3710 -1979 3762 -1970
rect 3710 -2013 3719 -1979
rect 3719 -2013 3753 -1979
rect 3753 -2013 3762 -1979
rect 3710 -2022 3762 -2013
rect 4004 -1806 4056 -1797
rect 4004 -1840 4013 -1806
rect 4013 -1840 4047 -1806
rect 4047 -1840 4056 -1806
rect 4004 -1849 4056 -1840
rect 4289 -1919 4341 -1867
rect 4289 -1991 4341 -1982
rect 4289 -2025 4298 -1991
rect 4298 -2025 4332 -1991
rect 4332 -2025 4341 -1991
rect 4289 -2034 4341 -2025
rect 4289 -2119 4341 -2110
rect 4289 -2153 4298 -2119
rect 4298 -2153 4332 -2119
rect 4332 -2153 4341 -2119
rect 4289 -2162 4341 -2153
rect 4289 -2239 4341 -2230
rect 4289 -2273 4298 -2239
rect 4298 -2273 4332 -2239
rect 4332 -2273 4341 -2239
rect 4289 -2282 4341 -2273
rect 4489 -1729 4541 -1720
rect 4489 -1763 4498 -1729
rect 4498 -1763 4532 -1729
rect 4532 -1763 4541 -1729
rect 4489 -1772 4541 -1763
rect 4601 -1849 4653 -1840
rect 4601 -1883 4610 -1849
rect 4610 -1883 4644 -1849
rect 4644 -1883 4653 -1849
rect 4601 -1892 4653 -1883
rect 4789 -1939 4841 -1930
rect 4789 -1973 4798 -1939
rect 4798 -1973 4832 -1939
rect 4832 -1973 4841 -1939
rect 4789 -1982 4841 -1973
rect 5769 -1729 5821 -1720
rect 5769 -1763 5778 -1729
rect 5778 -1763 5812 -1729
rect 5812 -1763 5821 -1729
rect 5769 -1772 5821 -1763
rect 6161 -1729 6213 -1720
rect 6161 -1763 6170 -1729
rect 6170 -1763 6204 -1729
rect 6204 -1763 6213 -1729
rect 6161 -1772 6213 -1763
rect 5889 -1839 5941 -1830
rect 5889 -1873 5898 -1839
rect 5898 -1873 5932 -1839
rect 5932 -1873 5941 -1839
rect 5889 -1882 5941 -1873
rect 6021 -1840 6073 -1831
rect 6021 -1874 6030 -1840
rect 6030 -1874 6064 -1840
rect 6064 -1874 6073 -1840
rect 6021 -1883 6073 -1874
rect 5769 -1939 5821 -1930
rect 5769 -1973 5778 -1939
rect 5778 -1973 5812 -1939
rect 5812 -1973 5821 -1939
rect 5769 -1982 5821 -1973
rect 5899 -2069 5951 -2017
rect 6383 -2026 6435 -2017
rect 6383 -2060 6392 -2026
rect 6392 -2060 6426 -2026
rect 6426 -2060 6435 -2026
rect 6383 -2069 6435 -2060
rect -69 -2659 -17 -2650
rect -69 -2693 -60 -2659
rect -60 -2693 -26 -2659
rect -26 -2693 -17 -2659
rect -69 -2702 -17 -2693
rect 4004 -2659 4056 -2650
rect 4004 -2693 4013 -2659
rect 4013 -2693 4047 -2659
rect 4047 -2693 4056 -2659
rect 4004 -2702 4056 -2693
rect 4201 -2659 4253 -2650
rect 4201 -2693 4210 -2659
rect 4210 -2693 4244 -2659
rect 4244 -2693 4253 -2659
rect 4201 -2702 4253 -2693
<< metal2 >>
rect 16 1244 56 1350
rect -5 1230 75 1244
rect -5 1178 9 1230
rect 61 1178 75 1230
rect -5 1164 75 1178
rect -783 1105 -703 1116
rect -783 1049 -771 1105
rect -715 1049 -703 1105
rect -783 1036 -703 1049
rect -897 370 -817 381
rect -897 314 -885 370
rect -829 314 -817 370
rect -897 301 -817 314
rect 387 184 427 1350
rect 455 1100 535 1114
rect 455 1048 469 1100
rect 521 1094 535 1100
rect 1715 1100 1795 1114
rect 1715 1094 1729 1100
rect 521 1054 1729 1094
rect 521 1048 535 1054
rect 455 1034 535 1048
rect 1715 1048 1729 1054
rect 1781 1048 1795 1100
rect 2795 1105 2875 1116
rect 2795 1049 2807 1105
rect 2863 1049 2875 1105
rect 1715 1034 1795 1048
rect 2507 1034 2587 1048
rect 2795 1036 2875 1049
rect 585 1000 665 1014
rect 585 948 599 1000
rect 651 994 665 1000
rect 1915 1000 1995 1014
rect 1915 994 1929 1000
rect 651 954 1929 994
rect 651 948 665 954
rect 585 934 665 948
rect 1915 948 1929 954
rect 1981 948 1995 1000
rect 2507 982 2521 1034
rect 2573 1008 2587 1034
rect 3983 1034 4063 1048
rect 3983 1008 3997 1034
rect 2573 982 3997 1008
rect 4049 982 4063 1034
rect 2507 968 4063 982
rect 1915 934 1995 948
rect 2507 933 2587 940
rect 2507 926 4063 933
rect 455 900 535 914
rect 455 848 469 900
rect 521 894 535 900
rect 2065 900 2145 914
rect 2065 894 2079 900
rect 521 854 2079 894
rect 521 848 535 854
rect 455 834 535 848
rect 2065 848 2079 854
rect 2131 848 2145 900
rect 2507 874 2521 926
rect 2573 919 4063 926
rect 2573 893 3997 919
rect 2573 874 2587 893
rect 2507 860 2587 874
rect 3983 867 3997 893
rect 4049 867 4063 919
rect 2065 834 2145 848
rect 2795 850 2875 864
rect 585 800 665 814
rect 585 748 599 800
rect 651 794 665 800
rect 1615 800 1695 814
rect 1615 794 1629 800
rect 651 754 1629 794
rect 651 748 665 754
rect 585 734 665 748
rect 1615 748 1629 754
rect 1681 748 1695 800
rect 2795 798 2809 850
rect 2861 844 2875 850
rect 3695 850 3775 864
rect 3983 853 4063 867
rect 3695 844 3709 850
rect 2861 804 3709 844
rect 2861 798 2875 804
rect 2795 784 2875 798
rect 3695 798 3709 804
rect 3761 798 3775 850
rect 3695 784 3775 798
rect 1615 734 1695 748
rect 2229 370 2309 381
rect 2229 314 2241 370
rect 2297 314 2309 370
rect 1815 290 1895 304
rect 2229 301 2309 314
rect 1815 238 1829 290
rect 1881 238 1895 290
rect 1815 224 1895 238
rect 367 170 447 184
rect 367 118 381 170
rect 433 118 447 170
rect 367 104 447 118
rect 387 -56 427 104
rect 367 -70 447 -56
rect 367 -122 381 -70
rect 433 -122 447 -70
rect 367 -136 447 -122
rect -669 -268 -589 -257
rect -669 -324 -657 -268
rect -601 -324 -589 -268
rect -669 -337 -589 -324
rect -555 -999 -475 -988
rect -555 -1055 -543 -999
rect -487 -1055 -475 -999
rect -555 -1068 -475 -1055
rect 387 -1276 427 -136
rect 1835 -176 1875 224
rect 1815 -190 1895 -176
rect 1815 -242 1829 -190
rect 1881 -242 1895 -190
rect 1815 -256 1895 -242
rect 2229 -268 2309 -257
rect 2229 -324 2241 -268
rect 2297 -324 2309 -268
rect 2229 -337 2309 -324
rect 2506 -341 2586 -327
rect 2506 -393 2520 -341
rect 2572 -346 2586 -341
rect 3983 -340 4063 -326
rect 3983 -346 3997 -340
rect 2572 -386 3997 -346
rect 2572 -393 2586 -386
rect 2506 -407 2586 -393
rect 3983 -392 3997 -386
rect 4049 -392 4063 -340
rect 3983 -406 4063 -392
rect 585 -700 665 -686
rect 585 -752 599 -700
rect 651 -706 665 -700
rect 1615 -700 1695 -686
rect 1615 -706 1629 -700
rect 651 -746 1629 -706
rect 651 -752 665 -746
rect 585 -766 665 -752
rect 1615 -752 1629 -746
rect 1681 -752 1695 -700
rect 1615 -766 1695 -752
rect 2795 -750 2875 -736
rect 455 -800 535 -786
rect 455 -852 469 -800
rect 521 -806 535 -800
rect 2065 -800 2145 -786
rect 2065 -806 2079 -800
rect 521 -846 2079 -806
rect 521 -852 535 -846
rect 455 -866 535 -852
rect 2065 -852 2079 -846
rect 2131 -852 2145 -800
rect 2795 -802 2809 -750
rect 2861 -756 2875 -750
rect 3695 -750 3775 -736
rect 3695 -756 3709 -750
rect 2861 -796 3709 -756
rect 2861 -802 2875 -796
rect 2795 -816 2875 -802
rect 3695 -802 3709 -796
rect 3761 -802 3775 -750
rect 3695 -816 3775 -802
rect 2065 -866 2145 -852
rect 585 -900 665 -886
rect 585 -952 599 -900
rect 651 -906 665 -900
rect 1915 -900 1995 -886
rect 1915 -906 1929 -900
rect 651 -946 1929 -906
rect 651 -952 665 -946
rect 585 -966 665 -952
rect 1915 -952 1929 -946
rect 1981 -952 1995 -900
rect 1915 -966 1995 -952
rect 2507 -900 2587 -886
rect 2507 -952 2521 -900
rect 2573 -906 2587 -900
rect 3695 -900 3775 -886
rect 3695 -906 3709 -900
rect 2573 -946 3709 -906
rect 2573 -952 2587 -946
rect 2507 -966 2587 -952
rect 3695 -952 3709 -946
rect 3761 -952 3775 -900
rect 3695 -966 3775 -952
rect 455 -1000 535 -986
rect 455 -1052 469 -1000
rect 521 -1006 535 -1000
rect 1715 -1000 1795 -986
rect 1715 -1006 1729 -1000
rect 521 -1046 1729 -1006
rect 521 -1052 535 -1046
rect 455 -1066 535 -1052
rect 1715 -1052 1729 -1046
rect 1781 -1052 1795 -1000
rect 1715 -1066 1795 -1052
rect 2795 -999 2875 -988
rect 2795 -1055 2807 -999
rect 2863 -1055 2875 -999
rect 2795 -1068 2875 -1055
rect -63 -1316 427 -1276
rect -63 -2636 -23 -1316
rect 5 -1401 85 -1387
rect 5 -1453 19 -1401
rect 71 -1407 85 -1401
rect 2015 -1401 2095 -1387
rect 2015 -1407 2029 -1401
rect 71 -1447 2029 -1407
rect 71 -1453 85 -1447
rect 5 -1467 85 -1453
rect 2015 -1453 2029 -1447
rect 2081 -1453 2095 -1401
rect 2015 -1467 2095 -1453
rect 5 -1521 85 -1507
rect 5 -1573 19 -1521
rect 71 -1527 85 -1521
rect 1865 -1521 1945 -1507
rect 1865 -1527 1879 -1521
rect 71 -1567 1879 -1527
rect 71 -1573 85 -1567
rect 5 -1587 85 -1573
rect 1865 -1573 1879 -1567
rect 1931 -1573 1945 -1521
rect 1865 -1587 1945 -1573
rect 5 -1641 85 -1627
rect 5 -1693 19 -1641
rect 71 -1647 85 -1641
rect 1715 -1641 1795 -1627
rect 1715 -1647 1729 -1641
rect 71 -1687 1729 -1647
rect 71 -1693 85 -1687
rect 5 -1707 85 -1693
rect 1715 -1693 1729 -1687
rect 1781 -1693 1795 -1641
rect 1715 -1707 1795 -1693
rect 5 -1761 85 -1747
rect 5 -1813 19 -1761
rect 71 -1767 85 -1761
rect 1565 -1761 1645 -1747
rect 1565 -1767 1579 -1761
rect 71 -1807 1579 -1767
rect 71 -1813 85 -1807
rect 5 -1827 85 -1813
rect 1565 -1813 1579 -1807
rect 1631 -1813 1645 -1761
rect 1565 -1827 1645 -1813
rect 3990 -1797 4070 -1783
rect 3990 -1849 4004 -1797
rect 4056 -1849 4070 -1797
rect 3990 -1863 4070 -1849
rect 2796 -1970 2876 -1956
rect 2796 -2022 2810 -1970
rect 2862 -1976 2876 -1970
rect 3696 -1970 3776 -1956
rect 3696 -1976 3710 -1970
rect 2862 -2016 3710 -1976
rect 2862 -2022 2876 -2016
rect 2796 -2036 2876 -2022
rect 3696 -2022 3710 -2016
rect 3762 -2022 3776 -1970
rect 3696 -2036 3776 -2022
rect 4010 -2636 4050 -1863
rect 4207 -2636 4247 1347
rect 4353 184 4393 1347
rect 4333 170 4413 184
rect 4333 118 4347 170
rect 4399 118 4413 170
rect 4333 104 4413 118
rect 4353 -56 4393 104
rect 4333 -70 4413 -56
rect 4333 -122 4347 -70
rect 4399 -122 4413 -70
rect 4333 -136 4413 -122
rect 4353 -1350 4393 -136
rect 4333 -1364 4413 -1350
rect 4333 -1416 4347 -1364
rect 4399 -1416 4413 -1364
rect 4333 -1430 4413 -1416
rect 4441 -1576 4481 1347
rect 4585 1244 4625 1346
rect 4565 1230 4645 1244
rect 4565 1178 4579 1230
rect 4631 1178 4645 1230
rect 4565 1164 4645 1178
rect 4675 1000 4755 1014
rect 4675 948 4689 1000
rect 4741 994 4755 1000
rect 5805 1000 5885 1014
rect 5805 994 5819 1000
rect 4741 954 5819 994
rect 4741 948 4755 954
rect 4675 934 4755 948
rect 5805 948 5819 954
rect 5871 948 5885 1000
rect 5805 934 5885 948
rect 4675 880 4755 894
rect 4675 828 4689 880
rect 4741 874 4755 880
rect 5655 880 5735 894
rect 5655 874 5669 880
rect 4741 834 5669 874
rect 4741 828 4755 834
rect 4675 814 4755 828
rect 5655 828 5669 834
rect 5721 828 5735 880
rect 5655 814 5735 828
rect 6008 609 6088 623
rect 6008 557 6022 609
rect 6074 604 6088 609
rect 6074 564 6206 604
rect 6074 557 6088 564
rect 6008 543 6088 557
rect 5905 290 5985 304
rect 5905 238 5919 290
rect 5971 238 5985 290
rect 5905 -190 5985 238
rect 5905 -242 5919 -190
rect 5971 -242 5985 -190
rect 5905 -256 5985 -242
rect 6008 -510 6088 -496
rect 6008 -562 6022 -510
rect 6074 -562 6088 -510
rect 6008 -576 6088 -562
rect 4675 -780 4755 -766
rect 4675 -832 4689 -780
rect 4741 -786 4755 -780
rect 5655 -780 5735 -766
rect 5655 -786 5669 -780
rect 4741 -826 5669 -786
rect 4741 -832 4755 -826
rect 4675 -846 4755 -832
rect 5655 -832 5669 -826
rect 5721 -832 5735 -780
rect 5655 -846 5735 -832
rect 4675 -900 4755 -886
rect 4675 -952 4689 -900
rect 4741 -906 4755 -900
rect 5805 -900 5885 -886
rect 5805 -906 5819 -900
rect 4741 -946 5819 -906
rect 4741 -952 4755 -946
rect 4675 -966 4755 -952
rect 5805 -952 5819 -946
rect 5871 -952 5885 -900
rect 5805 -966 5885 -952
rect 4421 -1590 4501 -1576
rect 4421 -1642 4435 -1590
rect 4487 -1642 4501 -1590
rect 4421 -1656 4501 -1642
rect 4475 -1720 4555 -1706
rect 4475 -1772 4489 -1720
rect 4541 -1726 4555 -1720
rect 5755 -1720 5835 -1706
rect 5755 -1726 5769 -1720
rect 4541 -1766 5769 -1726
rect 4541 -1772 4555 -1766
rect 4475 -1786 4555 -1772
rect 5755 -1772 5769 -1766
rect 5821 -1772 5835 -1720
rect 5755 -1786 5835 -1772
rect 4587 -1836 4667 -1826
rect 5875 -1830 5955 -1816
rect 6028 -1817 6068 -576
rect 6166 -1706 6206 564
rect 6369 -1396 6449 -1382
rect 6369 -1448 6383 -1396
rect 6435 -1448 6449 -1396
rect 6369 -1462 6449 -1448
rect 6147 -1720 6227 -1706
rect 6147 -1772 6161 -1720
rect 6213 -1772 6227 -1720
rect 6147 -1786 6227 -1772
rect 5875 -1836 5889 -1830
rect 4587 -1840 5889 -1836
rect 4275 -1867 4355 -1853
rect 4275 -1919 4289 -1867
rect 4341 -1893 4355 -1867
rect 4587 -1892 4601 -1840
rect 4653 -1876 5889 -1840
rect 4653 -1892 4667 -1876
rect 4341 -1919 4423 -1893
rect 4587 -1906 4667 -1892
rect 5875 -1882 5889 -1876
rect 5941 -1882 5955 -1830
rect 5875 -1896 5955 -1882
rect 6007 -1831 6087 -1817
rect 6007 -1883 6021 -1831
rect 6073 -1883 6087 -1831
rect 6007 -1897 6087 -1883
rect 4275 -1933 4423 -1919
rect 4383 -1936 4423 -1933
rect 4775 -1930 4855 -1916
rect 4775 -1936 4789 -1930
rect 4275 -1982 4355 -1968
rect 4383 -1976 4789 -1936
rect 4275 -2034 4289 -1982
rect 4341 -2008 4355 -1982
rect 4775 -1982 4789 -1976
rect 4841 -1936 4855 -1930
rect 5755 -1930 5835 -1916
rect 5755 -1936 5769 -1930
rect 4841 -1976 5769 -1936
rect 4841 -1982 4855 -1976
rect 4775 -1996 4855 -1982
rect 5755 -1982 5769 -1976
rect 5821 -1982 5835 -1930
rect 5755 -1996 5835 -1982
rect 6389 -2003 6429 -1462
rect 4341 -2024 4423 -2008
rect 5885 -2017 5965 -2003
rect 5885 -2024 5899 -2017
rect 4341 -2034 5899 -2024
rect 4275 -2048 5899 -2034
rect 4383 -2064 5899 -2048
rect 5885 -2069 5899 -2064
rect 5951 -2069 5965 -2017
rect 5885 -2083 5965 -2069
rect 6369 -2017 6449 -2003
rect 6369 -2069 6383 -2017
rect 6435 -2026 6449 -2017
rect 6435 -2066 6498 -2026
rect 6435 -2069 6449 -2066
rect 6369 -2083 6449 -2069
rect 4275 -2110 4355 -2096
rect 4275 -2162 4289 -2110
rect 4341 -2111 4355 -2110
rect 4341 -2151 6426 -2111
rect 4341 -2162 4355 -2151
rect 4275 -2176 4355 -2162
rect 4275 -2230 4355 -2216
rect 4275 -2282 4289 -2230
rect 4341 -2236 4355 -2230
rect 4341 -2276 6426 -2236
rect 4341 -2282 4355 -2276
rect 4275 -2296 4355 -2282
rect -83 -2650 -3 -2636
rect -83 -2702 -69 -2650
rect -17 -2702 -3 -2650
rect -83 -2716 -3 -2702
rect 3990 -2650 4070 -2636
rect 3990 -2702 4004 -2650
rect 4056 -2702 4070 -2650
rect 3990 -2716 4070 -2702
rect 4187 -2650 4267 -2636
rect 4187 -2702 4201 -2650
rect 4253 -2702 4267 -2650
rect 4187 -2716 4267 -2702
<< via2 >>
rect -771 1103 -715 1105
rect -771 1051 -769 1103
rect -769 1051 -717 1103
rect -717 1051 -715 1103
rect -771 1049 -715 1051
rect -885 368 -829 370
rect -885 316 -883 368
rect -883 316 -831 368
rect -831 316 -829 368
rect -885 314 -829 316
rect 2807 1103 2863 1105
rect 2807 1051 2809 1103
rect 2809 1051 2861 1103
rect 2861 1051 2863 1103
rect 2807 1049 2863 1051
rect 2241 368 2297 370
rect 2241 316 2243 368
rect 2243 316 2295 368
rect 2295 316 2297 368
rect 2241 314 2297 316
rect -657 -270 -601 -268
rect -657 -322 -655 -270
rect -655 -322 -603 -270
rect -603 -322 -601 -270
rect -657 -324 -601 -322
rect -543 -1001 -487 -999
rect -543 -1053 -541 -1001
rect -541 -1053 -489 -1001
rect -489 -1053 -487 -1001
rect -543 -1055 -487 -1053
rect 2241 -270 2297 -268
rect 2241 -322 2243 -270
rect 2243 -322 2295 -270
rect 2295 -322 2297 -270
rect 2241 -324 2297 -322
rect 2807 -1001 2863 -999
rect 2807 -1053 2809 -1001
rect 2809 -1053 2861 -1001
rect 2861 -1053 2863 -1001
rect 2807 -1055 2863 -1053
<< metal3 >>
rect -793 1106 -693 1126
rect 2785 1106 2885 1126
rect -793 1105 2885 1106
rect -793 1049 -771 1105
rect -715 1049 2807 1105
rect 2863 1049 2885 1105
rect -793 1046 2885 1049
rect -793 1026 -693 1046
rect 2785 1026 2885 1046
rect -907 372 -807 391
rect 2219 372 2319 391
rect -907 370 2319 372
rect -907 314 -885 370
rect -829 314 2241 370
rect 2297 314 2319 370
rect -907 312 2319 314
rect -907 291 -807 312
rect 2219 291 2319 312
rect -679 -266 -579 -247
rect 2219 -266 2319 -247
rect -679 -268 2319 -266
rect -679 -324 -657 -268
rect -601 -324 2241 -268
rect 2297 -324 2319 -268
rect -679 -326 2319 -324
rect -679 -347 -579 -326
rect 2219 -347 2319 -326
rect -565 -996 -465 -978
rect 2785 -996 2885 -978
rect -565 -999 2885 -996
rect -565 -1055 -543 -999
rect -487 -1055 2807 -999
rect 2863 -1055 2885 -999
rect -565 -1056 2885 -1055
rect -565 -1078 -465 -1056
rect 2785 -1078 2885 -1056
<< labels >>
flabel metal2 s 6395 -2267 6415 -2247 2 FreeSans 2000 0 0 0 s2
port 17 nsew
flabel metal2 s 6395 -2141 6415 -2121 2 FreeSans 2000 0 0 0 s2_bar
port 16 nsew
flabel metal2 s 4595 1320 4615 1340 2 FreeSans 2000 0 0 0 CLK2
port 15 nsew
flabel metal2 s 4451 1320 4471 1340 2 FreeSans 2000 0 0 0 CLK3
port 14 nsew
flabel metal2 s 4363 1320 4383 1340 2 FreeSans 2000 0 0 0 Dis2
port 13 nsew
flabel metal2 s 4217 1320 4237 1340 2 FreeSans 2000 0 0 0 Dis3
port 12 nsew
flabel metal2 s 397 1322 417 1342 2 FreeSans 2000 0 0 0 Dis1
port 11 nsew
flabel metal2 s 26 1325 46 1345 2 FreeSans 2000 0 0 0 CLK1
port 10 nsew
flabel metal1 s -317 960 -256 1020 2 FreeSans 3126 0 0 0 x3_bar
port 9 nsew
flabel metal1 s -431 1021 -370 1081 2 FreeSans 3126 0 0 0 x3
port 8 nsew
flabel metal1 s -546 960 -485 1020 2 FreeSans 3126 0 0 0 x2_bar
port 7 nsew
flabel metal1 s -659 1021 -598 1081 2 FreeSans 3126 0 0 0 x2
port 6 nsew
flabel metal1 s -773 959 -712 1019 2 FreeSans 3126 0 0 0 x1_bar
port 5 nsew
flabel metal1 s -887 1020 -826 1080 2 FreeSans 3126 0 0 0 x1
port 4 nsew
flabel metal1 s -1002 959 -941 1019 2 FreeSans 3126 0 0 0 x0_bar
port 3 nsew
flabel metal1 s -1115 1020 -1054 1080 2 FreeSans 3126 0 0 0 x0
port 2 nsew
flabel metal1 s -190 7 -156 41 2 FreeSans 2000 0 0 0 GND
port 1 nsew
rlabel locali 1005 -551 1045 -511 2 EESPFAL_XOR_v3_1/OUT
rlabel locali -55 -1036 -35 -1016 2 EESPFAL_XOR_v3_1/A
rlabel locali -55 -936 -35 -916 2 EESPFAL_XOR_v3_1/A_bar
rlabel locali -55 -836 -35 -816 2 EESPFAL_XOR_v3_1/B
rlabel locali -55 -736 -35 -716 2 EESPFAL_XOR_v3_1/B_bar
rlabel locali 855 -116 895 -76 2 EESPFAL_XOR_v3_1/Dis
rlabel metal1 1105 -676 1145 -636 2 EESPFAL_XOR_v3_1/OUT_bar
rlabel metal1 1055 4 1095 44 2 EESPFAL_XOR_v3_1/GND!
rlabel metal1 1055 -1176 1095 -1136 2 EESPFAL_XOR_v3_1/CLK
rlabel locali 1005 -2047 1045 -2007 4 EESPFAL_4in_NAND_0/OUT
rlabel locali -55 -1437 -35 -1417 4 EESPFAL_4in_NAND_0/A
rlabel locali -55 -1897 -35 -1877 4 EESPFAL_4in_NAND_0/A_bar
rlabel locali -55 -1557 -35 -1537 4 EESPFAL_4in_NAND_0/B
rlabel locali -55 -1997 -35 -1977 4 EESPFAL_4in_NAND_0/B_bar
rlabel locali -55 -1677 -35 -1657 4 EESPFAL_4in_NAND_0/C
rlabel locali -55 -2097 -35 -2077 4 EESPFAL_4in_NAND_0/C_bar
rlabel locali -55 -1797 -35 -1777 4 EESPFAL_4in_NAND_0/D
rlabel locali -55 -2197 -35 -2177 4 EESPFAL_4in_NAND_0/D_bar
rlabel locali 855 -2697 895 -2657 4 EESPFAL_4in_NAND_0/Dis
rlabel metal1 1105 -1907 1145 -1867 4 EESPFAL_4in_NAND_0/OUT_bar
rlabel metal1 1055 -2817 1095 -2777 4 EESPFAL_4in_NAND_0/GND!
rlabel metal1 1055 -1317 1095 -1277 4 EESPFAL_4in_NAND_0/CLK
rlabel locali 3215 -551 3255 -511 2 EESPFAL_INV4_0/OUT_bar
rlabel locali 3845 -796 3885 -756 2 EESPFAL_INV4_0/A
rlabel locali 2685 -556 2725 -516 2 EESPFAL_INV4_0/A_bar
rlabel locali 3065 -116 3105 -76 2 EESPFAL_INV4_0/Dis
rlabel metal1 3315 -676 3355 -636 2 EESPFAL_INV4_0/OUT
rlabel metal1 3265 4 3305 44 2 EESPFAL_INV4_0/GND!
rlabel metal1 3265 -1176 3305 -1136 2 EESPFAL_INV4_0/CLK
rlabel locali 3216 -2261 3256 -2221 4 EESPFAL_INV4_2/OUT_bar
rlabel locali 3846 -2016 3886 -1976 4 EESPFAL_INV4_2/A
rlabel locali 2686 -2256 2726 -2216 4 EESPFAL_INV4_2/A_bar
rlabel locali 3066 -2696 3106 -2656 4 EESPFAL_INV4_2/Dis
rlabel metal1 3316 -2136 3356 -2096 4 EESPFAL_INV4_2/OUT
rlabel metal1 3266 -2816 3306 -2776 4 EESPFAL_INV4_2/GND!
rlabel metal1 3266 -1636 3306 -1596 4 EESPFAL_INV4_2/CLK
rlabel locali 5095 -551 5135 -511 2 EESPFAL_NAND_v3_0/OUT
rlabel locali 4335 -936 4355 -916 2 EESPFAL_NAND_v3_0/A
rlabel locali 4335 -716 4355 -696 2 EESPFAL_NAND_v3_0/A_bar
rlabel locali 4335 -816 4355 -796 2 EESPFAL_NAND_v3_0/B
rlabel locali 4335 -616 4355 -596 2 EESPFAL_NAND_v3_0/B_bar
rlabel locali 4945 -116 4985 -76 2 EESPFAL_NAND_v3_0/Dis
rlabel metal1 5195 -676 5235 -636 2 EESPFAL_NAND_v3_0/OUT_bar
rlabel metal1 5145 4 5185 44 2 EESPFAL_NAND_v3_0/GND!
rlabel metal1 5145 -1176 5185 -1136 2 EESPFAL_NAND_v3_0/CLK
rlabel locali 5375 -2261 5415 -2221 6 EESPFAL_3in_NOR_v2_0/OUT
rlabel locali 6305 -1756 6325 -1736 6 EESPFAL_3in_NOR_v2_0/A
rlabel locali 6305 -2056 6325 -2036 6 EESPFAL_3in_NOR_v2_0/A_bar
rlabel locali 6305 -1866 6325 -1846 6 EESPFAL_3in_NOR_v2_0/B
rlabel locali 6305 -2176 6325 -2156 6 EESPFAL_3in_NOR_v2_0/B_bar
rlabel locali 6305 -1966 6325 -1946 6 EESPFAL_3in_NOR_v2_0/C
rlabel locali 6305 -2276 6325 -2256 6 EESPFAL_3in_NOR_v2_0/C_bar
rlabel locali 5525 -2696 5565 -2656 6 EESPFAL_3in_NOR_v2_0/Dis
rlabel metal1 5275 -2136 5315 -2096 6 EESPFAL_3in_NOR_v2_0/OUT_bar
rlabel metal1 5325 -2816 5365 -2776 6 EESPFAL_3in_NOR_v2_0/GND!
rlabel metal1 5325 -1636 5365 -1596 6 EESPFAL_3in_NOR_v2_0/CLK
rlabel locali 1005 559 1045 599 4 EESPFAL_XOR_v3_0/OUT
rlabel locali -55 1064 -35 1084 4 EESPFAL_XOR_v3_0/A
rlabel locali -55 964 -35 984 4 EESPFAL_XOR_v3_0/A_bar
rlabel locali -55 864 -35 884 4 EESPFAL_XOR_v3_0/B
rlabel locali -55 764 -35 784 4 EESPFAL_XOR_v3_0/B_bar
rlabel locali 855 124 895 164 4 EESPFAL_XOR_v3_0/Dis
rlabel metal1 1105 684 1145 724 4 EESPFAL_XOR_v3_0/OUT_bar
rlabel metal1 1055 4 1095 44 4 EESPFAL_XOR_v3_0/GND!
rlabel metal1 1055 1184 1095 1224 4 EESPFAL_XOR_v3_0/CLK
rlabel locali 3215 559 3255 599 4 EESPFAL_INV4_1/OUT_bar
rlabel locali 3845 804 3885 844 4 EESPFAL_INV4_1/A
rlabel locali 2685 564 2725 604 4 EESPFAL_INV4_1/A_bar
rlabel locali 3065 124 3105 164 4 EESPFAL_INV4_1/Dis
rlabel metal1 3315 684 3355 724 4 EESPFAL_INV4_1/OUT
rlabel metal1 3265 4 3305 44 4 EESPFAL_INV4_1/GND!
rlabel metal1 3265 1184 3305 1224 4 EESPFAL_INV4_1/CLK
rlabel locali 5095 559 5135 599 4 EESPFAL_NAND_v3_1/OUT
rlabel locali 4335 964 4355 984 4 EESPFAL_NAND_v3_1/A
rlabel locali 4335 744 4355 764 4 EESPFAL_NAND_v3_1/A_bar
rlabel locali 4335 844 4355 864 4 EESPFAL_NAND_v3_1/B
rlabel locali 4335 644 4355 664 4 EESPFAL_NAND_v3_1/B_bar
rlabel locali 4945 124 4985 164 4 EESPFAL_NAND_v3_1/Dis
rlabel metal1 5195 684 5235 724 4 EESPFAL_NAND_v3_1/OUT_bar
rlabel metal1 5145 4 5185 44 4 EESPFAL_NAND_v3_1/GND!
rlabel metal1 5145 1184 5185 1224 4 EESPFAL_NAND_v3_1/CLK
<< end >>
