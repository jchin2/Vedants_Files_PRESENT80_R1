magic
tech sky130A
magscale 1 2
timestamp 1671058898
<< poly >>
rect 778 1110 898 1140
rect 298 0 328 30
rect -50 -30 328 0
<< locali >>
rect -299 1261 1778 1284
rect -299 1227 -238 1261
rect -204 1227 -166 1261
rect -132 1227 -94 1261
rect -60 1227 -22 1261
rect 12 1227 50 1261
rect 84 1227 122 1261
rect 156 1227 194 1261
rect 228 1227 266 1261
rect 300 1227 338 1261
rect 372 1227 410 1261
rect 444 1227 482 1261
rect 516 1227 554 1261
rect 588 1227 626 1261
rect 660 1227 698 1261
rect 732 1227 770 1261
rect 804 1227 842 1261
rect 876 1227 914 1261
rect 948 1227 986 1261
rect 1020 1227 1058 1261
rect 1092 1227 1130 1261
rect 1164 1227 1202 1261
rect 1236 1227 1274 1261
rect 1308 1227 1346 1261
rect 1380 1227 1418 1261
rect 1452 1227 1490 1261
rect 1524 1227 1562 1261
rect 1596 1227 1634 1261
rect 1668 1227 1706 1261
rect 1740 1227 1778 1261
rect -299 1204 1778 1227
rect -130 380 -40 1204
rect 1308 1080 1776 1120
rect 218 -107 252 0
rect -260 -130 1751 -107
rect -260 -164 -199 -130
rect -165 -164 -127 -130
rect -93 -164 -55 -130
rect -21 -164 17 -130
rect 51 -164 89 -130
rect 123 -164 161 -130
rect 195 -164 233 -130
rect 267 -164 305 -130
rect 339 -164 377 -130
rect 411 -164 449 -130
rect 483 -164 521 -130
rect 555 -164 593 -130
rect 627 -164 665 -130
rect 699 -164 737 -130
rect 771 -164 809 -130
rect 843 -164 881 -130
rect 915 -164 953 -130
rect 987 -164 1025 -130
rect 1059 -131 1751 -130
rect 1059 -164 1097 -131
rect -260 -165 1097 -164
rect 1131 -165 1169 -131
rect 1203 -165 1241 -131
rect 1275 -165 1313 -131
rect 1347 -165 1385 -131
rect 1419 -165 1457 -131
rect 1491 -165 1529 -131
rect 1563 -165 1601 -131
rect 1635 -165 1673 -131
rect 1707 -165 1751 -131
rect -260 -187 1751 -165
<< viali >>
rect -238 1227 -204 1261
rect -166 1227 -132 1261
rect -94 1227 -60 1261
rect -22 1227 12 1261
rect 50 1227 84 1261
rect 122 1227 156 1261
rect 194 1227 228 1261
rect 266 1227 300 1261
rect 338 1227 372 1261
rect 410 1227 444 1261
rect 482 1227 516 1261
rect 554 1227 588 1261
rect 626 1227 660 1261
rect 698 1227 732 1261
rect 770 1227 804 1261
rect 842 1227 876 1261
rect 914 1227 948 1261
rect 986 1227 1020 1261
rect 1058 1227 1092 1261
rect 1130 1227 1164 1261
rect 1202 1227 1236 1261
rect 1274 1227 1308 1261
rect 1346 1227 1380 1261
rect 1418 1227 1452 1261
rect 1490 1227 1524 1261
rect 1562 1227 1596 1261
rect 1634 1227 1668 1261
rect 1706 1227 1740 1261
rect -199 -164 -165 -130
rect -127 -164 -93 -130
rect -55 -164 -21 -130
rect 17 -164 51 -130
rect 89 -164 123 -130
rect 161 -164 195 -130
rect 233 -164 267 -130
rect 305 -164 339 -130
rect 377 -164 411 -130
rect 449 -164 483 -130
rect 521 -164 555 -130
rect 593 -164 627 -130
rect 665 -164 699 -130
rect 737 -164 771 -130
rect 809 -164 843 -130
rect 881 -164 915 -130
rect 953 -164 987 -130
rect 1025 -164 1059 -130
rect 1097 -165 1131 -131
rect 1169 -165 1203 -131
rect 1241 -165 1275 -131
rect 1313 -165 1347 -131
rect 1385 -165 1419 -131
rect 1457 -165 1491 -131
rect 1529 -165 1563 -131
rect 1601 -165 1635 -131
rect 1673 -165 1707 -131
<< metal1 >>
rect -299 1261 1778 1294
rect -299 1227 -238 1261
rect -204 1227 -166 1261
rect -132 1227 -94 1261
rect -60 1227 -22 1261
rect 12 1227 50 1261
rect 84 1227 122 1261
rect 156 1227 194 1261
rect 228 1227 266 1261
rect 300 1227 338 1261
rect 372 1227 410 1261
rect 444 1227 482 1261
rect 516 1227 554 1261
rect 588 1227 626 1261
rect 660 1227 698 1261
rect 732 1227 770 1261
rect 804 1227 842 1261
rect 876 1227 914 1261
rect 948 1227 986 1261
rect 1020 1227 1058 1261
rect 1092 1227 1130 1261
rect 1164 1227 1202 1261
rect 1236 1227 1274 1261
rect 1308 1227 1346 1261
rect 1380 1227 1418 1261
rect 1452 1227 1490 1261
rect 1524 1227 1562 1261
rect 1596 1227 1634 1261
rect 1668 1227 1706 1261
rect 1740 1227 1778 1261
rect -299 1194 1778 1227
rect -260 -130 1751 -97
rect -260 -164 -199 -130
rect -165 -164 -127 -130
rect -93 -164 -55 -130
rect -21 -164 17 -130
rect 51 -164 89 -130
rect 123 -164 161 -130
rect 195 -164 233 -130
rect 267 -164 305 -130
rect 339 -164 377 -130
rect 411 -164 449 -130
rect 483 -164 521 -130
rect 555 -164 593 -130
rect 627 -164 665 -130
rect 699 -164 737 -130
rect 771 -164 809 -130
rect 843 -164 881 -130
rect 915 -164 953 -130
rect 987 -164 1025 -130
rect 1059 -131 1751 -130
rect 1059 -164 1097 -131
rect -260 -165 1097 -164
rect 1131 -165 1169 -131
rect 1203 -165 1241 -131
rect 1275 -165 1313 -131
rect 1347 -165 1385 -131
rect 1419 -165 1457 -131
rect 1491 -165 1529 -131
rect 1563 -165 1601 -131
rect 1635 -165 1673 -131
rect 1707 -165 1751 -131
rect -260 -197 1751 -165
use nmos_1v8_lvt_5p0_4finger  nmos_1v8_lvt_5p0_4finger_0
timestamp 1671058898
transform 1 0 1888 0 1 40
box -1136 -40 -364 1100
use nmos_1v8_lvt_5p0_body_4finger  nmos_1v8_lvt_5p0_body_4finger_0
timestamp 1671058898
transform 1 0 1288 0 1 40
box -1256 -40 -364 1100
use sky130_fd_pr__res_generic_po_RWRVR8  sky130_fd_pr__res_generic_po_RWRVR8_0
timestamp 1671058898
transform 1 0 -86 0 1 212
box -44 -242 44 242
<< labels >>
flabel metal1 s 664 -164 699 -130 2 FreeSans 5000 0 0 0 Ground
port 1 nsew
flabel metal1 s 626 1227 660 1261 2 FreeSans 5000 0 0 0 VDD
port 2 nsew
flabel locali s 746 -148 746 -148 2 FreeSans 5000 0 0 0 Ground
port 1 nsew
flabel locali s 1749 1090 1771 1110 2 FreeSans 5000 0 0 0 Mirror_out
port 3 nsew
<< end >>
