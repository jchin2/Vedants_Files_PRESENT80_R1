magic
tech sky130A
magscale 1 2
timestamp 1675786016
<< metal1 >>
rect -100 -13 -20 0
rect -100 -65 -86 -13
rect -34 -65 -20 -13
rect -100 -80 -20 -65
<< via1 >>
rect -86 -65 -34 -13
<< metal2 >>
rect -100 -11 -20 0
rect -100 -67 -88 -11
rect -32 -67 -20 -11
rect -100 -80 -20 -67
<< via2 >>
rect -88 -13 -32 -11
rect -88 -65 -86 -13
rect -86 -65 -34 -13
rect -34 -65 -32 -13
rect -88 -67 -32 -65
<< metal3 >>
rect -110 -11 -10 10
rect -110 -67 -88 -11
rect -32 -67 -10 -11
rect -110 -90 -10 -67
<< end >>
