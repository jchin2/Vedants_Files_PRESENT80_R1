* NGSPICE file created from INV_VP_VN.ext - technology: sky130A

.subckt INV_VP_VN A OUT VP VN
X0 OUT A VN VN sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X1 OUT A VP VP sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
.ends

