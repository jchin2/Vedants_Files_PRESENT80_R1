magic
tech sky130A
timestamp 1662787247
<< nwell >>
rect 65 160 315 475
<< nmos >>
rect 145 -25 160 125
rect 220 -25 235 125
<< pmos >>
rect 145 180 160 330
rect 220 180 235 330
<< ndiff >>
rect 85 90 145 125
rect 85 70 100 90
rect 120 70 145 90
rect 85 50 145 70
rect 85 30 100 50
rect 120 30 145 50
rect 85 10 145 30
rect 85 -10 100 10
rect 120 -10 145 10
rect 85 -25 145 -10
rect 160 90 220 125
rect 160 70 180 90
rect 200 70 220 90
rect 160 50 220 70
rect 160 30 180 50
rect 200 30 220 50
rect 160 10 220 30
rect 160 -10 180 10
rect 200 -10 220 10
rect 160 -25 220 -10
rect 235 90 295 125
rect 235 70 255 90
rect 275 70 295 90
rect 235 50 295 70
rect 235 30 255 50
rect 275 30 295 50
rect 235 10 295 30
rect 235 -10 255 10
rect 275 -10 295 10
rect 235 -25 295 -10
<< pdiff >>
rect 85 295 145 330
rect 85 275 100 295
rect 120 275 145 295
rect 85 255 145 275
rect 85 235 100 255
rect 120 235 145 255
rect 85 215 145 235
rect 85 195 100 215
rect 120 195 145 215
rect 85 180 145 195
rect 160 180 220 330
rect 235 295 295 330
rect 235 275 255 295
rect 275 275 295 295
rect 235 255 295 275
rect 235 235 255 255
rect 275 235 295 255
rect 235 215 295 235
rect 235 195 255 215
rect 275 195 295 215
rect 235 180 295 195
<< ndiffc >>
rect 100 70 120 90
rect 100 30 120 50
rect 100 -10 120 10
rect 180 70 200 90
rect 180 30 200 50
rect 180 -10 200 10
rect 255 70 275 90
rect 255 30 275 50
rect 255 -10 275 10
<< pdiffc >>
rect 100 275 120 295
rect 100 235 120 255
rect 100 195 120 215
rect 255 275 275 295
rect 255 235 275 255
rect 255 195 275 215
<< psubdiff >>
rect 85 -110 295 -95
rect 85 -130 100 -110
rect 120 -130 140 -110
rect 160 -130 180 -110
rect 200 -130 220 -110
rect 240 -130 260 -110
rect 280 -130 295 -110
rect 85 -145 295 -130
<< nsubdiff >>
rect 85 440 295 455
rect 85 420 100 440
rect 120 420 140 440
rect 160 420 180 440
rect 200 420 220 440
rect 240 420 260 440
rect 280 420 295 440
rect 85 405 295 420
<< psubdiffcont >>
rect 100 -130 120 -110
rect 140 -130 160 -110
rect 180 -130 200 -110
rect 220 -130 240 -110
rect 260 -130 280 -110
<< nsubdiffcont >>
rect 100 420 120 440
rect 140 420 160 440
rect 180 420 200 440
rect 220 420 240 440
rect 260 420 280 440
<< poly >>
rect 195 375 235 385
rect 195 355 205 375
rect 225 355 235 375
rect 195 345 235 355
rect 145 330 160 345
rect 220 330 235 345
rect 145 125 160 180
rect 220 125 235 180
rect 145 -40 160 -25
rect 120 -50 160 -40
rect 220 -45 235 -25
rect 120 -70 130 -50
rect 150 -70 160 -50
rect 120 -80 160 -70
<< polycont >>
rect 205 355 225 375
rect 130 -70 150 -50
<< locali >>
rect 85 440 295 450
rect 85 420 100 440
rect 120 420 140 440
rect 160 420 180 440
rect 200 420 220 440
rect 240 420 260 440
rect 280 420 295 440
rect 85 410 295 420
rect 195 375 235 385
rect 65 355 205 375
rect 225 355 235 375
rect 195 345 235 355
rect 90 295 130 310
rect 90 275 100 295
rect 120 275 130 295
rect 90 255 130 275
rect 90 235 100 255
rect 120 235 130 255
rect 90 215 130 235
rect 90 195 100 215
rect 120 195 130 215
rect 90 185 130 195
rect 245 295 285 310
rect 245 275 255 295
rect 275 275 285 295
rect 245 255 285 275
rect 245 235 255 255
rect 275 235 285 255
rect 245 215 285 235
rect 245 195 255 215
rect 275 195 285 215
rect 245 185 285 195
rect 245 145 265 185
rect 190 125 265 145
rect 190 105 210 125
rect 90 90 130 105
rect 90 70 100 90
rect 120 70 130 90
rect 90 50 130 70
rect 90 30 100 50
rect 120 30 130 50
rect 90 10 130 30
rect 90 -10 100 10
rect 120 -10 130 10
rect 90 -20 130 -10
rect 170 90 210 105
rect 170 70 180 90
rect 200 70 210 90
rect 170 50 210 70
rect 170 30 180 50
rect 200 30 210 50
rect 170 10 210 30
rect 170 -10 180 10
rect 200 -10 210 10
rect 170 -20 210 -10
rect 245 90 285 105
rect 245 70 255 90
rect 275 70 285 90
rect 245 50 285 70
rect 245 30 255 50
rect 275 30 285 50
rect 245 10 285 30
rect 245 -10 255 10
rect 275 -10 285 10
rect 245 -20 285 -10
rect 120 -50 160 -40
rect 65 -70 130 -50
rect 150 -70 160 -50
rect 190 -50 210 -20
rect 190 -70 315 -50
rect 120 -80 160 -70
rect 85 -110 295 -100
rect 85 -130 100 -110
rect 120 -130 140 -110
rect 160 -130 180 -110
rect 200 -130 220 -110
rect 240 -130 260 -110
rect 280 -130 295 -110
rect 85 -140 295 -130
<< viali >>
rect 100 420 120 440
rect 140 420 160 440
rect 180 420 200 440
rect 220 420 240 440
rect 260 420 280 440
rect 100 275 120 295
rect 100 235 120 255
rect 100 195 120 215
rect 100 70 120 90
rect 100 30 120 50
rect 100 -10 120 10
rect 255 70 275 90
rect 255 30 275 50
rect 255 -10 275 10
rect 100 -130 120 -110
rect 140 -130 160 -110
rect 180 -130 200 -110
rect 220 -130 240 -110
rect 260 -130 280 -110
<< metal1 >>
rect 65 440 315 455
rect 65 420 100 440
rect 120 420 140 440
rect 160 420 180 440
rect 200 420 220 440
rect 240 420 260 440
rect 280 420 315 440
rect 65 405 315 420
rect 90 295 130 405
rect 90 275 100 295
rect 120 275 130 295
rect 90 255 130 275
rect 90 235 100 255
rect 120 235 130 255
rect 90 215 130 235
rect 90 195 100 215
rect 120 195 130 215
rect 90 185 130 195
rect 90 90 130 105
rect 90 70 100 90
rect 120 70 130 90
rect 90 50 130 70
rect 90 30 100 50
rect 120 30 130 50
rect 90 10 130 30
rect 90 -10 100 10
rect 120 -10 130 10
rect 90 -20 130 -10
rect 245 90 285 105
rect 245 70 255 90
rect 275 70 285 90
rect 245 50 285 70
rect 245 30 255 50
rect 275 30 285 50
rect 245 10 285 30
rect 245 -10 255 10
rect 275 -10 285 10
rect 245 -20 285 -10
rect 100 -95 120 -20
rect 255 -95 275 -20
rect 65 -110 315 -95
rect 65 -130 100 -110
rect 120 -130 140 -110
rect 160 -130 180 -110
rect 200 -130 220 -110
rect 240 -130 260 -110
rect 280 -130 315 -110
rect 65 -145 315 -130
<< labels >>
rlabel metal1 65 -130 85 -110 7 GND!
port 5 w
rlabel metal1 65 420 85 440 7 VDD!
port 4 w
rlabel locali 295 -70 315 -50 3 OUT
port 3 e
rlabel locali 65 355 85 375 7 B
port 2 w
rlabel locali 65 -70 85 -50 7 A
port 1 w
<< end >>
