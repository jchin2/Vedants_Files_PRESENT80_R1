magic
tech sky130A
magscale 1 2
timestamp 1673382112
<< locali >>
rect -715 1054 -65 1094
rect 4315 1054 4585 1094
rect -601 954 -65 994
rect 2180 954 2555 994
rect -1171 854 -65 894
rect -1057 754 -65 794
rect 2180 654 2220 954
rect 4429 944 4585 984
rect 2408 834 2555 874
rect 4195 833 4471 873
rect 2254 734 2555 774
rect 2254 604 2294 734
rect 4195 724 4235 833
rect 4431 794 4471 833
rect 4431 754 4585 794
rect 2442 634 2555 674
rect 2215 564 2294 604
rect -255 -16 -65 64
rect 15 -116 385 -76
rect 2328 -437 2368 620
rect 2442 586 2482 634
rect 2021 -466 2368 -437
rect 1765 -477 2368 -466
rect 2402 546 2482 586
rect 1765 -506 2061 -477
rect 2402 -511 2442 546
rect 4349 530 4389 719
rect 6530 690 6554 716
rect -373 -556 385 -516
rect 2117 -551 2442 -511
rect 4279 490 4389 530
rect 4423 634 4585 674
rect 4279 -516 4319 490
rect 4423 456 4463 634
rect 2117 -636 2157 -551
rect 4235 -556 4319 -516
rect 4353 416 4463 456
rect 4501 534 4585 574
rect 6530 570 6556 597
rect 1765 -676 2157 -636
rect 2403 -626 2555 -586
rect -487 -796 385 -756
rect -943 -1306 -65 -1266
rect 2329 -1294 2369 -746
rect 2267 -1334 2369 -1294
rect -829 -1406 -65 -1366
rect -487 -1506 -65 -1466
rect -373 -1606 -65 -1566
rect 2267 -1666 2307 -1334
rect 2403 -1368 2443 -626
rect 4353 -636 4393 416
rect 4235 -676 4393 -636
rect 4501 -710 4541 534
rect 4269 -750 4541 -710
rect 2215 -1706 2307 -1666
rect 2341 -1408 2443 -1368
rect 2477 -826 2555 -786
rect 2215 -1796 2227 -1756
rect -255 -2376 -65 -2296
rect 2341 -2410 2381 -1408
rect 2477 -1442 2517 -826
rect 15 -2476 385 -2436
rect 1797 -2450 2381 -2410
rect 2415 -1482 2517 -1442
rect 1797 -2826 1837 -2450
rect 2415 -2484 2455 -1482
rect 1765 -2866 1837 -2826
rect 1871 -2524 2455 -2484
rect 2489 -1556 2705 -1516
rect -601 -2916 385 -2876
rect 1871 -2996 1911 -2524
rect 2489 -2580 2529 -1556
rect 4269 -1636 4309 -750
rect 4085 -1676 4309 -1636
rect 2263 -2620 2529 -2580
rect 2563 -1796 2705 -1756
rect 2563 -2673 2603 -1796
rect 4085 -1846 4266 -1806
rect 1765 -3036 1911 -2996
rect 2109 -2713 2603 -2673
rect -715 -3156 385 -3116
rect -373 -3656 85 -3616
rect -943 -3776 85 -3736
rect -653 -3846 -419 -3832
rect -1057 -3872 85 -3846
rect -1057 -3886 -619 -3872
rect -453 -3886 85 -3872
rect -487 -3966 85 -3926
rect 2109 -3996 2149 -2713
rect 3 -4020 85 -4006
rect -829 -4046 85 -4020
rect 2065 -4036 2149 -3996
rect -829 -4060 37 -4046
rect -1171 -4146 85 -4106
rect 2203 -4116 2243 -2827
rect 2065 -4156 2243 -4116
rect 15 -4596 85 -4556
rect -255 -4736 75 -4656
<< metal1 >>
rect -205 1154 -65 1254
rect 4171 1180 4220 1229
rect 6506 1179 6557 1228
rect -1251 -4086 -1171 1094
rect -1137 -3826 -1057 1094
rect -1023 -3716 -943 1094
rect -909 -3986 -829 1094
rect -795 -3096 -715 1094
rect -681 -2856 -601 1094
rect -567 -3906 -487 1094
rect -453 -3596 -373 1094
rect -345 -4736 -245 64
rect -205 -1106 -105 1154
rect 2348 700 2388 814
rect 4235 644 4275 1014
rect 4357 799 4397 987
rect 2215 -26 2555 74
rect 4235 -26 4575 74
rect 2369 -726 2477 -686
rect 2383 -948 2555 -908
rect -205 -1206 -65 -1106
rect -205 -3466 -105 -1206
rect 2383 -1775 2423 -948
rect 2307 -1815 2423 -1775
rect 2215 -2386 2705 -2286
rect 2203 -2747 2243 -2638
rect -205 -3566 75 -3466
<< via1 >>
rect 4149 238 4201 290
rect 4149 -242 4201 -190
<< metal2 >>
rect -65 -4516 15 1380
rect 2705 -2177 2785 1380
rect 4427 847 4505 887
rect 4135 290 4215 304
rect 4135 238 4149 290
rect 4201 238 4215 290
rect 4135 -190 4215 238
rect 4135 -242 4149 -190
rect 4201 -242 4215 -190
rect 4135 -256 4215 -242
rect 4427 -710 4467 847
rect 4693 184 4773 1380
rect 4286 -750 4467 -710
rect 4286 -1766 4326 -750
use EESPFAL_3in_NAND_v2  EESPFAL_3in_NAND_v2_0
timestamp 1501983338
transform 1 0 2705 0 1 -5146
box -2670 374 -590 1730
use EESPFAL_3in_NOR_v2  EESPFAL_3in_NOR_v2_0
timestamp 1501983338
transform 1 0 6875 0 1 -356
box -2340 304 -260 1660
use EESPFAL_INV4  EESPFAL_INV4_0
timestamp 1501983338
transform 1 0 3715 0 -1 694
box -3390 594 -1900 1950
use EESPFAL_INV4  EESPFAL_INV4_1
timestamp 1501983338
transform 1 0 6035 0 1 -3006
box -3390 594 -1900 1950
use EESPFAL_INV4  EESPFAL_INV4_2
timestamp 1501983338
transform 1 0 3715 0 -1 -1666
box -3390 594 -1900 1950
use EESPFAL_NAND_v3  EESPFAL_NAND_v3_0
timestamp 1501983338
transform 1 0 3464 0 1 628
box -949 -680 811 676
use EESPFAL_NAND_v3  EESPFAL_NAND_v3_1
timestamp 1501983338
transform 1 0 3464 0 -1 -580
box -949 -680 811 676
use EESPFAL_XOR_v3  EESPFAL_XOR_v3_0
timestamp 1501983338
transform 1 0 1225 0 1 -196
box -1330 144 1030 1500
use EESPFAL_XOR_v3  EESPFAL_XOR_v3_1
timestamp 1501983338
transform 1 0 1225 0 1 -2556
box -1330 144 1030 1500
use Li_via_M1  Li_via_M1_0
timestamp 1501983338
transform 1 0 4357 0 1 757
box -40 -38 40 42
use Li_via_M1  Li_via_M1_1
timestamp 1501983338
transform 1 0 4402 0 1 945
box -40 -38 40 42
use Li_via_M1  Li_via_M1_2
timestamp 1501983338
transform 1 0 4275 0 1 1052
box -40 -38 40 42
use Li_via_M1  Li_via_M1_3
timestamp 1501983338
transform 1 0 4275 0 1 602
box -40 -38 40 42
use Li_via_M1  Li_via_M1_4
timestamp 1501983338
transform 1 0 2368 0 1 852
box -40 -38 40 42
use Li_via_M1  Li_via_M1_5
timestamp 1501983338
transform 1 0 -1097 0 1 752
box -40 -38 40 42
use Li_via_M1  Li_via_M1_6
timestamp 1501983338
transform 1 0 -641 0 1 972
box -40 -38 40 42
use Li_via_M1  Li_via_M1_7
timestamp 1501983338
transform 1 0 -755 0 1 1052
box -40 -38 40 42
use Li_via_M1  Li_via_M1_8
timestamp 1501983338
transform 1 0 -1211 0 1 872
box -40 -38 40 42
use Li_via_M1  Li_via_M1_9
timestamp 1501983338
transform 1 0 2368 0 1 658
box -40 -38 40 42
use Li_via_M1  Li_via_M1_10
timestamp 1501983338
transform 1 0 -413 0 1 -558
box -40 -38 40 42
use Li_via_M1  Li_via_M1_11
timestamp 1501983338
transform 1 0 -295 0 1 22
box -40 -38 40 42
use Li_via_M1  Li_via_M1_12
timestamp 1501983338
transform 1 0 2329 0 1 -708
box -40 -38 40 42
use Li_via_M1  Li_via_M1_13
timestamp 1501983338
transform 1 0 2267 0 1 -1798
box -40 -38 40 42
use Li_via_M1  Li_via_M1_14
timestamp 1501983338
transform 1 0 2517 0 1 -708
box -40 -38 40 42
use Li_via_M1  Li_via_M1_15
timestamp 1501983338
transform 1 0 2595 0 1 -928
box -40 -38 40 42
use Li_via_M1  Li_via_M1_16
timestamp 1501983338
transform 1 0 -527 0 1 -798
box -40 -38 40 42
use Li_via_M1  Li_via_M1_17
timestamp 1501983338
transform 1 0 -983 0 1 -1308
box -40 -38 40 42
use Li_via_M1  Li_via_M1_18
timestamp 1501983338
transform 1 0 -869 0 1 -1408
box -40 -38 40 42
use Li_via_M1  Li_via_M1_19
timestamp 1501983338
transform 1 0 -527 0 1 -1508
box -40 -38 40 42
use Li_via_M1  Li_via_M1_20
timestamp 1501983338
transform 1 0 -413 0 1 -1608
box -40 -38 40 42
use Li_via_M1  Li_via_M1_21
timestamp 1501983338
transform 1 0 2223 0 1 -2789
box -40 -38 40 42
use Li_via_M1  Li_via_M1_22
timestamp 1501983338
transform 1 0 2223 0 1 -2601
box -40 -38 40 42
use Li_via_M1  Li_via_M1_23
timestamp 1501983338
transform 1 0 -641 0 1 -2898
box -40 -38 40 42
use Li_via_M1  Li_via_M1_24
timestamp 1501983338
transform 1 0 -755 0 1 -3138
box -40 -38 40 42
use Li_via_M1  Li_via_M1_25
timestamp 1501983338
transform 1 0 -295 0 1 -2338
box -40 -38 40 42
use Li_via_M1  Li_via_M1_26
timestamp 1501983338
transform 1 0 -983 0 1 -3758
box -40 -38 40 42
use Li_via_M1  Li_via_M1_27
timestamp 1501983338
transform 1 0 -869 0 1 -4022
box -40 -38 40 42
use Li_via_M1  Li_via_M1_28
timestamp 1501983338
transform 1 0 -1097 0 1 -3868
box -40 -38 40 42
use Li_via_M1  Li_via_M1_29
timestamp 1501983338
transform 1 0 -413 0 1 -3638
box -40 -38 40 42
use Li_via_M1  Li_via_M1_30
timestamp 1501983338
transform 1 0 -527 0 1 -3948
box -40 -38 40 42
use Li_via_M1  Li_via_M1_31
timestamp 1501983338
transform 1 0 -295 0 1 -4698
box -40 -38 40 42
use Li_via_M1  Li_via_M1_32
timestamp 1501983338
transform 1 0 -1211 0 1 -4128
box -40 -38 40 42
use Li_via_M2  Li_via_M2_0
timestamp 1501983338
transform 1 0 4733 0 1 142
box -40 -38 40 42
use Li_via_M2  Li_via_M2_1
timestamp 1501983338
transform 1 0 4306 0 1 -1808
box -40 -38 40 42
use Li_via_M2  Li_via_M2_2
timestamp 1501983338
transform 1 0 4545 0 1 866
box -40 -38 40 42
use Li_via_M2  Li_via_M2_3
timestamp 1501983338
transform 1 0 2745 0 1 142
box -40 -38 40 42
use Li_via_M2  Li_via_M2_4
timestamp 1501983338
transform 1 0 2745 0 1 -98
box -40 -38 40 42
use Li_via_M2  Li_via_M2_5
timestamp 1501983338
transform 1 0 -25 0 1 -108
box -40 -38 40 42
use Li_via_M2  Li_via_M2_6
timestamp 1501983338
transform 1 0 -25 0 1 142
box -40 -38 40 42
use Li_via_M2  Li_via_M2_7
timestamp 1501983338
transform 1 0 2745 0 1 -2219
box -40 -38 40 42
use Li_via_M2  Li_via_M2_8
timestamp 1501983338
transform 1 0 -25 0 1 -2218
box -40 -38 40 42
use Li_via_M2  Li_via_M2_9
timestamp 1501983338
transform 1 0 -25 0 1 -2468
box -40 -38 40 42
use Li_via_M2  Li_via_M2_10
timestamp 1501983338
transform 1 0 -25 0 1 -4558
box -40 -38 40 42
<< labels >>
flabel locali s 6530 690 6554 716 2 FreeSans 2000 0 0 0 s1_bar
port 1 nsew
flabel locali s 6530 570 6556 597 2 FreeSans 2000 0 0 0 s1
port 2 nsew
flabel metal1 s 6506 1179 6557 1228 2 FreeSans 2000 0 0 0 CLK3
port 3 nsew
flabel metal1 s -1241 1020 -1180 1080 2 FreeSans 2500 0 0 0 x0
port 4 nsew
flabel metal1 s -1128 959 -1067 1019 2 FreeSans 2500 0 0 0 x0_bar
port 5 nsew
flabel metal1 s -1013 1020 -952 1080 2 FreeSans 2500 0 0 0 x1
port 6 nsew
flabel metal1 s -899 959 -838 1019 2 FreeSans 2500 0 0 0 x1_bar
port 7 nsew
flabel metal1 s -785 1021 -724 1081 2 FreeSans 2500 0 0 0 x2
port 8 nsew
flabel metal1 s -672 960 -611 1020 2 FreeSans 2500 0 0 0 x2_bar
port 9 nsew
flabel metal1 s -557 1021 -496 1081 2 FreeSans 2500 0 0 0 x3
port 10 nsew
flabel metal1 s -443 960 -382 1020 2 FreeSans 2500 0 0 0 x3_bar
port 11 nsew
flabel metal1 s 4171 1180 4220 1229 2 FreeSans 2500 0 0 0 CLK2
port 12 nsew
flabel metal1 s -180 1176 -128 1230 2 FreeSans 2500 0 0 0 CLK1
port 13 nsew
flabel metal1 s -319 -1 -271 48 2 FreeSans 2500 0 0 0 GND
port 14 nsew
flabel locali s 2601 -808 2601 -808 2 FreeSans 2500 0 0 0 x2_bar_buff
port 15 nsew
flabel locali s 2597 -609 2597 -609 2 FreeSans 2500 0 0 0 x2_buff
port 16 nsew
flabel metal2 s 4708 1319 4759 1371 2 FreeSans 2000 0 0 0 Dis3
port 17 nsew
flabel metal2 s -50 1319 1 1367 2 FreeSans 2500 0 0 0 Dis1
port 18 nsew
flabel metal2 s 2720 1320 2772 1371 2 FreeSans 2500 0 0 0 Dis2
port 19 nsew
<< properties >>
string path 23.665 0.920 23.665 6.900 
<< end >>
