magic
tech sky130A
magscale 1 2
timestamp 1670967196
<< error_p >>
rect 17 -300 41 300
<< locali >>
rect -17 300 17 357
rect -17 -357 17 -300
<< rlocali >>
rect -17 -300 17 300
<< properties >>
string gencell sky130_fd_pr__res_generic_l1
string library sky130
string parameters w 0.17 l 3 m 1 nx 1 wmin 0.17 lmin 0.17 rho 12.8 val 225.882 dummy 0 dw 0.0 term 0.0 snake 1 roverlap 0
<< end >>
