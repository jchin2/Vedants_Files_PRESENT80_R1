magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect 184 552 217 585
<< l67d20 >>
rect 184 552 217 585
<< l66d20 >>
rect 187 555 214 582
<< l66d44 >>
rect 192 560 209 577
<< end >>
