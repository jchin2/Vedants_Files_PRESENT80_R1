magic
tech sky130A
timestamp 1671246442
<< pwell >>
rect -660 495 270 520
rect -658 -3 268 495
<< nmoslvt >>
rect -495 10 -480 505
rect -420 10 -405 505
rect -345 10 -330 505
rect -270 10 -255 505
rect -195 10 -180 505
rect -120 10 -105 505
rect -45 10 -30 505
rect 30 10 45 505
rect 105 10 120 505
rect 180 10 195 505
<< ndiff >>
rect -555 495 -495 505
rect -555 30 -535 495
rect -515 30 -495 495
rect -555 10 -495 30
rect -480 495 -420 505
rect -480 30 -460 495
rect -440 30 -420 495
rect -480 10 -420 30
rect -405 495 -345 505
rect -405 30 -385 495
rect -365 30 -345 495
rect -405 10 -345 30
rect -330 495 -270 505
rect -330 30 -310 495
rect -290 30 -270 495
rect -330 10 -270 30
rect -255 495 -195 505
rect -255 30 -235 495
rect -215 30 -195 495
rect -255 10 -195 30
rect -180 495 -120 505
rect -180 30 -160 495
rect -140 30 -120 495
rect -180 10 -120 30
rect -105 495 -45 505
rect -105 30 -85 495
rect -65 30 -45 495
rect -105 10 -45 30
rect -30 495 30 505
rect -30 30 -10 495
rect 10 30 30 495
rect -30 10 30 30
rect 45 495 105 505
rect 45 30 65 495
rect 85 30 105 495
rect 45 10 105 30
rect 120 495 180 505
rect 120 30 140 495
rect 160 30 180 495
rect 120 10 180 30
rect 195 495 255 505
rect 195 30 215 495
rect 235 30 255 495
rect 195 10 255 30
<< ndiffc >>
rect -535 30 -515 495
rect -460 30 -440 495
rect -385 30 -365 495
rect -310 30 -290 495
rect -235 30 -215 495
rect -160 30 -140 495
rect -85 30 -65 495
rect -10 30 10 495
rect 65 30 85 495
rect 140 30 160 495
rect 215 30 235 495
<< psubdiff >>
rect -645 495 -585 505
rect -645 30 -625 495
rect -605 30 -585 495
rect -645 10 -585 30
<< psubdiffcont >>
rect -625 30 -605 495
<< poly >>
rect -495 505 -480 520
rect -420 505 -405 520
rect -345 505 -330 520
rect -270 505 -255 520
rect -195 505 -180 520
rect -120 505 -105 520
rect -45 505 -30 520
rect 30 505 45 520
rect 105 505 120 520
rect 180 505 195 520
rect -495 -5 -480 10
rect -420 -5 -405 10
rect -345 -5 -330 10
rect -270 -5 -255 10
rect -195 -5 -180 10
rect -120 -5 -105 10
rect -45 -5 -30 10
rect 30 -5 45 10
rect 105 -5 120 10
rect 180 -5 195 10
<< locali >>
rect -635 30 -625 495
rect -605 30 -595 495
rect -635 20 -595 30
rect -545 30 -535 495
rect -515 30 -505 495
rect -545 20 -505 30
rect -470 30 -460 495
rect -440 30 -430 495
rect -470 20 -430 30
rect -395 30 -385 495
rect -365 30 -355 495
rect -395 20 -355 30
rect -320 30 -310 495
rect -290 30 -280 495
rect -320 20 -280 30
rect -245 30 -235 495
rect -215 30 -205 495
rect -245 20 -205 30
rect -170 30 -160 495
rect -140 30 -130 495
rect -170 20 -130 30
rect -95 30 -85 495
rect -65 30 -55 495
rect -95 20 -55 30
rect -20 30 -10 495
rect 10 30 20 495
rect -20 20 20 30
rect 55 30 65 495
rect 85 30 95 495
rect 55 20 95 30
rect 130 30 140 495
rect 160 30 170 495
rect 130 20 170 30
rect 205 30 215 495
rect 235 30 245 495
rect 205 20 245 30
<< end >>
