magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -2530 -2690 15070 14910
<< l71d20 >>
rect -130 140 -30 12410
rect 65 12410 12370 12510
rect 12570 5 12670 12350
rect -130 -290 12670 -190
rect -430 745 -330 12510
rect -430 12710 12675 12810
rect 12870 -290 12970 12650
rect -430 -590 12670 -490
rect -730 -290 -630 12810
rect -430 13010 12970 13110
rect -1030 -590 -930 13110
rect -1330 -890 -1230 13410
rect -1630 -1190 -1530 13710
rect -1930 -1490 -1830 14010
rect -2230 -1790 -2130 14310
rect -2530 -2090 -2430 14610
rect -430 13010 12670 13110
rect 13170 -290 13270 12810
rect -731 -890 12370 -790
rect 6170 -2690 14470 -2590
rect 13570 13610 13770 13710
rect 13770 13410 13870 13710
rect 14070 13710 14170 14010
rect 13870 13910 14070 14010
rect 14370 14010 14470 14310
rect 14170 14210 14370 14310
rect 14670 14310 14770 14610
rect 14470 14510 14670 14610
rect 14970 14610 15070 14910
rect 14770 14810 14970 14910
rect 12370 12410 12570 12510
rect 12570 12350 12670 12510
rect 13170 12805 13270 13010
rect 12970 13010 13270 13110
rect 12675 12710 12925 12810
rect 12870 12650 12970 12810
rect 13270 13310 13470 13410
rect 13470 13110 13570 13410
rect 13570 13610 13770 13710
rect 13770 13410 13870 13710
rect -1230 13610 -1030 13710
rect -1330 13410 -1230 13710
rect -1230 13610 -1030 13710
rect -1330 13410 -1230 13710
rect -1630 13710 -1530 14010
rect -1530 13910 -1330 14010
rect -1930 14010 -1830 14310
rect -1830 14210 -1630 14310
rect -2230 14310 -2130 14610
rect -2130 14510 -1930 14610
rect -2530 14610 -2430 14910
rect -2430 14810 -2230 14910
rect -430 12510 -330 12710
rect -730 12810 -630 13010
rect -730 13010 -430 13110
rect -130 12410 65 12510
rect -930 13310 -730 13410
rect -1030 13110 -930 13410
rect -1930 -1790 -1830 -1490
rect -1830 -1790 -1630 -1690
rect -2230 -2090 -2130 -1790
rect -2130 -2090 -1930 -1990
rect -2530 -2390 -2430 -2090
rect -2430 -2390 -2230 -2290
rect -630 -590 -430 -490
rect -730 -590 -630 -290
rect -130 10 -30 140
rect -30 10 165 110
rect -330 -290 -130 -190
rect -430 -290 -330 -135
rect -430 -135 -330 745
rect 165 10 6170 110
rect -930 -890 -730 -790
rect -1030 -890 -930 -590
rect -1230 -1190 -1030 -1090
rect -1330 -1190 -1230 -890
rect -1230 -1190 -1030 -1090
rect -1330 -1190 -1230 -890
rect -1630 -1490 -1530 -1190
rect -1530 -1490 -1330 -1390
rect 14670 -2390 14770 -2090
rect 14170 -2090 14370 -1990
rect 14370 -2090 14470 -1790
rect 13870 -1790 14070 -1690
rect 14070 -1790 14170 -1490
rect 13570 -1490 13770 -1390
rect 13770 -1490 13870 -1190
rect 13470 -1190 13570 -890
rect 13270 -1190 13470 -1090
rect 13470 -1190 13570 -890
rect 13270 -1190 13470 -1090
rect 13170 -890 13270 -590
rect 12970 -890 13170 -790
rect 12670 -590 12970 -490
rect 12570 -190 12670 5
rect 13170 -590 13270 -290
rect 12870 -490 12970 -290
rect 12370 -890 12970 -790
rect 12970 -1190 13270 -1090
rect 13270 -1490 13570 -1390
rect 13570 -1790 13870 -1690
rect 13870 -2090 14170 -1990
rect 14170 -2390 14470 -2290
rect 14770 -2690 14970 -2590
rect 14970 -2690 15070 -2390
rect 14470 -2690 14770 -2590
rect 14470 -2390 14670 -2290
rect -730 13310 13270 13410
rect -1030 13610 13570 13710
rect -1330 13910 13870 14010
rect -1630 14210 14170 14310
rect -1930 14510 14470 14610
rect -2230 14810 14770 14910
rect -2230 14810 14770 14910
rect -1930 14510 14470 14610
rect -1630 14210 14170 14310
rect -1330 13910 13870 14010
rect -1030 13610 13570 13710
rect -730 13310 13270 13410
rect 14970 -2390 15070 14610
rect 14670 -2090 14770 14310
rect 14370 -1790 14470 14010
rect 14070 -1490 14170 13710
rect 13770 -1190 13870 13410
rect 13470 -890 13570 13110
rect -1031 -1190 12970 -1090
rect -1331 -1490 13270 -1390
rect -1631 -1790 13570 -1690
rect -1931 -2090 13870 -1990
rect -2231 -2390 14170 -2290
<< end >>
