magic
tech sky130A
timestamp 1667345354
<< nwell >>
rect -1215 835 -35 930
rect -830 640 -420 835
<< nmos >>
rect -1135 385 -1120 535
rect -1060 385 -1045 535
rect -985 385 -970 535
rect -910 385 -895 535
rect -745 385 -730 535
rect -670 385 -655 535
rect -595 385 -580 535
rect -520 385 -505 535
rect -355 385 -340 535
rect -280 385 -265 535
rect -205 385 -190 535
rect -130 385 -115 535
<< pmos >>
rect -745 665 -730 815
rect -670 665 -655 815
rect -595 665 -580 815
rect -520 665 -505 815
<< ndiff >>
rect -1195 500 -1135 535
rect -1195 480 -1175 500
rect -1155 480 -1135 500
rect -1195 460 -1135 480
rect -1195 440 -1175 460
rect -1155 440 -1135 460
rect -1195 420 -1135 440
rect -1195 400 -1175 420
rect -1155 400 -1135 420
rect -1195 385 -1135 400
rect -1120 385 -1060 535
rect -1045 500 -985 535
rect -1045 480 -1025 500
rect -1005 480 -985 500
rect -1045 460 -985 480
rect -1045 440 -1025 460
rect -1005 440 -985 460
rect -1045 420 -985 440
rect -1045 400 -1025 420
rect -1005 400 -985 420
rect -1045 385 -985 400
rect -970 385 -910 535
rect -895 500 -835 535
rect -895 480 -875 500
rect -855 480 -835 500
rect -895 460 -835 480
rect -895 440 -875 460
rect -855 440 -835 460
rect -895 420 -835 440
rect -895 400 -875 420
rect -855 400 -835 420
rect -895 385 -835 400
rect -805 500 -745 535
rect -805 480 -785 500
rect -765 480 -745 500
rect -805 460 -745 480
rect -805 440 -785 460
rect -765 440 -745 460
rect -805 420 -745 440
rect -805 400 -785 420
rect -765 400 -745 420
rect -805 385 -745 400
rect -730 500 -670 535
rect -730 480 -710 500
rect -690 480 -670 500
rect -730 460 -670 480
rect -730 440 -710 460
rect -690 440 -670 460
rect -730 420 -670 440
rect -730 400 -710 420
rect -690 400 -670 420
rect -730 385 -670 400
rect -655 500 -595 535
rect -655 480 -635 500
rect -615 480 -595 500
rect -655 460 -595 480
rect -655 440 -635 460
rect -615 440 -595 460
rect -655 420 -595 440
rect -655 400 -635 420
rect -615 400 -595 420
rect -655 385 -595 400
rect -580 500 -520 535
rect -580 480 -560 500
rect -540 480 -520 500
rect -580 460 -520 480
rect -580 440 -560 460
rect -540 440 -520 460
rect -580 420 -520 440
rect -580 400 -560 420
rect -540 400 -520 420
rect -580 385 -520 400
rect -505 500 -445 535
rect -505 480 -485 500
rect -465 480 -445 500
rect -505 460 -445 480
rect -505 440 -485 460
rect -465 440 -445 460
rect -505 420 -445 440
rect -505 400 -485 420
rect -465 400 -445 420
rect -505 385 -445 400
rect -415 500 -355 535
rect -415 480 -395 500
rect -375 480 -355 500
rect -415 460 -355 480
rect -415 440 -395 460
rect -375 440 -355 460
rect -415 420 -355 440
rect -415 400 -395 420
rect -375 400 -355 420
rect -415 385 -355 400
rect -340 385 -280 535
rect -265 500 -205 535
rect -265 480 -245 500
rect -225 480 -205 500
rect -265 460 -205 480
rect -265 440 -245 460
rect -225 440 -205 460
rect -265 420 -205 440
rect -265 400 -245 420
rect -225 400 -205 420
rect -265 385 -205 400
rect -190 385 -130 535
rect -115 500 -55 535
rect -115 480 -95 500
rect -75 480 -55 500
rect -115 460 -55 480
rect -115 440 -95 460
rect -75 440 -55 460
rect -115 420 -55 440
rect -115 400 -95 420
rect -75 400 -55 420
rect -115 385 -55 400
<< pdiff >>
rect -805 780 -745 815
rect -805 760 -785 780
rect -765 760 -745 780
rect -805 740 -745 760
rect -805 720 -785 740
rect -765 720 -745 740
rect -805 700 -745 720
rect -805 680 -785 700
rect -765 680 -745 700
rect -805 665 -745 680
rect -730 780 -670 815
rect -730 760 -710 780
rect -690 760 -670 780
rect -730 740 -670 760
rect -730 720 -710 740
rect -690 720 -670 740
rect -730 700 -670 720
rect -730 680 -710 700
rect -690 680 -670 700
rect -730 665 -670 680
rect -655 780 -595 815
rect -655 760 -635 780
rect -615 760 -595 780
rect -655 740 -595 760
rect -655 720 -635 740
rect -615 720 -595 740
rect -655 700 -595 720
rect -655 680 -635 700
rect -615 680 -595 700
rect -655 665 -595 680
rect -580 780 -520 815
rect -580 760 -560 780
rect -540 760 -520 780
rect -580 740 -520 760
rect -580 720 -560 740
rect -540 720 -520 740
rect -580 700 -520 720
rect -580 680 -560 700
rect -540 680 -520 700
rect -580 665 -520 680
rect -505 780 -445 815
rect -505 760 -485 780
rect -465 760 -445 780
rect -505 740 -445 760
rect -505 720 -485 740
rect -465 720 -445 740
rect -505 700 -445 720
rect -505 680 -485 700
rect -465 680 -445 700
rect -505 665 -445 680
<< ndiffc >>
rect -1175 480 -1155 500
rect -1175 440 -1155 460
rect -1175 400 -1155 420
rect -1025 480 -1005 500
rect -1025 440 -1005 460
rect -1025 400 -1005 420
rect -875 480 -855 500
rect -875 440 -855 460
rect -875 400 -855 420
rect -785 480 -765 500
rect -785 440 -765 460
rect -785 400 -765 420
rect -710 480 -690 500
rect -710 440 -690 460
rect -710 400 -690 420
rect -635 480 -615 500
rect -635 440 -615 460
rect -635 400 -615 420
rect -560 480 -540 500
rect -560 440 -540 460
rect -560 400 -540 420
rect -485 480 -465 500
rect -485 440 -465 460
rect -485 400 -465 420
rect -395 480 -375 500
rect -395 440 -375 460
rect -395 400 -375 420
rect -245 480 -225 500
rect -245 440 -225 460
rect -245 400 -225 420
rect -95 480 -75 500
rect -95 440 -75 460
rect -95 400 -75 420
<< pdiffc >>
rect -785 760 -765 780
rect -785 720 -765 740
rect -785 680 -765 700
rect -710 760 -690 780
rect -710 720 -690 740
rect -710 680 -690 700
rect -635 760 -615 780
rect -635 720 -615 740
rect -635 680 -615 700
rect -560 760 -540 780
rect -560 720 -540 740
rect -560 680 -540 700
rect -485 760 -465 780
rect -485 720 -465 740
rect -485 680 -465 700
<< psubdiff >>
rect -1195 300 -55 315
rect -1195 280 -1155 300
rect -1135 280 -1115 300
rect -1095 280 -1075 300
rect -1055 280 -1035 300
rect -1015 280 -995 300
rect -975 280 -955 300
rect -935 280 -915 300
rect -895 280 -875 300
rect -855 280 -835 300
rect -815 280 -795 300
rect -775 280 -755 300
rect -735 280 -715 300
rect -695 280 -675 300
rect -655 280 -635 300
rect -615 280 -595 300
rect -575 280 -555 300
rect -535 280 -515 300
rect -495 280 -475 300
rect -455 280 -435 300
rect -415 280 -395 300
rect -375 280 -355 300
rect -335 280 -315 300
rect -295 280 -275 300
rect -255 280 -235 300
rect -215 280 -195 300
rect -175 280 -155 300
rect -135 280 -115 300
rect -95 280 -55 300
rect -1195 265 -55 280
<< nsubdiff >>
rect -1195 890 -55 905
rect -1195 870 -1155 890
rect -1135 870 -1115 890
rect -1095 870 -1075 890
rect -1055 870 -1035 890
rect -1015 870 -995 890
rect -975 870 -955 890
rect -935 870 -915 890
rect -895 870 -875 890
rect -855 870 -835 890
rect -815 870 -795 890
rect -775 870 -755 890
rect -735 870 -715 890
rect -695 870 -675 890
rect -655 870 -635 890
rect -615 870 -595 890
rect -575 870 -555 890
rect -535 870 -515 890
rect -495 870 -475 890
rect -455 870 -435 890
rect -415 870 -395 890
rect -375 870 -355 890
rect -335 870 -315 890
rect -295 870 -275 890
rect -255 870 -235 890
rect -215 870 -195 890
rect -175 870 -155 890
rect -135 870 -115 890
rect -95 870 -55 890
rect -1195 855 -55 870
<< psubdiffcont >>
rect -1155 280 -1135 300
rect -1115 280 -1095 300
rect -1075 280 -1055 300
rect -1035 280 -1015 300
rect -995 280 -975 300
rect -955 280 -935 300
rect -915 280 -895 300
rect -875 280 -855 300
rect -835 280 -815 300
rect -795 280 -775 300
rect -755 280 -735 300
rect -715 280 -695 300
rect -675 280 -655 300
rect -635 280 -615 300
rect -595 280 -575 300
rect -555 280 -535 300
rect -515 280 -495 300
rect -475 280 -455 300
rect -435 280 -415 300
rect -395 280 -375 300
rect -355 280 -335 300
rect -315 280 -295 300
rect -275 280 -255 300
rect -235 280 -215 300
rect -195 280 -175 300
rect -155 280 -135 300
rect -115 280 -95 300
<< nsubdiffcont >>
rect -1155 870 -1135 890
rect -1115 870 -1095 890
rect -1075 870 -1055 890
rect -1035 870 -1015 890
rect -995 870 -975 890
rect -955 870 -935 890
rect -915 870 -895 890
rect -875 870 -855 890
rect -835 870 -815 890
rect -795 870 -775 890
rect -755 870 -735 890
rect -715 870 -695 890
rect -675 870 -655 890
rect -635 870 -615 890
rect -595 870 -575 890
rect -555 870 -535 890
rect -515 870 -495 890
rect -475 870 -455 890
rect -435 870 -415 890
rect -395 870 -375 890
rect -355 870 -335 890
rect -315 870 -295 890
rect -275 870 -255 890
rect -235 870 -215 890
rect -195 870 -175 890
rect -155 870 -135 890
rect -115 870 -95 890
<< poly >>
rect -1000 825 -960 835
rect -1000 805 -990 825
rect -970 805 -960 825
rect -745 830 -655 845
rect -745 815 -730 830
rect -670 815 -655 830
rect -595 830 -505 845
rect -595 815 -580 830
rect -520 815 -505 830
rect -305 825 -265 835
rect -1000 795 -960 805
rect -1060 775 -1020 785
rect -1060 755 -1050 775
rect -1030 755 -1020 775
rect -1060 745 -1020 755
rect -1160 675 -1120 685
rect -1160 655 -1150 675
rect -1130 655 -1120 675
rect -1160 645 -1120 655
rect -1135 535 -1120 645
rect -1060 535 -1045 745
rect -985 535 -970 795
rect -935 725 -895 735
rect -935 705 -925 725
rect -905 705 -895 725
rect -935 695 -895 705
rect -910 535 -895 695
rect -305 805 -295 825
rect -275 805 -265 825
rect -305 795 -265 805
rect -355 675 -315 685
rect -745 650 -730 665
rect -670 590 -655 665
rect -595 650 -580 665
rect -520 650 -505 665
rect -355 655 -345 675
rect -325 655 -315 675
rect -620 640 -580 650
rect -620 620 -610 640
rect -590 620 -580 640
rect -620 610 -580 620
rect -670 580 -630 590
rect -670 560 -660 580
rect -640 560 -630 580
rect -670 550 -630 560
rect -745 535 -730 550
rect -670 535 -655 550
rect -595 535 -580 610
rect -355 645 -315 655
rect -520 535 -505 550
rect -355 535 -340 645
rect -280 535 -265 795
rect -205 775 -165 785
rect -205 755 -195 775
rect -175 755 -165 775
rect -205 745 -165 755
rect -205 535 -190 745
rect -130 725 -90 735
rect -130 705 -120 725
rect -100 705 -90 725
rect -130 695 -90 705
rect -130 535 -115 695
rect -1135 370 -1120 385
rect -1060 370 -1045 385
rect -985 370 -970 385
rect -910 370 -895 385
rect -745 370 -730 385
rect -670 370 -655 385
rect -595 370 -580 385
rect -520 370 -505 385
rect -355 370 -340 385
rect -745 360 -705 370
rect -745 340 -735 360
rect -715 340 -705 360
rect -745 330 -705 340
rect -545 360 -505 370
rect -280 365 -265 385
rect -205 365 -190 385
rect -130 365 -115 385
rect -545 340 -535 360
rect -515 340 -505 360
rect -545 330 -505 340
<< polycont >>
rect -990 805 -970 825
rect -1050 755 -1030 775
rect -1150 655 -1130 675
rect -925 705 -905 725
rect -295 805 -275 825
rect -345 655 -325 675
rect -610 620 -590 640
rect -660 560 -640 580
rect -195 755 -175 775
rect -120 705 -100 725
rect -735 340 -715 360
rect -535 340 -515 360
<< locali >>
rect -1195 890 -55 900
rect -1195 870 -1155 890
rect -1135 870 -1115 890
rect -1095 870 -1075 890
rect -1055 870 -1035 890
rect -1015 870 -995 890
rect -975 870 -955 890
rect -935 870 -915 890
rect -895 870 -875 890
rect -855 870 -835 890
rect -815 870 -795 890
rect -775 870 -755 890
rect -735 870 -715 890
rect -695 870 -675 890
rect -655 870 -635 890
rect -615 870 -595 890
rect -575 870 -555 890
rect -535 870 -515 890
rect -495 870 -475 890
rect -455 870 -435 890
rect -415 870 -395 890
rect -375 870 -355 890
rect -335 870 -315 890
rect -295 870 -275 890
rect -255 870 -235 890
rect -215 870 -195 890
rect -175 870 -155 890
rect -135 870 -115 890
rect -95 870 -55 890
rect -1195 860 -55 870
rect -1000 825 -960 835
rect -935 825 -895 835
rect -1195 805 -990 825
rect -970 805 -925 825
rect -905 805 -895 825
rect -1000 795 -960 805
rect -935 795 -895 805
rect -305 825 -265 835
rect -305 805 -295 825
rect -275 805 -265 825
rect -305 795 -265 805
rect -1060 775 -1020 785
rect -870 775 -830 785
rect -1195 755 -1050 775
rect -1030 755 -860 775
rect -840 755 -830 775
rect -1060 745 -1020 755
rect -870 745 -830 755
rect -795 780 -755 795
rect -795 760 -785 780
rect -765 760 -755 780
rect -795 740 -755 760
rect -935 725 -895 735
rect -1195 705 -925 725
rect -905 705 -895 725
rect -935 695 -895 705
rect -795 720 -785 740
rect -765 720 -755 740
rect -795 700 -755 720
rect -1160 675 -1120 685
rect -870 675 -830 685
rect -1195 655 -1150 675
rect -1130 655 -860 675
rect -840 655 -830 675
rect -795 680 -785 700
rect -765 680 -755 700
rect -795 670 -755 680
rect -720 780 -680 795
rect -720 760 -710 780
rect -690 760 -680 780
rect -720 740 -680 760
rect -720 720 -710 740
rect -690 720 -680 740
rect -720 700 -680 720
rect -720 680 -710 700
rect -690 680 -680 700
rect -720 665 -680 680
rect -645 780 -605 795
rect -645 760 -635 780
rect -615 760 -605 780
rect -645 740 -605 760
rect -645 720 -635 740
rect -615 720 -605 740
rect -645 700 -605 720
rect -645 680 -635 700
rect -615 680 -605 700
rect -645 670 -605 680
rect -570 780 -530 795
rect -570 760 -560 780
rect -540 760 -530 780
rect -570 740 -530 760
rect -570 720 -560 740
rect -540 720 -530 740
rect -570 700 -530 720
rect -570 680 -560 700
rect -540 680 -530 700
rect -570 665 -530 680
rect -495 780 -455 795
rect -495 760 -485 780
rect -465 760 -455 780
rect -495 740 -455 760
rect -205 775 -165 785
rect -205 755 -195 775
rect -175 755 -165 775
rect -205 745 -165 755
rect -495 720 -485 740
rect -465 720 -455 740
rect -495 700 -455 720
rect -495 680 -485 700
rect -465 680 -455 700
rect -130 725 -90 735
rect -130 705 -120 725
rect -100 705 -90 725
rect -130 695 -90 705
rect -495 670 -455 680
rect -355 675 -315 685
rect -1160 645 -1120 655
rect -870 645 -830 655
rect -710 640 -690 665
rect -620 640 -580 650
rect -710 620 -610 640
rect -590 620 -580 640
rect -710 555 -690 620
rect -620 610 -580 620
rect -1175 535 -690 555
rect -670 580 -630 590
rect -560 580 -540 665
rect -355 655 -345 675
rect -325 655 -315 675
rect -355 645 -315 655
rect -435 635 -395 645
rect -435 615 -425 635
rect -405 625 -395 635
rect -405 615 -55 625
rect -435 605 -55 615
rect -670 560 -660 580
rect -640 560 -55 580
rect -670 550 -630 560
rect -560 535 -540 560
rect -1175 515 -1155 535
rect -875 515 -855 535
rect -1185 500 -1145 515
rect -1185 480 -1175 500
rect -1155 480 -1145 500
rect -1185 460 -1145 480
rect -1185 440 -1175 460
rect -1155 440 -1145 460
rect -1185 420 -1145 440
rect -1185 400 -1175 420
rect -1155 400 -1145 420
rect -1185 390 -1145 400
rect -1035 500 -995 515
rect -1035 480 -1025 500
rect -1005 480 -995 500
rect -1035 460 -995 480
rect -1035 440 -1025 460
rect -1005 440 -995 460
rect -1035 420 -995 440
rect -1035 400 -1025 420
rect -1005 400 -995 420
rect -1035 390 -995 400
rect -885 500 -845 515
rect -885 480 -875 500
rect -855 480 -845 500
rect -885 460 -845 480
rect -885 440 -875 460
rect -855 440 -845 460
rect -885 420 -845 440
rect -885 400 -875 420
rect -855 400 -845 420
rect -885 390 -845 400
rect -795 500 -755 515
rect -795 480 -785 500
rect -765 480 -755 500
rect -795 460 -755 480
rect -795 440 -785 460
rect -765 440 -755 460
rect -795 420 -755 440
rect -795 400 -785 420
rect -765 400 -755 420
rect -795 390 -755 400
rect -720 500 -680 535
rect -720 480 -710 500
rect -690 480 -680 500
rect -720 460 -680 480
rect -720 440 -710 460
rect -690 440 -680 460
rect -720 420 -680 440
rect -720 400 -710 420
rect -690 400 -680 420
rect -720 390 -680 400
rect -645 500 -605 515
rect -645 480 -635 500
rect -615 480 -605 500
rect -645 460 -605 480
rect -645 440 -635 460
rect -615 440 -605 460
rect -645 420 -605 440
rect -645 400 -635 420
rect -615 400 -605 420
rect -645 390 -605 400
rect -570 500 -530 535
rect -395 515 -375 560
rect -95 515 -75 560
rect -570 480 -560 500
rect -540 480 -530 500
rect -570 460 -530 480
rect -570 440 -560 460
rect -540 440 -530 460
rect -570 420 -530 440
rect -570 400 -560 420
rect -540 400 -530 420
rect -570 390 -530 400
rect -495 500 -455 515
rect -495 480 -485 500
rect -465 480 -455 500
rect -495 460 -455 480
rect -495 440 -485 460
rect -465 440 -455 460
rect -495 420 -455 440
rect -495 400 -485 420
rect -465 400 -455 420
rect -495 390 -455 400
rect -405 500 -365 515
rect -405 480 -395 500
rect -375 480 -365 500
rect -405 460 -365 480
rect -405 440 -395 460
rect -375 440 -365 460
rect -405 420 -365 440
rect -405 400 -395 420
rect -375 400 -365 420
rect -405 390 -365 400
rect -255 500 -215 515
rect -255 480 -245 500
rect -225 480 -215 500
rect -255 460 -215 480
rect -255 440 -245 460
rect -225 440 -215 460
rect -255 420 -215 440
rect -255 400 -245 420
rect -225 400 -215 420
rect -255 390 -215 400
rect -105 500 -65 515
rect -105 480 -95 500
rect -75 480 -65 500
rect -105 460 -65 480
rect -105 440 -95 460
rect -75 440 -65 460
rect -105 420 -65 440
rect -105 400 -95 420
rect -75 400 -65 420
rect -105 390 -65 400
rect -745 360 -705 370
rect -545 360 -505 370
rect -1195 340 -735 360
rect -715 340 -535 360
rect -515 340 -505 360
rect -745 330 -705 340
rect -545 330 -505 340
rect -1195 300 -55 310
rect -1195 280 -1155 300
rect -1135 280 -1115 300
rect -1095 280 -1075 300
rect -1055 280 -1035 300
rect -1015 280 -995 300
rect -975 280 -955 300
rect -935 280 -915 300
rect -895 280 -875 300
rect -855 280 -835 300
rect -815 280 -795 300
rect -775 280 -755 300
rect -735 280 -715 300
rect -695 280 -675 300
rect -655 280 -635 300
rect -615 280 -595 300
rect -575 280 -555 300
rect -535 280 -515 300
rect -495 280 -475 300
rect -455 280 -435 300
rect -415 280 -395 300
rect -375 280 -355 300
rect -335 280 -315 300
rect -295 280 -275 300
rect -255 280 -235 300
rect -215 280 -195 300
rect -175 280 -155 300
rect -135 280 -115 300
rect -95 280 -55 300
rect -1195 270 -55 280
<< viali >>
rect -1155 870 -1135 890
rect -1115 870 -1095 890
rect -1075 870 -1055 890
rect -1035 870 -1015 890
rect -995 870 -975 890
rect -955 870 -935 890
rect -915 870 -895 890
rect -875 870 -855 890
rect -835 870 -815 890
rect -795 870 -775 890
rect -755 870 -735 890
rect -715 870 -695 890
rect -675 870 -655 890
rect -635 870 -615 890
rect -595 870 -575 890
rect -555 870 -535 890
rect -515 870 -495 890
rect -475 870 -455 890
rect -435 870 -415 890
rect -395 870 -375 890
rect -355 870 -335 890
rect -315 870 -295 890
rect -275 870 -255 890
rect -235 870 -215 890
rect -195 870 -175 890
rect -155 870 -135 890
rect -115 870 -95 890
rect -925 805 -905 825
rect -295 805 -275 825
rect -860 755 -840 775
rect -785 760 -765 780
rect -925 705 -905 725
rect -785 720 -765 740
rect -860 655 -840 675
rect -785 680 -765 700
rect -635 760 -615 780
rect -635 720 -615 740
rect -635 680 -615 700
rect -485 760 -465 780
rect -195 755 -175 775
rect -485 720 -465 740
rect -485 680 -465 700
rect -120 705 -100 725
rect -610 620 -590 640
rect -345 655 -325 675
rect -425 615 -405 635
rect -1025 480 -1005 500
rect -1025 440 -1005 460
rect -1025 400 -1005 420
rect -785 480 -765 500
rect -785 440 -765 460
rect -785 400 -765 420
rect -635 480 -615 500
rect -635 440 -615 460
rect -635 400 -615 420
rect -485 480 -465 500
rect -485 440 -465 460
rect -485 400 -465 420
rect -245 480 -225 500
rect -245 440 -225 460
rect -245 400 -225 420
rect -1155 280 -1135 300
rect -1115 280 -1095 300
rect -1075 280 -1055 300
rect -1035 280 -1015 300
rect -995 280 -975 300
rect -955 280 -935 300
rect -915 280 -895 300
rect -875 280 -855 300
rect -835 280 -815 300
rect -795 280 -775 300
rect -755 280 -735 300
rect -715 280 -695 300
rect -675 280 -655 300
rect -635 280 -615 300
rect -595 280 -575 300
rect -555 280 -535 300
rect -515 280 -495 300
rect -475 280 -455 300
rect -435 280 -415 300
rect -395 280 -375 300
rect -355 280 -335 300
rect -315 280 -295 300
rect -275 280 -255 300
rect -235 280 -215 300
rect -195 280 -175 300
rect -155 280 -135 300
rect -115 280 -95 300
<< metal1 >>
rect -1195 890 -55 905
rect -1195 870 -1155 890
rect -1135 870 -1115 890
rect -1095 870 -1075 890
rect -1055 870 -1035 890
rect -1015 870 -995 890
rect -975 870 -955 890
rect -935 870 -915 890
rect -895 870 -875 890
rect -855 870 -835 890
rect -815 870 -795 890
rect -775 870 -755 890
rect -735 870 -715 890
rect -695 870 -675 890
rect -655 870 -635 890
rect -615 870 -595 890
rect -575 870 -555 890
rect -535 870 -515 890
rect -495 870 -475 890
rect -455 870 -435 890
rect -415 870 -395 890
rect -375 870 -355 890
rect -335 870 -315 890
rect -295 870 -275 890
rect -255 870 -235 890
rect -215 870 -195 890
rect -175 870 -155 890
rect -135 870 -115 890
rect -95 870 -55 890
rect -1195 855 -55 870
rect -1025 515 -1005 855
rect -935 830 -895 835
rect -935 800 -930 830
rect -900 800 -895 830
rect -935 795 -895 800
rect -870 780 -830 785
rect -870 750 -865 780
rect -835 750 -830 780
rect -870 745 -830 750
rect -795 780 -755 855
rect -795 760 -785 780
rect -765 760 -755 780
rect -795 740 -755 760
rect -935 730 -895 735
rect -935 700 -930 730
rect -900 700 -895 730
rect -935 695 -895 700
rect -795 720 -785 740
rect -765 720 -755 740
rect -795 700 -755 720
rect -870 680 -830 685
rect -870 650 -865 680
rect -835 650 -830 680
rect -795 680 -785 700
rect -765 680 -755 700
rect -795 670 -755 680
rect -645 780 -605 855
rect -645 760 -635 780
rect -615 760 -605 780
rect -645 740 -605 760
rect -645 720 -635 740
rect -615 720 -605 740
rect -645 700 -605 720
rect -645 680 -635 700
rect -615 680 -605 700
rect -645 670 -605 680
rect -495 780 -455 855
rect -305 830 -265 835
rect -305 800 -300 830
rect -270 800 -265 830
rect -305 795 -265 800
rect -495 760 -485 780
rect -465 760 -455 780
rect -495 740 -455 760
rect -495 720 -485 740
rect -465 720 -455 740
rect -495 700 -455 720
rect -495 680 -485 700
rect -465 680 -455 700
rect -495 670 -455 680
rect -355 680 -315 685
rect -355 650 -350 680
rect -320 650 -315 680
rect -870 645 -830 650
rect -620 640 -580 650
rect -355 645 -315 650
rect -620 620 -610 640
rect -590 630 -580 640
rect -435 635 -395 645
rect -435 630 -425 635
rect -590 620 -425 630
rect -620 615 -425 620
rect -405 615 -395 635
rect -620 610 -395 615
rect -435 605 -395 610
rect -245 515 -225 855
rect -205 780 -165 785
rect -205 750 -200 780
rect -170 750 -165 780
rect -205 745 -165 750
rect -130 730 -90 735
rect -130 700 -125 730
rect -95 700 -90 730
rect -130 695 -90 700
rect -1035 500 -995 515
rect -1035 480 -1025 500
rect -1005 480 -995 500
rect -1035 460 -995 480
rect -1035 440 -1025 460
rect -1005 440 -995 460
rect -1035 420 -995 440
rect -1035 400 -1025 420
rect -1005 400 -995 420
rect -1035 390 -995 400
rect -795 500 -755 515
rect -795 480 -785 500
rect -765 480 -755 500
rect -795 460 -755 480
rect -795 440 -785 460
rect -765 440 -755 460
rect -795 420 -755 440
rect -795 400 -785 420
rect -765 400 -755 420
rect -795 390 -755 400
rect -645 500 -605 515
rect -645 480 -635 500
rect -615 480 -605 500
rect -645 460 -605 480
rect -645 440 -635 460
rect -615 440 -605 460
rect -645 420 -605 440
rect -645 400 -635 420
rect -615 400 -605 420
rect -645 390 -605 400
rect -495 500 -455 515
rect -495 480 -485 500
rect -465 480 -455 500
rect -495 460 -455 480
rect -495 440 -485 460
rect -465 440 -455 460
rect -495 420 -455 440
rect -495 400 -485 420
rect -465 400 -455 420
rect -495 390 -455 400
rect -255 500 -215 515
rect -255 480 -245 500
rect -225 480 -215 500
rect -255 460 -215 480
rect -255 440 -245 460
rect -225 440 -215 460
rect -255 420 -215 440
rect -255 400 -245 420
rect -225 400 -215 420
rect -255 390 -215 400
rect -785 315 -765 390
rect -635 315 -615 390
rect -485 315 -465 390
rect -1195 300 -55 315
rect -1195 280 -1155 300
rect -1135 280 -1115 300
rect -1095 280 -1075 300
rect -1055 280 -1035 300
rect -1015 280 -995 300
rect -975 280 -955 300
rect -935 280 -915 300
rect -895 280 -875 300
rect -855 280 -835 300
rect -815 280 -795 300
rect -775 280 -755 300
rect -735 280 -715 300
rect -695 280 -675 300
rect -655 280 -635 300
rect -615 280 -595 300
rect -575 280 -555 300
rect -535 280 -515 300
rect -495 280 -475 300
rect -455 280 -435 300
rect -415 280 -395 300
rect -375 280 -355 300
rect -335 280 -315 300
rect -295 280 -275 300
rect -255 280 -235 300
rect -215 280 -195 300
rect -175 280 -155 300
rect -135 280 -115 300
rect -95 280 -55 300
rect -1195 265 -55 280
<< via1 >>
rect -930 825 -900 830
rect -930 805 -925 825
rect -925 805 -905 825
rect -905 805 -900 825
rect -930 800 -900 805
rect -865 775 -835 780
rect -865 755 -860 775
rect -860 755 -840 775
rect -840 755 -835 775
rect -865 750 -835 755
rect -930 725 -900 730
rect -930 705 -925 725
rect -925 705 -905 725
rect -905 705 -900 725
rect -930 700 -900 705
rect -865 675 -835 680
rect -865 655 -860 675
rect -860 655 -840 675
rect -840 655 -835 675
rect -865 650 -835 655
rect -300 825 -270 830
rect -300 805 -295 825
rect -295 805 -275 825
rect -275 805 -270 825
rect -300 800 -270 805
rect -350 675 -320 680
rect -350 655 -345 675
rect -345 655 -325 675
rect -325 655 -320 675
rect -350 650 -320 655
rect -200 775 -170 780
rect -200 755 -195 775
rect -195 755 -175 775
rect -175 755 -170 775
rect -200 750 -170 755
rect -125 725 -95 730
rect -125 705 -120 725
rect -120 705 -100 725
rect -100 705 -95 725
rect -125 700 -95 705
<< metal2 >>
rect -935 830 -895 835
rect -935 800 -930 830
rect -900 825 -895 830
rect -305 830 -265 835
rect -305 825 -300 830
rect -900 805 -300 825
rect -900 800 -895 805
rect -935 795 -895 800
rect -305 800 -300 805
rect -270 800 -265 830
rect -305 795 -265 800
rect -870 780 -830 785
rect -870 750 -865 780
rect -835 775 -830 780
rect -205 780 -165 785
rect -205 775 -200 780
rect -835 755 -200 775
rect -835 750 -830 755
rect -870 745 -830 750
rect -205 750 -200 755
rect -170 750 -165 780
rect -205 745 -165 750
rect -935 730 -895 735
rect -935 700 -930 730
rect -900 725 -895 730
rect -130 730 -90 735
rect -130 725 -125 730
rect -900 705 -125 725
rect -900 700 -895 705
rect -935 695 -895 700
rect -130 700 -125 705
rect -95 700 -90 730
rect -130 695 -90 700
rect -870 680 -830 685
rect -870 650 -865 680
rect -835 675 -830 680
rect -355 680 -315 685
rect -355 675 -350 680
rect -835 655 -350 675
rect -835 650 -830 655
rect -870 645 -830 650
rect -355 650 -350 655
rect -320 650 -315 680
rect -355 645 -315 650
<< labels >>
rlabel metal1 -635 870 -615 890 7 CLK
port 9 w
rlabel locali -1190 660 -1180 670 7 B_bar
port 4 w
rlabel locali -1190 810 -1180 820 7 A
port 1 w
rlabel locali -1190 710 -1180 720 7 B
port 3 w
rlabel locali -1190 760 -1180 770 7 A_bar
port 2 w
rlabel viali -610 620 -590 640 7 OUT_bar
port 6 w
rlabel metal1 -635 280 -615 300 7 GND!
port 8 w
rlabel locali -735 340 -715 360 7 Dis
port 7 w
rlabel locali -660 560 -640 580 7 OUT
port 5 w
<< end >>
