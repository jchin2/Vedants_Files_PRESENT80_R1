* NGSPICE file created from EESPFAL_s1_flat.ext - technology: sky130A

.subckt EESPFAL_s1_flat GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar s1_bar s1 Dis1
+ Dis3 Dis2 CLK1 CLK2 CLK3
X0 a_n2159_n2753# x0_bar.t0 EESPFAL_INV4_0/A GND.t20 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X1 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar CLK2.t11 CLK2.t10 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X2 CLK1.t10 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar CLK1.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 EESPFAL_INV4_0/A EESPFAL_INV4_0/A_bar GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 GND.t59 EESPFAL_NAND_v3_0/A_bar.t6 EESPFAL_NAND_v3_0/A.t2 GND.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 GND.t40 EESPFAL_INV4_0/A EESPFAL_INV4_0/A_bar GND.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X6 EESPFAL_NAND_v3_1/B Dis1.t0 GND.t31 GND.t30 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_2081_n2754# EESPFAL_NAND_v3_1/OUT_bar a_1931_n2754# GND.t37 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X8 GND.t57 Dis2.t0 EESPFAL_NAND_v3_0/OUT GND.t56 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X9 a_n2160_67# x0_bar.t1 EESPFAL_NAND_v3_0/A_bar.t1 GND.t19 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X10 GND.t58 Dis2.t1 EESPFAL_NAND_v3_1/OUT GND.t56 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X11 CLK1.t50 EESPFAL_NAND_v3_1/A_bar.t6 EESPFAL_NAND_v3_1/A.t2 CLK1.t49 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK3.t4 EESPFAL_NAND_v3_0/OUT_bar.t6 a_2081_n2754# GND.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 EESPFAL_NAND_v3_1/A_bar.t3 x3.t0 a_n3420_n613# GND.t60 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X14 a_n3420_n613# x1.t0 CLK1.t23 GND.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_n1860_n613# x1_bar.t0 CLK1.t29 GND.t1 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X16 EESPFAL_NAND_v3_1/A.t0 EESPFAL_NAND_v3_1/A_bar.t7 GND.t83 GND.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 CLK2.t12 EESPFAL_INV4_0/A EESPFAL_3in_NOR_v2_0/C.t1 GND.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 GND.t51 Dis2.t2 EESPFAL_3in_NOR_v2_0/C.t0 GND.t50 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 GND.t55 EESPFAL_NAND_v3_1/A.t6 EESPFAL_NAND_v3_1/A_bar.t2 GND.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X20 GND.t14 Dis3.t0 s1_bar.t2 GND.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X21 s1.t2 s1_bar.t5 CLK3.t6 CLK3.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X22 EESPFAL_INV4_0/A_bar EESPFAL_INV4_0/A CLK1.t27 CLK1.t26 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X23 GND.t74 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X24 EESPFAL_3in_NOR_v2_0/C.t4 EESPFAL_3in_NOR_v2_0/C_bar.t5 GND.t63 GND.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X25 CLK2.t6 EESPFAL_NAND_v3_1/B_bar EESPFAL_NAND_v3_1/OUT_bar GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X26 EESPFAL_NAND_v3_0/OUT_bar.t0 Dis2.t3 GND.t53 GND.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X27 CLK1.t36 EESPFAL_NAND_v3_0/A.t6 EESPFAL_NAND_v3_0/A_bar.t2 CLK1.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X28 EESPFAL_NAND_v3_1/B x2_bar.t0 CLK1.t0 GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X29 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_1/OUT CLK2.t16 CLK2.t15 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X30 CLK1.t5 x2.t0 EESPFAL_NAND_v3_1/B_bar GND.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X31 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar CLK1.t45 CLK1.t44 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X32 a_n2009_n2753# x1.t1 a_n2159_n2753# GND.t34 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X33 a_n3420_67# x2.t1 CLK1.t6 GND.t8 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X34 CLK2.t30 EESPFAL_3in_NOR_v2_0/C.t5 EESPFAL_3in_NOR_v2_0/C_bar.t4 CLK2.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X35 CLK1.t32 EESPFAL_NAND_v3_0/A_bar.t7 EESPFAL_NAND_v3_0/A.t4 CLK1.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X36 GND.t33 Dis1.t1 EESPFAL_INV4_0/A GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X37 EESPFAL_3in_NOR_v2_0/C_bar.t3 EESPFAL_3in_NOR_v2_0/C.t6 CLK2.t26 CLK2.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X38 EESPFAL_INV4_0/A_bar x0.t0 CLK1.t48 GND.t82 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X39 CLK1.t12 x3_bar.t0 a_n2009_n2753# GND.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X40 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/B CLK1.t40 CLK1.t39 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X41 EESPFAL_NAND_v3_0/OUT_bar.t3 EESPFAL_NAND_v3_0/OUT CLK2.t24 CLK2.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X42 CLK1.t30 x1_bar.t1 a_n3720_n613# GND.t41 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X43 a_n3720_n613# x3_bar.t1 EESPFAL_NAND_v3_1/A_bar.t1 GND.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X44 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar CLK1.t20 CLK1.t19 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X45 EESPFAL_NAND_v3_1/A_bar.t4 Dis1.t2 GND.t64 GND.t45 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X46 GND.t87 s1_bar.t6 s1.t3 GND.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X47 EESPFAL_INV4_0/A EESPFAL_INV4_0/A_bar CLK1.t16 CLK1.t15 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X48 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar.t7 GND.t72 GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X49 CLK1.t4 x2.t2 a_n2160_67# GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X50 EESPFAL_NAND_v3_0/A_bar.t3 EESPFAL_NAND_v3_0/A.t7 GND.t70 GND.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X51 a_1910_n613# EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/OUT GND.t11 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X52 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_1/A_bar.t8 CLK2.t7 GND.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X53 s1_bar.t3 s1.t7 GND.t29 GND.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X54 CLK1.t25 EESPFAL_INV4_0/A EESPFAL_INV4_0/A_bar CLK1.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X55 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar.t8 CLK2.t1 CLK2.t0 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X56 a_1931_n2754# EESPFAL_3in_NOR_v2_0/C_bar.t6 s1_bar.t4 GND.t49 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X57 CLK1.t28 x1.t2 a_n2160_n613# GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X58 EESPFAL_NAND_v3_1/A_bar.t0 EESPFAL_NAND_v3_1/A.t7 CLK1.t3 CLK1.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X59 GND.t66 Dis1.t3 EESPFAL_NAND_v3_1/B_bar GND.t65 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X60 a_n3720_67# x0_bar.t2 EESPFAL_NAND_v3_0/A.t0 GND.t18 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X61 EESPFAL_NAND_v3_1/OUT_bar Dis2.t4 GND.t79 GND.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X62 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar GND.t75 GND.t9 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X63 CLK2.t20 EESPFAL_3in_NOR_v2_0/C_bar.t7 EESPFAL_3in_NOR_v2_0/C.t3 CLK2.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X64 EESPFAL_NAND_v3_0/OUT_bar.t5 EESPFAL_NAND_v3_0/A_bar.t8 CLK2.t31 GND.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X65 s1.t5 EESPFAL_3in_NOR_v2_0/C.t7 CLK3.t9 GND.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X66 CLK3.t1 s1.t8 s1_bar.t0 CLK3.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X67 a_n1860_67# x2_bar.t1 CLK1.t1 GND.t1 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X68 EESPFAL_3in_NOR_v2_0/C.t2 EESPFAL_3in_NOR_v2_0/C_bar.t8 CLK2.t18 CLK2.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X69 EESPFAL_INV4_0/A_bar x3.t1 CLK1.t33 GND.t61 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X70 EESPFAL_NAND_v3_0/A_bar.t4 EESPFAL_NAND_v3_0/A.t8 CLK1.t47 CLK1.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X71 CLK1.t11 x1_bar.t2 EESPFAL_INV4_0/A_bar GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X72 EESPFAL_NAND_v3_0/A.t1 Dis1.t4 GND.t46 GND.t45 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X73 CLK2.t9 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_1/OUT CLK2.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X74 EESPFAL_NAND_v3_1/B_bar EESPFAL_NAND_v3_1/B CLK1.t8 CLK1.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X75 CLK2.t28 EESPFAL_NAND_v3_0/A.t9 a_1910_67# GND.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X76 EESPFAL_NAND_v3_0/A.t5 x0.t1 a_n3420_67# GND.t60 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X77 CLK1.t18 EESPFAL_NAND_v3_1/B_bar EESPFAL_NAND_v3_1/B CLK1.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X78 EESPFAL_NAND_v3_0/A.t3 EESPFAL_NAND_v3_0/A_bar.t9 CLK1.t55 CLK1.t54 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X79 s1.t0 Dis3.t1 GND.t16 GND.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X80 EESPFAL_INV4_0/A_bar Dis1.t5 GND.t48 GND.t47 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X81 CLK1.t14 EESPFAL_INV4_0/A_bar EESPFAL_INV4_0/A CLK1.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X82 a_n2160_n613# x3_bar.t2 EESPFAL_NAND_v3_1/A.t4 GND.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X83 EESPFAL_NAND_v3_1/A.t1 EESPFAL_NAND_v3_1/A_bar.t9 CLK1.t22 CLK1.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X84 EESPFAL_NAND_v3_1/B_bar EESPFAL_NAND_v3_1/B GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X85 GND.t25 EESPFAL_NAND_v3_1/B_bar EESPFAL_NAND_v3_1/B GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X86 EESPFAL_NAND_v3_0/B_bar Dis1.t6 GND.t84 GND.t30 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X87 CLK2.t4 EESPFAL_NAND_v3_1/A.t8 a_1910_n613# GND.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X88 GND.t85 Dis1.t7 EESPFAL_NAND_v3_0/A_bar.t5 GND.t76 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X89 CLK2.t22 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar.t2 CLK2.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X90 GND.t44 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar GND.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X91 CLK1.t53 EESPFAL_NAND_v3_1/A.t9 EESPFAL_NAND_v3_1/A_bar.t5 CLK1.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X92 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar GND.t36 GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X93 a_1910_67# EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/OUT GND.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X94 GND.t68 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar.t1 GND.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X95 CLK1.t34 x3.t2 EESPFAL_NAND_v3_0/B GND.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X96 CLK1.t43 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/B CLK1.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X97 s1.t6 EESPFAL_NAND_v3_0/OUT CLK3.t8 GND.t67 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X98 CLK3.t11 s1_bar.t7 s1.t1 CLK3.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X99 GND.t4 EESPFAL_3in_NOR_v2_0/C.t8 EESPFAL_3in_NOR_v2_0/C_bar.t2 GND.t3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X100 GND.t77 Dis1.t8 EESPFAL_NAND_v3_1/A.t5 GND.t76 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X101 EESPFAL_3in_NOR_v2_0/C_bar.t1 EESPFAL_INV4_0/A_bar CLK2.t5 GND.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X102 EESPFAL_NAND_v3_1/A.t3 x3.t3 a_n1860_n613# GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X103 CLK3.t7 EESPFAL_NAND_v3_1/OUT s1.t4 GND.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X104 s1_bar.t1 s1.t9 CLK3.t3 CLK3.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X105 EESPFAL_3in_NOR_v2_0/C_bar.t0 Dis2.t5 GND.t81 GND.t80 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X106 CLK2.t3 EESPFAL_NAND_v3_0/OUT_bar.t9 EESPFAL_NAND_v3_0/OUT CLK2.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X107 GND.t78 Dis1.t9 EESPFAL_NAND_v3_0/B GND.t65 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X108 CLK1.t51 x2_bar.t2 a_n3720_67# GND.t41 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X109 CLK2.t27 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/OUT_bar.t4 GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X110 CLK2.t14 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar CLK2.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X111 EESPFAL_NAND_v3_0/B_bar x3_bar.t3 CLK1.t41 GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X112 EESPFAL_NAND_v3_0/A_bar.t0 x0.t2 a_n1860_67# GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X113 CLK1.t38 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar CLK1.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
R0 EESPFAL_3in_NAND_v2_0/C x0_bar.t0 904.039
R1 x0_bar.n0 x0_bar.t1 810.772
R2 x0_bar.n0 x0_bar.t2 694.566
R3 EESPFAL_3in_NAND_v2_0/C x0_bar.n1 325.825
R4 x0_bar.n1 x0_bar 278.57
R5 x0_bar x0_bar.n0 25.6
R6 x0_bar.n1 x0_bar 0.321
R7 GND.n405 GND.n404 341.085
R8 GND.n413 GND.n245 341.085
R9 GND.n415 GND.n414 341.085
R10 GND.n424 GND.n239 341.085
R11 GND.n425 GND.n424 341.085
R12 GND.n426 GND.n425 341.085
R13 GND.n437 GND.n233 341.085
R14 GND.n440 GND.n439 341.085
R15 GND.n450 GND.n449 341.085
R16 GND.n452 GND.n450 341.085
R17 GND.n452 GND.n451 341.085
R18 GND.n461 GND.n460 341.085
R19 GND.n463 GND.n462 341.085
R20 GND.n472 GND.n471 341.085
R21 GND.n311 GND.n310 341.085
R22 GND.n312 GND.n297 341.085
R23 GND.n321 GND.n297 341.085
R24 GND.n322 GND.n321 341.085
R25 GND.n324 GND.n323 341.085
R26 GND.n334 GND.n333 341.085
R27 GND.n343 GND.n284 341.085
R28 GND.n344 GND.n343 341.085
R29 GND.n345 GND.n344 341.085
R30 GND.n353 GND.n278 341.085
R31 GND.n365 GND.n364 341.085
R32 GND.n367 GND.n365 341.085
R33 GND.n367 GND.n366 341.085
R34 GND.n377 GND.n376 341.085
R35 GND.n387 GND.n260 341.085
R36 GND.n389 GND.n388 341.085
R37 GND.n389 GND.n254 341.085
R38 GND.n397 GND.n254 341.085
R39 GND.t19 GND.n239 319.767
R40 GND.n438 GND.t69 319.767
R41 GND.t54 GND.n438 319.767
R42 GND.n451 GND.t60 319.767
R43 GND.n312 GND.t11 319.767
R44 GND.n332 GND.t35 319.767
R45 GND.t43 GND.n332 319.767
R46 GND.n345 GND.t27 319.767
R47 GND.n364 GND.t7 319.767
R48 GND.n378 GND.t9 319.767
R49 GND.n378 GND.t24 319.767
R50 GND.t0 GND.n397 319.767
R51 GND.n414 GND.t6 277.131
R52 GND.t76 GND.n233 277.131
R53 GND.n439 GND.t45 277.131
R54 GND.t8 GND.n461 277.131
R55 GND.n310 GND.t5 277.131
R56 GND.n324 GND.t56 277.131
R57 GND.n334 GND.t52 277.131
R58 GND.t26 GND.n353 277.131
R59 GND.n376 GND.t65 277.131
R60 GND.t30 GND.n387 277.131
R61 GND.t1 GND.n245 234.496
R62 GND.n462 GND.t41 234.496
R63 GND.n95 GND.t67 192.984
R64 GND.n167 GND.t17 192.984
R65 GND.n7 GND.t71 192.984
R66 GND.n476 GND.t82 192.984
R67 GND.n404 GND.t2 191.86
R68 GND.t18 GND.n472 191.86
R69 GND.t2 GND.n403 158.378
R70 GND.n473 GND.t18 158.378
R71 GND.n403 GND.n250 157.6
R72 GND.n406 GND.n250 157.6
R73 GND.n406 GND.n246 157.6
R74 GND.n412 GND.n246 157.6
R75 GND.n412 GND.n244 157.6
R76 GND.n416 GND.n244 157.6
R77 GND.n416 GND.n240 157.6
R78 GND.n423 GND.n240 157.6
R79 GND.n423 GND.n238 157.6
R80 GND.n427 GND.n238 157.6
R81 GND.n427 GND.n234 157.6
R82 GND.n436 GND.n234 157.6
R83 GND.n436 GND.n232 157.6
R84 GND.n441 GND.n232 157.6
R85 GND.n441 GND.n229 157.6
R86 GND.n448 GND.n229 157.6
R87 GND.n448 GND.n228 157.6
R88 GND.n453 GND.n228 157.6
R89 GND.n453 GND.n224 157.6
R90 GND.n459 GND.n224 157.6
R91 GND.n459 GND.n223 157.6
R92 GND.n464 GND.n223 157.6
R93 GND.n464 GND.n218 157.6
R94 GND.n470 GND.n218 157.6
R95 GND.n470 GND.n217 157.6
R96 GND.n473 GND.n217 157.6
R97 GND.n309 GND.n303 157.6
R98 GND.n309 GND.n302 157.6
R99 GND.n313 GND.n302 157.6
R100 GND.n313 GND.n298 157.6
R101 GND.n320 GND.n298 157.6
R102 GND.n320 GND.n296 157.6
R103 GND.n325 GND.n296 157.6
R104 GND.n325 GND.n290 157.6
R105 GND.n331 GND.n290 157.6
R106 GND.n331 GND.n289 157.6
R107 GND.n335 GND.n289 157.6
R108 GND.n335 GND.n285 157.6
R109 GND.n342 GND.n285 157.6
R110 GND.n342 GND.n283 157.6
R111 GND.n346 GND.n283 157.6
R112 GND.n346 GND.n279 157.6
R113 GND.n352 GND.n279 157.6
R114 GND.n352 GND.n277 157.6
R115 GND.n363 GND.n273 157.6
R116 GND.n363 GND.n272 157.6
R117 GND.n368 GND.n272 157.6
R118 GND.n368 GND.n268 157.6
R119 GND.n375 GND.n268 157.6
R120 GND.n375 GND.n267 157.6
R121 GND.n379 GND.n267 157.6
R122 GND.n379 GND.n261 157.6
R123 GND.n386 GND.n261 157.6
R124 GND.n386 GND.n259 157.6
R125 GND.n390 GND.n259 157.6
R126 GND.n390 GND.n255 157.6
R127 GND.n396 GND.n255 157.6
R128 GND.n396 GND.n253 157.6
R129 GND.n306 GND.n305 118.661
R130 GND.n355 GND.n354 115.922
R131 GND.n358 GND.n357 115.922
R132 GND.n399 GND.n398 115.922
R133 GND.n120 GND.t50 111.486
R134 GND.n142 GND.t80 111.486
R135 GND.n15 GND.t37 111.486
R136 GND.n40 GND.t13 111.486
R137 GND.n62 GND.t15 111.486
R138 GND.n87 GND.t42 111.486
R139 GND.n175 GND.t34 111.486
R140 GND.n200 GND.t32 111.486
R141 GND.n509 GND.t47 111.486
R142 GND.n484 GND.t12 111.486
R143 GND.n405 GND.t1 106.589
R144 GND.n471 GND.t41 106.589
R145 GND.n305 GND.t5 70.155
R146 GND.n354 GND.t26 70.155
R147 GND.t6 GND.n413 63.953
R148 GND.n426 GND.t76 63.953
R149 GND.n449 GND.t45 63.953
R150 GND.n463 GND.t8 63.953
R151 GND.t56 GND.n322 63.953
R152 GND.t52 GND.n284 63.953
R153 GND.n366 GND.t65 63.953
R154 GND.n388 GND.t30 63.953
R155 GND.n475 GND 48.86
R156 GND.n159 GND.t21 44.336
R157 GND.n103 GND.t38 44.336
R158 GND.n128 GND.t62 37.162
R159 GND.n134 GND.t3 37.162
R160 GND.n23 GND.t49 37.162
R161 GND.n48 GND.t28 37.162
R162 GND.n54 GND.t86 37.162
R163 GND.n79 GND.t73 37.162
R164 GND.n183 GND.t20 37.162
R165 GND.n208 GND.t22 37.162
R166 GND.n517 GND.t39 37.162
R167 GND.n492 GND.t61 37.162
R168 GND GND.n474 31.565
R169 GND.n317 GND.t57 29.103
R170 GND.n339 GND.t53 29.103
R171 GND.n371 GND.t78 29.103
R172 GND.n257 GND.t84 29.103
R173 GND.n236 GND.t85 29.103
R174 GND.n445 GND.t46 29.103
R175 GND.n39 GND.t14 29.103
R176 GND.n66 GND.t16 29.103
R177 GND.n119 GND.t51 29.103
R178 GND.n146 GND.t81 29.103
R179 GND.n199 GND.t33 29.103
R180 GND.n508 GND.t48 29.103
R181 GND.n317 GND.t58 29.102
R182 GND.n339 GND.t79 29.102
R183 GND.n371 GND.t66 29.102
R184 GND.n257 GND.t31 29.102
R185 GND.n236 GND.t77 29.102
R186 GND.n445 GND.t64 29.102
R187 GND.n357 GND.t7 27.519
R188 GND.n398 GND.t0 27.519
R189 GND.n432 GND.t83 24
R190 GND.n432 GND.t55 24
R191 GND.n431 GND.t70 24
R192 GND.n431 GND.t59 24
R193 GND.n293 GND.t36 24
R194 GND.n293 GND.t44 24
R195 GND.n292 GND.t72 24
R196 GND.n292 GND.t68 24
R197 GND.n264 GND.t10 24
R198 GND.n264 GND.t25 24
R199 GND.n263 GND.t75 24
R200 GND.n263 GND.t74 24
R201 GND.n0 GND.t23 24
R202 GND.n0 GND.t40 24
R203 GND.n3 GND.t63 24
R204 GND.n3 GND.t4 24
R205 GND.n6 GND.t29 24
R206 GND.n6 GND.t87 24
R207 GND.n415 GND.t19 21.317
R208 GND.t69 GND.n437 21.317
R209 GND.n440 GND.t54 21.317
R210 GND.n460 GND.t60 21.317
R211 GND.t11 GND.n311 21.317
R212 GND.n323 GND.t35 21.317
R213 GND.n333 GND.t43 21.317
R214 GND.t27 GND.n278 21.317
R215 GND.t9 GND.n377 21.317
R216 GND.t24 GND.n260 21.317
R217 GND.n308 GND.n304 12.8
R218 GND.n308 GND.n301 12.8
R219 GND.n314 GND.n301 12.8
R220 GND.n314 GND.n299 12.8
R221 GND.n319 GND.n299 12.8
R222 GND.n319 GND.n295 12.8
R223 GND.n326 GND.n295 12.8
R224 GND.n326 GND.n291 12.8
R225 GND.n330 GND.n291 12.8
R226 GND.n330 GND.n288 12.8
R227 GND.n336 GND.n288 12.8
R228 GND.n336 GND.n286 12.8
R229 GND.n341 GND.n286 12.8
R230 GND.n341 GND.n282 12.8
R231 GND.n347 GND.n282 12.8
R232 GND.n347 GND.n280 12.8
R233 GND.n351 GND.n280 12.8
R234 GND.n351 GND.n276 12.8
R235 GND.n355 GND.n276 12.8
R236 GND.n358 GND.n274 12.8
R237 GND.n362 GND.n274 12.8
R238 GND.n362 GND.n271 12.8
R239 GND.n369 GND.n271 12.8
R240 GND.n369 GND.n269 12.8
R241 GND.n374 GND.n269 12.8
R242 GND.n374 GND.n266 12.8
R243 GND.n380 GND.n266 12.8
R244 GND.n380 GND.n262 12.8
R245 GND.n385 GND.n262 12.8
R246 GND.n385 GND.n258 12.8
R247 GND.n391 GND.n258 12.8
R248 GND.n391 GND.n256 12.8
R249 GND.n395 GND.n256 12.8
R250 GND.n395 GND.n252 12.8
R251 GND.n399 GND.n252 12.8
R252 GND.n402 GND.n249 12.8
R253 GND.n407 GND.n249 12.8
R254 GND.n407 GND.n247 12.8
R255 GND.n411 GND.n247 12.8
R256 GND.n411 GND.n243 12.8
R257 GND.n417 GND.n243 12.8
R258 GND.n417 GND.n241 12.8
R259 GND.n422 GND.n241 12.8
R260 GND.n422 GND.n237 12.8
R261 GND.n428 GND.n237 12.8
R262 GND.n428 GND.n235 12.8
R263 GND.n435 GND.n235 12.8
R264 GND.n435 GND.n231 12.8
R265 GND.n442 GND.n231 12.8
R266 GND.n442 GND.n230 12.8
R267 GND.n447 GND.n230 12.8
R268 GND.n447 GND.n227 12.8
R269 GND.n454 GND.n227 12.8
R270 GND.n454 GND.n225 12.8
R271 GND.n458 GND.n225 12.8
R272 GND.n458 GND.n222 12.8
R273 GND.n465 GND.n222 12.8
R274 GND.n465 GND.n219 12.8
R275 GND.n469 GND.n219 12.8
R276 GND.n469 GND.n220 12.8
R277 GND.n136 GND.n133 12.8
R278 GND.n56 GND.n53 12.8
R279 GND.n304 GND.n303 9.154
R280 GND.n274 GND.n273 9.154
R281 GND.n363 GND.n362 9.154
R282 GND.n364 GND.n363 9.154
R283 GND.n272 GND.n271 9.154
R284 GND.n365 GND.n272 9.154
R285 GND.n369 GND.n368 9.154
R286 GND.n368 GND.n367 9.154
R287 GND.n269 GND.n268 9.154
R288 GND.n366 GND.n268 9.154
R289 GND.n375 GND.n374 9.154
R290 GND.n376 GND.n375 9.154
R291 GND.n267 GND.n266 9.154
R292 GND.n377 GND.n267 9.154
R293 GND.n380 GND.n379 9.154
R294 GND.n379 GND.n378 9.154
R295 GND.n262 GND.n261 9.154
R296 GND.n261 GND.n260 9.154
R297 GND.n386 GND.n385 9.154
R298 GND.n387 GND.n386 9.154
R299 GND.n259 GND.n258 9.154
R300 GND.n388 GND.n259 9.154
R301 GND.n391 GND.n390 9.154
R302 GND.n390 GND.n389 9.154
R303 GND.n256 GND.n255 9.154
R304 GND.n255 GND.n254 9.154
R305 GND.n396 GND.n395 9.154
R306 GND.n397 GND.n396 9.154
R307 GND.n253 GND.n252 9.154
R308 GND.n309 GND.n308 9.154
R309 GND.n310 GND.n309 9.154
R310 GND.n302 GND.n301 9.154
R311 GND.n311 GND.n302 9.154
R312 GND.n314 GND.n313 9.154
R313 GND.n313 GND.n312 9.154
R314 GND.n299 GND.n298 9.154
R315 GND.n298 GND.n297 9.154
R316 GND.n320 GND.n319 9.154
R317 GND.n321 GND.n320 9.154
R318 GND.n296 GND.n295 9.154
R319 GND.n322 GND.n296 9.154
R320 GND.n326 GND.n325 9.154
R321 GND.n325 GND.n324 9.154
R322 GND.n291 GND.n290 9.154
R323 GND.n323 GND.n290 9.154
R324 GND.n331 GND.n330 9.154
R325 GND.n332 GND.n331 9.154
R326 GND.n289 GND.n288 9.154
R327 GND.n333 GND.n289 9.154
R328 GND.n336 GND.n335 9.154
R329 GND.n335 GND.n334 9.154
R330 GND.n286 GND.n285 9.154
R331 GND.n285 GND.n284 9.154
R332 GND.n342 GND.n341 9.154
R333 GND.n343 GND.n342 9.154
R334 GND.n283 GND.n282 9.154
R335 GND.n344 GND.n283 9.154
R336 GND.n347 GND.n346 9.154
R337 GND.n346 GND.n345 9.154
R338 GND.n280 GND.n279 9.154
R339 GND.n279 GND.n278 9.154
R340 GND.n352 GND.n351 9.154
R341 GND.n353 GND.n352 9.154
R342 GND.n277 GND.n276 9.154
R343 GND.n250 GND.n249 9.154
R344 GND.n404 GND.n250 9.154
R345 GND.n407 GND.n406 9.154
R346 GND.n406 GND.n405 9.154
R347 GND.n247 GND.n246 9.154
R348 GND.n246 GND.n245 9.154
R349 GND.n412 GND.n411 9.154
R350 GND.n413 GND.n412 9.154
R351 GND.n244 GND.n243 9.154
R352 GND.n414 GND.n244 9.154
R353 GND.n417 GND.n416 9.154
R354 GND.n416 GND.n415 9.154
R355 GND.n241 GND.n240 9.154
R356 GND.n240 GND.n239 9.154
R357 GND.n423 GND.n422 9.154
R358 GND.n424 GND.n423 9.154
R359 GND.n238 GND.n237 9.154
R360 GND.n425 GND.n238 9.154
R361 GND.n428 GND.n427 9.154
R362 GND.n427 GND.n426 9.154
R363 GND.n235 GND.n234 9.154
R364 GND.n234 GND.n233 9.154
R365 GND.n436 GND.n435 9.154
R366 GND.n437 GND.n436 9.154
R367 GND.n232 GND.n231 9.154
R368 GND.n438 GND.n232 9.154
R369 GND.n442 GND.n441 9.154
R370 GND.n441 GND.n440 9.154
R371 GND.n230 GND.n229 9.154
R372 GND.n439 GND.n229 9.154
R373 GND.n448 GND.n447 9.154
R374 GND.n449 GND.n448 9.154
R375 GND.n228 GND.n227 9.154
R376 GND.n450 GND.n228 9.154
R377 GND.n454 GND.n453 9.154
R378 GND.n453 GND.n452 9.154
R379 GND.n225 GND.n224 9.154
R380 GND.n451 GND.n224 9.154
R381 GND.n459 GND.n458 9.154
R382 GND.n460 GND.n459 9.154
R383 GND.n223 GND.n222 9.154
R384 GND.n461 GND.n223 9.154
R385 GND.n465 GND.n464 9.154
R386 GND.n464 GND.n463 9.154
R387 GND.n219 GND.n218 9.154
R388 GND.n462 GND.n218 9.154
R389 GND.n470 GND.n469 9.154
R390 GND.n471 GND.n470 9.154
R391 GND.n220 GND.n217 9.154
R392 GND.n472 GND.n217 9.154
R393 GND.n474 GND.n473 9.154
R394 GND.n403 GND.n402 9.154
R395 GND.n9 GND.n8 9.154
R396 GND.n13 GND.n12 9.154
R397 GND.n12 GND.n11 9.154
R398 GND.n17 GND.n16 9.154
R399 GND.n16 GND.n15 9.154
R400 GND.n21 GND.n20 9.154
R401 GND.n20 GND.n19 9.154
R402 GND.n25 GND.n24 9.154
R403 GND.n24 GND.n23 9.154
R404 GND.n29 GND.n28 9.154
R405 GND.n28 GND.n27 9.154
R406 GND.n33 GND.n32 9.154
R407 GND.n32 GND.n31 9.154
R408 GND.n37 GND.n36 9.154
R409 GND.n36 GND.n35 9.154
R410 GND.n42 GND.n41 9.154
R411 GND.n41 GND.n40 9.154
R412 GND.n46 GND.n45 9.154
R413 GND.n45 GND.n44 9.154
R414 GND.n50 GND.n49 9.154
R415 GND.n49 GND.n48 9.154
R416 GND.n53 GND.n5 9.154
R417 GND.n5 GND.n4 9.154
R418 GND.n56 GND.n55 9.154
R419 GND.n55 GND.n54 9.154
R420 GND.n60 GND.n59 9.154
R421 GND.n59 GND.n58 9.154
R422 GND.n64 GND.n63 9.154
R423 GND.n63 GND.n62 9.154
R424 GND.n69 GND.n68 9.154
R425 GND.n68 GND.n67 9.154
R426 GND.n73 GND.n72 9.154
R427 GND.n72 GND.n71 9.154
R428 GND.n77 GND.n76 9.154
R429 GND.n76 GND.n75 9.154
R430 GND.n81 GND.n80 9.154
R431 GND.n80 GND.n79 9.154
R432 GND.n85 GND.n84 9.154
R433 GND.n84 GND.n83 9.154
R434 GND.n89 GND.n88 9.154
R435 GND.n88 GND.n87 9.154
R436 GND.n93 GND.n92 9.154
R437 GND.n92 GND.n91 9.154
R438 GND.n97 GND.n96 9.154
R439 GND.n105 GND.n104 9.154
R440 GND.n109 GND.n108 9.154
R441 GND.n108 GND.n107 9.154
R442 GND.n113 GND.n112 9.154
R443 GND.n112 GND.n111 9.154
R444 GND.n117 GND.n116 9.154
R445 GND.n116 GND.n115 9.154
R446 GND.n122 GND.n121 9.154
R447 GND.n121 GND.n120 9.154
R448 GND.n126 GND.n125 9.154
R449 GND.n125 GND.n124 9.154
R450 GND.n130 GND.n129 9.154
R451 GND.n129 GND.n128 9.154
R452 GND.n133 GND.n2 9.154
R453 GND.n2 GND.n1 9.154
R454 GND.n136 GND.n135 9.154
R455 GND.n135 GND.n134 9.154
R456 GND.n140 GND.n139 9.154
R457 GND.n139 GND.n138 9.154
R458 GND.n144 GND.n143 9.154
R459 GND.n143 GND.n142 9.154
R460 GND.n149 GND.n148 9.154
R461 GND.n148 GND.n147 9.154
R462 GND.n153 GND.n152 9.154
R463 GND.n152 GND.n151 9.154
R464 GND.n157 GND.n156 9.154
R465 GND.n156 GND.n155 9.154
R466 GND.n161 GND.n160 9.154
R467 GND.n169 GND.n168 9.154
R468 GND.n173 GND.n172 9.154
R469 GND.n172 GND.n171 9.154
R470 GND.n177 GND.n176 9.154
R471 GND.n176 GND.n175 9.154
R472 GND.n181 GND.n180 9.154
R473 GND.n180 GND.n179 9.154
R474 GND.n185 GND.n184 9.154
R475 GND.n184 GND.n183 9.154
R476 GND.n189 GND.n188 9.154
R477 GND.n188 GND.n187 9.154
R478 GND.n193 GND.n192 9.154
R479 GND.n192 GND.n191 9.154
R480 GND.n197 GND.n196 9.154
R481 GND.n196 GND.n195 9.154
R482 GND.n202 GND.n201 9.154
R483 GND.n201 GND.n200 9.154
R484 GND.n206 GND.n205 9.154
R485 GND.n205 GND.n204 9.154
R486 GND.n210 GND.n209 9.154
R487 GND.n209 GND.n208 9.154
R488 GND.n214 GND.n213 9.154
R489 GND.n213 GND.n212 9.154
R490 GND.n519 GND.n518 9.154
R491 GND.n518 GND.n517 9.154
R492 GND.n515 GND.n514 9.154
R493 GND.n514 GND.n513 9.154
R494 GND.n511 GND.n510 9.154
R495 GND.n510 GND.n509 9.154
R496 GND.n506 GND.n505 9.154
R497 GND.n505 GND.n504 9.154
R498 GND.n502 GND.n501 9.154
R499 GND.n501 GND.n500 9.154
R500 GND.n498 GND.n497 9.154
R501 GND.n497 GND.n496 9.154
R502 GND.n494 GND.n493 9.154
R503 GND.n493 GND.n492 9.154
R504 GND.n490 GND.n489 9.154
R505 GND.n489 GND.n488 9.154
R506 GND.n486 GND.n485 9.154
R507 GND.n485 GND.n484 9.154
R508 GND.n482 GND.n481 9.154
R509 GND.n481 GND.n480 9.154
R510 GND.n478 GND.n477 9.154
R511 GND.n433 GND.n432 5.103
R512 GND.n433 GND.n431 5.103
R513 GND.n329 GND.n293 5.103
R514 GND.n329 GND.n292 5.103
R515 GND.n381 GND.n264 5.103
R516 GND.n381 GND.n263 5.103
R517 GND.n215 GND.n0 5.103
R518 GND.n132 GND.n3 5.103
R519 GND.n52 GND.n6 5.103
R520 GND.n400 GND.n399 4.65
R521 GND.n360 GND.n274 4.65
R522 GND.n362 GND.n361 4.65
R523 GND.n271 GND.n270 4.65
R524 GND.n370 GND.n369 4.65
R525 GND.n372 GND.n269 4.65
R526 GND.n374 GND.n373 4.65
R527 GND.n266 GND.n265 4.65
R528 GND.n381 GND.n380 4.65
R529 GND.n382 GND.n262 4.65
R530 GND.n385 GND.n384 4.65
R531 GND.n383 GND.n258 4.65
R532 GND.n392 GND.n391 4.65
R533 GND.n393 GND.n256 4.65
R534 GND.n395 GND.n394 4.65
R535 GND.n252 GND.n251 4.65
R536 GND.n359 GND.n358 4.65
R537 GND.n356 GND.n355 4.65
R538 GND.n308 GND.n307 4.65
R539 GND.n301 GND.n300 4.65
R540 GND.n315 GND.n314 4.65
R541 GND.n316 GND.n299 4.65
R542 GND.n319 GND.n318 4.65
R543 GND.n295 GND.n294 4.65
R544 GND.n327 GND.n326 4.65
R545 GND.n328 GND.n291 4.65
R546 GND.n330 GND.n329 4.65
R547 GND.n288 GND.n287 4.65
R548 GND.n337 GND.n336 4.65
R549 GND.n338 GND.n286 4.65
R550 GND.n341 GND.n340 4.65
R551 GND.n282 GND.n281 4.65
R552 GND.n348 GND.n347 4.65
R553 GND.n349 GND.n280 4.65
R554 GND.n351 GND.n350 4.65
R555 GND.n276 GND.n275 4.65
R556 GND.n249 GND.n248 4.65
R557 GND.n408 GND.n407 4.65
R558 GND.n409 GND.n247 4.65
R559 GND.n411 GND.n410 4.65
R560 GND.n243 GND.n242 4.65
R561 GND.n418 GND.n417 4.65
R562 GND.n419 GND.n241 4.65
R563 GND.n422 GND.n421 4.65
R564 GND.n420 GND.n237 4.65
R565 GND.n429 GND.n428 4.65
R566 GND.n430 GND.n235 4.65
R567 GND.n435 GND.n434 4.65
R568 GND.n433 GND.n231 4.65
R569 GND.n443 GND.n442 4.65
R570 GND.n444 GND.n230 4.65
R571 GND.n447 GND.n446 4.65
R572 GND.n227 GND.n226 4.65
R573 GND.n455 GND.n454 4.65
R574 GND.n456 GND.n225 4.65
R575 GND.n458 GND.n457 4.65
R576 GND.n222 GND.n221 4.65
R577 GND.n466 GND.n465 4.65
R578 GND.n467 GND.n219 4.65
R579 GND.n469 GND.n468 4.65
R580 GND.n402 GND.n401 4.65
R581 GND.n14 GND.n13 4.65
R582 GND.n18 GND.n17 4.65
R583 GND.n22 GND.n21 4.65
R584 GND.n26 GND.n25 4.65
R585 GND.n30 GND.n29 4.65
R586 GND.n34 GND.n33 4.65
R587 GND.n38 GND.n37 4.65
R588 GND.n43 GND.n42 4.65
R589 GND.n47 GND.n46 4.65
R590 GND.n51 GND.n50 4.65
R591 GND.n53 GND.n52 4.65
R592 GND.n57 GND.n56 4.65
R593 GND.n61 GND.n60 4.65
R594 GND.n65 GND.n64 4.65
R595 GND.n70 GND.n69 4.65
R596 GND.n74 GND.n73 4.65
R597 GND.n78 GND.n77 4.65
R598 GND.n82 GND.n81 4.65
R599 GND.n86 GND.n85 4.65
R600 GND.n90 GND.n89 4.65
R601 GND.n94 GND.n93 4.65
R602 GND.n98 GND.n97 4.65
R603 GND.n100 GND.n99 4.65
R604 GND.n102 GND.n101 4.65
R605 GND.n106 GND.n105 4.65
R606 GND.n110 GND.n109 4.65
R607 GND.n114 GND.n113 4.65
R608 GND.n118 GND.n117 4.65
R609 GND.n123 GND.n122 4.65
R610 GND.n127 GND.n126 4.65
R611 GND.n131 GND.n130 4.65
R612 GND.n133 GND.n132 4.65
R613 GND.n137 GND.n136 4.65
R614 GND.n141 GND.n140 4.65
R615 GND.n145 GND.n144 4.65
R616 GND.n150 GND.n149 4.65
R617 GND.n154 GND.n153 4.65
R618 GND.n158 GND.n157 4.65
R619 GND.n162 GND.n161 4.65
R620 GND.n164 GND.n163 4.65
R621 GND.n166 GND.n165 4.65
R622 GND.n170 GND.n169 4.65
R623 GND.n174 GND.n173 4.65
R624 GND.n178 GND.n177 4.65
R625 GND.n182 GND.n181 4.65
R626 GND.n186 GND.n185 4.65
R627 GND.n190 GND.n189 4.65
R628 GND.n194 GND.n193 4.65
R629 GND.n198 GND.n197 4.65
R630 GND.n203 GND.n202 4.65
R631 GND.n207 GND.n206 4.65
R632 GND.n211 GND.n210 4.65
R633 GND.n215 GND.n214 4.65
R634 GND.n520 GND.n519 4.65
R635 GND.n516 GND.n515 4.65
R636 GND.n512 GND.n511 4.65
R637 GND.n507 GND.n506 4.65
R638 GND.n503 GND.n502 4.65
R639 GND.n499 GND.n498 4.65
R640 GND.n495 GND.n494 4.65
R641 GND.n491 GND.n490 4.65
R642 GND.n487 GND.n486 4.65
R643 GND.n483 GND.n482 4.65
R644 GND.n305 GND.n303 2.791
R645 GND.n357 GND.n273 2.791
R646 GND.n398 GND.n253 2.791
R647 GND.n354 GND.n277 2.791
R648 GND.n474 GND.n216 2.739
R649 GND.n479 GND.n475 2.739
R650 GND.n10 GND.n9 2.682
R651 GND.n306 GND.n304 2.682
R652 GND.n220 GND.n216 2.682
R653 GND.n479 GND.n478 2.682
R654 GND.n8 GND.n7 1.873
R655 GND.n104 GND.n103 1.873
R656 GND.n477 GND.n476 1.873
R657 GND.n96 GND.n95 1.873
R658 GND.n160 GND.n159 1.873
R659 GND.n168 GND.n167 1.873
R660 GND.n14 GND.n10 1.096
R661 GND.n307 GND.n306 1.095
R662 GND.n468 GND.n216 1.095
R663 GND.n483 GND.n479 1.095
R664 GND.n401 GND.n400 0.637
R665 GND.n166 GND.n164 0.562
R666 GND.n359 GND.n356 0.55
R667 GND.n102 GND.n100 0.55
R668 GND.n307 GND.n300 0.1
R669 GND.n315 GND.n300 0.1
R670 GND.n316 GND.n315 0.1
R671 GND.n318 GND.n316 0.1
R672 GND.n327 GND.n294 0.1
R673 GND.n328 GND.n327 0.1
R674 GND.n329 GND.n328 0.1
R675 GND.n337 GND.n287 0.1
R676 GND.n338 GND.n337 0.1
R677 GND.n340 GND.n281 0.1
R678 GND.n348 GND.n281 0.1
R679 GND.n349 GND.n348 0.1
R680 GND.n350 GND.n349 0.1
R681 GND.n350 GND.n275 0.1
R682 GND.n356 GND.n275 0.1
R683 GND.n360 GND.n359 0.1
R684 GND.n361 GND.n360 0.1
R685 GND.n361 GND.n270 0.1
R686 GND.n370 GND.n270 0.1
R687 GND.n373 GND.n372 0.1
R688 GND.n373 GND.n265 0.1
R689 GND.n381 GND.n265 0.1
R690 GND.n384 GND.n382 0.1
R691 GND.n384 GND.n383 0.1
R692 GND.n393 GND.n392 0.1
R693 GND.n394 GND.n393 0.1
R694 GND.n394 GND.n251 0.1
R695 GND.n400 GND.n251 0.1
R696 GND.n401 GND.n248 0.1
R697 GND.n408 GND.n248 0.1
R698 GND.n409 GND.n408 0.1
R699 GND.n410 GND.n409 0.1
R700 GND.n410 GND.n242 0.1
R701 GND.n418 GND.n242 0.1
R702 GND.n419 GND.n418 0.1
R703 GND.n421 GND.n419 0.1
R704 GND.n421 GND.n420 0.1
R705 GND.n430 GND.n429 0.1
R706 GND.n434 GND.n430 0.1
R707 GND.n434 GND.n433 0.1
R708 GND.n444 GND.n443 0.1
R709 GND.n446 GND.n444 0.1
R710 GND.n455 GND.n226 0.1
R711 GND.n456 GND.n455 0.1
R712 GND.n457 GND.n456 0.1
R713 GND.n457 GND.n221 0.1
R714 GND.n466 GND.n221 0.1
R715 GND.n467 GND.n466 0.1
R716 GND.n468 GND.n467 0.1
R717 GND.n18 GND.n14 0.1
R718 GND.n22 GND.n18 0.1
R719 GND.n26 GND.n22 0.1
R720 GND.n30 GND.n26 0.1
R721 GND.n34 GND.n30 0.1
R722 GND.n38 GND.n34 0.1
R723 GND.n47 GND.n43 0.1
R724 GND.n51 GND.n47 0.1
R725 GND.n52 GND.n51 0.1
R726 GND.n61 GND.n57 0.1
R727 GND.n65 GND.n61 0.1
R728 GND.n74 GND.n70 0.1
R729 GND.n78 GND.n74 0.1
R730 GND.n82 GND.n78 0.1
R731 GND.n86 GND.n82 0.1
R732 GND.n90 GND.n86 0.1
R733 GND.n94 GND.n90 0.1
R734 GND.n98 GND.n94 0.1
R735 GND.n100 GND.n98 0.1
R736 GND.n106 GND.n102 0.1
R737 GND.n110 GND.n106 0.1
R738 GND.n114 GND.n110 0.1
R739 GND.n118 GND.n114 0.1
R740 GND.n127 GND.n123 0.1
R741 GND.n131 GND.n127 0.1
R742 GND.n132 GND.n131 0.1
R743 GND.n141 GND.n137 0.1
R744 GND.n145 GND.n141 0.1
R745 GND.n154 GND.n150 0.1
R746 GND.n158 GND.n154 0.1
R747 GND.n162 GND.n158 0.1
R748 GND.n164 GND.n162 0.1
R749 GND.n170 GND.n166 0.1
R750 GND.n174 GND.n170 0.1
R751 GND.n178 GND.n174 0.1
R752 GND.n182 GND.n178 0.1
R753 GND.n186 GND.n182 0.1
R754 GND.n190 GND.n186 0.1
R755 GND.n194 GND.n190 0.1
R756 GND.n198 GND.n194 0.1
R757 GND.n207 GND.n203 0.1
R758 GND.n211 GND.n207 0.1
R759 GND.n215 GND.n211 0.1
R760 GND.n520 GND.n516 0.1
R761 GND.n516 GND.n512 0.1
R762 GND.n507 GND.n503 0.1
R763 GND.n503 GND.n499 0.1
R764 GND.n499 GND.n495 0.1
R765 GND.n495 GND.n491 0.1
R766 GND.n491 GND.n487 0.1
R767 GND.n487 GND.n483 0.1
R768 GND.n317 GND.n294 0.075
R769 GND GND.n287 0.075
R770 GND.n339 GND.n338 0.075
R771 GND.n372 GND.n371 0.075
R772 GND.n382 EESPFAL_INV4_2/GND 0.075
R773 GND.n383 GND.n257 0.075
R774 GND.n429 GND.n236 0.075
R775 GND.n443 EESPFAL_XOR_v3_0/GND 0.075
R776 GND.n446 GND.n445 0.075
R777 GND.n43 GND.n39 0.075
R778 GND.n57 EESPFAL_3in_NOR_v2_0/GND 0.075
R779 GND.n66 GND.n65 0.075
R780 GND.n123 GND.n119 0.075
R781 GND.n137 EESPFAL_INV4_0/GND 0.075
R782 GND.n146 GND.n145 0.075
R783 GND.n203 GND.n199 0.075
R784 EESPFAL_3in_NAND_v2_0/GND GND.n520 0.075
R785 GND.n512 GND.n508 0.075
R786 GND.n318 GND.n317 0.025
R787 GND.n329 GND 0.025
R788 GND.n340 GND.n339 0.025
R789 GND.n371 GND.n370 0.025
R790 EESPFAL_INV4_2/GND GND.n381 0.025
R791 GND.n392 GND.n257 0.025
R792 GND.n420 GND.n236 0.025
R793 GND.n433 EESPFAL_XOR_v3_0/GND 0.025
R794 GND.n445 GND.n226 0.025
R795 GND.n39 GND.n38 0.025
R796 GND.n52 EESPFAL_3in_NOR_v2_0/GND 0.025
R797 GND.n70 GND.n66 0.025
R798 GND.n119 GND.n118 0.025
R799 GND.n132 EESPFAL_INV4_0/GND 0.025
R800 GND.n150 GND.n146 0.025
R801 GND.n199 GND.n198 0.025
R802 EESPFAL_3in_NAND_v2_0/GND GND.n215 0.025
R803 GND.n508 GND.n507 0.025
R804 CLK2.n132 CLK2.t9 44.338
R805 CLK2.n103 CLK2.t16 44.338
R806 CLK2.n240 CLK2.t24 44.337
R807 CLK2.n197 CLK2.t3 44.337
R808 CLK2.n29 CLK2.t26 44.337
R809 CLK2.n58 CLK2.t20 44.337
R810 CLK2.n0 CLK2.t1 39.4
R811 CLK2.n0 CLK2.t22 39.4
R812 CLK2.n6 CLK2.t11 39.4
R813 CLK2.n6 CLK2.t14 39.4
R814 CLK2.n10 CLK2.t18 39.4
R815 CLK2.n10 CLK2.t30 39.4
R816 CLK2.n12 CLK2.t5 29.712
R817 CLK2.n75 CLK2.t12 29.712
R818 CLK2.n198 CLK2.t2 24.568
R819 CLK2.n241 CLK2.t23 24.568
R820 CLK2.n128 CLK2.t8 24.568
R821 CLK2.n104 CLK2.t15 24.568
R822 CLK2.n54 CLK2.t19 24.568
R823 CLK2.n30 CLK2.t25 24.568
R824 CLK2.n214 CLK2.t31 24
R825 CLK2.n214 CLK2.t27 24
R826 CLK2.n161 CLK2.t4 24
R827 CLK2.n7 CLK2.t7 24
R828 CLK2.n7 CLK2.t6 24
R829 CLK2.n1 CLK2.t28 24
R830 CLK2.n118 CLK2.n115 12.8
R831 CLK2.n44 CLK2.n41 12.8
R832 CLK2.n155 CLK2.n154 8.855
R833 CLK2.n73 CLK2.n72 8.855
R834 CLK2.n69 CLK2.n68 8.855
R835 CLK2.n68 CLK2.n67 8.855
R836 CLK2.n65 CLK2.n64 8.855
R837 CLK2.n64 CLK2.n63 8.855
R838 CLK2.n61 CLK2.n60 8.855
R839 CLK2.n60 CLK2.n59 8.855
R840 CLK2.n56 CLK2.n55 8.855
R841 CLK2.n55 CLK2.n54 8.855
R842 CLK2.n52 CLK2.n51 8.855
R843 CLK2.n51 CLK2.n50 8.855
R844 CLK2.n48 CLK2.n47 8.855
R845 CLK2.n47 CLK2.n46 8.855
R846 CLK2.n44 CLK2.n43 8.855
R847 CLK2.n43 CLK2.n42 8.855
R848 CLK2.n41 CLK2.n40 8.855
R849 CLK2.n40 CLK2.n39 8.855
R850 CLK2.n36 CLK2.n35 8.855
R851 CLK2.n35 CLK2.n34 8.855
R852 CLK2.n32 CLK2.n31 8.855
R853 CLK2.n31 CLK2.n30 8.855
R854 CLK2.n27 CLK2.n26 8.855
R855 CLK2.n26 CLK2.n25 8.855
R856 CLK2.n23 CLK2.n22 8.855
R857 CLK2.n22 CLK2.n21 8.855
R858 CLK2.n19 CLK2.n18 8.855
R859 CLK2.n18 CLK2.n17 8.855
R860 CLK2.n15 CLK2.n14 8.855
R861 CLK2.n151 CLK2.n150 8.855
R862 CLK2.n150 CLK2.n149 8.855
R863 CLK2.n147 CLK2.n146 8.855
R864 CLK2.n146 CLK2.n145 8.855
R865 CLK2.n143 CLK2.n142 8.855
R866 CLK2.n142 CLK2.n141 8.855
R867 CLK2.n139 CLK2.n138 8.855
R868 CLK2.n138 CLK2.n137 8.855
R869 CLK2.n135 CLK2.n134 8.855
R870 CLK2.n134 CLK2.n133 8.855
R871 CLK2.n130 CLK2.n129 8.855
R872 CLK2.n129 CLK2.n128 8.855
R873 CLK2.n126 CLK2.n125 8.855
R874 CLK2.n125 CLK2.n124 8.855
R875 CLK2.n122 CLK2.n121 8.855
R876 CLK2.n121 CLK2.n120 8.855
R877 CLK2.n118 CLK2.n117 8.855
R878 CLK2.n117 CLK2.n116 8.855
R879 CLK2.n115 CLK2.n114 8.855
R880 CLK2.n114 CLK2.n113 8.855
R881 CLK2.n110 CLK2.n109 8.855
R882 CLK2.n109 CLK2.n108 8.855
R883 CLK2.n106 CLK2.n105 8.855
R884 CLK2.n105 CLK2.n104 8.855
R885 CLK2.n101 CLK2.n100 8.855
R886 CLK2.n100 CLK2.n99 8.855
R887 CLK2.n97 CLK2.n96 8.855
R888 CLK2.n96 CLK2.n95 8.855
R889 CLK2.n93 CLK2.n92 8.855
R890 CLK2.n92 CLK2.n91 8.855
R891 CLK2.n89 CLK2.n88 8.855
R892 CLK2.n88 CLK2.n87 8.855
R893 CLK2.n84 CLK2.n83 8.855
R894 CLK2.n83 CLK2.n82 8.855
R895 CLK2.n80 CLK2.n79 8.855
R896 CLK2.n175 CLK2.n174 8.855
R897 CLK2.n179 CLK2.n178 8.855
R898 CLK2.n178 CLK2.n177 8.855
R899 CLK2.n183 CLK2.n182 8.855
R900 CLK2.n182 CLK2.n181 8.855
R901 CLK2.n187 CLK2.n186 8.855
R902 CLK2.n186 CLK2.n185 8.855
R903 CLK2.n191 CLK2.n190 8.855
R904 CLK2.n190 CLK2.n189 8.855
R905 CLK2.n195 CLK2.n194 8.855
R906 CLK2.n194 CLK2.n193 8.855
R907 CLK2.n200 CLK2.n199 8.855
R908 CLK2.n199 CLK2.n198 8.855
R909 CLK2.n204 CLK2.n203 8.855
R910 CLK2.n203 CLK2.n202 8.855
R911 CLK2.n208 CLK2.n207 8.855
R912 CLK2.n207 CLK2.n206 8.855
R913 CLK2.n212 CLK2.n211 8.855
R914 CLK2.n211 CLK2.n210 8.855
R915 CLK2.n251 CLK2.n250 8.855
R916 CLK2.n250 CLK2.n249 8.855
R917 CLK2.n247 CLK2.n246 8.855
R918 CLK2.n246 CLK2.n245 8.855
R919 CLK2.n243 CLK2.n242 8.855
R920 CLK2.n242 CLK2.n241 8.855
R921 CLK2.n238 CLK2.n237 8.855
R922 CLK2.n237 CLK2.n236 8.855
R923 CLK2.n234 CLK2.n233 8.855
R924 CLK2.n233 CLK2.n232 8.855
R925 CLK2.n230 CLK2.n229 8.855
R926 CLK2.n229 CLK2.n228 8.855
R927 CLK2.n226 CLK2.n225 8.855
R928 CLK2.n225 CLK2.n224 8.855
R929 CLK2.n221 CLK2.n220 8.855
R930 CLK2.n220 CLK2.n219 8.855
R931 CLK2.n217 CLK2.n216 8.855
R932 CLK2.n167 CLK2.n2 8.365
R933 CLK2.n206 CLK2.t0 8.189
R934 CLK2.n249 CLK2.t21 8.189
R935 CLK2.n120 CLK2.t10 8.189
R936 CLK2.n113 CLK2.t13 8.189
R937 CLK2.n46 CLK2.t17 8.189
R938 CLK2.n39 CLK2.t29 8.189
R939 CLK2.n223 CLK2.n214 6.776
R940 CLK2.n86 CLK2.n7 6.776
R941 CLK2.n163 CLK2.n162 6.754
R942 CLK2.n213 CLK2.n0 4.938
R943 CLK2.n119 CLK2.n6 4.938
R944 CLK2.n45 CLK2.n10 4.938
R945 CLK2.n157 CLK2.n5 4.675
R946 CLK2.n12 CLK2.n11 4.662
R947 CLK2.n74 CLK2.n73 4.65
R948 CLK2.n70 CLK2.n69 4.65
R949 CLK2.n66 CLK2.n65 4.65
R950 CLK2.n62 CLK2.n61 4.65
R951 CLK2.n57 CLK2.n56 4.65
R952 CLK2.n53 CLK2.n52 4.65
R953 CLK2.n49 CLK2.n48 4.65
R954 CLK2.n45 CLK2.n44 4.65
R955 CLK2.n41 CLK2.n38 4.65
R956 CLK2.n37 CLK2.n36 4.65
R957 CLK2.n33 CLK2.n32 4.65
R958 CLK2.n28 CLK2.n27 4.65
R959 CLK2.n24 CLK2.n23 4.65
R960 CLK2.n20 CLK2.n19 4.65
R961 CLK2.n16 CLK2.n15 4.65
R962 CLK2.n76 CLK2.n9 4.65
R963 CLK2.n77 CLK2.n8 4.65
R964 CLK2.n156 CLK2.n155 4.65
R965 CLK2.n152 CLK2.n151 4.65
R966 CLK2.n148 CLK2.n147 4.65
R967 CLK2.n144 CLK2.n143 4.65
R968 CLK2.n140 CLK2.n139 4.65
R969 CLK2.n136 CLK2.n135 4.65
R970 CLK2.n131 CLK2.n130 4.65
R971 CLK2.n127 CLK2.n126 4.65
R972 CLK2.n123 CLK2.n122 4.65
R973 CLK2.n119 CLK2.n118 4.65
R974 CLK2.n115 CLK2.n112 4.65
R975 CLK2.n111 CLK2.n110 4.65
R976 CLK2.n107 CLK2.n106 4.65
R977 CLK2.n102 CLK2.n101 4.65
R978 CLK2.n98 CLK2.n97 4.65
R979 CLK2.n94 CLK2.n93 4.65
R980 CLK2.n90 CLK2.n89 4.65
R981 CLK2.n85 CLK2.n84 4.65
R982 CLK2.n81 CLK2.n80 4.65
R983 CLK2.n160 CLK2.n4 4.65
R984 CLK2.n159 CLK2.n158 4.65
R985 CLK2.n166 CLK2.n165 4.65
R986 CLK2.n176 CLK2.n175 4.65
R987 CLK2.n180 CLK2.n179 4.65
R988 CLK2.n184 CLK2.n183 4.65
R989 CLK2.n188 CLK2.n187 4.65
R990 CLK2.n192 CLK2.n191 4.65
R991 CLK2.n196 CLK2.n195 4.65
R992 CLK2.n201 CLK2.n200 4.65
R993 CLK2.n205 CLK2.n204 4.65
R994 CLK2.n209 CLK2.n208 4.65
R995 CLK2.n213 CLK2.n212 4.65
R996 CLK2.n252 CLK2.n251 4.65
R997 CLK2.n248 CLK2.n247 4.65
R998 CLK2.n244 CLK2.n243 4.65
R999 CLK2.n239 CLK2.n238 4.65
R1000 CLK2.n235 CLK2.n234 4.65
R1001 CLK2.n231 CLK2.n230 4.65
R1002 CLK2.n227 CLK2.n226 4.65
R1003 CLK2.n222 CLK2.n221 4.65
R1004 CLK2.n164 CLK2.n3 3.039
R1005 CLK2.n170 CLK2.n169 3.033
R1006 CLK2.n218 CLK2.n217 2.682
R1007 CLK2.n162 CLK2.n161 2.57
R1008 CLK2.n2 CLK2.n1 2.57
R1009 CLK2.n164 CLK2.n163 2.224
R1010 CLK2.n159 CLK2.n157 2.203
R1011 CLK2.n171 CLK2.n167 2.203
R1012 CLK2.n174 CLK2.n173 1.655
R1013 CLK2.n154 CLK2.n153 1.655
R1014 CLK2.n72 CLK2.n71 1.655
R1015 CLK2.n14 CLK2.n13 1.655
R1016 CLK2.n79 CLK2.n78 1.655
R1017 CLK2.n216 CLK2.n215 1.655
R1018 CLK2.n222 CLK2.n218 1.095
R1019 CLK2.n77 CLK2.n76 1.047
R1020 CLK2.n170 CLK2.n168 0.898
R1021 CLK2.n168 CLK2 0.155
R1022 CLK2.n160 CLK2.n159 0.125
R1023 CLK2.n167 CLK2.n166 0.125
R1024 CLK2.n166 CLK2.n164 0.12
R1025 CLK2.n163 CLK2.n160 0.119
R1026 CLK2.n74 CLK2.n70 0.1
R1027 CLK2.n70 CLK2.n66 0.1
R1028 CLK2.n66 CLK2.n62 0.1
R1029 CLK2.n57 CLK2.n53 0.1
R1030 CLK2.n53 CLK2.n49 0.1
R1031 CLK2.n49 CLK2.n45 0.1
R1032 CLK2.n38 CLK2.n37 0.1
R1033 CLK2.n37 CLK2.n33 0.1
R1034 CLK2.n28 CLK2.n24 0.1
R1035 CLK2.n24 CLK2.n20 0.1
R1036 CLK2.n20 CLK2.n16 0.1
R1037 CLK2.n156 CLK2.n152 0.1
R1038 CLK2.n152 CLK2.n148 0.1
R1039 CLK2.n148 CLK2.n144 0.1
R1040 CLK2.n144 CLK2.n140 0.1
R1041 CLK2.n140 CLK2.n136 0.1
R1042 CLK2.n131 CLK2.n127 0.1
R1043 CLK2.n127 CLK2.n123 0.1
R1044 CLK2.n123 CLK2.n119 0.1
R1045 CLK2.n112 CLK2.n111 0.1
R1046 CLK2.n111 CLK2.n107 0.1
R1047 CLK2.n102 CLK2.n98 0.1
R1048 CLK2.n98 CLK2.n94 0.1
R1049 CLK2.n94 CLK2.n90 0.1
R1050 CLK2.n85 CLK2.n81 0.1
R1051 CLK2.n81 CLK2.n77 0.1
R1052 CLK2.n180 CLK2.n176 0.1
R1053 CLK2.n184 CLK2.n180 0.1
R1054 CLK2.n188 CLK2.n184 0.1
R1055 CLK2.n192 CLK2.n188 0.1
R1056 CLK2.n196 CLK2.n192 0.1
R1057 CLK2.n205 CLK2.n201 0.1
R1058 CLK2.n209 CLK2.n205 0.1
R1059 CLK2.n213 CLK2.n209 0.1
R1060 CLK2.n252 CLK2.n248 0.1
R1061 CLK2.n248 CLK2.n244 0.1
R1062 CLK2.n239 CLK2.n235 0.1
R1063 CLK2.n235 CLK2.n231 0.1
R1064 CLK2.n231 CLK2.n227 0.1
R1065 CLK2.n75 CLK2.n74 0.087
R1066 CLK2.n16 CLK2.n12 0.087
R1067 CLK2.n90 CLK2.n86 0.087
R1068 CLK2.n227 CLK2.n223 0.087
R1069 CLK2.n58 CLK2.n57 0.075
R1070 CLK2.n38 EESPFAL_INV4_0/CLK 0.075
R1071 CLK2.n33 CLK2.n29 0.075
R1072 CLK2.n157 CLK2.n156 0.075
R1073 CLK2.n132 CLK2.n131 0.075
R1074 CLK2.n112 EESPFAL_NAND_v3_1/CLK 0.075
R1075 CLK2.n107 CLK2.n103 0.075
R1076 CLK2.n201 CLK2.n197 0.075
R1077 CLK2 CLK2.n252 0.075
R1078 CLK2.n244 CLK2.n240 0.075
R1079 CLK2.n176 CLK2.n172 0.072
R1080 CLK2.n62 CLK2.n58 0.025
R1081 CLK2.n45 EESPFAL_INV4_0/CLK 0.025
R1082 CLK2.n29 CLK2.n28 0.025
R1083 CLK2.n136 CLK2.n132 0.025
R1084 CLK2.n119 EESPFAL_NAND_v3_1/CLK 0.025
R1085 CLK2.n103 CLK2.n102 0.025
R1086 CLK2.n171 CLK2.n170 0.025
R1087 CLK2.n197 CLK2.n196 0.025
R1088 CLK2 CLK2.n213 0.025
R1089 CLK2.n240 CLK2.n239 0.025
R1090 CLK2.n76 CLK2.n75 0.012
R1091 CLK2.n86 CLK2.n85 0.012
R1092 CLK2.n223 CLK2.n222 0.012
R1093 CLK2.n172 CLK2.n171 0.002
R1094 CLK1.n21 CLK1.t10 44.338
R1095 CLK1.n50 CLK1.t20 44.338
R1096 CLK1.n109 CLK1.t50 44.338
R1097 CLK1.n461 CLK1.t3 44.338
R1098 CLK1.n267 CLK1.t55 44.337
R1099 CLK1.n240 CLK1.t36 44.337
R1100 CLK1.n181 CLK1.t40 44.337
R1101 CLK1.n154 CLK1.t43 44.337
R1102 CLK1.n380 CLK1.t27 44.337
R1103 CLK1.n351 CLK1.t14 44.337
R1104 CLK1.n131 CLK1.t47 39.4
R1105 CLK1.n131 CLK1.t32 39.4
R1106 CLK1.n135 CLK1.t45 39.4
R1107 CLK1.n135 CLK1.t38 39.4
R1108 CLK1.n316 CLK1.t16 39.4
R1109 CLK1.n316 CLK1.t25 39.4
R1110 CLK1.n0 CLK1.t22 39.4
R1111 CLK1.n0 CLK1.t53 39.4
R1112 CLK1.n2 CLK1.t8 39.4
R1113 CLK1.n2 CLK1.t18 39.4
R1114 CLK1.n414 CLK1.t48 30.775
R1115 CLK1.n318 CLK1.t12 30.775
R1116 CLK1.n4 CLK1.t5 29.713
R1117 CLK1.n67 CLK1.t0 29.713
R1118 CLK1.n198 CLK1.t41 29.712
R1119 CLK1.n137 CLK1.t34 29.712
R1120 CLK1.n241 CLK1.t35 24.568
R1121 CLK1.n263 CLK1.t54 24.568
R1122 CLK1.n155 CLK1.t42 24.568
R1123 CLK1.n177 CLK1.t39 24.568
R1124 CLK1.n352 CLK1.t13 24.568
R1125 CLK1.n376 CLK1.t26 24.568
R1126 CLK1.n110 CLK1.t49 24.568
R1127 CLK1.n462 CLK1.t2 24.568
R1128 CLK1.n22 CLK1.t9 24.568
R1129 CLK1.n46 CLK1.t19 24.568
R1130 CLK1.n128 CLK1.t6 24
R1131 CLK1.n128 CLK1.t51 24
R1132 CLK1.n132 CLK1.t1 24
R1133 CLK1.n132 CLK1.t4 24
R1134 CLK1.n315 CLK1.t33 24
R1135 CLK1.n315 CLK1.t11 24
R1136 CLK1.n1 CLK1.t29 24
R1137 CLK1.n1 CLK1.t28 24
R1138 CLK1.n126 CLK1.t23 24
R1139 CLK1.n126 CLK1.t30 24
R1140 CLK1.n257 CLK1.n254 12.8
R1141 CLK1.n171 CLK1.n168 12.8
R1142 CLK1.n370 CLK1.n367 12.8
R1143 CLK1.n40 CLK1.n37 12.8
R1144 CLK1.n140 CLK1.n139 8.855
R1145 CLK1.n144 CLK1.n143 8.855
R1146 CLK1.n143 CLK1.n142 8.855
R1147 CLK1.n148 CLK1.n147 8.855
R1148 CLK1.n147 CLK1.n146 8.855
R1149 CLK1.n152 CLK1.n151 8.855
R1150 CLK1.n151 CLK1.n150 8.855
R1151 CLK1.n157 CLK1.n156 8.855
R1152 CLK1.n156 CLK1.n155 8.855
R1153 CLK1.n161 CLK1.n160 8.855
R1154 CLK1.n160 CLK1.n159 8.855
R1155 CLK1.n165 CLK1.n164 8.855
R1156 CLK1.n164 CLK1.n163 8.855
R1157 CLK1.n168 CLK1.n134 8.855
R1158 CLK1.n134 CLK1.n133 8.855
R1159 CLK1.n171 CLK1.n170 8.855
R1160 CLK1.n170 CLK1.n169 8.855
R1161 CLK1.n175 CLK1.n174 8.855
R1162 CLK1.n174 CLK1.n173 8.855
R1163 CLK1.n179 CLK1.n178 8.855
R1164 CLK1.n178 CLK1.n177 8.855
R1165 CLK1.n184 CLK1.n183 8.855
R1166 CLK1.n183 CLK1.n182 8.855
R1167 CLK1.n188 CLK1.n187 8.855
R1168 CLK1.n187 CLK1.n186 8.855
R1169 CLK1.n192 CLK1.n191 8.855
R1170 CLK1.n191 CLK1.n190 8.855
R1171 CLK1.n196 CLK1.n195 8.855
R1172 CLK1.n205 CLK1.n204 8.855
R1173 CLK1.n209 CLK1.n208 8.855
R1174 CLK1.n208 CLK1.n207 8.855
R1175 CLK1.n213 CLK1.n212 8.855
R1176 CLK1.n212 CLK1.n211 8.855
R1177 CLK1.n218 CLK1.n217 8.855
R1178 CLK1.n217 CLK1.n216 8.855
R1179 CLK1.n222 CLK1.n221 8.855
R1180 CLK1.n221 CLK1.n220 8.855
R1181 CLK1.n226 CLK1.n225 8.855
R1182 CLK1.n225 CLK1.n224 8.855
R1183 CLK1.n230 CLK1.n229 8.855
R1184 CLK1.n229 CLK1.n228 8.855
R1185 CLK1.n234 CLK1.n233 8.855
R1186 CLK1.n233 CLK1.n232 8.855
R1187 CLK1.n238 CLK1.n237 8.855
R1188 CLK1.n237 CLK1.n236 8.855
R1189 CLK1.n243 CLK1.n242 8.855
R1190 CLK1.n242 CLK1.n241 8.855
R1191 CLK1.n247 CLK1.n246 8.855
R1192 CLK1.n246 CLK1.n245 8.855
R1193 CLK1.n251 CLK1.n250 8.855
R1194 CLK1.n250 CLK1.n249 8.855
R1195 CLK1.n254 CLK1.n130 8.855
R1196 CLK1.n130 CLK1.n129 8.855
R1197 CLK1.n257 CLK1.n256 8.855
R1198 CLK1.n256 CLK1.n255 8.855
R1199 CLK1.n261 CLK1.n260 8.855
R1200 CLK1.n260 CLK1.n259 8.855
R1201 CLK1.n265 CLK1.n264 8.855
R1202 CLK1.n264 CLK1.n263 8.855
R1203 CLK1.n270 CLK1.n269 8.855
R1204 CLK1.n269 CLK1.n268 8.855
R1205 CLK1.n274 CLK1.n273 8.855
R1206 CLK1.n273 CLK1.n272 8.855
R1207 CLK1.n278 CLK1.n277 8.855
R1208 CLK1.n277 CLK1.n276 8.855
R1209 CLK1.n282 CLK1.n281 8.855
R1210 CLK1.n281 CLK1.n280 8.855
R1211 CLK1.n286 CLK1.n285 8.855
R1212 CLK1.n285 CLK1.n284 8.855
R1213 CLK1.n290 CLK1.n289 8.855
R1214 CLK1.n289 CLK1.n288 8.855
R1215 CLK1.n295 CLK1.n294 8.855
R1216 CLK1.n294 CLK1.n293 8.855
R1217 CLK1.n299 CLK1.n298 8.855
R1218 CLK1.n298 CLK1.n297 8.855
R1219 CLK1.n303 CLK1.n302 8.855
R1220 CLK1.n321 CLK1.n320 8.855
R1221 CLK1.n325 CLK1.n324 8.855
R1222 CLK1.n324 CLK1.n323 8.855
R1223 CLK1.n329 CLK1.n328 8.855
R1224 CLK1.n328 CLK1.n327 8.855
R1225 CLK1.n333 CLK1.n332 8.855
R1226 CLK1.n332 CLK1.n331 8.855
R1227 CLK1.n337 CLK1.n336 8.855
R1228 CLK1.n336 CLK1.n335 8.855
R1229 CLK1.n341 CLK1.n340 8.855
R1230 CLK1.n340 CLK1.n339 8.855
R1231 CLK1.n345 CLK1.n344 8.855
R1232 CLK1.n344 CLK1.n343 8.855
R1233 CLK1.n349 CLK1.n348 8.855
R1234 CLK1.n348 CLK1.n347 8.855
R1235 CLK1.n354 CLK1.n353 8.855
R1236 CLK1.n353 CLK1.n352 8.855
R1237 CLK1.n358 CLK1.n357 8.855
R1238 CLK1.n357 CLK1.n356 8.855
R1239 CLK1.n362 CLK1.n361 8.855
R1240 CLK1.n361 CLK1.n360 8.855
R1241 CLK1.n367 CLK1.n366 8.855
R1242 CLK1.n366 CLK1.n365 8.855
R1243 CLK1.n370 CLK1.n369 8.855
R1244 CLK1.n369 CLK1.n368 8.855
R1245 CLK1.n374 CLK1.n373 8.855
R1246 CLK1.n373 CLK1.n372 8.855
R1247 CLK1.n378 CLK1.n377 8.855
R1248 CLK1.n377 CLK1.n376 8.855
R1249 CLK1.n383 CLK1.n382 8.855
R1250 CLK1.n382 CLK1.n381 8.855
R1251 CLK1.n387 CLK1.n386 8.855
R1252 CLK1.n386 CLK1.n385 8.855
R1253 CLK1.n391 CLK1.n390 8.855
R1254 CLK1.n390 CLK1.n389 8.855
R1255 CLK1.n395 CLK1.n394 8.855
R1256 CLK1.n394 CLK1.n393 8.855
R1257 CLK1.n400 CLK1.n399 8.855
R1258 CLK1.n399 CLK1.n398 8.855
R1259 CLK1.n404 CLK1.n403 8.855
R1260 CLK1.n403 CLK1.n402 8.855
R1261 CLK1.n408 CLK1.n407 8.855
R1262 CLK1.n407 CLK1.n406 8.855
R1263 CLK1.n412 CLK1.n411 8.855
R1264 CLK1.n7 CLK1.n6 8.855
R1265 CLK1.n11 CLK1.n10 8.855
R1266 CLK1.n10 CLK1.n9 8.855
R1267 CLK1.n15 CLK1.n14 8.855
R1268 CLK1.n14 CLK1.n13 8.855
R1269 CLK1.n19 CLK1.n18 8.855
R1270 CLK1.n18 CLK1.n17 8.855
R1271 CLK1.n24 CLK1.n23 8.855
R1272 CLK1.n23 CLK1.n22 8.855
R1273 CLK1.n28 CLK1.n27 8.855
R1274 CLK1.n27 CLK1.n26 8.855
R1275 CLK1.n32 CLK1.n31 8.855
R1276 CLK1.n31 CLK1.n30 8.855
R1277 CLK1.n37 CLK1.n36 8.855
R1278 CLK1.n36 CLK1.n35 8.855
R1279 CLK1.n40 CLK1.n39 8.855
R1280 CLK1.n39 CLK1.n38 8.855
R1281 CLK1.n44 CLK1.n43 8.855
R1282 CLK1.n43 CLK1.n42 8.855
R1283 CLK1.n48 CLK1.n47 8.855
R1284 CLK1.n47 CLK1.n46 8.855
R1285 CLK1.n53 CLK1.n52 8.855
R1286 CLK1.n52 CLK1.n51 8.855
R1287 CLK1.n57 CLK1.n56 8.855
R1288 CLK1.n56 CLK1.n55 8.855
R1289 CLK1.n61 CLK1.n60 8.855
R1290 CLK1.n60 CLK1.n59 8.855
R1291 CLK1.n65 CLK1.n64 8.855
R1292 CLK1.n74 CLK1.n73 8.855
R1293 CLK1.n78 CLK1.n77 8.855
R1294 CLK1.n77 CLK1.n76 8.855
R1295 CLK1.n82 CLK1.n81 8.855
R1296 CLK1.n81 CLK1.n80 8.855
R1297 CLK1.n87 CLK1.n86 8.855
R1298 CLK1.n86 CLK1.n85 8.855
R1299 CLK1.n91 CLK1.n90 8.855
R1300 CLK1.n90 CLK1.n89 8.855
R1301 CLK1.n95 CLK1.n94 8.855
R1302 CLK1.n94 CLK1.n93 8.855
R1303 CLK1.n99 CLK1.n98 8.855
R1304 CLK1.n98 CLK1.n97 8.855
R1305 CLK1.n103 CLK1.n102 8.855
R1306 CLK1.n102 CLK1.n101 8.855
R1307 CLK1.n107 CLK1.n106 8.855
R1308 CLK1.n106 CLK1.n105 8.855
R1309 CLK1.n112 CLK1.n111 8.855
R1310 CLK1.n111 CLK1.n110 8.855
R1311 CLK1.n116 CLK1.n115 8.855
R1312 CLK1.n115 CLK1.n114 8.855
R1313 CLK1.n120 CLK1.n119 8.855
R1314 CLK1.n119 CLK1.n118 8.855
R1315 CLK1.n124 CLK1.n123 8.855
R1316 CLK1.n123 CLK1.n122 8.855
R1317 CLK1.n472 CLK1.n471 8.855
R1318 CLK1.n471 CLK1.n470 8.855
R1319 CLK1.n468 CLK1.n467 8.855
R1320 CLK1.n467 CLK1.n466 8.855
R1321 CLK1.n464 CLK1.n463 8.855
R1322 CLK1.n463 CLK1.n462 8.855
R1323 CLK1.n459 CLK1.n458 8.855
R1324 CLK1.n458 CLK1.n457 8.855
R1325 CLK1.n455 CLK1.n454 8.855
R1326 CLK1.n454 CLK1.n453 8.855
R1327 CLK1.n451 CLK1.n450 8.855
R1328 CLK1.n450 CLK1.n449 8.855
R1329 CLK1.n447 CLK1.n446 8.855
R1330 CLK1.n446 CLK1.n445 8.855
R1331 CLK1.n443 CLK1.n442 8.855
R1332 CLK1.n442 CLK1.n441 8.855
R1333 CLK1.n439 CLK1.n438 8.855
R1334 CLK1.n438 CLK1.n437 8.855
R1335 CLK1.n434 CLK1.n433 8.855
R1336 CLK1.n433 CLK1.n432 8.855
R1337 CLK1.n430 CLK1.n429 8.855
R1338 CLK1.n429 CLK1.n428 8.855
R1339 CLK1.n426 CLK1.n425 8.855
R1340 CLK1.n249 CLK1.t46 8.189
R1341 CLK1.n255 CLK1.t31 8.189
R1342 CLK1.n163 CLK1.t44 8.189
R1343 CLK1.n169 CLK1.t37 8.189
R1344 CLK1.n360 CLK1.t15 8.189
R1345 CLK1.n368 CLK1.t24 8.189
R1346 CLK1.n118 CLK1.t21 8.189
R1347 CLK1.n470 CLK1.t52 8.189
R1348 CLK1.n30 CLK1.t7 8.189
R1349 CLK1.n38 CLK1.t17 8.189
R1350 CLK1.n292 CLK1.n128 6.776
R1351 CLK1.n215 CLK1.n132 6.776
R1352 CLK1.n397 CLK1.n315 6.776
R1353 CLK1.n84 CLK1.n1 6.776
R1354 CLK1.n436 CLK1.n126 6.776
R1355 CLK1.n253 CLK1.n131 4.938
R1356 CLK1.n167 CLK1.n135 4.938
R1357 CLK1.n364 CLK1.n316 4.938
R1358 CLK1.n125 CLK1.n0 4.938
R1359 CLK1.n34 CLK1.n2 4.938
R1360 CLK1.n318 CLK1.n317 4.687
R1361 CLK1.n137 CLK1.n136 4.662
R1362 CLK1.n4 CLK1.n3 4.662
R1363 CLK1.n141 CLK1.n140 4.65
R1364 CLK1.n145 CLK1.n144 4.65
R1365 CLK1.n149 CLK1.n148 4.65
R1366 CLK1.n153 CLK1.n152 4.65
R1367 CLK1.n158 CLK1.n157 4.65
R1368 CLK1.n162 CLK1.n161 4.65
R1369 CLK1.n166 CLK1.n165 4.65
R1370 CLK1.n168 CLK1.n167 4.65
R1371 CLK1.n172 CLK1.n171 4.65
R1372 CLK1.n176 CLK1.n175 4.65
R1373 CLK1.n180 CLK1.n179 4.65
R1374 CLK1.n185 CLK1.n184 4.65
R1375 CLK1.n189 CLK1.n188 4.65
R1376 CLK1.n193 CLK1.n192 4.65
R1377 CLK1.n197 CLK1.n196 4.65
R1378 CLK1.n200 CLK1.n199 4.65
R1379 CLK1.n202 CLK1.n201 4.65
R1380 CLK1.n206 CLK1.n205 4.65
R1381 CLK1.n210 CLK1.n209 4.65
R1382 CLK1.n214 CLK1.n213 4.65
R1383 CLK1.n219 CLK1.n218 4.65
R1384 CLK1.n223 CLK1.n222 4.65
R1385 CLK1.n227 CLK1.n226 4.65
R1386 CLK1.n231 CLK1.n230 4.65
R1387 CLK1.n235 CLK1.n234 4.65
R1388 CLK1.n239 CLK1.n238 4.65
R1389 CLK1.n244 CLK1.n243 4.65
R1390 CLK1.n248 CLK1.n247 4.65
R1391 CLK1.n252 CLK1.n251 4.65
R1392 CLK1.n254 CLK1.n253 4.65
R1393 CLK1.n258 CLK1.n257 4.65
R1394 CLK1.n262 CLK1.n261 4.65
R1395 CLK1.n266 CLK1.n265 4.65
R1396 CLK1.n271 CLK1.n270 4.65
R1397 CLK1.n275 CLK1.n274 4.65
R1398 CLK1.n279 CLK1.n278 4.65
R1399 CLK1.n283 CLK1.n282 4.65
R1400 CLK1.n287 CLK1.n286 4.65
R1401 CLK1.n291 CLK1.n290 4.65
R1402 CLK1.n296 CLK1.n295 4.65
R1403 CLK1.n300 CLK1.n299 4.65
R1404 CLK1.n304 CLK1.n303 4.65
R1405 CLK1.n322 CLK1.n321 4.65
R1406 CLK1.n326 CLK1.n325 4.65
R1407 CLK1.n330 CLK1.n329 4.65
R1408 CLK1.n334 CLK1.n333 4.65
R1409 CLK1.n338 CLK1.n337 4.65
R1410 CLK1.n342 CLK1.n341 4.65
R1411 CLK1.n346 CLK1.n345 4.65
R1412 CLK1.n350 CLK1.n349 4.65
R1413 CLK1.n355 CLK1.n354 4.65
R1414 CLK1.n359 CLK1.n358 4.65
R1415 CLK1.n363 CLK1.n362 4.65
R1416 CLK1.n367 CLK1.n364 4.65
R1417 CLK1.n371 CLK1.n370 4.65
R1418 CLK1.n375 CLK1.n374 4.65
R1419 CLK1.n379 CLK1.n378 4.65
R1420 CLK1.n384 CLK1.n383 4.65
R1421 CLK1.n388 CLK1.n387 4.65
R1422 CLK1.n392 CLK1.n391 4.65
R1423 CLK1.n396 CLK1.n395 4.65
R1424 CLK1.n401 CLK1.n400 4.65
R1425 CLK1.n405 CLK1.n404 4.65
R1426 CLK1.n409 CLK1.n408 4.65
R1427 CLK1.n413 CLK1.n412 4.65
R1428 CLK1.n416 CLK1.n415 4.65
R1429 CLK1.n8 CLK1.n7 4.65
R1430 CLK1.n12 CLK1.n11 4.65
R1431 CLK1.n16 CLK1.n15 4.65
R1432 CLK1.n20 CLK1.n19 4.65
R1433 CLK1.n25 CLK1.n24 4.65
R1434 CLK1.n29 CLK1.n28 4.65
R1435 CLK1.n33 CLK1.n32 4.65
R1436 CLK1.n37 CLK1.n34 4.65
R1437 CLK1.n41 CLK1.n40 4.65
R1438 CLK1.n45 CLK1.n44 4.65
R1439 CLK1.n49 CLK1.n48 4.65
R1440 CLK1.n54 CLK1.n53 4.65
R1441 CLK1.n58 CLK1.n57 4.65
R1442 CLK1.n62 CLK1.n61 4.65
R1443 CLK1.n66 CLK1.n65 4.65
R1444 CLK1.n69 CLK1.n68 4.65
R1445 CLK1.n71 CLK1.n70 4.65
R1446 CLK1.n75 CLK1.n74 4.65
R1447 CLK1.n79 CLK1.n78 4.65
R1448 CLK1.n83 CLK1.n82 4.65
R1449 CLK1.n88 CLK1.n87 4.65
R1450 CLK1.n92 CLK1.n91 4.65
R1451 CLK1.n96 CLK1.n95 4.65
R1452 CLK1.n100 CLK1.n99 4.65
R1453 CLK1.n104 CLK1.n103 4.65
R1454 CLK1.n108 CLK1.n107 4.65
R1455 CLK1.n113 CLK1.n112 4.65
R1456 CLK1.n117 CLK1.n116 4.65
R1457 CLK1.n121 CLK1.n120 4.65
R1458 CLK1.n125 CLK1.n124 4.65
R1459 CLK1.n473 CLK1.n472 4.65
R1460 CLK1.n469 CLK1.n468 4.65
R1461 CLK1.n465 CLK1.n464 4.65
R1462 CLK1.n460 CLK1.n459 4.65
R1463 CLK1.n456 CLK1.n455 4.65
R1464 CLK1.n452 CLK1.n451 4.65
R1465 CLK1.n448 CLK1.n447 4.65
R1466 CLK1.n444 CLK1.n443 4.65
R1467 CLK1.n440 CLK1.n439 4.65
R1468 CLK1.n435 CLK1.n434 4.65
R1469 CLK1.n431 CLK1.n430 4.65
R1470 CLK1.n427 CLK1.n426 4.65
R1471 CLK1.n313 CLK1.n312 3.635
R1472 CLK1.n308 CLK1.n307 3.563
R1473 CLK1.n422 CLK1.n421 3.563
R1474 CLK1.n417 CLK1.n416 3.067
R1475 CLK1.n314 CLK1.n313 2.245
R1476 CLK1.n419 CLK1.n418 2.245
R1477 CLK1.n139 CLK1.n138 1.655
R1478 CLK1.n204 CLK1.n203 1.655
R1479 CLK1.n320 CLK1.n319 1.655
R1480 CLK1.n6 CLK1.n5 1.655
R1481 CLK1.n73 CLK1.n72 1.655
R1482 CLK1.n195 CLK1.n194 1.655
R1483 CLK1.n302 CLK1.n301 1.655
R1484 CLK1.n411 CLK1.n410 1.655
R1485 CLK1.n64 CLK1.n63 1.655
R1486 CLK1.n425 CLK1.n424 1.655
R1487 CLK1.n311 CLK1.n310 1.498
R1488 CLK1.n307 CLK1.n306 1.44
R1489 CLK1.n421 CLK1.n420 1.44
R1490 CLK1.n202 CLK1.n200 0.637
R1491 CLK1.n71 CLK1.n69 0.637
R1492 CLK1.n127 CLK1 0.125
R1493 CLK1.n145 CLK1.n141 0.1
R1494 CLK1.n149 CLK1.n145 0.1
R1495 CLK1.n153 CLK1.n149 0.1
R1496 CLK1.n162 CLK1.n158 0.1
R1497 CLK1.n166 CLK1.n162 0.1
R1498 CLK1.n167 CLK1.n166 0.1
R1499 CLK1.n176 CLK1.n172 0.1
R1500 CLK1.n180 CLK1.n176 0.1
R1501 CLK1.n189 CLK1.n185 0.1
R1502 CLK1.n193 CLK1.n189 0.1
R1503 CLK1.n197 CLK1.n193 0.1
R1504 CLK1.n206 CLK1.n202 0.1
R1505 CLK1.n210 CLK1.n206 0.1
R1506 CLK1.n214 CLK1.n210 0.1
R1507 CLK1.n223 CLK1.n219 0.1
R1508 CLK1.n227 CLK1.n223 0.1
R1509 CLK1.n231 CLK1.n227 0.1
R1510 CLK1.n235 CLK1.n231 0.1
R1511 CLK1.n239 CLK1.n235 0.1
R1512 CLK1.n248 CLK1.n244 0.1
R1513 CLK1.n252 CLK1.n248 0.1
R1514 CLK1.n253 CLK1.n252 0.1
R1515 CLK1.n262 CLK1.n258 0.1
R1516 CLK1.n266 CLK1.n262 0.1
R1517 CLK1.n275 CLK1.n271 0.1
R1518 CLK1.n279 CLK1.n275 0.1
R1519 CLK1.n283 CLK1.n279 0.1
R1520 CLK1.n287 CLK1.n283 0.1
R1521 CLK1.n291 CLK1.n287 0.1
R1522 CLK1.n300 CLK1.n296 0.1
R1523 CLK1.n304 CLK1.n300 0.1
R1524 CLK1.n326 CLK1.n322 0.1
R1525 CLK1.n330 CLK1.n326 0.1
R1526 CLK1.n334 CLK1.n330 0.1
R1527 CLK1.n338 CLK1.n334 0.1
R1528 CLK1.n342 CLK1.n338 0.1
R1529 CLK1.n346 CLK1.n342 0.1
R1530 CLK1.n350 CLK1.n346 0.1
R1531 CLK1.n359 CLK1.n355 0.1
R1532 CLK1.n363 CLK1.n359 0.1
R1533 CLK1.n364 CLK1.n363 0.1
R1534 CLK1.n375 CLK1.n371 0.1
R1535 CLK1.n379 CLK1.n375 0.1
R1536 CLK1.n388 CLK1.n384 0.1
R1537 CLK1.n392 CLK1.n388 0.1
R1538 CLK1.n396 CLK1.n392 0.1
R1539 CLK1.n405 CLK1.n401 0.1
R1540 CLK1.n409 CLK1.n405 0.1
R1541 CLK1.n413 CLK1.n409 0.1
R1542 CLK1.n12 CLK1.n8 0.1
R1543 CLK1.n16 CLK1.n12 0.1
R1544 CLK1.n20 CLK1.n16 0.1
R1545 CLK1.n29 CLK1.n25 0.1
R1546 CLK1.n33 CLK1.n29 0.1
R1547 CLK1.n34 CLK1.n33 0.1
R1548 CLK1.n45 CLK1.n41 0.1
R1549 CLK1.n49 CLK1.n45 0.1
R1550 CLK1.n58 CLK1.n54 0.1
R1551 CLK1.n62 CLK1.n58 0.1
R1552 CLK1.n66 CLK1.n62 0.1
R1553 CLK1.n75 CLK1.n71 0.1
R1554 CLK1.n79 CLK1.n75 0.1
R1555 CLK1.n83 CLK1.n79 0.1
R1556 CLK1.n92 CLK1.n88 0.1
R1557 CLK1.n96 CLK1.n92 0.1
R1558 CLK1.n100 CLK1.n96 0.1
R1559 CLK1.n104 CLK1.n100 0.1
R1560 CLK1.n108 CLK1.n104 0.1
R1561 CLK1.n117 CLK1.n113 0.1
R1562 CLK1.n121 CLK1.n117 0.1
R1563 CLK1.n125 CLK1.n121 0.1
R1564 CLK1.n473 CLK1.n469 0.1
R1565 CLK1.n469 CLK1.n465 0.1
R1566 CLK1.n460 CLK1.n456 0.1
R1567 CLK1.n456 CLK1.n452 0.1
R1568 CLK1.n452 CLK1.n448 0.1
R1569 CLK1.n448 CLK1.n444 0.1
R1570 CLK1.n444 CLK1.n440 0.1
R1571 CLK1.n435 CLK1.n431 0.1
R1572 CLK1.n431 CLK1.n427 0.1
R1573 CLK1.n305 CLK1.n304 0.088
R1574 CLK1.n427 CLK1.n423 0.088
R1575 CLK1.n141 CLK1.n137 0.087
R1576 CLK1.n198 CLK1.n197 0.087
R1577 CLK1.n397 CLK1.n396 0.087
R1578 CLK1.n8 CLK1.n4 0.087
R1579 CLK1.n67 CLK1.n66 0.087
R1580 CLK1.n158 CLK1.n154 0.075
R1581 CLK1.n172 CLK1 0.075
R1582 CLK1.n181 CLK1.n180 0.075
R1583 CLK1.n219 CLK1.n215 0.075
R1584 CLK1.n244 CLK1.n240 0.075
R1585 CLK1.n258 EESPFAL_XOR_v3_0/CLK 0.075
R1586 CLK1.n267 CLK1.n266 0.075
R1587 CLK1.n292 CLK1.n291 0.075
R1588 CLK1.n355 CLK1.n351 0.075
R1589 CLK1.n371 EESPFAL_3in_NAND_v2_0/CLK 0.075
R1590 CLK1.n380 CLK1.n379 0.075
R1591 CLK1.n25 CLK1.n21 0.075
R1592 CLK1.n41 EESPFAL_INV4_1/CLK 0.075
R1593 CLK1.n50 CLK1.n49 0.075
R1594 CLK1.n88 CLK1.n84 0.075
R1595 CLK1.n113 CLK1.n109 0.075
R1596 EESPFAL_XOR_v3_1/CLK CLK1.n473 0.075
R1597 CLK1.n465 CLK1.n461 0.075
R1598 CLK1.n440 CLK1.n436 0.075
R1599 CLK1.n322 CLK1.n318 0.062
R1600 CLK1.n414 CLK1.n413 0.062
R1601 CLK1.n416 CLK1.n414 0.037
R1602 CLK1.n418 CLK1.n417 0.034
R1603 CLK1.n312 CLK1.n311 0.033
R1604 CLK1.n311 CLK1.n127 0.032
R1605 CLK1.n154 CLK1.n153 0.025
R1606 CLK1.n167 CLK1 0.025
R1607 CLK1.n185 CLK1.n181 0.025
R1608 CLK1.n215 CLK1.n214 0.025
R1609 CLK1.n240 CLK1.n239 0.025
R1610 CLK1.n253 EESPFAL_XOR_v3_0/CLK 0.025
R1611 CLK1.n271 CLK1.n267 0.025
R1612 CLK1.n296 CLK1.n292 0.025
R1613 CLK1.n351 CLK1.n350 0.025
R1614 CLK1.n364 EESPFAL_3in_NAND_v2_0/CLK 0.025
R1615 CLK1.n384 CLK1.n380 0.025
R1616 CLK1.n21 CLK1.n20 0.025
R1617 CLK1.n34 EESPFAL_INV4_1/CLK 0.025
R1618 CLK1.n54 CLK1.n50 0.025
R1619 CLK1.n84 CLK1.n83 0.025
R1620 CLK1.n109 CLK1.n108 0.025
R1621 EESPFAL_XOR_v3_1/CLK CLK1.n125 0.025
R1622 CLK1.n461 CLK1.n460 0.025
R1623 CLK1.n436 CLK1.n435 0.025
R1624 CLK1.n310 CLK1.n308 0.019
R1625 CLK1.n308 CLK1.n305 0.018
R1626 CLK1.n423 CLK1.n422 0.018
R1627 CLK1.n422 CLK1.n419 0.015
R1628 CLK1.n200 CLK1.n198 0.012
R1629 CLK1.n401 CLK1.n397 0.012
R1630 CLK1.n69 CLK1.n67 0.012
R1631 CLK1.n419 CLK1.n314 0.011
R1632 CLK1.n310 CLK1.n309 0.007
R1633 EESPFAL_NAND_v3_0/A_bar.t7 EESPFAL_NAND_v3_0/A_bar.t9 819.4
R1634 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/A_bar.t8 736.033
R1635 EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_NAND_v3_0/A_bar.t7 514.133
R1636 EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_NAND_v3_0/A_bar.t6 305.266
R1637 EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_NAND_v3_0/A_bar.n5 192
R1638 EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_NAND_v3_0/A_bar.n0 166.734
R1639 EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_NAND_v3_0/A_bar.n4 105.6
R1640 EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_NAND_v3_0/A_bar.t0 97.939
R1641 EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_NAND_v3_0/A_bar.t1 97.937
R1642 EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_NAND_v3_0/A_bar.n2 76
R1643 EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_NAND_v3_0/A_bar.n1 73.937
R1644 EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_NAND_v3_0/A_bar.n3 57.6
R1645 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/A_bar.n6 56.157
R1646 EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_NAND_v3_0/A_bar.t2 39.4
R1647 EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_NAND_v3_0/A_bar.t4 39.4
R1648 EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_NAND_v3_0/A_bar.t5 24
R1649 EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_NAND_v3_0/A_bar.t3 24
R1650 EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_XOR_v3_0/OUT 3.2
R1651 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/A.t9 1074.82
R1652 EESPFAL_NAND_v3_0/A.t8 EESPFAL_NAND_v3_0/A.t6 819.4
R1653 EESPFAL_NAND_v3_0/A.n5 EESPFAL_NAND_v3_0/A.t7 506.1
R1654 EESPFAL_XOR_v3_0/OUT_bar EESPFAL_NAND_v3_0/A 442.013
R1655 EESPFAL_NAND_v3_0/A.n5 EESPFAL_NAND_v3_0/A.t8 313.3
R1656 EESPFAL_NAND_v3_0/A.n1 EESPFAL_NAND_v3_0/A.t0 273.936
R1657 EESPFAL_NAND_v3_0/A.n4 EESPFAL_NAND_v3_0/A.n3 128.335
R1658 EESPFAL_NAND_v3_0/A.n2 EESPFAL_NAND_v3_0/A.n1 105.6
R1659 EESPFAL_NAND_v3_0/A.n1 EESPFAL_NAND_v3_0/A.t5 81.937
R1660 EESPFAL_NAND_v3_0/A.n2 EESPFAL_NAND_v3_0/A.n0 57.937
R1661 EESPFAL_NAND_v3_0/A.n6 EESPFAL_NAND_v3_0/A.n4 57.6
R1662 EESPFAL_NAND_v3_0/A.n4 EESPFAL_NAND_v3_0/A.n2 41.6
R1663 EESPFAL_NAND_v3_0/A.n3 EESPFAL_NAND_v3_0/A.t4 39.4
R1664 EESPFAL_NAND_v3_0/A.n3 EESPFAL_NAND_v3_0/A.t3 39.4
R1665 EESPFAL_NAND_v3_0/A.n0 EESPFAL_NAND_v3_0/A.t2 24
R1666 EESPFAL_NAND_v3_0/A.n0 EESPFAL_NAND_v3_0/A.t1 24
R1667 EESPFAL_NAND_v3_0/A.n6 EESPFAL_NAND_v3_0/A.n5 8.764
R1668 EESPFAL_XOR_v3_0/OUT_bar EESPFAL_NAND_v3_0/A.n6 4.65
R1669 Dis1.n5 Dis1 556.8
R1670 Dis1.n2 EESPFAL_INV4_1/Dis 556.8
R1671 Dis1.n4 Dis1.t9 504.5
R1672 Dis1.n1 Dis1.t3 504.5
R1673 Dis1.n0 Dis1.t1 504.5
R1674 Dis1.n6 Dis1.t4 389.3
R1675 Dis1.n5 Dis1.t7 389.3
R1676 Dis1.n4 Dis1.t6 389.3
R1677 Dis1.n3 Dis1.t2 389.3
R1678 Dis1.n2 Dis1.t8 389.3
R1679 Dis1.n1 Dis1.t0 389.3
R1680 Dis1.n0 Dis1.t5 389.3
R1681 EESPFAL_3in_NAND_v2_0/Dis Dis1.n8 235.714
R1682 Dis1.n7 EESPFAL_XOR_v3_0/Dis 227.457
R1683 Dis1.n8 EESPFAL_XOR_v3_1/Dis 227.456
R1684 Dis1.n6 Dis1.n5 115.2
R1685 Dis1.n3 Dis1.n2 115.2
R1686 Dis1.n7 Dis1 3.587
R1687 Dis1 Dis1.n4 3.2
R1688 EESPFAL_XOR_v3_0/Dis Dis1.n6 3.2
R1689 EESPFAL_INV4_1/Dis Dis1.n1 3.2
R1690 EESPFAL_XOR_v3_1/Dis Dis1.n3 3.2
R1691 EESPFAL_3in_NAND_v2_0/Dis Dis1.n0 3.2
R1692 Dis1.n8 Dis1.n7 0.625
R1693 Dis2.n4 Dis2.n3 532.126
R1694 Dis2.n1 Dis2.t0 504.5
R1695 Dis2.n0 Dis2.t1 504.5
R1696 Dis2.n1 Dis2.t3 389.3
R1697 Dis2.n0 Dis2.t4 389.3
R1698 Dis2.n4 Dis2.t2 389.3
R1699 Dis2.n5 Dis2.t5 389.3
R1700 Dis2.n2 Dis2 177.217
R1701 Dis2.n3 EESPFAL_NAND_v3_1/Dis 177.216
R1702 Dis2.n5 Dis2.n4 115.2
R1703 Dis2.n2 Dis2 3.605
R1704 Dis2 Dis2.n1 3.2
R1705 EESPFAL_NAND_v3_1/Dis Dis2.n0 3.2
R1706 EESPFAL_INV4_0/Dis Dis2.n5 3.2
R1707 Dis2.n3 Dis2.n2 0.621
R1708 EESPFAL_NAND_v3_1/A_bar.t9 EESPFAL_NAND_v3_1/A_bar.t6 819.4
R1709 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/A_bar.t8 736.033
R1710 EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_NAND_v3_1/A_bar.t7 506.1
R1711 EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_NAND_v3_1/A_bar.t9 313.3
R1712 EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_NAND_v3_1/A_bar.t1 273.937
R1713 EESPFAL_XOR_v3_1/OUT_bar EESPFAL_NAND_v3_1/A_bar 266.318
R1714 EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_NAND_v3_1/A_bar.n0 128.334
R1715 EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_NAND_v3_1/A_bar.n2 105.6
R1716 EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_NAND_v3_1/A_bar.t3 81.937
R1717 EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_NAND_v3_1/A_bar.n1 57.937
R1718 EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_NAND_v3_1/A_bar.n4 57.6
R1719 EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_NAND_v3_1/A_bar.n3 41.6
R1720 EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_NAND_v3_1/A_bar.t5 39.4
R1721 EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_NAND_v3_1/A_bar.t0 39.4
R1722 EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_NAND_v3_1/A_bar.t2 24
R1723 EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_NAND_v3_1/A_bar.t4 24
R1724 EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_NAND_v3_1/A_bar.n5 8.764
R1725 EESPFAL_XOR_v3_1/OUT_bar EESPFAL_NAND_v3_1/A_bar.n6 4.65
R1726 EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/A.t8 1074.82
R1727 EESPFAL_NAND_v3_1/A.t9 EESPFAL_NAND_v3_1/A.t7 819.4
R1728 EESPFAL_NAND_v3_1/A.n1 EESPFAL_NAND_v3_1/A.t9 514.133
R1729 EESPFAL_NAND_v3_1/A.n1 EESPFAL_NAND_v3_1/A.t6 305.266
R1730 EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/A.n6 260.333
R1731 EESPFAL_NAND_v3_1/A.n6 EESPFAL_NAND_v3_1/A.n5 192
R1732 EESPFAL_NAND_v3_1/A.n4 EESPFAL_NAND_v3_1/A.n3 166.736
R1733 EESPFAL_NAND_v3_1/A.n5 EESPFAL_NAND_v3_1/A.n4 105.6
R1734 EESPFAL_NAND_v3_1/A.n6 EESPFAL_NAND_v3_1/A.t3 97.937
R1735 EESPFAL_NAND_v3_1/A.n5 EESPFAL_NAND_v3_1/A.t4 97.937
R1736 EESPFAL_NAND_v3_1/A.n2 EESPFAL_NAND_v3_1/A.n1 76
R1737 EESPFAL_NAND_v3_1/A.n4 EESPFAL_NAND_v3_1/A.n0 73.937
R1738 EESPFAL_NAND_v3_1/A.n4 EESPFAL_NAND_v3_1/A.n2 57.6
R1739 EESPFAL_NAND_v3_1/A.n3 EESPFAL_NAND_v3_1/A.t2 39.4
R1740 EESPFAL_NAND_v3_1/A.n3 EESPFAL_NAND_v3_1/A.t1 39.4
R1741 EESPFAL_NAND_v3_1/A.n0 EESPFAL_NAND_v3_1/A.t5 24
R1742 EESPFAL_NAND_v3_1/A.n0 EESPFAL_NAND_v3_1/A.t0 24
R1743 EESPFAL_NAND_v3_1/A.n2 EESPFAL_XOR_v3_1/OUT 3.2
R1744 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_3in_NOR_v2_0/A_bar 922.56
R1745 EESPFAL_NAND_v3_0/OUT_bar.t8 EESPFAL_NAND_v3_0/OUT_bar.t9 819.4
R1746 EESPFAL_3in_NOR_v2_0/A_bar EESPFAL_NAND_v3_0/OUT_bar.t6 684.833
R1747 EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_NAND_v3_0/OUT_bar.t7 506.1
R1748 EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_NAND_v3_0/OUT_bar.t8 313.3
R1749 EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_NAND_v3_0/OUT_bar.t4 177.936
R1750 EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_NAND_v3_0/OUT_bar.n3 128.335
R1751 EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_NAND_v3_0/OUT_bar.n1 105.6
R1752 EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_NAND_v3_0/OUT_bar.t5 81.937
R1753 EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_NAND_v3_0/OUT_bar.n0 58.265
R1754 EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_NAND_v3_0/OUT_bar.n4 57.6
R1755 EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_NAND_v3_0/OUT_bar.n2 41.6
R1756 EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_NAND_v3_0/OUT_bar.t2 39.4
R1757 EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_NAND_v3_0/OUT_bar.t3 39.4
R1758 EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_NAND_v3_0/OUT_bar.t1 24
R1759 EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_NAND_v3_0/OUT_bar.t0 24
R1760 EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_NAND_v3_0/OUT_bar.n5 8.764
R1761 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_NAND_v3_0/OUT_bar.n6 4.65
R1762 CLK3.n89 CLK3.t6 44.337
R1763 CLK3.n35 CLK3.t1 44.337
R1764 CLK3.n0 CLK3.t3 39.4
R1765 CLK3.n0 CLK3.t11 39.4
R1766 CLK3.n55 CLK3.t8 30.775
R1767 CLK3.n2 CLK3.t4 30.775
R1768 CLK3.n36 CLK3.t0 24.568
R1769 CLK3.n90 CLK3.t5 24.568
R1770 CLK3.n52 CLK3.t9 24
R1771 CLK3.n52 CLK3.t7 24
R1772 CLK3.n54 CLK3 9.841
R1773 CLK3.n5 CLK3.n4 8.855
R1774 CLK3.n9 CLK3.n8 8.855
R1775 CLK3.n8 CLK3.n7 8.855
R1776 CLK3.n13 CLK3.n12 8.855
R1777 CLK3.n12 CLK3.n11 8.855
R1778 CLK3.n17 CLK3.n16 8.855
R1779 CLK3.n16 CLK3.n15 8.855
R1780 CLK3.n21 CLK3.n20 8.855
R1781 CLK3.n20 CLK3.n19 8.855
R1782 CLK3.n25 CLK3.n24 8.855
R1783 CLK3.n24 CLK3.n23 8.855
R1784 CLK3.n29 CLK3.n28 8.855
R1785 CLK3.n28 CLK3.n27 8.855
R1786 CLK3.n33 CLK3.n32 8.855
R1787 CLK3.n32 CLK3.n31 8.855
R1788 CLK3.n38 CLK3.n37 8.855
R1789 CLK3.n37 CLK3.n36 8.855
R1790 CLK3.n42 CLK3.n41 8.855
R1791 CLK3.n41 CLK3.n40 8.855
R1792 CLK3.n46 CLK3.n45 8.855
R1793 CLK3.n45 CLK3.n44 8.855
R1794 CLK3.n50 CLK3.n49 8.855
R1795 CLK3.n49 CLK3.n48 8.855
R1796 CLK3.n100 CLK3.n99 8.855
R1797 CLK3.n99 CLK3.n98 8.855
R1798 CLK3.n96 CLK3.n95 8.855
R1799 CLK3.n95 CLK3.n94 8.855
R1800 CLK3.n92 CLK3.n91 8.855
R1801 CLK3.n91 CLK3.n90 8.855
R1802 CLK3.n87 CLK3.n86 8.855
R1803 CLK3.n86 CLK3.n85 8.855
R1804 CLK3.n83 CLK3.n82 8.855
R1805 CLK3.n82 CLK3.n81 8.855
R1806 CLK3.n79 CLK3.n78 8.855
R1807 CLK3.n78 CLK3.n77 8.855
R1808 CLK3.n75 CLK3.n74 8.855
R1809 CLK3.n74 CLK3.n73 8.855
R1810 CLK3.n70 CLK3.n69 8.855
R1811 CLK3.n69 CLK3.n68 8.855
R1812 CLK3.n66 CLK3.n65 8.855
R1813 CLK3.n65 CLK3.n64 8.855
R1814 CLK3.n62 CLK3.n61 8.855
R1815 CLK3.n61 CLK3.n60 8.855
R1816 CLK3.n58 CLK3.n57 8.855
R1817 CLK3.n44 CLK3.t2 8.189
R1818 CLK3.n98 CLK3.t10 8.189
R1819 CLK3.n72 CLK3.n52 6.776
R1820 CLK3.n51 CLK3.n0 4.938
R1821 CLK3.n2 CLK3.n1 4.687
R1822 CLK3.n6 CLK3.n5 4.65
R1823 CLK3.n10 CLK3.n9 4.65
R1824 CLK3.n14 CLK3.n13 4.65
R1825 CLK3.n18 CLK3.n17 4.65
R1826 CLK3.n22 CLK3.n21 4.65
R1827 CLK3.n26 CLK3.n25 4.65
R1828 CLK3.n30 CLK3.n29 4.65
R1829 CLK3.n34 CLK3.n33 4.65
R1830 CLK3.n39 CLK3.n38 4.65
R1831 CLK3.n43 CLK3.n42 4.65
R1832 CLK3.n47 CLK3.n46 4.65
R1833 CLK3.n51 CLK3.n50 4.65
R1834 CLK3.n101 CLK3.n100 4.65
R1835 CLK3.n97 CLK3.n96 4.65
R1836 CLK3.n93 CLK3.n92 4.65
R1837 CLK3.n88 CLK3.n87 4.65
R1838 CLK3.n84 CLK3.n83 4.65
R1839 CLK3.n80 CLK3.n79 4.65
R1840 CLK3.n76 CLK3.n75 4.65
R1841 CLK3.n71 CLK3.n70 4.65
R1842 CLK3.n67 CLK3.n66 4.65
R1843 CLK3.n63 CLK3.n62 4.65
R1844 CLK3.n59 CLK3.n58 4.65
R1845 CLK3.n54 CLK3.n53 3.038
R1846 CLK3.n4 CLK3.n3 1.655
R1847 CLK3.n57 CLK3.n56 1.655
R1848 CLK3.n10 CLK3.n6 0.1
R1849 CLK3.n14 CLK3.n10 0.1
R1850 CLK3.n18 CLK3.n14 0.1
R1851 CLK3.n22 CLK3.n18 0.1
R1852 CLK3.n26 CLK3.n22 0.1
R1853 CLK3.n30 CLK3.n26 0.1
R1854 CLK3.n34 CLK3.n30 0.1
R1855 CLK3.n43 CLK3.n39 0.1
R1856 CLK3.n47 CLK3.n43 0.1
R1857 CLK3.n51 CLK3.n47 0.1
R1858 CLK3.n101 CLK3.n97 0.1
R1859 CLK3.n97 CLK3.n93 0.1
R1860 CLK3.n88 CLK3.n84 0.1
R1861 CLK3.n84 CLK3.n80 0.1
R1862 CLK3.n80 CLK3.n76 0.1
R1863 CLK3.n71 CLK3.n67 0.1
R1864 CLK3.n67 CLK3.n63 0.1
R1865 CLK3.n63 CLK3.n59 0.1
R1866 CLK3.n76 CLK3.n72 0.087
R1867 CLK3.n39 CLK3.n35 0.075
R1868 CLK3 CLK3.n101 0.075
R1869 CLK3.n93 CLK3.n89 0.075
R1870 CLK3.n6 CLK3.n2 0.062
R1871 CLK3.n59 CLK3.n55 0.062
R1872 CLK3.n55 CLK3.n54 0.034
R1873 CLK3.n35 CLK3.n34 0.025
R1874 CLK3 CLK3.n51 0.025
R1875 CLK3.n89 CLK3.n88 0.025
R1876 CLK3.n72 CLK3.n71 0.012
R1877 x3.n0 x3.t3 800.452
R1878 x3.n0 x3.t0 787.997
R1879 x3 x3.t2 778.1
R1880 EESPFAL_3in_NAND_v2_0/A_bar x3.t1 696.166
R1881 EESPFAL_XOR_v3_1/B x3.n0 169.6
R1882 x3.n1 EESPFAL_3in_NAND_v2_0/A_bar 146.405
R1883 EESPFAL_XOR_v3_1/B x3.n1 96.17
R1884 x3.n1 x3 2.854
R1885 x1.n0 x1.t0 1176.57
R1886 x1.n0 x1.t2 1149.49
R1887 EESPFAL_3in_NAND_v2_0/B x1.t1 1106.75
R1888 EESPFAL_3in_NAND_v2_0/B x1.n1 291.644
R1889 x1.n1 x1 242.09
R1890 x1 x1.n0 128
R1891 x1.n1 x1 3.228
R1892 x1_bar.n0 x1_bar.t0 1069.04
R1893 x1_bar.n0 x1_bar.t1 1015.9
R1894 EESPFAL_3in_NAND_v2_0/B_bar x1_bar.t2 604.112
R1895 EESPFAL_3in_NAND_v2_0/B_bar x1_bar.n1 255.773
R1896 x1_bar.n1 x1_bar 205.61
R1897 x1_bar x1_bar.n0 89.6
R1898 x1_bar.n1 x1_bar 2.945
R1899 EESPFAL_3in_NOR_v2_0/C.t5 EESPFAL_3in_NOR_v2_0/C.t6 819.4
R1900 EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_3in_NOR_v2_0/C.t7 775.706
R1901 EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_3in_NOR_v2_0/C.t5 514.133
R1902 EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_3in_NOR_v2_0/C.t8 305.266
R1903 EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_3in_NOR_v2_0/C.n0 166.734
R1904 EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_3in_NOR_v2_0/C 163.511
R1905 EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_3in_NOR_v2_0/C.n2 102.4
R1906 EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_3in_NOR_v2_0/C.n1 88.255
R1907 EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_3in_NOR_v2_0/C.t1 81.937
R1908 EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_3in_NOR_v2_0/C.n6 76
R1909 EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_3in_NOR_v2_0/C.n5 57.6
R1910 EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_3in_NOR_v2_0/C.n3 51.539
R1911 EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_3in_NOR_v2_0/C.t3 39.4
R1912 EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_3in_NOR_v2_0/C.t2 39.4
R1913 EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_3in_NOR_v2_0/C.t0 24
R1914 EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_3in_NOR_v2_0/C.t4 24
R1915 EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_3in_NOR_v2_0/C.n4 6.4
R1916 EESPFAL_INV4_0/OUT_bar EESPFAL_3in_NOR_v2_0/C.n7 3.2
R1917 Dis3 Dis3.t0 392.5
R1918 Dis3.n0 Dis3.t1 389.3
R1919 Dis3.n0 Dis3 297.494
R1920 Dis3 Dis3.n0 112
R1921 s1_bar.t7 s1_bar.t5 819.4
R1922 s1_bar.n4 s1_bar.t6 506.1
R1923 s1_bar.n4 s1_bar.t7 313.3
R1924 s1_bar.n2 s1_bar.t4 181.136
R1925 s1_bar.n3 s1_bar.n0 128.334
R1926 s1_bar.n2 s1_bar.n1 57.937
R1927 s1_bar.n5 s1_bar.n3 57.6
R1928 s1_bar.n3 s1_bar.n2 41.6
R1929 s1_bar.n0 s1_bar.t0 39.4
R1930 s1_bar.n0 s1_bar.t1 39.4
R1931 s1_bar.n1 s1_bar.t2 24
R1932 s1_bar.n1 s1_bar.t3 24
R1933 s1_bar.n5 s1_bar.n4 8.764
R1934 s1_bar s1_bar.n5 4.681
R1935 s1.t9 s1.t8 819.4
R1936 s1.n3 s1.t9 514.133
R1937 s1.n3 s1.t7 305.266
R1938 s1.n4 s1.n1 166.734
R1939 s1.n5 s1.n4 105.6
R1940 s1.n5 s1.t5 97.937
R1941 s1.n6 s1.n5 96
R1942 s1 s1.n6 83.684
R1943 s1 s1.n3 79.2
R1944 s1.n4 s1.n2 73.937
R1945 s1.n6 s1.n0 73.937
R1946 s1.n4 s1 54.4
R1947 s1.n1 s1.t1 39.4
R1948 s1.n1 s1.t2 39.4
R1949 s1.n2 s1.t3 24
R1950 s1.n2 s1.t0 24
R1951 s1.n0 s1.t4 24
R1952 s1.n0 s1.t6 24
R1953 EESPFAL_3in_NOR_v2_0/C_bar.t8 EESPFAL_3in_NOR_v2_0/C_bar.t7 819.4
R1954 EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_3in_NOR_v2_0/C_bar.t5 506.1
R1955 EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_3in_NOR_v2_0/C_bar.t8 313.3
R1956 EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_3in_NOR_v2_0/C_bar.t6 305.997
R1957 EESPFAL_INV4_0/OUT EESPFAL_3in_NOR_v2_0/C_bar.n0 206.179
R1958 EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_3in_NOR_v2_0/C_bar.t1 187.536
R1959 EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_3in_NOR_v2_0/C_bar.n3 128.335
R1960 EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_3in_NOR_v2_0/C_bar 115.2
R1961 EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_3in_NOR_v2_0/C_bar.n1 57.937
R1962 EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_3in_NOR_v2_0/C_bar.n4 57.6
R1963 EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_3in_NOR_v2_0/C_bar.n2 41.6
R1964 EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_3in_NOR_v2_0/C_bar.t4 39.4
R1965 EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_3in_NOR_v2_0/C_bar.t3 39.4
R1966 EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_3in_NOR_v2_0/C_bar.t2 24
R1967 EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_3in_NOR_v2_0/C_bar.t0 24
R1968 EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_3in_NOR_v2_0/C_bar.n5 8.764
R1969 EESPFAL_INV4_0/OUT EESPFAL_3in_NOR_v2_0/C_bar.n6 4.65
R1970 x2_bar.n0 x2_bar.t1 1069.04
R1971 x2_bar.n0 x2_bar.t2 1015.9
R1972 EESPFAL_INV4_1/A_bar x2_bar.t0 392.5
R1973 EESPFAL_INV4_1/A_bar x2_bar 184.698
R1974 x2_bar x2_bar.n0 89.6
R1975 x2.n0 x2.t1 1176.57
R1976 x2.n0 x2.t2 1149.49
R1977 EESPFAL_INV4_1/A x2.t0 778.1
R1978 x2 x2.n0 128
R1979 EESPFAL_INV4_1/A x2 44.3
R1980 x0.n0 x0.t2 800.452
R1981 x0.n0 x0.t1 787.997
R1982 EESPFAL_3in_NAND_v2_0/C_bar x0.t0 430.966
R1983 EESPFAL_3in_NAND_v2_0/C_bar x0.n1 368.182
R1984 x0.n1 x0 315.05
R1985 x0 x0.n0 169.6
R1986 x0.n1 x0 0.228
R1987 EESPFAL_3in_NAND_v2_0/A x3_bar.t0 1271.5
R1988 x3_bar.n0 x3_bar.t2 810.772
R1989 x3_bar.n0 x3_bar.t1 694.566
R1990 x3_bar x3_bar.t3 392.5
R1991 x3_bar.n1 x3_bar 179.639
R1992 x3_bar.n2 EESPFAL_3in_NAND_v2_0/A 109.588
R1993 EESPFAL_XOR_v3_1/B_bar x3_bar.n2 59.69
R1994 EESPFAL_XOR_v3_1/B_bar x3_bar.n0 25.6
R1995 x3_bar.n2 x3_bar.n1 1.69
R1996 x3_bar.n1 x3_bar 0.912
C0 x2 a_n3420_n613# 0.00fF
C1 EESPFAL_NAND_v3_1/B a_n1860_n613# 0.00fF
C2 EESPFAL_NAND_v3_0/B CLK1 0.70fF
C3 EESPFAL_INV4_0/A_bar x2_bar 0.00fF
C4 EESPFAL_NAND_v3_0/B x3_bar 0.01fF
C5 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_1/A 0.00fF
C6 Dis2 CLK1 0.08fF
C7 a_n3720_67# x3 0.00fF
C8 Dis2 EESPFAL_NAND_v3_1/A 0.04fF
C9 a_n1860_n613# Dis1 0.00fF
C10 a_1910_n613# EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C11 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/A 3.15fF
C12 a_n1860_n613# EESPFAL_NAND_v3_1/A_bar 0.00fF
C13 EESPFAL_INV4_0/A_bar x0 0.01fF
C14 EESPFAL_3in_NOR_v2_0/C CLK3 0.50fF
C15 x1 CLK2 0.03fF
C16 a_n3720_67# x2_bar 0.00fF
C17 EESPFAL_NAND_v3_0/A x1_bar 0.01fF
C18 EESPFAL_NAND_v3_0/A_bar CLK3 0.01fF
C19 s1 EESPFAL_NAND_v3_1/B_bar 0.00fF
C20 EESPFAL_NAND_v3_0/B_bar x2 0.02fF
C21 a_n3720_67# x0 0.00fF
C22 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_NAND_v3_1/B_bar 0.00fF
C23 EESPFAL_INV4_0/A_bar CLK2 0.08fF
C24 x1_bar a_n3420_n613# 0.00fF
C25 a_n2160_67# x0_bar 0.00fF
C26 a_n3420_67# EESPFAL_NAND_v3_0/A 0.01fF
C27 EESPFAL_3in_NOR_v2_0/C_bar Dis2 0.23fF
C28 a_n1860_n613# x3 0.00fF
C29 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/A_bar 0.38fF
C30 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/A 0.99fF
C31 EESPFAL_NAND_v3_1/B EESPFAL_INV4_0/A 0.01fF
C32 EESPFAL_NAND_v3_1/OUT a_1910_n613# 0.01fF
C33 s1 EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C34 Dis2 EESPFAL_NAND_v3_0/A 0.02fF
C35 s1_bar CLK2 0.26fF
C36 a_n2160_67# CLK1 0.02fF
C37 a_n2160_67# x3_bar 0.01fF
C38 x2_bar a_n1860_n613# 0.01fF
C39 a_n2160_67# EESPFAL_NAND_v3_1/A 0.00fF
C40 EESPFAL_INV4_0/A Dis1 0.11fF
C41 EESPFAL_NAND_v3_0/B CLK3 0.01fF
C42 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/OUT_bar 0.14fF
C43 EESPFAL_INV4_0/A EESPFAL_NAND_v3_1/A_bar 0.01fF
C44 s1_bar EESPFAL_NAND_v3_0/OUT 0.07fF
C45 Dis2 CLK3 1.29fF
C46 a_n1860_n613# x0 0.00fF
C47 EESPFAL_NAND_v3_1/OUT_bar Dis1 0.00fF
C48 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_1/A_bar 0.05fF
C49 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/B_bar 0.01fF
C50 x1 x2 0.28fF
C51 EESPFAL_INV4_0/A a_n2009_n2753# 0.01fF
C52 x1 a_n2160_n613# 0.00fF
C53 s1_bar a_2081_n2754# 0.00fF
C54 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar 0.55fF
C55 EESPFAL_3in_NOR_v2_0/C x1 0.00fF
C56 EESPFAL_INV4_0/A_bar x2 0.04fF
C57 EESPFAL_NAND_v3_1/OUT_bar a_1910_67# 0.00fF
C58 Dis3 EESPFAL_NAND_v3_1/B_bar 0.04fF
C59 Dis2 EESPFAL_NAND_v3_0/B_bar 0.02fF
C60 a_1910_n613# EESPFAL_NAND_v3_1/A 0.01fF
C61 s1 EESPFAL_NAND_v3_1/OUT 0.06fF
C62 EESPFAL_NAND_v3_0/A_bar x1 0.00fF
C63 EESPFAL_INV4_0/A x3 0.02fF
C64 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_0/OUT_bar 0.09fF
C65 EESPFAL_NAND_v3_1/B Dis1 0.16fF
C66 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/A_bar 0.36fF
C67 a_n3720_67# x2 0.00fF
C68 a_n2160_67# EESPFAL_NAND_v3_0/A 0.00fF
C69 x1_bar x1 5.71fF
C70 EESPFAL_INV4_0/A_bar EESPFAL_3in_NOR_v2_0/C 0.01fF
C71 x2_bar EESPFAL_INV4_0/A 0.00fF
C72 Dis1 EESPFAL_NAND_v3_1/A_bar 0.32fF
C73 CLK1 EESPFAL_NAND_v3_1/B_bar 0.70fF
C74 x3_bar EESPFAL_NAND_v3_1/B_bar 0.00fF
C75 EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/B_bar 0.03fF
C76 s1 Dis3 0.41fF
C77 EESPFAL_INV4_0/A x0 0.00fF
C78 a_n3720_n613# Dis1 0.02fF
C79 Dis3 EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C80 a_n3720_n613# EESPFAL_NAND_v3_1/A_bar 0.01fF
C81 a_n1860_67# CLK1 0.02fF
C82 a_n3420_67# x1 0.00fF
C83 a_n1860_67# x3_bar 0.01fF
C84 a_n1860_67# EESPFAL_NAND_v3_1/A 0.00fF
C85 EESPFAL_INV4_0/A_bar x1_bar 0.08fF
C86 s1_bar EESPFAL_3in_NOR_v2_0/C 0.12fF
C87 a_n3720_67# EESPFAL_NAND_v3_0/A_bar 0.00fF
C88 EESPFAL_3in_NOR_v2_0/C_bar a_1910_n613# 0.00fF
C89 a_n2159_n2753# x0_bar 0.00fF
C90 s1 EESPFAL_NAND_v3_1/A 0.02fF
C91 EESPFAL_INV4_0/A CLK2 0.72fF
C92 EESPFAL_NAND_v3_1/B x3 0.03fF
C93 EESPFAL_NAND_v3_0/A a_1910_n613# 0.00fF
C94 CLK1 EESPFAL_NAND_v3_0/OUT_bar 0.05fF
C95 a_n3720_67# x1_bar 0.00fF
C96 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_NAND_v3_1/A 0.01fF
C97 a_n2160_67# EESPFAL_NAND_v3_0/B_bar 0.00fF
C98 a_n1860_n613# x2 0.00fF
C99 x3 Dis1 0.18fF
C100 EESPFAL_NAND_v3_1/OUT_bar CLK2 1.23fF
C101 x3 EESPFAL_NAND_v3_1/A_bar 0.10fF
C102 EESPFAL_NAND_v3_0/OUT EESPFAL_INV4_0/A 0.01fF
C103 EESPFAL_NAND_v3_1/B x2_bar 0.04fF
C104 a_1910_n613# CLK3 0.00fF
C105 EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_NAND_v3_1/B_bar 0.01fF
C106 a_n2159_n2753# CLK1 0.02fF
C107 x3_bar a_n2159_n2753# 0.00fF
C108 x2_bar Dis1 0.23fF
C109 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_0/OUT 0.09fF
C110 x3 a_n3720_n613# 0.00fF
C111 s1 a_1931_n2754# 0.01fF
C112 x2_bar EESPFAL_NAND_v3_1/A_bar 0.12fF
C113 x3 a_n2009_n2753# 0.00fF
C114 EESPFAL_INV4_0/A_bar Dis2 0.01fF
C115 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/B_bar 0.00fF
C116 EESPFAL_NAND_v3_1/OUT Dis3 0.02fF
C117 Dis1 x0 0.08fF
C118 EESPFAL_NAND_v3_1/A_bar x0 0.01fF
C119 CLK3 EESPFAL_NAND_v3_1/B_bar 0.02fF
C120 x2_bar a_n3720_n613# 0.01fF
C121 EESPFAL_NAND_v3_0/A_bar a_n1860_n613# 0.00fF
C122 a_n1860_67# EESPFAL_NAND_v3_0/A 0.00fF
C123 EESPFAL_NAND_v3_1/OUT_bar a_2081_n2754# 0.00fF
C124 s1 EESPFAL_3in_NOR_v2_0/C_bar 0.08fF
C125 a_n3720_n613# x0 0.00fF
C126 EESPFAL_NAND_v3_1/B CLK2 0.47fF
C127 s1_bar Dis2 0.01fF
C128 EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_NAND_v3_0/OUT_bar 0.02fF
C129 a_n1860_n613# x1_bar 0.00fF
C130 EESPFAL_NAND_v3_1/OUT CLK1 0.01fF
C131 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/A 0.07fF
C132 CLK2 Dis1 0.01fF
C133 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/OUT_bar 0.06fF
C134 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_0/OUT 0.03fF
C135 CLK2 EESPFAL_NAND_v3_1/A_bar 0.10fF
C136 a_n2160_67# x1 0.00fF
C137 EESPFAL_3in_NOR_v2_0/C_bar a_n2159_n2753# 0.00fF
C138 s1 CLK3 1.06fF
C139 x2_bar x3 3.66fF
C140 EESPFAL_INV4_0/A x2 0.05fF
C141 EESPFAL_NAND_v3_0/OUT Dis1 0.00fF
C142 CLK3 EESPFAL_NAND_v3_0/OUT_bar 0.13fF
C143 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_1/A_bar 0.00fF
C144 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_1/B_bar 0.02fF
C145 a_n2009_n2753# CLK2 0.00fF
C146 CLK1 x0_bar 0.72fF
C147 x3 x0 0.09fF
C148 x3_bar x0_bar 0.18fF
C149 EESPFAL_NAND_v3_1/A x0_bar 0.02fF
C150 Dis3 CLK1 0.26fF
C151 EESPFAL_NAND_v3_1/OUT_bar x2 0.00fF
C152 x3_bar Dis3 0.00fF
C153 Dis3 EESPFAL_NAND_v3_1/A 0.08fF
C154 EESPFAL_NAND_v3_1/OUT a_1931_n2754# 0.00fF
C155 a_1910_67# CLK2 0.02fF
C156 a_n1860_67# EESPFAL_NAND_v3_0/B_bar 0.00fF
C157 EESPFAL_3in_NOR_v2_0/C EESPFAL_INV4_0/A 0.07fF
C158 x2_bar x0 1.81fF
C159 EESPFAL_NAND_v3_0/OUT a_1910_67# 0.01fF
C160 EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_NAND_v3_1/OUT 0.08fF
C161 EESPFAL_3in_NOR_v2_0/C EESPFAL_NAND_v3_1/OUT_bar 0.04fF
C162 x3_bar CLK1 2.40fF
C163 x3 CLK2 0.02fF
C164 x3_bar EESPFAL_NAND_v3_1/A 0.13fF
C165 CLK1 EESPFAL_NAND_v3_1/A 1.43fF
C166 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/OUT_bar 0.09fF
C167 Dis3 a_1931_n2754# 0.00fF
C168 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_0/A 0.00fF
C169 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_0/A_bar 0.00fF
C170 EESPFAL_INV4_0/A x1_bar 0.01fF
C171 EESPFAL_NAND_v3_0/OUT x3 0.00fF
C172 x2_bar CLK2 0.01fF
C173 EESPFAL_NAND_v3_1/B x2 0.33fF
C174 EESPFAL_NAND_v3_1/OUT CLK3 0.76fF
C175 EESPFAL_3in_NOR_v2_0/C_bar x0_bar 0.00fF
C176 x2 Dis1 0.16fF
C177 EESPFAL_NAND_v3_1/B a_n2160_n613# 0.00fF
C178 EESPFAL_3in_NOR_v2_0/C_bar Dis3 0.18fF
C179 x1 EESPFAL_NAND_v3_1/B_bar 0.00fF
C180 x2 EESPFAL_NAND_v3_1/A_bar 1.05fF
C181 a_1931_n2754# EESPFAL_NAND_v3_1/A 0.00fF
C182 EESPFAL_NAND_v3_0/A x0_bar 0.31fF
C183 EESPFAL_NAND_v3_0/A Dis3 0.08fF
C184 a_n2160_n613# Dis1 0.00fF
C185 EESPFAL_3in_NOR_v2_0/C EESPFAL_NAND_v3_1/B 0.01fF
C186 a_n2160_n613# EESPFAL_NAND_v3_1/A_bar 0.00fF
C187 x2 a_n3720_n613# 0.00fF
C188 a_n2009_n2753# x2 0.00fF
C189 EESPFAL_3in_NOR_v2_0/C Dis1 0.00fF
C190 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_0/A_bar 0.00fF
C191 Dis3 CLK3 1.19fF
C192 EESPFAL_3in_NOR_v2_0/C_bar x3_bar 0.01fF
C193 EESPFAL_3in_NOR_v2_0/C_bar CLK1 0.16fF
C194 a_n3420_n613# x0_bar 0.00fF
C195 EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_NAND_v3_1/A 0.03fF
C196 EESPFAL_3in_NOR_v2_0/C EESPFAL_NAND_v3_1/A_bar 0.00fF
C197 Dis2 EESPFAL_INV4_0/A 0.04fF
C198 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_0/B 0.02fF
C199 EESPFAL_NAND_v3_0/A_bar Dis1 0.29fF
C200 EESPFAL_NAND_v3_0/A x3_bar 0.15fF
C201 EESPFAL_NAND_v3_0/A CLK1 1.45fF
C202 EESPFAL_NAND_v3_1/B x1_bar 0.00fF
C203 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/A 0.02fF
C204 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_1/A_bar 0.02fF
C205 Dis2 EESPFAL_NAND_v3_1/OUT_bar 0.31fF
C206 EESPFAL_NAND_v3_0/OUT CLK2 0.97fF
C207 EESPFAL_3in_NOR_v2_0/C a_n2009_n2753# 0.00fF
C208 x1_bar Dis1 0.08fF
C209 CLK1 CLK3 0.04fF
C210 x1_bar EESPFAL_NAND_v3_1/A_bar 0.06fF
C211 x3_bar CLK3 0.00fF
C212 CLK3 EESPFAL_NAND_v3_1/A 0.20fF
C213 x3 x2 0.34fF
C214 CLK1 a_n3420_n613# 0.02fF
C215 s1_bar EESPFAL_NAND_v3_1/B_bar 0.00fF
C216 a_n3420_n613# EESPFAL_NAND_v3_1/A 0.00fF
C217 EESPFAL_3in_NOR_v2_0/C_bar a_1931_n2754# 0.00fF
C218 x3_bar a_n3420_n613# 0.01fF
C219 a_n2159_n2753# x1 0.01fF
C220 s1 EESPFAL_INV4_0/A_bar 0.00fF
C221 EESPFAL_NAND_v3_0/B_bar x0_bar 0.00fF
C222 x3 a_n2160_n613# 0.00fF
C223 x1_bar a_n3720_n613# 0.00fF
C224 EESPFAL_NAND_v3_0/B_bar Dis3 0.05fF
C225 CLK2 a_2081_n2754# 0.00fF
C226 a_n2009_n2753# x1_bar 0.00fF
C227 x2_bar x2 6.02fF
C228 a_n3420_67# Dis1 0.01fF
C229 a_n3420_67# EESPFAL_NAND_v3_1/A_bar 0.00fF
C230 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_0/B 0.03fF
C231 x2 x0 0.23fF
C232 x2_bar a_n2160_n613# 0.01fF
C233 EESPFAL_NAND_v3_0/OUT a_2081_n2754# 0.00fF
C234 CLK3 a_1931_n2754# 0.01fF
C235 Dis2 EESPFAL_NAND_v3_1/B 0.06fF
C236 EESPFAL_INV4_0/A_bar a_n2159_n2753# 0.00fF
C237 EESPFAL_NAND_v3_0/A_bar x3 0.98fF
C238 s1_bar s1 2.14fF
C239 EESPFAL_NAND_v3_0/B Dis1 0.10fF
C240 EESPFAL_NAND_v3_0/B_bar x3_bar 0.04fF
C241 EESPFAL_NAND_v3_0/B_bar CLK1 1.03fF
C242 a_n2160_n613# x0 0.00fF
C243 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_1/A 0.00fF
C244 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_1/A_bar 0.00fF
C245 Dis2 Dis1 0.03fF
C246 s1_bar EESPFAL_NAND_v3_0/OUT_bar 0.05fF
C247 Dis2 EESPFAL_NAND_v3_1/A_bar 0.02fF
C248 x3 x1_bar 2.32fF
C249 a_n1860_n613# EESPFAL_NAND_v3_1/B_bar 0.00fF
C250 EESPFAL_NAND_v3_0/A_bar x2_bar 0.07fF
C251 EESPFAL_3in_NOR_v2_0/C_bar CLK3 0.32fF
C252 CLK2 x2 0.15fF
C253 EESPFAL_NAND_v3_0/A_bar x0 0.07fF
C254 x2_bar x1_bar 0.08fF
C255 EESPFAL_NAND_v3_0/A CLK3 0.01fF
C256 EESPFAL_NAND_v3_0/A a_n3420_n613# 0.00fF
C257 a_n3420_67# x3 0.01fF
C258 Dis2 a_1910_67# 0.00fF
C259 x1 x0_bar 5.56fF
C260 x1_bar x0 0.56fF
C261 EESPFAL_3in_NOR_v2_0/C CLK2 1.06fF
C262 EESPFAL_NAND_v3_0/B x3 0.08fF
C263 a_n3420_67# x2_bar 0.00fF
C264 EESPFAL_NAND_v3_0/A_bar CLK2 0.09fF
C265 EESPFAL_3in_NOR_v2_0/C EESPFAL_NAND_v3_0/OUT 0.10fF
C266 Dis2 x3 0.00fF
C267 a_n3420_67# x0 0.00fF
C268 EESPFAL_INV4_0/A_bar x0_bar 0.15fF
C269 s1_bar EESPFAL_NAND_v3_1/OUT 0.11fF
C270 x1 CLK1 1.79fF
C271 x1 EESPFAL_NAND_v3_1/A 0.05fF
C272 EESPFAL_INV4_0/A_bar Dis3 0.00fF
C273 EESPFAL_NAND_v3_0/B x2_bar 0.00fF
C274 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/A_bar 0.01fF
C275 x3_bar x1 1.29fF
C276 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/A 0.03fF
C277 EESPFAL_NAND_v3_1/OUT_bar a_1910_n613# 0.00fF
C278 a_n2160_67# Dis1 0.00fF
C279 a_n2160_67# EESPFAL_NAND_v3_1/A_bar 0.00fF
C280 EESPFAL_NAND_v3_0/B x0 0.01fF
C281 EESPFAL_3in_NOR_v2_0/C a_2081_n2754# 0.00fF
C282 EESPFAL_NAND_v3_0/B_bar CLK3 0.02fF
C283 EESPFAL_INV4_0/A EESPFAL_NAND_v3_1/B_bar 0.01fF
C284 a_n3720_67# x0_bar 0.00fF
C285 EESPFAL_INV4_0/A_bar x3_bar 0.06fF
C286 EESPFAL_INV4_0/A_bar CLK1 1.42fF
C287 EESPFAL_INV4_0/A_bar EESPFAL_NAND_v3_1/A 0.01fF
C288 s1_bar Dis3 0.28fF
C289 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_1/B_bar 0.12fF
C290 EESPFAL_NAND_v3_0/B CLK2 0.38fF
C291 x2 a_n2160_n613# 0.00fF
C292 Dis2 CLK2 1.30fF
C293 a_n3720_67# CLK1 0.01fF
C294 a_n3720_67# x3_bar 0.01fF
C295 s1 EESPFAL_INV4_0/A 0.00fF
C296 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/OUT 0.07fF
C297 s1_bar EESPFAL_NAND_v3_1/A 0.03fF
C298 EESPFAL_3in_NOR_v2_0/C_bar x1 0.00fF
C299 EESPFAL_3in_NOR_v2_0/C x2 0.00fF
C300 Dis2 EESPFAL_NAND_v3_0/OUT 0.16fF
C301 a_n2160_67# x3 0.00fF
C302 s1 EESPFAL_NAND_v3_1/OUT_bar 0.02fF
C303 EESPFAL_NAND_v3_0/A x1 0.01fF
C304 EESPFAL_NAND_v3_0/A_bar x2 0.04fF
C305 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_0/OUT_bar 1.02fF
C306 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar 0.49fF
C307 EESPFAL_INV4_0/A a_n2159_n2753# 0.01fF
C308 a_n2160_67# x2_bar 0.00fF
C309 EESPFAL_NAND_v3_0/A_bar a_n2160_n613# 0.00fF
C310 x1_bar x2 2.72fF
C311 EESPFAL_INV4_0/A_bar EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C312 Dis1 EESPFAL_NAND_v3_1/B_bar 0.09fF
C313 x1 a_n3420_n613# 0.00fF
C314 s1_bar a_1931_n2754# 0.00fF
C315 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/B_bar 0.21fF
C316 a_n2160_67# x0 0.00fF
C317 x1_bar a_n2160_n613# 0.00fF
C318 a_n1860_67# Dis1 0.00fF
C319 a_n1860_n613# CLK1 0.02fF
C320 a_n1860_n613# x3_bar 0.00fF
C321 a_n1860_n613# EESPFAL_NAND_v3_1/A 0.01fF
C322 a_n1860_67# EESPFAL_NAND_v3_1/A_bar 0.00fF
C323 a_n3420_67# x2 0.00fF
C324 s1 EESPFAL_NAND_v3_1/B 0.00fF
C325 s1_bar EESPFAL_3in_NOR_v2_0/C_bar 1.83fF
C326 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_0/OUT_bar 0.02fF
C327 a_n3720_67# EESPFAL_NAND_v3_0/A 0.01fF
C328 EESPFAL_NAND_v3_0/A_bar x1_bar 0.00fF
C329 EESPFAL_NAND_v3_1/OUT EESPFAL_INV4_0/A 0.00fF
C330 s1 EESPFAL_NAND_v3_1/A_bar 0.00fF
C331 EESPFAL_NAND_v3_0/B x2 0.02fF
C332 EESPFAL_NAND_v3_0/OUT_bar Dis1 0.00fF
C333 Dis2 x2 0.00fF
C334 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_NAND_v3_1/A_bar 0.00fF
C335 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar 0.66fF
C336 x3 EESPFAL_NAND_v3_1/B_bar 0.02fF
C337 s1_bar CLK3 1.19fF
C338 a_n3420_67# EESPFAL_NAND_v3_0/A_bar 0.00fF
C339 a_n2159_n2753# Dis1 0.00fF
C340 EESPFAL_INV4_0/A x0_bar 0.08fF
C341 EESPFAL_INV4_0/A Dis3 0.00fF
C342 EESPFAL_3in_NOR_v2_0/C Dis2 0.41fF
C343 x2_bar EESPFAL_NAND_v3_1/B_bar 0.01fF
C344 a_n1860_67# x3 0.00fF
C345 a_1910_67# EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C346 a_n3420_67# x1_bar 0.00fF
C347 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/A_bar 0.31fF
C348 EESPFAL_NAND_v3_1/OUT_bar Dis3 0.01fF
C349 Dis2 EESPFAL_NAND_v3_0/A_bar 0.02fF
C350 a_1910_n613# CLK2 0.02fF
C351 EESPFAL_NAND_v3_0/A a_n1860_n613# 0.00fF
C352 a_n1860_67# x2_bar 0.01fF
C353 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/OUT 0.08fF
C354 EESPFAL_INV4_0/A x3_bar 0.04fF
C355 EESPFAL_INV4_0/A CLK1 1.05fF
C356 EESPFAL_INV4_0/A EESPFAL_NAND_v3_1/A 0.06fF
C357 x3 EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C358 EESPFAL_NAND_v3_0/OUT a_1910_n613# 0.01fF
C359 a_n1860_67# x0 0.00fF
C360 EESPFAL_NAND_v3_1/OUT Dis1 0.00fF
C361 EESPFAL_NAND_v3_1/OUT_bar CLK1 0.05fF
C362 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/A_bar 0.01fF
C363 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_1/A 0.07fF
C364 CLK2 EESPFAL_NAND_v3_1/B_bar 0.12fF
C365 x3 a_n2159_n2753# 0.00fF
C366 a_n2160_67# x2 0.00fF
C367 EESPFAL_NAND_v3_1/B Dis3 0.04fF
C368 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_1/B_bar 0.00fF
C369 Dis1 x0_bar 0.12fF
C370 EESPFAL_INV4_0/A_bar x1 0.08fF
C371 EESPFAL_NAND_v3_1/A_bar x0_bar 0.03fF
C372 Dis3 Dis1 0.02fF
C373 EESPFAL_NAND_v3_1/OUT a_1910_67# 0.00fF
C374 Dis3 EESPFAL_NAND_v3_1/A_bar 0.08fF
C375 Dis2 EESPFAL_NAND_v3_0/B 0.05fF
C376 s1 CLK2 0.11fF
C377 a_n3720_n613# x0_bar 0.00fF
C378 EESPFAL_NAND_v3_1/B CLK1 0.88fF
C379 EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_INV4_0/A 0.34fF
C380 EESPFAL_NAND_v3_1/B x3_bar 0.00fF
C381 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/A 0.98fF
C382 CLK2 EESPFAL_NAND_v3_0/OUT_bar 1.19fF
C383 a_n3720_67# x1 0.00fF
C384 a_n2160_67# EESPFAL_NAND_v3_0/A_bar 0.01fF
C385 CLK1 Dis1 3.35fF
C386 s1 EESPFAL_NAND_v3_0/OUT 0.05fF
C387 x3_bar Dis1 0.29fF
C388 EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_NAND_v3_1/OUT_bar 0.22fF
C389 Dis1 EESPFAL_NAND_v3_1/A 0.28fF
C390 CLK1 EESPFAL_NAND_v3_1/A_bar 1.68fF
C391 EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/A_bar 3.23fF
C392 x3_bar EESPFAL_NAND_v3_1/A_bar 0.38fF
C393 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar 0.87fF
C394 a_n2160_67# x1_bar 0.00fF
C395 a_n2159_n2753# CLK2 0.00fF
C396 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_0/A 0.00fF
C397 EESPFAL_INV4_0/A CLK3 0.01fF
C398 CLK1 a_n3720_n613# 0.01fF
C399 x3_bar a_n3720_n613# 0.01fF
C400 a_n3720_n613# EESPFAL_NAND_v3_1/A 0.00fF
C401 a_n2009_n2753# CLK1 0.02fF
C402 x3_bar a_n2009_n2753# 0.01fF
C403 x3 x0_bar 0.77fF
C404 s1 a_2081_n2754# 0.01fF
C405 EESPFAL_NAND_v3_1/OUT_bar CLK3 0.38fF
C406 x3 Dis3 0.01fF
C407 EESPFAL_NAND_v3_0/OUT_bar a_2081_n2754# 0.00fF
C408 EESPFAL_3in_NOR_v2_0/C a_1910_n613# 0.00fF
C409 x2 EESPFAL_NAND_v3_1/B_bar 0.07fF
C410 a_1910_67# EESPFAL_NAND_v3_1/A 0.00fF
C411 x2_bar x0_bar 0.18fF
C412 x2_bar Dis3 0.00fF
C413 EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_NAND_v3_1/B 0.01fF
C414 x0_bar x0 5.73fF
C415 a_n1860_67# x2 0.00fF
C416 x3 CLK1 1.85fF
C417 x3 x3_bar 5.75fF
C418 EESPFAL_NAND_v3_1/OUT CLK2 0.94fF
C419 x3 EESPFAL_NAND_v3_1/A 0.07fF
C420 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_0/A 0.00fF
C421 EESPFAL_3in_NOR_v2_0/C_bar Dis1 0.00fF
C422 EESPFAL_3in_NOR_v2_0/C EESPFAL_NAND_v3_1/B_bar 0.01fF
C423 EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_NAND_v3_1/A_bar 0.00fF
C424 EESPFAL_NAND_v3_0/A Dis1 0.32fF
C425 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_0/OUT 1.64fF
C426 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_0/B_bar 0.00fF
C427 x2_bar CLK1 1.21fF
C428 x2_bar x3_bar 0.41fF
C429 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_1/B_bar 0.00fF
C430 x2_bar EESPFAL_NAND_v3_1/A 0.21fF
C431 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/A_bar 0.02fF
C432 EESPFAL_NAND_v3_1/B CLK3 0.05fF
C433 EESPFAL_3in_NOR_v2_0/C_bar a_n2009_n2753# 0.00fF
C434 CLK2 x0_bar 0.01fF
C435 CLK1 x0 0.49fF
C436 CLK3 Dis1 0.00fF
C437 x3_bar x0 0.09fF
C438 EESPFAL_NAND_v3_1/A x0 0.01fF
C439 Dis3 CLK2 0.18fF
C440 x1_bar EESPFAL_NAND_v3_1/B_bar 0.00fF
C441 EESPFAL_NAND_v3_0/A a_n3720_n613# 0.00fF
C442 CLK3 EESPFAL_NAND_v3_1/A_bar 0.03fF
C443 a_n3420_n613# Dis1 0.01fF
C444 a_n1860_67# EESPFAL_NAND_v3_0/A_bar 0.01fF
C445 a_n3420_n613# EESPFAL_NAND_v3_1/A_bar 0.01fF
C446 EESPFAL_NAND_v3_1/OUT a_2081_n2754# 0.00fF
C447 s1 EESPFAL_3in_NOR_v2_0/C 0.08fF
C448 a_n2159_n2753# x2 0.00fF
C449 EESPFAL_NAND_v3_0/OUT Dis3 0.03fF
C450 EESPFAL_NAND_v3_0/A a_1910_67# 0.01fF
C451 EESPFAL_3in_NOR_v2_0/C EESPFAL_NAND_v3_0/OUT_bar 0.10fF
C452 a_n1860_67# x1_bar 0.00fF
C453 Dis2 a_1910_n613# 0.00fF
C454 CLK1 CLK2 1.29fF
C455 x3_bar CLK2 0.07fF
C456 CLK2 EESPFAL_NAND_v3_1/A 0.95fF
C457 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/OUT_bar 0.05fF
C458 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_0/B_bar 0.01fF
C459 a_1910_67# CLK3 0.00fF
C460 EESPFAL_3in_NOR_v2_0/C a_n2159_n2753# 0.00fF
C461 EESPFAL_NAND_v3_0/A x3 0.27fF
C462 EESPFAL_INV4_0/A x1 0.04fF
C463 EESPFAL_NAND_v3_0/B_bar Dis1 0.17fF
C464 Dis3 a_2081_n2754# 0.00fF
C465 EESPFAL_NAND_v3_0/OUT CLK1 0.01fF
C466 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_1/B_bar 0.02fF
C467 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_1/A 0.07fF
C468 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_1/A_bar 0.00fF
C469 Dis2 EESPFAL_NAND_v3_1/B_bar 0.03fF
C470 x3 CLK3 0.00fF
C471 EESPFAL_NAND_v3_1/OUT x2 0.00fF
C472 EESPFAL_NAND_v3_0/A x2_bar 0.13fF
C473 x3 a_n3420_n613# 0.01fF
C474 CLK2 a_1931_n2754# 0.00fF
C475 a_n1860_67# EESPFAL_NAND_v3_0/B 0.00fF
C476 a_n2159_n2753# x1_bar 0.00fF
C477 EESPFAL_NAND_v3_0/A x0 0.09fF
C478 EESPFAL_INV4_0/A_bar EESPFAL_INV4_0/A 0.73fF
C479 x2_bar CLK3 0.00fF
C480 x2_bar a_n3420_n613# 0.01fF
C481 EESPFAL_NAND_v3_0/OUT a_1931_n2754# 0.00fF
C482 EESPFAL_3in_NOR_v2_0/C EESPFAL_NAND_v3_1/OUT 1.45fF
C483 x2 x0_bar 0.13fF
C484 s1 Dis2 0.02fF
C485 EESPFAL_3in_NOR_v2_0/C_bar CLK2 0.91fF
C486 Dis3 x2 0.01fF
C487 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/OUT_bar 0.15fF
C488 a_n3420_n613# x0 0.00fF
C489 Dis2 EESPFAL_NAND_v3_0/OUT_bar 0.32fF
C490 a_n2160_n613# x0_bar 0.00fF
C491 EESPFAL_NAND_v3_0/B_bar x3 0.33fF
C492 s1_bar EESPFAL_INV4_0/A 0.00fF
C493 EESPFAL_NAND_v3_0/A CLK2 0.66fF
C494 EESPFAL_NAND_v3_1/B x1 0.00fF
C495 EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_NAND_v3_0/OUT 0.01fF
C496 EESPFAL_3in_NOR_v2_0/C x0_bar 0.00fF
C497 x1 Dis1 0.08fF
C498 s1_bar EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C499 EESPFAL_3in_NOR_v2_0/C Dis3 0.18fF
C500 EESPFAL_NAND_v3_0/B_bar x2_bar 0.00fF
C501 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/A 0.04fF
C502 x3_bar x2 0.18fF
C503 x1 EESPFAL_NAND_v3_1/A_bar 0.06fF
C504 CLK1 x2 2.78fF
C505 CLK2 CLK3 0.97fF
C506 x2 EESPFAL_NAND_v3_1/A 0.26fF
C507 EESPFAL_NAND_v3_0/A_bar x0_bar 0.07fF
C508 EESPFAL_NAND_v3_0/A_bar Dis3 0.08fF
C509 EESPFAL_NAND_v3_0/B_bar x0 0.01fF
C510 CLK1 a_n2160_n613# 0.02fF
C511 x3_bar a_n2160_n613# 0.01fF
C512 a_n2160_n613# EESPFAL_NAND_v3_1/A 0.01fF
C513 EESPFAL_3in_NOR_v2_0/C_bar a_2081_n2754# 0.00fF
C514 EESPFAL_NAND_v3_0/OUT CLK3 1.16fF
C515 x1 a_n3720_n613# 0.00fF
C516 x1_bar x0_bar 0.13fF
C517 EESPFAL_INV4_0/A_bar Dis1 0.27fF
C518 EESPFAL_3in_NOR_v2_0/C CLK1 0.11fF
C519 EESPFAL_3in_NOR_v2_0/C x3_bar 0.01fF
C520 EESPFAL_3in_NOR_v2_0/C EESPFAL_NAND_v3_1/A 0.03fF
C521 EESPFAL_INV4_0/A_bar EESPFAL_NAND_v3_1/A_bar 0.02fF
C522 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_0/B 0.02fF
C523 EESPFAL_NAND_v3_0/A_bar CLK1 1.20fF
C524 EESPFAL_NAND_v3_0/A_bar x3_bar 0.23fF
C525 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_1/A 0.02fF
C526 CLK3 a_2081_n2754# 0.01fF
C527 Dis2 EESPFAL_NAND_v3_1/OUT 0.13fF
C528 EESPFAL_NAND_v3_0/B_bar CLK2 0.04fF
C529 s1_bar EESPFAL_NAND_v3_1/B 0.01fF
C530 EESPFAL_INV4_0/A_bar a_n2009_n2753# 0.00fF
C531 a_n3720_67# Dis1 0.02fF
C532 a_n3420_67# x0_bar 0.00fF
C533 a_n3720_67# EESPFAL_NAND_v3_1/A_bar 0.00fF
C534 x1_bar CLK1 0.88fF
C535 x3_bar x1_bar 0.17fF
C536 x3 x1 0.20fF
C537 x1_bar EESPFAL_NAND_v3_1/A 0.06fF
C538 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/OUT 0.00fF
C539 EESPFAL_3in_NOR_v2_0/C_bar x2 0.01fF
C540 s1_bar EESPFAL_NAND_v3_1/A_bar 0.00fF
C541 EESPFAL_3in_NOR_v2_0/C a_1931_n2754# 0.00fF
C542 EESPFAL_NAND_v3_0/B x0_bar 0.00fF
C543 EESPFAL_NAND_v3_0/B Dis3 0.05fF
C544 x2_bar x1 0.08fF
C545 EESPFAL_NAND_v3_0/A x2 0.07fF
C546 Dis2 Dis3 0.59fF
C547 a_n3420_67# CLK1 0.01fF
C548 a_n3420_67# x3_bar 0.01fF
C549 EESPFAL_INV4_0/A_bar x3 0.08fF
C550 x1 x0 0.04fF
C551 EESPFAL_NAND_v3_0/A a_n2160_n613# 0.00fF
C552 CLK3 x2 0.00fF
C553 EESPFAL_3in_NOR_v2_0/C EESPFAL_3in_NOR_v2_0/C_bar 2.13fF
C554 a_2081_n2754# GND 0.02fF
C555 a_1931_n2754# GND 0.02fF
C556 Dis3 GND 4.02fF
C557 a_n2009_n2753# GND 0.02fF
C558 a_n2159_n2753# GND 0.02fF
C559 s1 GND 1.76fF
C560 s1_bar GND 1.71fF
C561 EESPFAL_3in_NOR_v2_0/C_bar GND 1.26fF $ **FLOATING
C562 EESPFAL_3in_NOR_v2_0/C GND 1.22fF $ **FLOATING
C563 EESPFAL_INV4_0/A_bar GND 1.23fF
C564 EESPFAL_INV4_0/A GND 1.36fF
C565 a_1910_n613# GND 0.02fF
C566 a_n1860_n613# GND 0.01fF
C567 a_n2160_n613# GND 0.01fF
C568 a_n3420_n613# GND 0.01fF
C569 a_n3720_n613# GND 0.01fF
C570 EESPFAL_NAND_v3_1/OUT_bar GND 1.49fF
C571 EESPFAL_NAND_v3_1/OUT GND 1.14fF
C572 EESPFAL_NAND_v3_1/B GND 1.21fF
C573 EESPFAL_NAND_v3_1/B_bar GND 1.11fF
C574 EESPFAL_NAND_v3_1/A_bar GND 2.41fF $ **FLOATING
C575 EESPFAL_NAND_v3_1/A GND 2.46fF $ **FLOATING
C576 x1 GND 3.15fF
C577 x1_bar GND 3.01fF
C578 a_1910_67# GND 0.02fF
C579 a_n1860_67# GND 0.01fF
C580 a_n2160_67# GND 0.01fF
C581 a_n3420_67# GND 0.01fF
C582 a_n3720_67# GND 0.01fF
C583 Dis2 GND 4.83fF
C584 x3_bar GND 4.95fF
C585 x3 GND 8.10fF
C586 Dis1 GND 8.94fF
C587 EESPFAL_NAND_v3_0/OUT_bar GND 2.58fF $ **FLOATING
C588 EESPFAL_NAND_v3_0/OUT GND 1.78fF
C589 EESPFAL_NAND_v3_0/B_bar GND 1.17fF
C590 EESPFAL_NAND_v3_0/B GND 1.35fF
C591 x0 GND 2.65fF
C592 x0_bar GND 2.48fF
C593 x2_bar GND 5.37fF
C594 EESPFAL_NAND_v3_0/A GND 2.99fF $ **FLOATING
C595 EESPFAL_NAND_v3_0/A_bar GND 1.95fF $ **FLOATING
C596 x2 GND 9.30fF
C597 CLK3 GND 3.69fF
C598 CLK2 GND 9.52fF
C599 CLK1 GND 17.65fF
C600 x3_bar.t2 GND 0.44fF
C601 x3_bar.t1 GND 0.15fF
C602 x3_bar.n0 GND 1.46fF $ **FLOATING
C603 x3_bar.t3 GND 0.12fF
C604 x3_bar.n1 GND 3.72fF $ **FLOATING
C605 x3_bar.t0 GND 0.38fF
C606 EESPFAL_3in_NAND_v2_0/A GND 1.68fF $ **FLOATING
C607 x3_bar.n2 GND 3.28fF $ **FLOATING
C608 EESPFAL_XOR_v3_1/B_bar GND 0.09fF $ **FLOATING
C609 x0.t0 GND 0.12fF
C610 x0.t1 GND 0.14fF
C611 x0.t2 GND 0.15fF
C612 x0.n0 GND 1.75fF $ **FLOATING
C613 x0.n1 GND 4.59fF $ **FLOATING
C614 EESPFAL_3in_NAND_v2_0/C_bar GND 0.53fF $ **FLOATING
C615 x2.t0 GND 0.16fF
C616 x2.t2 GND 0.23fF
C617 x2.t1 GND 0.20fF
C618 x2.n0 GND 1.75fF $ **FLOATING
C619 EESPFAL_INV4_1/A GND 1.30fF $ **FLOATING
C620 x2_bar.t0 GND 0.23fF
C621 x2_bar.t1 GND 0.65fF
C622 x2_bar.t2 GND 0.37fF
C623 x2_bar.n0 GND 3.46fF $ **FLOATING
C624 EESPFAL_INV4_1/A_bar GND 0.82fF $ **FLOATING
C625 EESPFAL_INV4_0/OUT GND 0.23fF $ **FLOATING
C626 EESPFAL_3in_NOR_v2_0/C_bar.t6 GND 0.03fF
C627 EESPFAL_3in_NOR_v2_0/C_bar.n0 GND 0.63fF $ **FLOATING
C628 EESPFAL_3in_NOR_v2_0/C_bar.t2 GND 0.04fF
C629 EESPFAL_3in_NOR_v2_0/C_bar.t0 GND 0.04fF
C630 EESPFAL_3in_NOR_v2_0/C_bar.n1 GND 0.13fF $ **FLOATING
C631 EESPFAL_3in_NOR_v2_0/C_bar.t1 GND 0.25fF
C632 EESPFAL_3in_NOR_v2_0/C_bar.n2 GND 0.17fF $ **FLOATING
C633 EESPFAL_3in_NOR_v2_0/C_bar.t4 GND 0.04fF
C634 EESPFAL_3in_NOR_v2_0/C_bar.t3 GND 0.04fF
C635 EESPFAL_3in_NOR_v2_0/C_bar.n3 GND 0.11fF $ **FLOATING
C636 EESPFAL_3in_NOR_v2_0/C_bar.n4 GND 0.12fF $ **FLOATING
C637 EESPFAL_3in_NOR_v2_0/C_bar.t7 GND 0.06fF
C638 EESPFAL_3in_NOR_v2_0/C_bar.t8 GND 0.05fF
C639 EESPFAL_3in_NOR_v2_0/C_bar.t5 GND 0.04fF
C640 EESPFAL_3in_NOR_v2_0/C_bar.n5 GND 0.06fF $ **FLOATING
C641 EESPFAL_3in_NOR_v2_0/C_bar.n6 GND 0.04fF $ **FLOATING
C642 s1.t4 GND 0.04fF
C643 s1.t6 GND 0.04fF
C644 s1.n0 GND 0.15fF $ **FLOATING
C645 s1.t5 GND 0.19fF
C646 s1.t1 GND 0.04fF
C647 s1.t2 GND 0.04fF
C648 s1.n1 GND 0.14fF $ **FLOATING
C649 s1.t3 GND 0.04fF
C650 s1.t0 GND 0.04fF
C651 s1.n2 GND 0.15fF $ **FLOATING
C652 s1.t8 GND 0.06fF
C653 s1.t9 GND 0.06fF
C654 s1.t7 GND 0.03fF
C655 s1.n3 GND 0.06fF $ **FLOATING
C656 s1.n4 GND 0.20fF $ **FLOATING
C657 s1.n5 GND 0.17fF $ **FLOATING
C658 s1.n6 GND 0.14fF $ **FLOATING
C659 s1_bar.t0 GND 0.05fF
C660 s1_bar.t1 GND 0.05fF
C661 s1_bar.n0 GND 0.12fF $ **FLOATING
C662 s1_bar.t2 GND 0.05fF
C663 s1_bar.t3 GND 0.05fF
C664 s1_bar.n1 GND 0.14fF $ **FLOATING
C665 s1_bar.t4 GND 0.27fF
C666 s1_bar.n2 GND 0.19fF $ **FLOATING
C667 s1_bar.n3 GND 0.13fF $ **FLOATING
C668 s1_bar.t5 GND 0.06fF
C669 s1_bar.t7 GND 0.06fF
C670 s1_bar.t6 GND 0.04fF
C671 s1_bar.n4 GND 0.07fF $ **FLOATING
C672 s1_bar.n5 GND 0.05fF $ **FLOATING
C673 Dis3.t0 GND 0.08fF
C674 Dis3.t1 GND 0.08fF
C675 Dis3.n0 GND 0.40fF $ **FLOATING
C676 EESPFAL_3in_NOR_v2_0/C.t3 GND 0.04fF
C677 EESPFAL_3in_NOR_v2_0/C.t2 GND 0.04fF
C678 EESPFAL_3in_NOR_v2_0/C.n0 GND 0.13fF $ **FLOATING
C679 EESPFAL_3in_NOR_v2_0/C.t1 GND 0.16fF
C680 EESPFAL_3in_NOR_v2_0/C.t7 GND 0.05fF
C681 EESPFAL_3in_NOR_v2_0/C.n1 GND 0.77fF $ **FLOATING
C682 EESPFAL_3in_NOR_v2_0/C.n2 GND 0.18fF $ **FLOATING
C683 EESPFAL_3in_NOR_v2_0/C.t0 GND 0.04fF
C684 EESPFAL_3in_NOR_v2_0/C.t4 GND 0.04fF
C685 EESPFAL_3in_NOR_v2_0/C.n3 GND 0.12fF $ **FLOATING
C686 EESPFAL_3in_NOR_v2_0/C.n4 GND 0.11fF $ **FLOATING
C687 EESPFAL_3in_NOR_v2_0/C.n5 GND 0.11fF $ **FLOATING
C688 EESPFAL_3in_NOR_v2_0/C.t6 GND 0.06fF
C689 EESPFAL_3in_NOR_v2_0/C.t5 GND 0.06fF
C690 EESPFAL_3in_NOR_v2_0/C.t8 GND 0.03fF
C691 EESPFAL_3in_NOR_v2_0/C.n6 GND 0.06fF $ **FLOATING
C692 EESPFAL_3in_NOR_v2_0/C.n7 GND 0.03fF $ **FLOATING
C693 EESPFAL_INV4_0/OUT_bar GND 0.01fF $ **FLOATING
C694 x1_bar.t2 GND 0.22fF
C695 x1_bar.t0 GND 0.44fF
C696 x1_bar.t1 GND 0.25fF
C697 x1_bar.n0 GND 2.34fF $ **FLOATING
C698 x1_bar.n1 GND 4.88fF $ **FLOATING
C699 EESPFAL_3in_NAND_v2_0/B_bar GND 0.71fF $ **FLOATING
C700 x1.t1 GND 0.46fF
C701 x1.t2 GND 0.28fF
C702 x1.t0 GND 0.24fF
C703 x1.n0 GND 2.12fF $ **FLOATING
C704 x1.n1 GND 4.42fF $ **FLOATING
C705 EESPFAL_3in_NAND_v2_0/B GND 1.92fF $ **FLOATING
C706 x3.t3 GND 0.18fF
C707 x3.t0 GND 0.17fF
C708 x3.n0 GND 2.07fF $ **FLOATING
C709 x3.t2 GND 0.18fF
C710 x3.t1 GND 0.22fF
C711 EESPFAL_3in_NAND_v2_0/A_bar GND 0.61fF $ **FLOATING
C712 x3.n1 GND 4.00fF $ **FLOATING
C713 EESPFAL_XOR_v3_1/B GND 0.26fF $ **FLOATING
C714 CLK3.t3 GND 0.02fF
C715 CLK3.t11 GND 0.02fF
C716 CLK3.n0 GND 0.05fF $ **FLOATING
C717 CLK3.t1 GND 0.02fF
C718 CLK3.t4 GND 0.04fF
C719 CLK3.n1 GND 0.06fF $ **FLOATING
C720 CLK3.n2 GND 0.17fF $ **FLOATING
C721 CLK3.n3 GND 0.03fF $ **FLOATING
C722 CLK3.n4 GND 0.01fF $ **FLOATING
C723 CLK3.n5 GND 0.01fF $ **FLOATING
C724 CLK3.n6 GND 0.01fF $ **FLOATING
C725 CLK3.n7 GND 0.03fF $ **FLOATING
C726 CLK3.n8 GND 0.01fF $ **FLOATING
C727 CLK3.n9 GND 0.01fF $ **FLOATING
C728 CLK3.n10 GND 0.01fF $ **FLOATING
C729 CLK3.n11 GND 0.03fF $ **FLOATING
C730 CLK3.n12 GND 0.01fF $ **FLOATING
C731 CLK3.n13 GND 0.01fF $ **FLOATING
C732 CLK3.n14 GND 0.01fF $ **FLOATING
C733 CLK3.n15 GND 0.03fF $ **FLOATING
C734 CLK3.n16 GND 0.01fF $ **FLOATING
C735 CLK3.n17 GND 0.01fF $ **FLOATING
C736 CLK3.n18 GND 0.01fF $ **FLOATING
C737 CLK3.n19 GND 0.03fF $ **FLOATING
C738 CLK3.n20 GND 0.01fF $ **FLOATING
C739 CLK3.n21 GND 0.01fF $ **FLOATING
C740 CLK3.n22 GND 0.01fF $ **FLOATING
C741 CLK3.n23 GND 0.03fF $ **FLOATING
C742 CLK3.n24 GND 0.01fF $ **FLOATING
C743 CLK3.n25 GND 0.01fF $ **FLOATING
C744 CLK3.n26 GND 0.01fF $ **FLOATING
C745 CLK3.n27 GND 0.06fF $ **FLOATING
C746 CLK3.n28 GND 0.01fF $ **FLOATING
C747 CLK3.n29 GND 0.01fF $ **FLOATING
C748 CLK3.n30 GND 0.01fF $ **FLOATING
C749 CLK3.n31 GND 0.08fF $ **FLOATING
C750 CLK3.n32 GND 0.01fF $ **FLOATING
C751 CLK3.n33 GND 0.01fF $ **FLOATING
C752 CLK3.n34 GND 0.01fF $ **FLOATING
C753 CLK3.n35 GND 0.14fF $ **FLOATING
C754 CLK3.t0 GND 0.04fF
C755 CLK3.n36 GND 0.05fF $ **FLOATING
C756 CLK3.n37 GND 0.01fF $ **FLOATING
C757 CLK3.n38 GND 0.01fF $ **FLOATING
C758 CLK3.n39 GND 0.01fF $ **FLOATING
C759 CLK3.n40 GND 0.08fF $ **FLOATING
C760 CLK3.n41 GND 0.01fF $ **FLOATING
C761 CLK3.n42 GND 0.01fF $ **FLOATING
C762 CLK3.n43 GND 0.01fF $ **FLOATING
C763 CLK3.t2 GND 0.04fF
C764 CLK3.n44 GND 0.04fF $ **FLOATING
C765 CLK3.n45 GND 0.01fF $ **FLOATING
C766 CLK3.n46 GND 0.01fF $ **FLOATING
C767 CLK3.n47 GND 0.01fF $ **FLOATING
C768 CLK3.n48 GND 0.08fF $ **FLOATING
C769 CLK3.n49 GND 0.01fF $ **FLOATING
C770 CLK3.n50 GND 0.01fF $ **FLOATING
C771 CLK3.n51 GND 0.08fF $ **FLOATING
C772 CLK3.t6 GND 0.02fF
C773 CLK3.t9 GND 0.02fF
C774 CLK3.t7 GND 0.02fF
C775 CLK3.n52 GND 0.07fF $ **FLOATING
C776 CLK3.t8 GND 0.04fF
C777 CLK3.n53 GND 0.06fF $ **FLOATING
C778 CLK3.n54 GND 0.12fF $ **FLOATING
C779 CLK3.n55 GND 0.16fF $ **FLOATING
C780 CLK3.n56 GND 0.03fF $ **FLOATING
C781 CLK3.n57 GND 0.01fF $ **FLOATING
C782 CLK3.n58 GND 0.01fF $ **FLOATING
C783 CLK3.n59 GND 0.01fF $ **FLOATING
C784 CLK3.n60 GND 0.03fF $ **FLOATING
C785 CLK3.n61 GND 0.01fF $ **FLOATING
C786 CLK3.n62 GND 0.01fF $ **FLOATING
C787 CLK3.n63 GND 0.01fF $ **FLOATING
C788 CLK3.n64 GND 0.03fF $ **FLOATING
C789 CLK3.n65 GND 0.01fF $ **FLOATING
C790 CLK3.n66 GND 0.01fF $ **FLOATING
C791 CLK3.n67 GND 0.01fF $ **FLOATING
C792 CLK3.n68 GND 0.03fF $ **FLOATING
C793 CLK3.n69 GND 0.01fF $ **FLOATING
C794 CLK3.n70 GND 0.01fF $ **FLOATING
C795 CLK3.n71 GND 0.01fF $ **FLOATING
C796 CLK3.n72 GND 0.09fF $ **FLOATING
C797 CLK3.n73 GND 0.03fF $ **FLOATING
C798 CLK3.n74 GND 0.01fF $ **FLOATING
C799 CLK3.n75 GND 0.01fF $ **FLOATING
C800 CLK3.n76 GND 0.01fF $ **FLOATING
C801 CLK3.n77 GND 0.03fF $ **FLOATING
C802 CLK3.n78 GND 0.01fF $ **FLOATING
C803 CLK3.n79 GND 0.01fF $ **FLOATING
C804 CLK3.n80 GND 0.01fF $ **FLOATING
C805 CLK3.n81 GND 0.06fF $ **FLOATING
C806 CLK3.n82 GND 0.01fF $ **FLOATING
C807 CLK3.n83 GND 0.01fF $ **FLOATING
C808 CLK3.n84 GND 0.01fF $ **FLOATING
C809 CLK3.n85 GND 0.08fF $ **FLOATING
C810 CLK3.n86 GND 0.01fF $ **FLOATING
C811 CLK3.n87 GND 0.01fF $ **FLOATING
C812 CLK3.n88 GND 0.01fF $ **FLOATING
C813 CLK3.n89 GND 0.14fF $ **FLOATING
C814 CLK3.t5 GND 0.04fF
C815 CLK3.n90 GND 0.05fF $ **FLOATING
C816 CLK3.n91 GND 0.01fF $ **FLOATING
C817 CLK3.n92 GND 0.01fF $ **FLOATING
C818 CLK3.n93 GND 0.01fF $ **FLOATING
C819 CLK3.n94 GND 0.08fF $ **FLOATING
C820 CLK3.n95 GND 0.01fF $ **FLOATING
C821 CLK3.n96 GND 0.01fF $ **FLOATING
C822 CLK3.n97 GND 0.01fF $ **FLOATING
C823 CLK3.t10 GND 0.04fF
C824 CLK3.n98 GND 0.04fF $ **FLOATING
C825 CLK3.n99 GND 0.01fF $ **FLOATING
C826 CLK3.n100 GND 0.01fF $ **FLOATING
C827 CLK3.n101 GND 0.01fF $ **FLOATING
C828 EESPFAL_NAND_v3_0/OUT_bar.t6 GND 0.04fF
C829 EESPFAL_3in_NOR_v2_0/A_bar GND 0.54fF $ **FLOATING
C830 EESPFAL_NAND_v3_0/OUT_bar.t1 GND 0.04fF
C831 EESPFAL_NAND_v3_0/OUT_bar.t0 GND 0.04fF
C832 EESPFAL_NAND_v3_0/OUT_bar.n0 GND 0.11fF $ **FLOATING
C833 EESPFAL_NAND_v3_0/OUT_bar.t5 GND 0.14fF
C834 EESPFAL_NAND_v3_0/OUT_bar.t4 GND 0.20fF
C835 EESPFAL_NAND_v3_0/OUT_bar.n1 GND 0.20fF $ **FLOATING
C836 EESPFAL_NAND_v3_0/OUT_bar.n2 GND 0.09fF $ **FLOATING
C837 EESPFAL_NAND_v3_0/OUT_bar.t2 GND 0.04fF
C838 EESPFAL_NAND_v3_0/OUT_bar.t3 GND 0.04fF
C839 EESPFAL_NAND_v3_0/OUT_bar.n3 GND 0.09fF $ **FLOATING
C840 EESPFAL_NAND_v3_0/OUT_bar.n4 GND 0.10fF $ **FLOATING
C841 EESPFAL_NAND_v3_0/OUT_bar.t9 GND 0.05fF
C842 EESPFAL_NAND_v3_0/OUT_bar.t8 GND 0.04fF
C843 EESPFAL_NAND_v3_0/OUT_bar.t7 GND 0.03fF
C844 EESPFAL_NAND_v3_0/OUT_bar.n5 GND 0.05fF $ **FLOATING
C845 EESPFAL_NAND_v3_0/OUT_bar.n6 GND 0.04fF $ **FLOATING
C846 EESPFAL_NAND_v3_1/A.t8 GND 0.13fF
C847 EESPFAL_NAND_v3_1/A.t3 GND 0.21fF
C848 EESPFAL_NAND_v3_1/A.t4 GND 0.21fF
C849 EESPFAL_NAND_v3_1/A.t5 GND 0.05fF
C850 EESPFAL_NAND_v3_1/A.t0 GND 0.05fF
C851 EESPFAL_NAND_v3_1/A.n0 GND 0.16fF $ **FLOATING
C852 EESPFAL_NAND_v3_1/A.t6 GND 0.04fF
C853 EESPFAL_NAND_v3_1/A.t7 GND 0.06fF
C854 EESPFAL_NAND_v3_1/A.t9 GND 0.07fF
C855 EESPFAL_NAND_v3_1/A.n1 GND 0.07fF $ **FLOATING
C856 EESPFAL_XOR_v3_1/OUT GND 0.01fF $ **FLOATING
C857 EESPFAL_NAND_v3_1/A.n2 GND 0.04fF $ **FLOATING
C858 EESPFAL_NAND_v3_1/A.t2 GND 0.05fF
C859 EESPFAL_NAND_v3_1/A.t1 GND 0.05fF
C860 EESPFAL_NAND_v3_1/A.n3 GND 0.15fF $ **FLOATING
C861 EESPFAL_NAND_v3_1/A.n4 GND 0.22fF $ **FLOATING
C862 EESPFAL_NAND_v3_1/A.n5 GND 0.22fF $ **FLOATING
C863 EESPFAL_NAND_v3_1/A.n6 GND 0.31fF $ **FLOATING
C864 EESPFAL_XOR_v3_1/OUT_bar GND 0.32fF $ **FLOATING
C865 EESPFAL_NAND_v3_1/A_bar.t8 GND 0.07fF
C866 EESPFAL_NAND_v3_1/A_bar.t5 GND 0.05fF
C867 EESPFAL_NAND_v3_1/A_bar.t0 GND 0.05fF
C868 EESPFAL_NAND_v3_1/A_bar.n0 GND 0.13fF $ **FLOATING
C869 EESPFAL_NAND_v3_1/A_bar.t2 GND 0.05fF
C870 EESPFAL_NAND_v3_1/A_bar.t4 GND 0.05fF
C871 EESPFAL_NAND_v3_1/A_bar.n1 GND 0.16fF $ **FLOATING
C872 EESPFAL_NAND_v3_1/A_bar.t3 GND 0.20fF
C873 EESPFAL_NAND_v3_1/A_bar.t1 GND 0.34fF
C874 EESPFAL_NAND_v3_1/A_bar.n2 GND 0.30fF $ **FLOATING
C875 EESPFAL_NAND_v3_1/A_bar.n3 GND 0.13fF $ **FLOATING
C876 EESPFAL_NAND_v3_1/A_bar.n4 GND 0.14fF $ **FLOATING
C877 EESPFAL_NAND_v3_1/A_bar.t7 GND 0.05fF
C878 EESPFAL_NAND_v3_1/A_bar.t6 GND 0.07fF
C879 EESPFAL_NAND_v3_1/A_bar.t9 GND 0.06fF
C880 EESPFAL_NAND_v3_1/A_bar.n5 GND 0.07fF $ **FLOATING
C881 EESPFAL_NAND_v3_1/A_bar.n6 GND 0.05fF $ **FLOATING
C882 Dis2.t1 GND 0.12fF
C883 Dis2.t4 GND 0.08fF
C884 Dis2.n0 GND 0.31fF $ **FLOATING
C885 EESPFAL_NAND_v3_1/Dis GND 0.13fF $ **FLOATING
C886 Dis2.t0 GND 0.12fF
C887 Dis2.t3 GND 0.08fF
C888 Dis2.n1 GND 0.31fF $ **FLOATING
C889 Dis2.n2 GND 0.51fF $ **FLOATING
C890 Dis2.n3 GND 1.52fF $ **FLOATING
C891 Dis2.t2 GND 0.08fF
C892 Dis2.n4 GND 0.76fF $ **FLOATING
C893 Dis2.t5 GND 0.08fF
C894 Dis2.n5 GND 0.17fF $ **FLOATING
C895 EESPFAL_INV4_0/Dis GND -0.15fF $ **FLOATING
C896 Dis1.t1 GND 0.21fF
C897 Dis1.t5 GND 0.14fF
C898 Dis1.n0 GND 0.53fF $ **FLOATING
C899 Dis1.t3 GND 0.21fF
C900 Dis1.t0 GND 0.14fF
C901 Dis1.n1 GND 0.53fF $ **FLOATING
C902 EESPFAL_INV4_1/Dis GND 0.60fF $ **FLOATING
C903 Dis1.t8 GND 0.14fF
C904 Dis1.n2 GND 0.87fF $ **FLOATING
C905 Dis1.t2 GND 0.14fF
C906 Dis1.n3 GND 0.28fF $ **FLOATING
C907 EESPFAL_XOR_v3_1/Dis GND 0.26fF $ **FLOATING
C908 Dis1.t9 GND 0.21fF
C909 Dis1.t6 GND 0.14fF
C910 Dis1.n4 GND 0.53fF $ **FLOATING
C911 Dis1.t7 GND 0.14fF
C912 Dis1.n5 GND 0.87fF $ **FLOATING
C913 Dis1.t4 GND 0.14fF
C914 Dis1.n6 GND 0.28fF $ **FLOATING
C915 EESPFAL_XOR_v3_0/Dis GND 0.26fF $ **FLOATING
C916 Dis1.n7 GND 0.83fF $ **FLOATING
C917 Dis1.n8 GND 2.57fF $ **FLOATING
C918 EESPFAL_3in_NAND_v2_0/Dis GND 0.31fF $ **FLOATING
C919 EESPFAL_XOR_v3_0/OUT_bar GND 0.30fF $ **FLOATING
C920 EESPFAL_NAND_v3_0/A.t9 GND 0.12fF
C921 EESPFAL_NAND_v3_0/A.t2 GND 0.04fF
C922 EESPFAL_NAND_v3_0/A.t1 GND 0.04fF
C923 EESPFAL_NAND_v3_0/A.n0 GND 0.13fF $ **FLOATING
C924 EESPFAL_NAND_v3_0/A.t5 GND 0.17fF
C925 EESPFAL_NAND_v3_0/A.t0 GND 0.29fF
C926 EESPFAL_NAND_v3_0/A.n1 GND 0.26fF $ **FLOATING
C927 EESPFAL_NAND_v3_0/A.n2 GND 0.11fF $ **FLOATING
C928 EESPFAL_NAND_v3_0/A.t4 GND 0.04fF
C929 EESPFAL_NAND_v3_0/A.t3 GND 0.04fF
C930 EESPFAL_NAND_v3_0/A.n3 GND 0.11fF $ **FLOATING
C931 EESPFAL_NAND_v3_0/A.n4 GND 0.12fF $ **FLOATING
C932 EESPFAL_NAND_v3_0/A.t6 GND 0.06fF
C933 EESPFAL_NAND_v3_0/A.t8 GND 0.05fF
C934 EESPFAL_NAND_v3_0/A.t7 GND 0.04fF
C935 EESPFAL_NAND_v3_0/A.n5 GND 0.06fF $ **FLOATING
C936 EESPFAL_NAND_v3_0/A.n6 GND 0.04fF $ **FLOATING
C937 EESPFAL_NAND_v3_0/A_bar.t8 GND 0.08fF
C938 EESPFAL_NAND_v3_0/A_bar.t1 GND 0.24fF
C939 EESPFAL_NAND_v3_0/A_bar.t2 GND 0.05fF
C940 EESPFAL_NAND_v3_0/A_bar.t4 GND 0.05fF
C941 EESPFAL_NAND_v3_0/A_bar.n0 GND 0.17fF $ **FLOATING
C942 EESPFAL_NAND_v3_0/A_bar.t5 GND 0.05fF
C943 EESPFAL_NAND_v3_0/A_bar.t3 GND 0.05fF
C944 EESPFAL_NAND_v3_0/A_bar.n1 GND 0.18fF $ **FLOATING
C945 EESPFAL_NAND_v3_0/A_bar.t9 GND 0.07fF
C946 EESPFAL_NAND_v3_0/A_bar.t7 GND 0.08fF
C947 EESPFAL_NAND_v3_0/A_bar.t6 GND 0.04fF
C948 EESPFAL_NAND_v3_0/A_bar.n2 GND 0.08fF $ **FLOATING
C949 EESPFAL_XOR_v3_0/OUT GND 0.01fF $ **FLOATING
C950 EESPFAL_NAND_v3_0/A_bar.n3 GND 0.04fF $ **FLOATING
C951 EESPFAL_NAND_v3_0/A_bar.n4 GND 0.24fF $ **FLOATING
C952 EESPFAL_NAND_v3_0/A_bar.n5 GND 0.24fF $ **FLOATING
C953 EESPFAL_NAND_v3_0/A_bar.t0 GND 0.24fF
C954 EESPFAL_NAND_v3_0/A_bar.n6 GND 0.52fF $ **FLOATING
C955 CLK1.t22 GND 0.03fF
C956 CLK1.t53 GND 0.03fF
C957 CLK1.n0 GND 0.08fF $ **FLOATING
C958 CLK1.t50 GND 0.04fF
C959 CLK1.t29 GND 0.03fF
C960 CLK1.t28 GND 0.03fF
C961 CLK1.n1 GND 0.12fF $ **FLOATING
C962 CLK1.t0 GND 0.05fF
C963 CLK1.t20 GND 0.04fF
C964 EESPFAL_INV4_1/CLK GND 0.01fF $ **FLOATING
C965 CLK1.t8 GND 0.03fF
C966 CLK1.t18 GND 0.03fF
C967 CLK1.n2 GND 0.08fF $ **FLOATING
C968 CLK1.t10 GND 0.04fF
C969 CLK1.t5 GND 0.05fF
C970 CLK1.n3 GND 0.11fF $ **FLOATING
C971 CLK1.n4 GND 0.36fF $ **FLOATING
C972 CLK1.n5 GND 0.06fF $ **FLOATING
C973 CLK1.n6 GND 0.02fF $ **FLOATING
C974 CLK1.n7 GND 0.02fF $ **FLOATING
C975 CLK1.n8 GND 0.02fF $ **FLOATING
C976 CLK1.n9 GND 0.04fF $ **FLOATING
C977 CLK1.n10 GND 0.02fF $ **FLOATING
C978 CLK1.n11 GND 0.02fF $ **FLOATING
C979 CLK1.n12 GND 0.02fF $ **FLOATING
C980 CLK1.n13 GND 0.10fF $ **FLOATING
C981 CLK1.n14 GND 0.02fF $ **FLOATING
C982 CLK1.n15 GND 0.02fF $ **FLOATING
C983 CLK1.n16 GND 0.02fF $ **FLOATING
C984 CLK1.n17 GND 0.14fF $ **FLOATING
C985 CLK1.n18 GND 0.02fF $ **FLOATING
C986 CLK1.n19 GND 0.02fF $ **FLOATING
C987 CLK1.n20 GND 0.01fF $ **FLOATING
C988 CLK1.n21 GND 0.22fF $ **FLOATING
C989 CLK1.t9 GND 0.07fF
C990 CLK1.n22 GND 0.08fF $ **FLOATING
C991 CLK1.n23 GND 0.02fF $ **FLOATING
C992 CLK1.n24 GND 0.02fF $ **FLOATING
C993 CLK1.n25 GND 0.02fF $ **FLOATING
C994 CLK1.n26 GND 0.12fF $ **FLOATING
C995 CLK1.n27 GND 0.02fF $ **FLOATING
C996 CLK1.n28 GND 0.02fF $ **FLOATING
C997 CLK1.n29 GND 0.02fF $ **FLOATING
C998 CLK1.t7 GND 0.07fF
C999 CLK1.n30 GND 0.07fF $ **FLOATING
C1000 CLK1.n31 GND 0.02fF $ **FLOATING
C1001 CLK1.n32 GND 0.02fF $ **FLOATING
C1002 CLK1.n33 GND 0.02fF $ **FLOATING
C1003 CLK1.n34 GND 0.13fF $ **FLOATING
C1004 CLK1.n35 GND 0.13fF $ **FLOATING
C1005 CLK1.n36 GND 0.02fF $ **FLOATING
C1006 CLK1.n37 GND 0.02fF $ **FLOATING
C1007 CLK1.t17 GND 0.07fF
C1008 CLK1.n38 GND 0.07fF $ **FLOATING
C1009 CLK1.n39 GND 0.02fF $ **FLOATING
C1010 CLK1.n40 GND 0.02fF $ **FLOATING
C1011 CLK1.n41 GND 0.02fF $ **FLOATING
C1012 CLK1.n42 GND 0.12fF $ **FLOATING
C1013 CLK1.n43 GND 0.02fF $ **FLOATING
C1014 CLK1.n44 GND 0.02fF $ **FLOATING
C1015 CLK1.n45 GND 0.02fF $ **FLOATING
C1016 CLK1.t19 GND 0.07fF
C1017 CLK1.n46 GND 0.08fF $ **FLOATING
C1018 CLK1.n47 GND 0.02fF $ **FLOATING
C1019 CLK1.n48 GND 0.02fF $ **FLOATING
C1020 CLK1.n49 GND 0.02fF $ **FLOATING
C1021 CLK1.n50 GND 0.22fF $ **FLOATING
C1022 CLK1.n51 GND 0.14fF $ **FLOATING
C1023 CLK1.n52 GND 0.02fF $ **FLOATING
C1024 CLK1.n53 GND 0.02fF $ **FLOATING
C1025 CLK1.n54 GND 0.01fF $ **FLOATING
C1026 CLK1.n55 GND 0.10fF $ **FLOATING
C1027 CLK1.n56 GND 0.02fF $ **FLOATING
C1028 CLK1.n57 GND 0.02fF $ **FLOATING
C1029 CLK1.n58 GND 0.02fF $ **FLOATING
C1030 CLK1.n59 GND 0.04fF $ **FLOATING
C1031 CLK1.n60 GND 0.02fF $ **FLOATING
C1032 CLK1.n61 GND 0.02fF $ **FLOATING
C1033 CLK1.n62 GND 0.02fF $ **FLOATING
C1034 CLK1.n63 GND 0.06fF $ **FLOATING
C1035 CLK1.n64 GND 0.02fF $ **FLOATING
C1036 CLK1.n65 GND 0.02fF $ **FLOATING
C1037 CLK1.n66 GND 0.02fF $ **FLOATING
C1038 CLK1.n67 GND 0.34fF $ **FLOATING
C1039 CLK1.n68 GND 0.12fF $ **FLOATING
C1040 CLK1.n69 GND 0.08fF $ **FLOATING
C1041 CLK1.n70 GND 0.16fF $ **FLOATING
C1042 CLK1.n71 GND 0.09fF $ **FLOATING
C1043 CLK1.n72 GND 0.06fF $ **FLOATING
C1044 CLK1.n73 GND 0.02fF $ **FLOATING
C1045 CLK1.n74 GND 0.02fF $ **FLOATING
C1046 CLK1.n75 GND 0.02fF $ **FLOATING
C1047 CLK1.n76 GND 0.05fF $ **FLOATING
C1048 CLK1.n77 GND 0.02fF $ **FLOATING
C1049 CLK1.n78 GND 0.02fF $ **FLOATING
C1050 CLK1.n79 GND 0.02fF $ **FLOATING
C1051 CLK1.n80 GND 0.04fF $ **FLOATING
C1052 CLK1.n81 GND 0.02fF $ **FLOATING
C1053 CLK1.n82 GND 0.02fF $ **FLOATING
C1054 CLK1.n83 GND 0.01fF $ **FLOATING
C1055 CLK1.n84 GND 0.14fF $ **FLOATING
C1056 CLK1.n85 GND 0.04fF $ **FLOATING
C1057 CLK1.n86 GND 0.02fF $ **FLOATING
C1058 CLK1.n87 GND 0.02fF $ **FLOATING
C1059 CLK1.n88 GND 0.02fF $ **FLOATING
C1060 CLK1.n89 GND 0.04fF $ **FLOATING
C1061 CLK1.n90 GND 0.02fF $ **FLOATING
C1062 CLK1.n91 GND 0.02fF $ **FLOATING
C1063 CLK1.n92 GND 0.02fF $ **FLOATING
C1064 CLK1.n93 GND 0.04fF $ **FLOATING
C1065 CLK1.n94 GND 0.02fF $ **FLOATING
C1066 CLK1.n95 GND 0.02fF $ **FLOATING
C1067 CLK1.n96 GND 0.02fF $ **FLOATING
C1068 CLK1.n97 GND 0.04fF $ **FLOATING
C1069 CLK1.n98 GND 0.02fF $ **FLOATING
C1070 CLK1.n99 GND 0.02fF $ **FLOATING
C1071 CLK1.n100 GND 0.02fF $ **FLOATING
C1072 CLK1.n101 GND 0.10fF $ **FLOATING
C1073 CLK1.n102 GND 0.02fF $ **FLOATING
C1074 CLK1.n103 GND 0.02fF $ **FLOATING
C1075 CLK1.n104 GND 0.02fF $ **FLOATING
C1076 CLK1.n105 GND 0.14fF $ **FLOATING
C1077 CLK1.n106 GND 0.02fF $ **FLOATING
C1078 CLK1.n107 GND 0.02fF $ **FLOATING
C1079 CLK1.n108 GND 0.01fF $ **FLOATING
C1080 CLK1.n109 GND 0.22fF $ **FLOATING
C1081 CLK1.t49 GND 0.07fF
C1082 CLK1.n110 GND 0.08fF $ **FLOATING
C1083 CLK1.n111 GND 0.02fF $ **FLOATING
C1084 CLK1.n112 GND 0.02fF $ **FLOATING
C1085 CLK1.n113 GND 0.02fF $ **FLOATING
C1086 CLK1.n114 GND 0.12fF $ **FLOATING
C1087 CLK1.n115 GND 0.02fF $ **FLOATING
C1088 CLK1.n116 GND 0.02fF $ **FLOATING
C1089 CLK1.n117 GND 0.02fF $ **FLOATING
C1090 CLK1.t21 GND 0.07fF
C1091 CLK1.n118 GND 0.07fF $ **FLOATING
C1092 CLK1.n119 GND 0.02fF $ **FLOATING
C1093 CLK1.n120 GND 0.02fF $ **FLOATING
C1094 CLK1.n121 GND 0.02fF $ **FLOATING
C1095 CLK1.n122 GND 0.13fF $ **FLOATING
C1096 CLK1.n123 GND 0.02fF $ **FLOATING
C1097 CLK1.n124 GND 0.02fF $ **FLOATING
C1098 CLK1.n125 GND 0.13fF $ **FLOATING
C1099 CLK1.t3 GND 0.04fF
C1100 CLK1.t23 GND 0.03fF
C1101 CLK1.t30 GND 0.03fF
C1102 CLK1.n126 GND 0.12fF $ **FLOATING
C1103 CLK1.n127 GND 0.01fF $ **FLOATING
C1104 CLK1.t6 GND 0.03fF
C1105 CLK1.t51 GND 0.03fF
C1106 CLK1.n128 GND 0.12fF $ **FLOATING
C1107 CLK1.t55 GND 0.04fF
C1108 EESPFAL_XOR_v3_0/CLK GND 0.01fF $ **FLOATING
C1109 CLK1.n129 GND 0.13fF $ **FLOATING
C1110 CLK1.n130 GND 0.02fF $ **FLOATING
C1111 CLK1.t47 GND 0.03fF
C1112 CLK1.t32 GND 0.03fF
C1113 CLK1.n131 GND 0.08fF $ **FLOATING
C1114 CLK1.t36 GND 0.04fF
C1115 CLK1.t1 GND 0.03fF
C1116 CLK1.t4 GND 0.03fF
C1117 CLK1.n132 GND 0.12fF $ **FLOATING
C1118 CLK1.t41 GND 0.05fF
C1119 CLK1.t40 GND 0.04fF
C1120 CLK1.n133 GND 0.13fF $ **FLOATING
C1121 CLK1.n134 GND 0.02fF $ **FLOATING
C1122 CLK1.t45 GND 0.03fF
C1123 CLK1.t38 GND 0.03fF
C1124 CLK1.n135 GND 0.08fF $ **FLOATING
C1125 CLK1.t43 GND 0.04fF
C1126 CLK1.t34 GND 0.05fF
C1127 CLK1.n136 GND 0.11fF $ **FLOATING
C1128 CLK1.n137 GND 0.36fF $ **FLOATING
C1129 CLK1.n138 GND 0.06fF $ **FLOATING
C1130 CLK1.n139 GND 0.02fF $ **FLOATING
C1131 CLK1.n140 GND 0.02fF $ **FLOATING
C1132 CLK1.n141 GND 0.02fF $ **FLOATING
C1133 CLK1.n142 GND 0.04fF $ **FLOATING
C1134 CLK1.n143 GND 0.02fF $ **FLOATING
C1135 CLK1.n144 GND 0.02fF $ **FLOATING
C1136 CLK1.n145 GND 0.02fF $ **FLOATING
C1137 CLK1.n146 GND 0.10fF $ **FLOATING
C1138 CLK1.n147 GND 0.02fF $ **FLOATING
C1139 CLK1.n148 GND 0.02fF $ **FLOATING
C1140 CLK1.n149 GND 0.02fF $ **FLOATING
C1141 CLK1.n150 GND 0.14fF $ **FLOATING
C1142 CLK1.n151 GND 0.02fF $ **FLOATING
C1143 CLK1.n152 GND 0.02fF $ **FLOATING
C1144 CLK1.n153 GND 0.01fF $ **FLOATING
C1145 CLK1.n154 GND 0.22fF $ **FLOATING
C1146 CLK1.t42 GND 0.07fF
C1147 CLK1.n155 GND 0.08fF $ **FLOATING
C1148 CLK1.n156 GND 0.02fF $ **FLOATING
C1149 CLK1.n157 GND 0.02fF $ **FLOATING
C1150 CLK1.n158 GND 0.02fF $ **FLOATING
C1151 CLK1.n159 GND 0.12fF $ **FLOATING
C1152 CLK1.n160 GND 0.02fF $ **FLOATING
C1153 CLK1.n161 GND 0.02fF $ **FLOATING
C1154 CLK1.n162 GND 0.02fF $ **FLOATING
C1155 CLK1.t44 GND 0.07fF
C1156 CLK1.n163 GND 0.07fF $ **FLOATING
C1157 CLK1.n164 GND 0.02fF $ **FLOATING
C1158 CLK1.n165 GND 0.02fF $ **FLOATING
C1159 CLK1.n166 GND 0.02fF $ **FLOATING
C1160 CLK1.n167 GND 0.13fF $ **FLOATING
C1161 CLK1.n168 GND 0.02fF $ **FLOATING
C1162 CLK1.t37 GND 0.07fF
C1163 CLK1.n169 GND 0.07fF $ **FLOATING
C1164 CLK1.n170 GND 0.02fF $ **FLOATING
C1165 CLK1.n171 GND 0.02fF $ **FLOATING
C1166 CLK1.n172 GND 0.02fF $ **FLOATING
C1167 CLK1.n173 GND 0.12fF $ **FLOATING
C1168 CLK1.n174 GND 0.02fF $ **FLOATING
C1169 CLK1.n175 GND 0.02fF $ **FLOATING
C1170 CLK1.n176 GND 0.02fF $ **FLOATING
C1171 CLK1.t39 GND 0.07fF
C1172 CLK1.n177 GND 0.08fF $ **FLOATING
C1173 CLK1.n178 GND 0.02fF $ **FLOATING
C1174 CLK1.n179 GND 0.02fF $ **FLOATING
C1175 CLK1.n180 GND 0.02fF $ **FLOATING
C1176 CLK1.n181 GND 0.22fF $ **FLOATING
C1177 CLK1.n182 GND 0.14fF $ **FLOATING
C1178 CLK1.n183 GND 0.02fF $ **FLOATING
C1179 CLK1.n184 GND 0.02fF $ **FLOATING
C1180 CLK1.n185 GND 0.01fF $ **FLOATING
C1181 CLK1.n186 GND 0.10fF $ **FLOATING
C1182 CLK1.n187 GND 0.02fF $ **FLOATING
C1183 CLK1.n188 GND 0.02fF $ **FLOATING
C1184 CLK1.n189 GND 0.02fF $ **FLOATING
C1185 CLK1.n190 GND 0.04fF $ **FLOATING
C1186 CLK1.n191 GND 0.02fF $ **FLOATING
C1187 CLK1.n192 GND 0.02fF $ **FLOATING
C1188 CLK1.n193 GND 0.02fF $ **FLOATING
C1189 CLK1.n194 GND 0.06fF $ **FLOATING
C1190 CLK1.n195 GND 0.02fF $ **FLOATING
C1191 CLK1.n196 GND 0.02fF $ **FLOATING
C1192 CLK1.n197 GND 0.02fF $ **FLOATING
C1193 CLK1.n198 GND 0.34fF $ **FLOATING
C1194 CLK1.n199 GND 0.12fF $ **FLOATING
C1195 CLK1.n200 GND 0.08fF $ **FLOATING
C1196 CLK1.n201 GND 0.16fF $ **FLOATING
C1197 CLK1.n202 GND 0.09fF $ **FLOATING
C1198 CLK1.n203 GND 0.06fF $ **FLOATING
C1199 CLK1.n204 GND 0.02fF $ **FLOATING
C1200 CLK1.n205 GND 0.02fF $ **FLOATING
C1201 CLK1.n206 GND 0.02fF $ **FLOATING
C1202 CLK1.n207 GND 0.05fF $ **FLOATING
C1203 CLK1.n208 GND 0.02fF $ **FLOATING
C1204 CLK1.n209 GND 0.02fF $ **FLOATING
C1205 CLK1.n210 GND 0.02fF $ **FLOATING
C1206 CLK1.n211 GND 0.04fF $ **FLOATING
C1207 CLK1.n212 GND 0.02fF $ **FLOATING
C1208 CLK1.n213 GND 0.02fF $ **FLOATING
C1209 CLK1.n214 GND 0.01fF $ **FLOATING
C1210 CLK1.n215 GND 0.14fF $ **FLOATING
C1211 CLK1.n216 GND 0.04fF $ **FLOATING
C1212 CLK1.n217 GND 0.02fF $ **FLOATING
C1213 CLK1.n218 GND 0.02fF $ **FLOATING
C1214 CLK1.n219 GND 0.02fF $ **FLOATING
C1215 CLK1.n220 GND 0.04fF $ **FLOATING
C1216 CLK1.n221 GND 0.02fF $ **FLOATING
C1217 CLK1.n222 GND 0.02fF $ **FLOATING
C1218 CLK1.n223 GND 0.02fF $ **FLOATING
C1219 CLK1.n224 GND 0.04fF $ **FLOATING
C1220 CLK1.n225 GND 0.02fF $ **FLOATING
C1221 CLK1.n226 GND 0.02fF $ **FLOATING
C1222 CLK1.n227 GND 0.02fF $ **FLOATING
C1223 CLK1.n228 GND 0.04fF $ **FLOATING
C1224 CLK1.n229 GND 0.02fF $ **FLOATING
C1225 CLK1.n230 GND 0.02fF $ **FLOATING
C1226 CLK1.n231 GND 0.02fF $ **FLOATING
C1227 CLK1.n232 GND 0.10fF $ **FLOATING
C1228 CLK1.n233 GND 0.02fF $ **FLOATING
C1229 CLK1.n234 GND 0.02fF $ **FLOATING
C1230 CLK1.n235 GND 0.02fF $ **FLOATING
C1231 CLK1.n236 GND 0.14fF $ **FLOATING
C1232 CLK1.n237 GND 0.02fF $ **FLOATING
C1233 CLK1.n238 GND 0.02fF $ **FLOATING
C1234 CLK1.n239 GND 0.01fF $ **FLOATING
C1235 CLK1.n240 GND 0.22fF $ **FLOATING
C1236 CLK1.t35 GND 0.07fF
C1237 CLK1.n241 GND 0.08fF $ **FLOATING
C1238 CLK1.n242 GND 0.02fF $ **FLOATING
C1239 CLK1.n243 GND 0.02fF $ **FLOATING
C1240 CLK1.n244 GND 0.02fF $ **FLOATING
C1241 CLK1.n245 GND 0.12fF $ **FLOATING
C1242 CLK1.n246 GND 0.02fF $ **FLOATING
C1243 CLK1.n247 GND 0.02fF $ **FLOATING
C1244 CLK1.n248 GND 0.02fF $ **FLOATING
C1245 CLK1.t46 GND 0.07fF
C1246 CLK1.n249 GND 0.07fF $ **FLOATING
C1247 CLK1.n250 GND 0.02fF $ **FLOATING
C1248 CLK1.n251 GND 0.02fF $ **FLOATING
C1249 CLK1.n252 GND 0.02fF $ **FLOATING
C1250 CLK1.n253 GND 0.13fF $ **FLOATING
C1251 CLK1.n254 GND 0.02fF $ **FLOATING
C1252 CLK1.t31 GND 0.07fF
C1253 CLK1.n255 GND 0.07fF $ **FLOATING
C1254 CLK1.n256 GND 0.02fF $ **FLOATING
C1255 CLK1.n257 GND 0.02fF $ **FLOATING
C1256 CLK1.n258 GND 0.02fF $ **FLOATING
C1257 CLK1.n259 GND 0.12fF $ **FLOATING
C1258 CLK1.n260 GND 0.02fF $ **FLOATING
C1259 CLK1.n261 GND 0.02fF $ **FLOATING
C1260 CLK1.n262 GND 0.02fF $ **FLOATING
C1261 CLK1.t54 GND 0.07fF
C1262 CLK1.n263 GND 0.08fF $ **FLOATING
C1263 CLK1.n264 GND 0.02fF $ **FLOATING
C1264 CLK1.n265 GND 0.02fF $ **FLOATING
C1265 CLK1.n266 GND 0.02fF $ **FLOATING
C1266 CLK1.n267 GND 0.22fF $ **FLOATING
C1267 CLK1.n268 GND 0.14fF $ **FLOATING
C1268 CLK1.n269 GND 0.02fF $ **FLOATING
C1269 CLK1.n270 GND 0.02fF $ **FLOATING
C1270 CLK1.n271 GND 0.01fF $ **FLOATING
C1271 CLK1.n272 GND 0.10fF $ **FLOATING
C1272 CLK1.n273 GND 0.02fF $ **FLOATING
C1273 CLK1.n274 GND 0.02fF $ **FLOATING
C1274 CLK1.n275 GND 0.02fF $ **FLOATING
C1275 CLK1.n276 GND 0.04fF $ **FLOATING
C1276 CLK1.n277 GND 0.02fF $ **FLOATING
C1277 CLK1.n278 GND 0.02fF $ **FLOATING
C1278 CLK1.n279 GND 0.02fF $ **FLOATING
C1279 CLK1.n280 GND 0.04fF $ **FLOATING
C1280 CLK1.n281 GND 0.02fF $ **FLOATING
C1281 CLK1.n282 GND 0.02fF $ **FLOATING
C1282 CLK1.n283 GND 0.02fF $ **FLOATING
C1283 CLK1.n284 GND 0.04fF $ **FLOATING
C1284 CLK1.n285 GND 0.02fF $ **FLOATING
C1285 CLK1.n286 GND 0.02fF $ **FLOATING
C1286 CLK1.n287 GND 0.02fF $ **FLOATING
C1287 CLK1.n288 GND 0.04fF $ **FLOATING
C1288 CLK1.n289 GND 0.02fF $ **FLOATING
C1289 CLK1.n290 GND 0.02fF $ **FLOATING
C1290 CLK1.n291 GND 0.02fF $ **FLOATING
C1291 CLK1.n292 GND 0.14fF $ **FLOATING
C1292 CLK1.n293 GND 0.04fF $ **FLOATING
C1293 CLK1.n294 GND 0.02fF $ **FLOATING
C1294 CLK1.n295 GND 0.02fF $ **FLOATING
C1295 CLK1.n296 GND 0.01fF $ **FLOATING
C1296 CLK1.n297 GND 0.05fF $ **FLOATING
C1297 CLK1.n298 GND 0.02fF $ **FLOATING
C1298 CLK1.n299 GND 0.02fF $ **FLOATING
C1299 CLK1.n300 GND 0.02fF $ **FLOATING
C1300 CLK1.n301 GND 0.06fF $ **FLOATING
C1301 CLK1.n302 GND 0.02fF $ **FLOATING
C1302 CLK1.n303 GND 0.02fF $ **FLOATING
C1303 CLK1.n304 GND 0.02fF $ **FLOATING
C1304 CLK1.n305 GND 0.01fF $ **FLOATING
C1305 CLK1.n306 GND 0.01fF $ **FLOATING
C1306 CLK1.n307 GND 0.14fF $ **FLOATING
C1307 CLK1.n308 GND 0.01fF $ **FLOATING
C1308 CLK1.n309 GND 0.02fF $ **FLOATING
C1309 CLK1.n310 GND 0.00fF $ **FLOATING
C1310 CLK1.n311 GND 0.01fF $ **FLOATING
C1311 CLK1.n312 GND 0.28fF $ **FLOATING
C1312 CLK1.n313 GND 0.27fF $ **FLOATING
C1313 CLK1.n314 GND 0.02fF $ **FLOATING
C1314 CLK1.t48 GND 0.06fF
C1315 CLK1.t33 GND 0.03fF
C1316 CLK1.t11 GND 0.03fF
C1317 CLK1.n315 GND 0.12fF $ **FLOATING
C1318 CLK1.t27 GND 0.04fF
C1319 EESPFAL_3in_NAND_v2_0/CLK GND 0.01fF $ **FLOATING
C1320 CLK1.t16 GND 0.03fF
C1321 CLK1.t25 GND 0.03fF
C1322 CLK1.n316 GND 0.08fF $ **FLOATING
C1323 CLK1.t14 GND 0.04fF
C1324 CLK1.t12 GND 0.06fF
C1325 CLK1.n317 GND 0.10fF $ **FLOATING
C1326 CLK1.n318 GND 0.27fF $ **FLOATING
C1327 CLK1.n319 GND 0.05fF $ **FLOATING
C1328 CLK1.n320 GND 0.02fF $ **FLOATING
C1329 CLK1.n321 GND 0.02fF $ **FLOATING
C1330 CLK1.n322 GND 0.02fF $ **FLOATING
C1331 CLK1.n323 GND 0.05fF $ **FLOATING
C1332 CLK1.n324 GND 0.02fF $ **FLOATING
C1333 CLK1.n325 GND 0.02fF $ **FLOATING
C1334 CLK1.n326 GND 0.02fF $ **FLOATING
C1335 CLK1.n327 GND 0.04fF $ **FLOATING
C1336 CLK1.n328 GND 0.02fF $ **FLOATING
C1337 CLK1.n329 GND 0.02fF $ **FLOATING
C1338 CLK1.n330 GND 0.02fF $ **FLOATING
C1339 CLK1.n331 GND 0.04fF $ **FLOATING
C1340 CLK1.n332 GND 0.02fF $ **FLOATING
C1341 CLK1.n333 GND 0.02fF $ **FLOATING
C1342 CLK1.n334 GND 0.02fF $ **FLOATING
C1343 CLK1.n335 GND 0.04fF $ **FLOATING
C1344 CLK1.n336 GND 0.02fF $ **FLOATING
C1345 CLK1.n337 GND 0.02fF $ **FLOATING
C1346 CLK1.n338 GND 0.02fF $ **FLOATING
C1347 CLK1.n339 GND 0.04fF $ **FLOATING
C1348 CLK1.n340 GND 0.02fF $ **FLOATING
C1349 CLK1.n341 GND 0.02fF $ **FLOATING
C1350 CLK1.n342 GND 0.02fF $ **FLOATING
C1351 CLK1.n343 GND 0.10fF $ **FLOATING
C1352 CLK1.n344 GND 0.02fF $ **FLOATING
C1353 CLK1.n345 GND 0.02fF $ **FLOATING
C1354 CLK1.n346 GND 0.02fF $ **FLOATING
C1355 CLK1.n347 GND 0.14fF $ **FLOATING
C1356 CLK1.n348 GND 0.02fF $ **FLOATING
C1357 CLK1.n349 GND 0.02fF $ **FLOATING
C1358 CLK1.n350 GND 0.01fF $ **FLOATING
C1359 CLK1.n351 GND 0.22fF $ **FLOATING
C1360 CLK1.t13 GND 0.07fF
C1361 CLK1.n352 GND 0.08fF $ **FLOATING
C1362 CLK1.n353 GND 0.02fF $ **FLOATING
C1363 CLK1.n354 GND 0.02fF $ **FLOATING
C1364 CLK1.n355 GND 0.02fF $ **FLOATING
C1365 CLK1.n356 GND 0.12fF $ **FLOATING
C1366 CLK1.n357 GND 0.02fF $ **FLOATING
C1367 CLK1.n358 GND 0.02fF $ **FLOATING
C1368 CLK1.n359 GND 0.02fF $ **FLOATING
C1369 CLK1.t15 GND 0.07fF
C1370 CLK1.n360 GND 0.07fF $ **FLOATING
C1371 CLK1.n361 GND 0.02fF $ **FLOATING
C1372 CLK1.n362 GND 0.02fF $ **FLOATING
C1373 CLK1.n363 GND 0.02fF $ **FLOATING
C1374 CLK1.n364 GND 0.13fF $ **FLOATING
C1375 CLK1.n365 GND 0.13fF $ **FLOATING
C1376 CLK1.n366 GND 0.02fF $ **FLOATING
C1377 CLK1.n367 GND 0.02fF $ **FLOATING
C1378 CLK1.t24 GND 0.07fF
C1379 CLK1.n368 GND 0.07fF $ **FLOATING
C1380 CLK1.n369 GND 0.02fF $ **FLOATING
C1381 CLK1.n370 GND 0.02fF $ **FLOATING
C1382 CLK1.n371 GND 0.02fF $ **FLOATING
C1383 CLK1.n372 GND 0.12fF $ **FLOATING
C1384 CLK1.n373 GND 0.02fF $ **FLOATING
C1385 CLK1.n374 GND 0.02fF $ **FLOATING
C1386 CLK1.n375 GND 0.02fF $ **FLOATING
C1387 CLK1.t26 GND 0.07fF
C1388 CLK1.n376 GND 0.08fF $ **FLOATING
C1389 CLK1.n377 GND 0.02fF $ **FLOATING
C1390 CLK1.n378 GND 0.02fF $ **FLOATING
C1391 CLK1.n379 GND 0.02fF $ **FLOATING
C1392 CLK1.n380 GND 0.22fF $ **FLOATING
C1393 CLK1.n381 GND 0.14fF $ **FLOATING
C1394 CLK1.n382 GND 0.02fF $ **FLOATING
C1395 CLK1.n383 GND 0.02fF $ **FLOATING
C1396 CLK1.n384 GND 0.01fF $ **FLOATING
C1397 CLK1.n385 GND 0.10fF $ **FLOATING
C1398 CLK1.n386 GND 0.02fF $ **FLOATING
C1399 CLK1.n387 GND 0.02fF $ **FLOATING
C1400 CLK1.n388 GND 0.02fF $ **FLOATING
C1401 CLK1.n389 GND 0.04fF $ **FLOATING
C1402 CLK1.n390 GND 0.02fF $ **FLOATING
C1403 CLK1.n391 GND 0.02fF $ **FLOATING
C1404 CLK1.n392 GND 0.02fF $ **FLOATING
C1405 CLK1.n393 GND 0.04fF $ **FLOATING
C1406 CLK1.n394 GND 0.02fF $ **FLOATING
C1407 CLK1.n395 GND 0.02fF $ **FLOATING
C1408 CLK1.n396 GND 0.02fF $ **FLOATING
C1409 CLK1.n397 GND 0.14fF $ **FLOATING
C1410 CLK1.n398 GND 0.04fF $ **FLOATING
C1411 CLK1.n399 GND 0.02fF $ **FLOATING
C1412 CLK1.n400 GND 0.02fF $ **FLOATING
C1413 CLK1.n401 GND 0.01fF $ **FLOATING
C1414 CLK1.n402 GND 0.04fF $ **FLOATING
C1415 CLK1.n403 GND 0.02fF $ **FLOATING
C1416 CLK1.n404 GND 0.02fF $ **FLOATING
C1417 CLK1.n405 GND 0.02fF $ **FLOATING
C1418 CLK1.n406 GND 0.05fF $ **FLOATING
C1419 CLK1.n407 GND 0.02fF $ **FLOATING
C1420 CLK1.n408 GND 0.02fF $ **FLOATING
C1421 CLK1.n409 GND 0.02fF $ **FLOATING
C1422 CLK1.n410 GND 0.05fF $ **FLOATING
C1423 CLK1.n411 GND 0.02fF $ **FLOATING
C1424 CLK1.n412 GND 0.02fF $ **FLOATING
C1425 CLK1.n413 GND 0.02fF $ **FLOATING
C1426 CLK1.n414 GND 0.26fF $ **FLOATING
C1427 CLK1.n415 GND 0.10fF $ **FLOATING
C1428 CLK1.n416 GND 0.06fF $ **FLOATING
C1429 CLK1.n417 GND 0.10fF $ **FLOATING
C1430 CLK1.n418 GND 0.01fF $ **FLOATING
C1431 CLK1.n419 GND 0.00fF $ **FLOATING
C1432 CLK1.n420 GND 0.01fF $ **FLOATING
C1433 CLK1.n421 GND 0.14fF $ **FLOATING
C1434 CLK1.n422 GND 0.01fF $ **FLOATING
C1435 CLK1.n423 GND 0.01fF $ **FLOATING
C1436 CLK1.n424 GND 0.06fF $ **FLOATING
C1437 CLK1.n425 GND 0.02fF $ **FLOATING
C1438 CLK1.n426 GND 0.02fF $ **FLOATING
C1439 CLK1.n427 GND 0.02fF $ **FLOATING
C1440 CLK1.n428 GND 0.05fF $ **FLOATING
C1441 CLK1.n429 GND 0.02fF $ **FLOATING
C1442 CLK1.n430 GND 0.02fF $ **FLOATING
C1443 CLK1.n431 GND 0.02fF $ **FLOATING
C1444 CLK1.n432 GND 0.04fF $ **FLOATING
C1445 CLK1.n433 GND 0.02fF $ **FLOATING
C1446 CLK1.n434 GND 0.02fF $ **FLOATING
C1447 CLK1.n435 GND 0.01fF $ **FLOATING
C1448 CLK1.n436 GND 0.14fF $ **FLOATING
C1449 CLK1.n437 GND 0.04fF $ **FLOATING
C1450 CLK1.n438 GND 0.02fF $ **FLOATING
C1451 CLK1.n439 GND 0.02fF $ **FLOATING
C1452 CLK1.n440 GND 0.02fF $ **FLOATING
C1453 CLK1.n441 GND 0.04fF $ **FLOATING
C1454 CLK1.n442 GND 0.02fF $ **FLOATING
C1455 CLK1.n443 GND 0.02fF $ **FLOATING
C1456 CLK1.n444 GND 0.02fF $ **FLOATING
C1457 CLK1.n445 GND 0.04fF $ **FLOATING
C1458 CLK1.n446 GND 0.02fF $ **FLOATING
C1459 CLK1.n447 GND 0.02fF $ **FLOATING
C1460 CLK1.n448 GND 0.02fF $ **FLOATING
C1461 CLK1.n449 GND 0.04fF $ **FLOATING
C1462 CLK1.n450 GND 0.02fF $ **FLOATING
C1463 CLK1.n451 GND 0.02fF $ **FLOATING
C1464 CLK1.n452 GND 0.02fF $ **FLOATING
C1465 CLK1.n453 GND 0.10fF $ **FLOATING
C1466 CLK1.n454 GND 0.02fF $ **FLOATING
C1467 CLK1.n455 GND 0.02fF $ **FLOATING
C1468 CLK1.n456 GND 0.02fF $ **FLOATING
C1469 CLK1.n457 GND 0.14fF $ **FLOATING
C1470 CLK1.n458 GND 0.02fF $ **FLOATING
C1471 CLK1.n459 GND 0.02fF $ **FLOATING
C1472 CLK1.n460 GND 0.01fF $ **FLOATING
C1473 CLK1.n461 GND 0.22fF $ **FLOATING
C1474 CLK1.t2 GND 0.07fF
C1475 CLK1.n462 GND 0.08fF $ **FLOATING
C1476 CLK1.n463 GND 0.02fF $ **FLOATING
C1477 CLK1.n464 GND 0.02fF $ **FLOATING
C1478 CLK1.n465 GND 0.02fF $ **FLOATING
C1479 CLK1.n466 GND 0.12fF $ **FLOATING
C1480 CLK1.n467 GND 0.02fF $ **FLOATING
C1481 CLK1.n468 GND 0.02fF $ **FLOATING
C1482 CLK1.n469 GND 0.02fF $ **FLOATING
C1483 CLK1.t52 GND 0.07fF
C1484 CLK1.n470 GND 0.07fF $ **FLOATING
C1485 CLK1.n471 GND 0.02fF $ **FLOATING
C1486 CLK1.n472 GND 0.02fF $ **FLOATING
C1487 CLK1.n473 GND 0.02fF $ **FLOATING
C1488 EESPFAL_XOR_v3_1/CLK GND 0.01fF $ **FLOATING
C1489 CLK2.t1 GND 0.02fF
C1490 CLK2.t22 GND 0.02fF
C1491 CLK2.n0 GND 0.05fF $ **FLOATING
C1492 CLK2.t3 GND 0.03fF
C1493 CLK2.t28 GND 0.02fF
C1494 CLK2.n1 GND 0.05fF $ **FLOATING
C1495 CLK2.n2 GND 0.01fF $ **FLOATING
C1496 CLK2.n3 GND 0.01fF $ **FLOATING
C1497 CLK2.n4 GND 0.01fF $ **FLOATING
C1498 CLK2.n5 GND 0.07fF $ **FLOATING
C1499 CLK2.t9 GND 0.03fF
C1500 CLK2.t11 GND 0.02fF
C1501 CLK2.t14 GND 0.02fF
C1502 CLK2.n6 GND 0.05fF $ **FLOATING
C1503 EESPFAL_NAND_v3_1/CLK GND 0.01fF $ **FLOATING
C1504 CLK2.t16 GND 0.03fF
C1505 CLK2.t7 GND 0.02fF
C1506 CLK2.t6 GND 0.02fF
C1507 CLK2.n7 GND 0.08fF $ **FLOATING
C1508 CLK2.n8 GND 0.07fF $ **FLOATING
C1509 CLK2.n9 GND 0.08fF $ **FLOATING
C1510 CLK2.t12 GND 0.04fF
C1511 CLK2.t20 GND 0.03fF
C1512 CLK2.t18 GND 0.02fF
C1513 CLK2.t30 GND 0.02fF
C1514 CLK2.n10 GND 0.05fF $ **FLOATING
C1515 EESPFAL_INV4_0/CLK GND 0.01fF $ **FLOATING
C1516 CLK2.t26 GND 0.03fF
C1517 CLK2.t5 GND 0.04fF
C1518 CLK2.n11 GND 0.08fF $ **FLOATING
C1519 CLK2.n12 GND 0.24fF $ **FLOATING
C1520 CLK2.n13 GND 0.04fF $ **FLOATING
C1521 CLK2.n14 GND 0.02fF $ **FLOATING
C1522 CLK2.n15 GND 0.01fF $ **FLOATING
C1523 CLK2.n16 GND 0.01fF $ **FLOATING
C1524 CLK2.n17 GND 0.03fF $ **FLOATING
C1525 CLK2.n18 GND 0.02fF $ **FLOATING
C1526 CLK2.n19 GND 0.01fF $ **FLOATING
C1527 CLK2.n20 GND 0.02fF $ **FLOATING
C1528 CLK2.n21 GND 0.07fF $ **FLOATING
C1529 CLK2.n22 GND 0.02fF $ **FLOATING
C1530 CLK2.n23 GND 0.01fF $ **FLOATING
C1531 CLK2.n24 GND 0.02fF $ **FLOATING
C1532 CLK2.n25 GND 0.09fF $ **FLOATING
C1533 CLK2.n26 GND 0.02fF $ **FLOATING
C1534 CLK2.n27 GND 0.01fF $ **FLOATING
C1535 CLK2.n28 GND 0.01fF $ **FLOATING
C1536 CLK2.n29 GND 0.15fF $ **FLOATING
C1537 CLK2.t25 GND 0.05fF
C1538 CLK2.n30 GND 0.05fF $ **FLOATING
C1539 CLK2.n31 GND 0.02fF $ **FLOATING
C1540 CLK2.n32 GND 0.01fF $ **FLOATING
C1541 CLK2.n33 GND 0.01fF $ **FLOATING
C1542 CLK2.n34 GND 0.08fF $ **FLOATING
C1543 CLK2.n35 GND 0.02fF $ **FLOATING
C1544 CLK2.n36 GND 0.01fF $ **FLOATING
C1545 CLK2.n37 GND 0.02fF $ **FLOATING
C1546 CLK2.n38 GND 0.01fF $ **FLOATING
C1547 CLK2.t29 GND 0.05fF
C1548 CLK2.n39 GND 0.05fF $ **FLOATING
C1549 CLK2.n40 GND 0.02fF $ **FLOATING
C1550 CLK2.n41 GND 0.01fF $ **FLOATING
C1551 CLK2.n42 GND 0.09fF $ **FLOATING
C1552 CLK2.n43 GND 0.02fF $ **FLOATING
C1553 CLK2.n44 GND 0.01fF $ **FLOATING
C1554 CLK2.n45 GND 0.09fF $ **FLOATING
C1555 CLK2.t17 GND 0.05fF
C1556 CLK2.n46 GND 0.05fF $ **FLOATING
C1557 CLK2.n47 GND 0.02fF $ **FLOATING
C1558 CLK2.n48 GND 0.01fF $ **FLOATING
C1559 CLK2.n49 GND 0.02fF $ **FLOATING
C1560 CLK2.n50 GND 0.08fF $ **FLOATING
C1561 CLK2.n51 GND 0.02fF $ **FLOATING
C1562 CLK2.n52 GND 0.01fF $ **FLOATING
C1563 CLK2.n53 GND 0.02fF $ **FLOATING
C1564 CLK2.t19 GND 0.05fF
C1565 CLK2.n54 GND 0.05fF $ **FLOATING
C1566 CLK2.n55 GND 0.02fF $ **FLOATING
C1567 CLK2.n56 GND 0.01fF $ **FLOATING
C1568 CLK2.n57 GND 0.01fF $ **FLOATING
C1569 CLK2.n58 GND 0.15fF $ **FLOATING
C1570 CLK2.n59 GND 0.09fF $ **FLOATING
C1571 CLK2.n60 GND 0.02fF $ **FLOATING
C1572 CLK2.n61 GND 0.01fF $ **FLOATING
C1573 CLK2.n62 GND 0.01fF $ **FLOATING
C1574 CLK2.n63 GND 0.07fF $ **FLOATING
C1575 CLK2.n64 GND 0.02fF $ **FLOATING
C1576 CLK2.n65 GND 0.01fF $ **FLOATING
C1577 CLK2.n66 GND 0.02fF $ **FLOATING
C1578 CLK2.n67 GND 0.03fF $ **FLOATING
C1579 CLK2.n68 GND 0.02fF $ **FLOATING
C1580 CLK2.n69 GND 0.01fF $ **FLOATING
C1581 CLK2.n70 GND 0.02fF $ **FLOATING
C1582 CLK2.n71 GND 0.04fF $ **FLOATING
C1583 CLK2.n72 GND 0.02fF $ **FLOATING
C1584 CLK2.n73 GND 0.01fF $ **FLOATING
C1585 CLK2.n74 GND 0.01fF $ **FLOATING
C1586 CLK2.n75 GND 0.23fF $ **FLOATING
C1587 CLK2.n76 GND 0.11fF $ **FLOATING
C1588 CLK2.n77 GND 0.10fF $ **FLOATING
C1589 CLK2.n78 GND 0.04fF $ **FLOATING
C1590 CLK2.n79 GND 0.02fF $ **FLOATING
C1591 CLK2.n80 GND 0.01fF $ **FLOATING
C1592 CLK2.n81 GND 0.02fF $ **FLOATING
C1593 CLK2.n82 GND 0.03fF $ **FLOATING
C1594 CLK2.n83 GND 0.02fF $ **FLOATING
C1595 CLK2.n84 GND 0.01fF $ **FLOATING
C1596 CLK2.n85 GND 0.01fF $ **FLOATING
C1597 CLK2.n86 GND 0.10fF $ **FLOATING
C1598 CLK2.n87 GND 0.03fF $ **FLOATING
C1599 CLK2.n88 GND 0.02fF $ **FLOATING
C1600 CLK2.n89 GND 0.01fF $ **FLOATING
C1601 CLK2.n90 GND 0.01fF $ **FLOATING
C1602 CLK2.n91 GND 0.03fF $ **FLOATING
C1603 CLK2.n92 GND 0.02fF $ **FLOATING
C1604 CLK2.n93 GND 0.01fF $ **FLOATING
C1605 CLK2.n94 GND 0.02fF $ **FLOATING
C1606 CLK2.n95 GND 0.07fF $ **FLOATING
C1607 CLK2.n96 GND 0.02fF $ **FLOATING
C1608 CLK2.n97 GND 0.01fF $ **FLOATING
C1609 CLK2.n98 GND 0.02fF $ **FLOATING
C1610 CLK2.n99 GND 0.09fF $ **FLOATING
C1611 CLK2.n100 GND 0.02fF $ **FLOATING
C1612 CLK2.n101 GND 0.01fF $ **FLOATING
C1613 CLK2.n102 GND 0.01fF $ **FLOATING
C1614 CLK2.n103 GND 0.15fF $ **FLOATING
C1615 CLK2.t15 GND 0.05fF
C1616 CLK2.n104 GND 0.05fF $ **FLOATING
C1617 CLK2.n105 GND 0.02fF $ **FLOATING
C1618 CLK2.n106 GND 0.01fF $ **FLOATING
C1619 CLK2.n107 GND 0.01fF $ **FLOATING
C1620 CLK2.n108 GND 0.08fF $ **FLOATING
C1621 CLK2.n109 GND 0.02fF $ **FLOATING
C1622 CLK2.n110 GND 0.01fF $ **FLOATING
C1623 CLK2.n111 GND 0.02fF $ **FLOATING
C1624 CLK2.n112 GND 0.01fF $ **FLOATING
C1625 CLK2.t13 GND 0.05fF
C1626 CLK2.n113 GND 0.05fF $ **FLOATING
C1627 CLK2.n114 GND 0.02fF $ **FLOATING
C1628 CLK2.n115 GND 0.01fF $ **FLOATING
C1629 CLK2.n116 GND 0.09fF $ **FLOATING
C1630 CLK2.n117 GND 0.02fF $ **FLOATING
C1631 CLK2.n118 GND 0.01fF $ **FLOATING
C1632 CLK2.n119 GND 0.09fF $ **FLOATING
C1633 CLK2.t10 GND 0.05fF
C1634 CLK2.n120 GND 0.05fF $ **FLOATING
C1635 CLK2.n121 GND 0.02fF $ **FLOATING
C1636 CLK2.n122 GND 0.01fF $ **FLOATING
C1637 CLK2.n123 GND 0.02fF $ **FLOATING
C1638 CLK2.n124 GND 0.08fF $ **FLOATING
C1639 CLK2.n125 GND 0.02fF $ **FLOATING
C1640 CLK2.n126 GND 0.01fF $ **FLOATING
C1641 CLK2.n127 GND 0.02fF $ **FLOATING
C1642 CLK2.t8 GND 0.05fF
C1643 CLK2.n128 GND 0.05fF $ **FLOATING
C1644 CLK2.n129 GND 0.02fF $ **FLOATING
C1645 CLK2.n130 GND 0.01fF $ **FLOATING
C1646 CLK2.n131 GND 0.01fF $ **FLOATING
C1647 CLK2.n132 GND 0.15fF $ **FLOATING
C1648 CLK2.n133 GND 0.09fF $ **FLOATING
C1649 CLK2.n134 GND 0.02fF $ **FLOATING
C1650 CLK2.n135 GND 0.01fF $ **FLOATING
C1651 CLK2.n136 GND 0.01fF $ **FLOATING
C1652 CLK2.n137 GND 0.07fF $ **FLOATING
C1653 CLK2.n138 GND 0.02fF $ **FLOATING
C1654 CLK2.n139 GND 0.01fF $ **FLOATING
C1655 CLK2.n140 GND 0.02fF $ **FLOATING
C1656 CLK2.n141 GND 0.03fF $ **FLOATING
C1657 CLK2.n142 GND 0.02fF $ **FLOATING
C1658 CLK2.n143 GND 0.01fF $ **FLOATING
C1659 CLK2.n144 GND 0.02fF $ **FLOATING
C1660 CLK2.n145 GND 0.03fF $ **FLOATING
C1661 CLK2.n146 GND 0.02fF $ **FLOATING
C1662 CLK2.n147 GND 0.01fF $ **FLOATING
C1663 CLK2.n148 GND 0.02fF $ **FLOATING
C1664 CLK2.n149 GND 0.03fF $ **FLOATING
C1665 CLK2.n150 GND 0.02fF $ **FLOATING
C1666 CLK2.n151 GND 0.01fF $ **FLOATING
C1667 CLK2.n152 GND 0.02fF $ **FLOATING
C1668 CLK2.n153 GND 0.04fF $ **FLOATING
C1669 CLK2.n154 GND 0.02fF $ **FLOATING
C1670 CLK2.n155 GND 0.01fF $ **FLOATING
C1671 CLK2.n156 GND 0.01fF $ **FLOATING
C1672 CLK2.n157 GND 0.05fF $ **FLOATING
C1673 CLK2.n158 GND 0.01fF $ **FLOATING
C1674 CLK2.n159 GND 0.04fF $ **FLOATING
C1675 CLK2.n160 GND 0.01fF $ **FLOATING
C1676 CLK2.t4 GND 0.02fF
C1677 CLK2.n161 GND 0.05fF $ **FLOATING
C1678 CLK2.n162 GND 0.01fF $ **FLOATING
C1679 CLK2.n163 GND 0.06fF $ **FLOATING
C1680 CLK2.n164 GND 0.06fF $ **FLOATING
C1681 CLK2.n165 GND 0.01fF $ **FLOATING
C1682 CLK2.n166 GND 0.01fF $ **FLOATING
C1683 CLK2.n167 GND 0.05fF $ **FLOATING
C1684 CLK2.n168 GND 0.01fF $ **FLOATING
C1685 CLK2.n169 GND 0.07fF $ **FLOATING
C1686 CLK2.n170 GND 0.01fF $ **FLOATING
C1687 CLK2.n171 GND 0.03fF $ **FLOATING
C1688 CLK2.n172 GND 0.01fF $ **FLOATING
C1689 CLK2.n173 GND 0.04fF $ **FLOATING
C1690 CLK2.n174 GND 0.02fF $ **FLOATING
C1691 CLK2.n175 GND 0.01fF $ **FLOATING
C1692 CLK2.n176 GND 0.01fF $ **FLOATING
C1693 CLK2.n177 GND 0.03fF $ **FLOATING
C1694 CLK2.n178 GND 0.02fF $ **FLOATING
C1695 CLK2.n179 GND 0.01fF $ **FLOATING
C1696 CLK2.n180 GND 0.02fF $ **FLOATING
C1697 CLK2.n181 GND 0.03fF $ **FLOATING
C1698 CLK2.n182 GND 0.02fF $ **FLOATING
C1699 CLK2.n183 GND 0.01fF $ **FLOATING
C1700 CLK2.n184 GND 0.02fF $ **FLOATING
C1701 CLK2.n185 GND 0.03fF $ **FLOATING
C1702 CLK2.n186 GND 0.02fF $ **FLOATING
C1703 CLK2.n187 GND 0.01fF $ **FLOATING
C1704 CLK2.n188 GND 0.02fF $ **FLOATING
C1705 CLK2.n189 GND 0.07fF $ **FLOATING
C1706 CLK2.n190 GND 0.02fF $ **FLOATING
C1707 CLK2.n191 GND 0.01fF $ **FLOATING
C1708 CLK2.n192 GND 0.02fF $ **FLOATING
C1709 CLK2.n193 GND 0.09fF $ **FLOATING
C1710 CLK2.n194 GND 0.02fF $ **FLOATING
C1711 CLK2.n195 GND 0.01fF $ **FLOATING
C1712 CLK2.n196 GND 0.01fF $ **FLOATING
C1713 CLK2.n197 GND 0.15fF $ **FLOATING
C1714 CLK2.t2 GND 0.05fF
C1715 CLK2.n198 GND 0.05fF $ **FLOATING
C1716 CLK2.n199 GND 0.02fF $ **FLOATING
C1717 CLK2.n200 GND 0.01fF $ **FLOATING
C1718 CLK2.n201 GND 0.01fF $ **FLOATING
C1719 CLK2.n202 GND 0.08fF $ **FLOATING
C1720 CLK2.n203 GND 0.02fF $ **FLOATING
C1721 CLK2.n204 GND 0.01fF $ **FLOATING
C1722 CLK2.n205 GND 0.02fF $ **FLOATING
C1723 CLK2.t0 GND 0.05fF
C1724 CLK2.n206 GND 0.05fF $ **FLOATING
C1725 CLK2.n207 GND 0.02fF $ **FLOATING
C1726 CLK2.n208 GND 0.01fF $ **FLOATING
C1727 CLK2.n209 GND 0.02fF $ **FLOATING
C1728 CLK2.n210 GND 0.09fF $ **FLOATING
C1729 CLK2.n211 GND 0.02fF $ **FLOATING
C1730 CLK2.n212 GND 0.01fF $ **FLOATING
C1731 CLK2.n213 GND 0.09fF $ **FLOATING
C1732 CLK2.t24 GND 0.03fF
C1733 CLK2.t31 GND 0.02fF
C1734 CLK2.t27 GND 0.02fF
C1735 CLK2.n214 GND 0.08fF $ **FLOATING
C1736 CLK2.n215 GND 0.04fF $ **FLOATING
C1737 CLK2.n216 GND 0.02fF $ **FLOATING
C1738 CLK2.n217 GND 0.01fF $ **FLOATING
C1739 CLK2.n218 GND 0.07fF $ **FLOATING
C1740 CLK2.n219 GND 0.03fF $ **FLOATING
C1741 CLK2.n220 GND 0.02fF $ **FLOATING
C1742 CLK2.n221 GND 0.01fF $ **FLOATING
C1743 CLK2.n222 GND 0.04fF $ **FLOATING
C1744 CLK2.n223 GND 0.10fF $ **FLOATING
C1745 CLK2.n224 GND 0.03fF $ **FLOATING
C1746 CLK2.n225 GND 0.02fF $ **FLOATING
C1747 CLK2.n226 GND 0.01fF $ **FLOATING
C1748 CLK2.n227 GND 0.01fF $ **FLOATING
C1749 CLK2.n228 GND 0.03fF $ **FLOATING
C1750 CLK2.n229 GND 0.02fF $ **FLOATING
C1751 CLK2.n230 GND 0.01fF $ **FLOATING
C1752 CLK2.n231 GND 0.02fF $ **FLOATING
C1753 CLK2.n232 GND 0.07fF $ **FLOATING
C1754 CLK2.n233 GND 0.02fF $ **FLOATING
C1755 CLK2.n234 GND 0.01fF $ **FLOATING
C1756 CLK2.n235 GND 0.02fF $ **FLOATING
C1757 CLK2.n236 GND 0.09fF $ **FLOATING
C1758 CLK2.n237 GND 0.02fF $ **FLOATING
C1759 CLK2.n238 GND 0.01fF $ **FLOATING
C1760 CLK2.n239 GND 0.01fF $ **FLOATING
C1761 CLK2.n240 GND 0.15fF $ **FLOATING
C1762 CLK2.t23 GND 0.05fF
C1763 CLK2.n241 GND 0.05fF $ **FLOATING
C1764 CLK2.n242 GND 0.02fF $ **FLOATING
C1765 CLK2.n243 GND 0.01fF $ **FLOATING
C1766 CLK2.n244 GND 0.01fF $ **FLOATING
C1767 CLK2.n245 GND 0.08fF $ **FLOATING
C1768 CLK2.n246 GND 0.02fF $ **FLOATING
C1769 CLK2.n247 GND 0.01fF $ **FLOATING
C1770 CLK2.n248 GND 0.02fF $ **FLOATING
C1771 CLK2.t21 GND 0.05fF
C1772 CLK2.n249 GND 0.05fF $ **FLOATING
C1773 CLK2.n250 GND 0.02fF $ **FLOATING
C1774 CLK2.n251 GND 0.01fF $ **FLOATING
C1775 CLK2.n252 GND 0.01fF $ **FLOATING
C1776 x0_bar.t0 GND 0.47fF
C1777 x0_bar.t1 GND 0.53fF
C1778 x0_bar.t2 GND 0.18fF
C1779 x0_bar.n0 GND 1.75fF $ **FLOATING
C1780 x0_bar.n1 GND 5.78fF $ **FLOATING
C1781 EESPFAL_3in_NAND_v2_0/C GND 1.93fF $ **FLOATING
.ends

