* NGSPICE file created from EESPFAL_64bitwidth_PRESENT80_R1.ext - technology: sky130A

.subckt EESPFAL_XOR_v3 OUT_bar GND OUT A A_bar B B_bar Dis CLK
X0 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X2 a_n840_410# A CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=7.5e+12p ps=3.22e+07u w=1.5e+06u l=150000u
X3 a_n1140_410# B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_420_410# B_bar OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X5 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X7 a_720_410# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar B a_n840_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 CLK A_bar a_n1140_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK A a_420_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 OUT B a_720_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_4in_XOR EESPFAL_XOR_v3_3/GND x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar
+ x2 x2_bar k2 k2_bar x3 x3_bar k3 k3_bar XOR0_bar XOR0 XOR1_bar XOR1 XOR2_bar XOR2
+ XOR3_bar XOR3 CLK Dis
XEESPFAL_XOR_v3_0 XOR0_bar EESPFAL_XOR_v3_3/GND XOR0 x0 x0_bar k0 k0_bar Dis CLK EESPFAL_XOR_v3
XEESPFAL_XOR_v3_1 XOR1_bar EESPFAL_XOR_v3_3/GND XOR1 x1 x1_bar k1 k1_bar Dis CLK EESPFAL_XOR_v3
XEESPFAL_XOR_v3_2 XOR2_bar EESPFAL_XOR_v3_3/GND XOR2 x2 x2_bar k2 k2_bar Dis CLK EESPFAL_XOR_v3
XEESPFAL_XOR_v3_3 XOR3_bar EESPFAL_XOR_v3_3/GND XOR3 x3 x3_bar k3 k3_bar Dis CLK EESPFAL_XOR_v3
.ends

.subckt EESPFAL_3in_NAND_v2 OUT_bar GND OUT A A_bar B B_bar C C_bar Dis CLK
X0 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u M=2
X1 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X2 a_n910_640# B a_n1060_640# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X4 CLK B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=7.7e+12p pd=3.36e+07u as=0p ps=0u w=1.5e+06u l=150000u
X5 CLK A a_n910_640# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n1060_640# C OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 OUT_bar A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 OUT_bar C_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_INV4 OUT GND OUT_bar A A_bar Dis CLK
X0 OUT A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=5.25e+12p ps=2.32e+07u w=1.5e+06u l=150000u
X1 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X2 GND Dis OUT_bar GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X3 GND OUT_bar OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X5 OUT_bar OUT GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 CLK A OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT Dis GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_3in_NOR_v2 OUT_bar GND OUT A A_bar B B_bar C C_bar Dis CLK
X0 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 OUT B CLK GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=7.7e+12p ps=3.36e+07u w=1.5e+06u l=150000u
X2 OUT_bar OUT CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X3 a_n1990_570# B_bar a_n2140_570# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X4 CLK A OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X6 CLK C OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n2140_570# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 OUT_bar C_bar a_n1990_570# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_NAND_v3 OUT_bar GND OUT A A_bar B B_bar Dis CLK
X0 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X2 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X3 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X5 OUT_bar A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6e+12p ps=2.62e+07u w=1.5e+06u l=150000u
X6 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_501_n414# B OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 CLK A a_501_n414# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 CLK B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_s3 EESPFAL_INV4_2/GND x0 x1 x2 x2_bar x3 x3_bar s3_bar s3 Dis1 Dis3
+ Dis2 x0_bar CLK2 x1_bar CLK1 CLK3 EESPFAL_XOR_v3_0/OUT
XEESPFAL_3in_NAND_v2_0 EESPFAL_INV4_2/A_bar EESPFAL_INV4_2/GND EESPFAL_INV4_2/A x2_bar
+ x2 x0 x0_bar x3 x3_bar Dis1 CLK1 EESPFAL_3in_NAND_v2
XEESPFAL_INV4_0 EESPFAL_INV4_0/OUT EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/B x3_bar x3
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_INV4_1 EESPFAL_INV4_1/OUT EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/B x1 x1_bar
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_INV4_2 EESPFAL_INV4_2/OUT EESPFAL_INV4_2/GND EESPFAL_INV4_2/OUT_bar EESPFAL_INV4_2/A
+ EESPFAL_INV4_2/A_bar Dis2 CLK2 EESPFAL_INV4
XEESPFAL_XOR_v3_0 EESPFAL_NAND_v3_0/A EESPFAL_INV4_2/GND EESPFAL_XOR_v3_0/OUT x1 x1_bar
+ x0 x0_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_XOR_v3_1 EESPFAL_NAND_v3_1/A_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/A x2
+ x2_bar x3 x3_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_3in_NOR_v2_0 s3_bar EESPFAL_INV4_2/GND s3 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar
+ EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_2/OUT_bar EESPFAL_INV4_2/OUT
+ Dis3 CLK3 EESPFAL_3in_NOR_v2
XEESPFAL_NAND_v3_0 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/OUT
+ EESPFAL_NAND_v3_0/A EESPFAL_XOR_v3_0/OUT EESPFAL_NAND_v3_0/B EESPFAL_INV4_0/OUT
+ Dis2 CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_1 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/OUT
+ EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/B EESPFAL_INV4_1/OUT
+ Dis2 CLK2 EESPFAL_NAND_v3
.ends

.subckt EESPFAL_s1 EESPFAL_INV4_2/GND x0 x0_bar x1 x2 x2_bar x3 s1_bar s1 Dis1 Dis3
+ Dis2 x3_bar x1_bar CLK2 CLK1 CLK3
XEESPFAL_3in_NAND_v2_0 EESPFAL_INV4_2/A_bar EESPFAL_INV4_2/GND EESPFAL_INV4_2/A x3_bar
+ x3 x1 x1_bar x0_bar x0 Dis1 CLK1 EESPFAL_3in_NAND_v2
XEESPFAL_INV4_0 EESPFAL_INV4_0/OUT EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/B x3 x3_bar
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_INV4_1 EESPFAL_INV4_1/OUT EESPFAL_INV4_2/GND EESPFAL_INV4_1/OUT_bar x2 x2_bar
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_INV4_2 EESPFAL_INV4_2/OUT EESPFAL_INV4_2/GND EESPFAL_INV4_2/OUT_bar EESPFAL_INV4_2/A
+ EESPFAL_INV4_2/A_bar Dis2 CLK2 EESPFAL_INV4
XEESPFAL_XOR_v3_0 EESPFAL_NAND_v3_0/A EESPFAL_INV4_2/GND EESPFAL_XOR_v3_0/OUT x2 x2_bar
+ x0 x0_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_XOR_v3_1 EESPFAL_NAND_v3_1/A_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/A x1
+ x1_bar x3 x3_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_3in_NOR_v2_0 s1_bar EESPFAL_INV4_2/GND s1 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar
+ EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_2/OUT_bar EESPFAL_INV4_2/OUT
+ Dis3 CLK3 EESPFAL_3in_NOR_v2
XEESPFAL_NAND_v3_0 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/OUT
+ EESPFAL_NAND_v3_0/A EESPFAL_XOR_v3_0/OUT EESPFAL_NAND_v3_0/B EESPFAL_INV4_0/OUT
+ Dis2 CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_1 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/OUT
+ EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/A_bar EESPFAL_INV4_1/OUT EESPFAL_INV4_1/OUT_bar
+ Dis2 CLK2 EESPFAL_NAND_v3
.ends

.subckt EESPFAL_4in_NAND OUT_bar GND OUT A A_bar B B_bar C C_bar D D_bar Dis CLK
X0 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=3.6e+12p pd=1.68e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X1 CLK B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=8.5e+12p pd=3.68e+07u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n1040_180# B a_n1190_180# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 OUT_bar OUT CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u M=2
X4 CLK D_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n1340_180# D OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT_bar A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar C_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X11 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK A a_n1040_180# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_n1190_180# C a_n1340_180# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_s2 x0 x1 x1_bar x2 x2_bar x3 x3_bar Dis3 Dis2 CLK2 s2_bar s2 CLK1
+ x0_bar EESPFAL_INV4_2/GND CLK3 Dis1
XEESPFAL_4in_NAND_0 EESPFAL_INV4_1/A_bar EESPFAL_INV4_2/GND EESPFAL_INV4_1/A x3_bar
+ x3 x1 x1_bar x0 x0_bar x2 x2_bar Dis1 CLK1 EESPFAL_4in_NAND
XEESPFAL_INV4_0 EESPFAL_INV4_0/OUT EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/B x1_bar x1
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_INV4_1 EESPFAL_INV4_1/OUT EESPFAL_INV4_2/GND EESPFAL_INV4_1/OUT_bar EESPFAL_INV4_1/A
+ EESPFAL_INV4_1/A_bar Dis2 CLK2 EESPFAL_INV4
XEESPFAL_INV4_2 EESPFAL_INV4_2/OUT EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/B x2_bar x2
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_XOR_v3_0 EESPFAL_NAND_v3_0/A EESPFAL_INV4_2/GND EESPFAL_XOR_v3_0/OUT x3 x3_bar
+ x2 x2_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_XOR_v3_1 EESPFAL_NAND_v3_1/A_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/A x1
+ x1_bar x0 x0_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_3in_NOR_v2_0 s2_bar EESPFAL_INV4_2/GND s2 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar
+ EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_1/OUT_bar EESPFAL_INV4_1/OUT
+ Dis3 CLK3 EESPFAL_3in_NOR_v2
XEESPFAL_NAND_v3_0 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/OUT
+ EESPFAL_NAND_v3_0/A EESPFAL_XOR_v3_0/OUT EESPFAL_NAND_v3_0/B EESPFAL_INV4_0/OUT
+ Dis2 CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_1 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/OUT
+ EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/B EESPFAL_INV4_2/OUT
+ Dis2 CLK2 EESPFAL_NAND_v3
.ends

.subckt EESPFAL_NOR_v3 OUT_bar GND OUT A A_bar B B_bar Dis CLK
X0 a_n1820_550# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=6e+12p ps=2.62e+07u w=1.5e+06u l=150000u
X1 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X2 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u M=2
X3 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X4 OUT_bar B_bar a_n1820_550# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X6 OUT A CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 CLK B OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_s0 EESPFAL_XOR_v3_0/GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar Dis1
+ Dis2 Dis3 s0 s0_bar CLK3 CLK2 CLK1
XEESPFAL_XOR_v3_0 EESPFAL_NAND_v3_1/A EESPFAL_XOR_v3_0/GND EESPFAL_NAND_v3_0/A x0
+ x0_bar x3 x3_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_NOR_v3_0 s0_bar EESPFAL_XOR_v3_0/GND s0 EESPFAL_NOR_v3_0/A EESPFAL_NOR_v3_0/A_bar
+ EESPFAL_NOR_v3_0/B EESPFAL_NOR_v3_0/B_bar Dis3 CLK3 EESPFAL_NOR_v3
XEESPFAL_NOR_v3_1 EESPFAL_NAND_v3_0/B_bar EESPFAL_XOR_v3_0/GND EESPFAL_NAND_v3_0/B
+ x1 x1_bar x2_bar x2 Dis1 CLK1 EESPFAL_NOR_v3
XEESPFAL_NAND_v3_0 EESPFAL_NOR_v3_0/A_bar EESPFAL_XOR_v3_0/GND EESPFAL_NOR_v3_0/A
+ EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar
+ Dis2 CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_1 EESPFAL_NOR_v3_0/B_bar EESPFAL_XOR_v3_0/GND EESPFAL_NOR_v3_0/B
+ EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar
+ Dis2 CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_2 EESPFAL_NAND_v3_1/B_bar EESPFAL_XOR_v3_0/GND EESPFAL_NAND_v3_1/B
+ x2 x2_bar x1_bar x1 Dis1 CLK1 EESPFAL_NAND_v3
.ends

.subckt EESPFAL_Sbox x0 x1 x2_bar Dis1 Dis2 Dis3 s0 s0_bar s1 s2 s2_bar s3_bar s3
+ s1_bar CLK2 CLK3 CLK1 x3_bar x3 x2 EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT EESPFAL_s3_0/EESPFAL_INV4_2/GND
+ x0_bar x1_bar
XEESPFAL_s3_0 EESPFAL_s3_0/EESPFAL_INV4_2/GND x0 x1 x2 x2_bar x3 x3_bar s3_bar s3
+ Dis1 Dis3 Dis2 x0_bar CLK2 x1_bar CLK1 CLK3 EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT EESPFAL_s3
XEESPFAL_s1_0 EESPFAL_s3_0/EESPFAL_INV4_2/GND x0 x0_bar x1 x2 x2_bar x3 s1_bar s1
+ Dis1 Dis3 Dis2 x3_bar x1_bar CLK2 CLK1 CLK3 EESPFAL_s1
XEESPFAL_s2_0 x0 x1 x1_bar x2 x2_bar x3 x3_bar Dis3 Dis2 CLK2 s2_bar s2 CLK1 x0_bar
+ EESPFAL_s3_0/EESPFAL_INV4_2/GND CLK3 Dis1 EESPFAL_s2
XEESPFAL_s0_0 EESPFAL_s3_0/EESPFAL_INV4_2/GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar
+ Dis1 Dis2 Dis3 s0 s0_bar CLK3 CLK2 CLK1 EESPFAL_s0
.ends

.subckt EESPFAL_PRESENT_R1 x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar x2 x2_bar k2 k2_bar
+ x3 x3_bar k3 k3_bar s0 s0_bar Dis0 Dis1 s3_bar s3 s1 Dis3 CLK0 s2_bar CLK2 s1_bar
+ s2 CLK3 Dis2 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/GND CLK1
XEESPFAL_4in_XOR_0 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/GND x0 x0_bar k0 k0_bar x1 x1_bar
+ k1 k1_bar x2 x2_bar k2 k2_bar x3 x3_bar k3 k3_bar EESPFAL_Sbox_0/x0_bar EESPFAL_Sbox_0/x0
+ EESPFAL_Sbox_0/x1_bar EESPFAL_Sbox_0/x1 EESPFAL_Sbox_0/x2_bar EESPFAL_Sbox_0/x2
+ EESPFAL_Sbox_0/x3_bar EESPFAL_Sbox_0/x3 CLK0 Dis0 EESPFAL_4in_XOR
XEESPFAL_Sbox_0 EESPFAL_Sbox_0/x0 EESPFAL_Sbox_0/x1 EESPFAL_Sbox_0/x2_bar Dis1 Dis2
+ Dis3 s0 s0_bar s1 s2 s2_bar s3_bar s3 s1_bar CLK2 CLK3 CLK1 EESPFAL_Sbox_0/x3_bar
+ EESPFAL_Sbox_0/x3 EESPFAL_Sbox_0/x2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT
+ EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/GND EESPFAL_Sbox_0/x0_bar EESPFAL_Sbox_0/x1_bar
+ EESPFAL_Sbox
.ends

.subckt EESPFAL_64bitwidth_PRESENT80_R1 GND k3_bar x3_bar x0 x0_bar k0 k0_bar x1 k1_bar
+ k1 k2 k2_bar x2 x2_bar k3 x3 k4 k5 k6 k7 k4_bar k5_bar k6_bar k7_bar x4 x5 x6 x7
+ x4_bar x5_bar x6_bar x7_bar x14 k15_bar k14_bar k13_bar k12_bar x13 x12 x12_bar
+ x13_bar x15 k12 x15_bar x14_bar k15 k14 k13 x8_bar x9_bar k8 x10_bar k9 x11_bar
+ k10 k11 x11 x10 x9 x8 k8_bar k11_bar k10_bar k9_bar x17 x16 k18_bar k17_bar k16_bar
+ k17 k16 k19 k18 k19_bar x16_bar x17_bar x18_bar x19_bar x18 x19 x21_bar x22_bar
+ x23_bar k20_bar x20_bar k21_bar k22_bar k23_bar k22 k21 k20 k23 x20 x21 x22 x23
+ x25 x24_bar x24 k24_bar k25_bar k26_bar x25_bar x26_bar k25 k24 k26 x26 x27 x27_bar
+ k27 k27_bar k30 k30_bar x29_bar k29_bar x28 k28_bar x28_bar x29 k31 k31_bar x30_bar
+ x31_bar k29 x30 k28 x31 x1_bar k34 k35 x32 x33 x34 x35 x35_bar x34_bar x33_bar x32_bar
+ k33 k32 k32_bar k35_bar k33_bar k34_bar x38 k38_bar k39_bar x39 k38 x37 x36 k39
+ k36 k37_bar k36_bar x39_bar x38_bar x36_bar x37_bar k37 x41_bar x40_bar x43 x42
+ x41 k40_bar x40 k41_bar k42_bar k40 k43_bar k41 k42 k43 x42_bar x43_bar k47_bar
+ k46_bar k45_bar k44_bar x44 x47 x47_bar k47 x46 k46 k45 k44 x44_bar x45_bar x46_bar
+ x45 x51_bar x50_bar k51_bar k49 k48 x50 k48_bar x49 x48_bar x48 x49_bar k50_bar
+ x51 k50 k49_bar k51 x54 k55_bar x55 k55 x54_bar x55_bar k54_bar x52 k53 k52 x53_bar
+ x53 k53_bar k52_bar k54 x52_bar k60 k62 k63 k62_bar k60_bar k61_bar x63 k63_bar
+ x60 x61 x60_bar x63_bar x61_bar k61 x62 x62_bar k58 x56_bar x59 k57 k59_bar k56_bar
+ k58_bar x58_bar x56 x58 k56 x59_bar x57_bar x57 k59 k57_bar Dis0 CLK1 Dis1 CLK3
+ Dis2 CLK2 Dis3 s12 s13 s14 s12_bar s13_bar s14_bar s16 s17 s18 s19 s16_bar s17_bar
+ s18_bar s19_bar s22 s23 s20 s21 s20_bar s21_bar s22_bar s23_bar s24 s25 s26 s27
+ s24_bar s26_bar s27_bar s28 s29 s30 s31 s28_bar s29_bar s30_bar s31_bar s0 s1 s2
+ s3 s4 s6 s7 s8 s9 s10 s0_bar s1_bar s2_bar s3_bar s4_bar s6_bar s7_bar s8_bar s9_bar
+ s10_bar s5_bar s5 s11 s15 s11_bar s15_bar s25_bar CLK0 s35 s35_bar s52 s53 s54 s55
+ s56 s57 s58 s59 s60 s61 s62 s63 s40_bar s41_bar s42_bar s43_bar s44_bar s45_bar
+ s46_bar s47_bar s48_bar s49_bar s50_bar s51_bar s52_bar s53_bar s54_bar s55_bar
+ s56_bar s57_bar s58_bar s59_bar s60_bar s61_bar s62_bar s63_bar s33 s34 s32_bar
+ s33_bar s34_bar s37 s38 s39 s37_bar s38_bar s39_bar s32 s36_bar s36 s40 s41 s42
+ s43 s44 s45 s46 s47 s48 s49 s50 s51
XEESPFAL_PRESENT_R1_0 x60 x60_bar k60 k60_bar x61 x61_bar k61 k61_bar x62 x62_bar
+ k62 k62_bar x63 x63_bar k63 k63_bar s60 s60_bar Dis0 Dis1 s63_bar s63 s61 Dis3 CLK0
+ s62_bar CLK2 s61_bar s62 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_1 x52 x52_bar k52 k52_bar x53 x53_bar k53 k53_bar x54 x54_bar
+ k54 k54_bar x55 x55_bar k55 k55_bar s52 s52_bar Dis0 Dis1 s55_bar s55 s53 Dis3 CLK0
+ s54_bar CLK2 s53_bar s54 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_3 x48 x48_bar k48 k48_bar x49 x49_bar k49 k49_bar x50 x50_bar
+ k50 k50_bar x51 x51_bar k51 k51_bar s48 s48_bar Dis0 Dis1 s51_bar s51 s49 Dis3 CLK0
+ s50_bar CLK2 s49_bar s50 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_2 x56 x56_bar k56 k56_bar x57 x57_bar k57 k57_bar x58 x58_bar
+ k58 k58_bar x59 x59_bar k59 k59_bar s56 s56_bar Dis0 Dis1 s59_bar s59 s57 Dis3 CLK0
+ s58_bar CLK2 s57_bar s58 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_4 x44 x44_bar k44 k44_bar x45 x45_bar k45 k45_bar x46 x46_bar
+ k46 k46_bar x47 x47_bar k47 k47_bar s44 s44_bar Dis0 Dis1 s47_bar s47 s45 Dis3 CLK0
+ s46_bar CLK2 s45_bar s46 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_5 x40 x40_bar k40 k40_bar x41 x41_bar k41 k41_bar x42 x42_bar
+ k42 k42_bar x43 x43_bar k43 k43_bar s40 s40_bar Dis0 Dis1 s43_bar s43 s41 Dis3 CLK0
+ s42_bar CLK2 s41_bar s42 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_6 x32 x32_bar k32 k32_bar x33 x33_bar k33 k33_bar x34 x34_bar
+ k34 k34_bar x35 x35_bar k35 k35_bar s32 s32_bar Dis0 Dis1 s35_bar s35 s33 Dis3 CLK0
+ s34_bar CLK2 s33_bar s34 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_7 x36 x36_bar k36 k36_bar x37 x37_bar k37 k37_bar x38 x38_bar
+ k38 k38_bar x39 x39_bar k39 k39_bar s36 s36_bar Dis0 Dis1 s39_bar s39 s37 Dis3 CLK0
+ s38_bar CLK2 s37_bar s38 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_8 x28 x28_bar k28 k28_bar x29 x29_bar k29 k29_bar x30 x30_bar
+ k30 k30_bar x31 x31_bar k31 k31_bar s28 s28_bar Dis0 Dis1 s31_bar s31 s29 Dis3 CLK0
+ s30_bar CLK2 s29_bar s30 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_9 x24 x24_bar k24 k24_bar x25 x25_bar k25 k25_bar x26 x26_bar
+ k26 k26_bar x27 x27_bar k27 k27_bar s24 s24_bar Dis0 Dis1 s27_bar s27 s25 Dis3 CLK0
+ s26_bar CLK2 s25_bar s26 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_10 x20 x20_bar k20 k20_bar x21 x21_bar k21 k21_bar x22 x22_bar
+ k22 k22_bar x23 x23_bar k23 k23_bar s20 s20_bar Dis0 Dis1 s23_bar s23 s21 Dis3 CLK0
+ s22_bar CLK2 s21_bar s22 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_11 x16 x16_bar k16 k16_bar x17 x17_bar k17 k17_bar x18 x18_bar
+ k18 k18_bar x19 x19_bar k19 k19_bar s16 s16_bar Dis0 Dis1 s19_bar s19 s17 Dis3 CLK0
+ s18_bar CLK2 s17_bar s18 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_12 x4 x4_bar k4 k4_bar x5 x5_bar k5 k5_bar x6 x6_bar k6 k6_bar
+ x7 x7_bar k7 k7_bar s4 s4_bar Dis0 Dis1 s7_bar s7 s5 Dis3 CLK0 s6_bar CLK2 s5_bar
+ s6 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_13 x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar x2 x2_bar k2 k2_bar
+ x3 x3_bar k3 k3_bar s0 s0_bar Dis0 Dis1 s3_bar s3 s1 Dis3 CLK0 s2_bar CLK2 s1_bar
+ s2 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_14 x12 x12_bar k12 k12_bar x13 x13_bar k13 k13_bar x14 x14_bar
+ k14 k14_bar x15 x15_bar k15 k15_bar s12 s12_bar Dis0 Dis1 s15_bar s15 s13 Dis3 CLK0
+ s14_bar CLK2 s13_bar s14 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
XEESPFAL_PRESENT_R1_15 x8 x8_bar k8 k8_bar x9 x9_bar k9 k9_bar x10 x10_bar k10 k10_bar
+ x11 x11_bar k11 k11_bar s8 s8_bar Dis0 Dis1 s11_bar s11 s9 Dis3 CLK0 s10_bar CLK2
+ s9_bar s10 CLK3 Dis2 GND CLK1 EESPFAL_PRESENT_R1
.ends

