magic
tech sky130A
timestamp 1664857990
<< nwell >>
rect -885 795 20 885
rect -575 430 -305 795
<< nmos >>
rect -795 175 -780 325
rect -720 175 -705 325
rect -555 175 -540 325
rect -480 175 -465 325
rect -405 175 -390 325
rect -330 175 -315 325
rect -165 175 -150 325
rect -90 175 -75 325
<< pmos >>
rect -480 455 -465 755
rect -405 455 -390 755
<< ndiff >>
rect -855 290 -795 325
rect -855 270 -835 290
rect -815 270 -795 290
rect -855 250 -795 270
rect -855 230 -835 250
rect -815 230 -795 250
rect -855 210 -795 230
rect -855 190 -835 210
rect -815 190 -795 210
rect -855 175 -795 190
rect -780 175 -720 325
rect -705 290 -645 325
rect -705 270 -685 290
rect -665 270 -645 290
rect -705 250 -645 270
rect -705 230 -685 250
rect -665 230 -645 250
rect -705 210 -645 230
rect -705 190 -685 210
rect -665 190 -645 210
rect -705 175 -645 190
rect -615 290 -555 325
rect -615 270 -595 290
rect -575 270 -555 290
rect -615 250 -555 270
rect -615 230 -595 250
rect -575 230 -555 250
rect -615 210 -555 230
rect -615 190 -595 210
rect -575 190 -555 210
rect -615 175 -555 190
rect -540 290 -480 325
rect -540 270 -520 290
rect -500 270 -480 290
rect -540 250 -480 270
rect -540 230 -520 250
rect -500 230 -480 250
rect -540 210 -480 230
rect -540 190 -520 210
rect -500 190 -480 210
rect -540 175 -480 190
rect -465 290 -405 325
rect -465 270 -445 290
rect -425 270 -405 290
rect -465 250 -405 270
rect -465 230 -445 250
rect -425 230 -405 250
rect -465 210 -405 230
rect -465 190 -445 210
rect -425 190 -405 210
rect -465 175 -405 190
rect -390 290 -330 325
rect -390 270 -370 290
rect -350 270 -330 290
rect -390 250 -330 270
rect -390 230 -370 250
rect -350 230 -330 250
rect -390 210 -330 230
rect -390 190 -370 210
rect -350 190 -330 210
rect -390 175 -330 190
rect -315 290 -255 325
rect -315 270 -295 290
rect -275 270 -255 290
rect -315 250 -255 270
rect -315 230 -295 250
rect -275 230 -255 250
rect -315 210 -255 230
rect -315 190 -295 210
rect -275 190 -255 210
rect -315 175 -255 190
rect -225 290 -165 325
rect -225 270 -205 290
rect -185 270 -165 290
rect -225 250 -165 270
rect -225 230 -205 250
rect -185 230 -165 250
rect -225 210 -165 230
rect -225 190 -205 210
rect -185 190 -165 210
rect -225 175 -165 190
rect -150 290 -90 325
rect -150 270 -130 290
rect -110 270 -90 290
rect -150 250 -90 270
rect -150 230 -130 250
rect -110 230 -90 250
rect -150 210 -90 230
rect -150 190 -130 210
rect -110 190 -90 210
rect -150 175 -90 190
rect -75 290 -15 325
rect -75 270 -55 290
rect -35 270 -15 290
rect -75 250 -15 270
rect -75 230 -55 250
rect -35 230 -15 250
rect -75 210 -15 230
rect -75 190 -55 210
rect -35 190 -15 210
rect -75 175 -15 190
<< pdiff >>
rect -540 730 -480 755
rect -540 710 -520 730
rect -500 710 -480 730
rect -540 690 -480 710
rect -540 670 -520 690
rect -500 670 -480 690
rect -540 650 -480 670
rect -540 630 -520 650
rect -500 630 -480 650
rect -540 610 -480 630
rect -540 590 -520 610
rect -500 590 -480 610
rect -540 570 -480 590
rect -540 550 -520 570
rect -500 550 -480 570
rect -540 530 -480 550
rect -540 510 -520 530
rect -500 510 -480 530
rect -540 490 -480 510
rect -540 470 -520 490
rect -500 470 -480 490
rect -540 455 -480 470
rect -465 730 -405 755
rect -465 710 -445 730
rect -425 710 -405 730
rect -465 690 -405 710
rect -465 670 -445 690
rect -425 670 -405 690
rect -465 650 -405 670
rect -465 630 -445 650
rect -425 630 -405 650
rect -465 610 -405 630
rect -465 590 -445 610
rect -425 590 -405 610
rect -465 570 -405 590
rect -465 550 -445 570
rect -425 550 -405 570
rect -465 530 -405 550
rect -465 510 -445 530
rect -425 510 -405 530
rect -465 490 -405 510
rect -465 470 -445 490
rect -425 470 -405 490
rect -465 455 -405 470
rect -390 730 -330 755
rect -390 710 -370 730
rect -350 710 -330 730
rect -390 690 -330 710
rect -390 670 -370 690
rect -350 670 -330 690
rect -390 650 -330 670
rect -390 630 -370 650
rect -350 630 -330 650
rect -390 610 -330 630
rect -390 590 -370 610
rect -350 590 -330 610
rect -390 570 -330 590
rect -390 550 -370 570
rect -350 550 -330 570
rect -390 530 -330 550
rect -390 510 -370 530
rect -350 510 -330 530
rect -390 490 -330 510
rect -390 470 -370 490
rect -350 470 -330 490
rect -390 455 -330 470
<< ndiffc >>
rect -835 270 -815 290
rect -835 230 -815 250
rect -835 190 -815 210
rect -685 270 -665 290
rect -685 230 -665 250
rect -685 190 -665 210
rect -595 270 -575 290
rect -595 230 -575 250
rect -595 190 -575 210
rect -520 270 -500 290
rect -520 230 -500 250
rect -520 190 -500 210
rect -445 270 -425 290
rect -445 230 -425 250
rect -445 190 -425 210
rect -370 270 -350 290
rect -370 230 -350 250
rect -370 190 -350 210
rect -295 270 -275 290
rect -295 230 -275 250
rect -295 190 -275 210
rect -205 270 -185 290
rect -205 230 -185 250
rect -205 190 -185 210
rect -130 270 -110 290
rect -130 230 -110 250
rect -130 190 -110 210
rect -55 270 -35 290
rect -55 230 -35 250
rect -55 190 -35 210
<< pdiffc >>
rect -520 710 -500 730
rect -520 670 -500 690
rect -520 630 -500 650
rect -520 590 -500 610
rect -520 550 -500 570
rect -520 510 -500 530
rect -520 470 -500 490
rect -445 710 -425 730
rect -445 670 -425 690
rect -445 630 -425 650
rect -445 590 -425 610
rect -445 550 -425 570
rect -445 510 -425 530
rect -445 470 -425 490
rect -370 710 -350 730
rect -370 670 -350 690
rect -370 630 -350 650
rect -370 590 -350 610
rect -370 550 -350 570
rect -370 510 -350 530
rect -370 470 -350 490
<< psubdiff >>
rect -865 -130 0 -115
rect -865 -150 -845 -130
rect -825 -150 -805 -130
rect -785 -150 -765 -130
rect -745 -150 -725 -130
rect -705 -150 -685 -130
rect -665 -150 -645 -130
rect -625 -150 -605 -130
rect -585 -150 -565 -130
rect -545 -150 -525 -130
rect -505 -150 -485 -130
rect -465 -150 -445 -130
rect -425 -150 -405 -130
rect -385 -150 -365 -130
rect -345 -150 -325 -130
rect -305 -150 -285 -130
rect -265 -150 -245 -130
rect -225 -150 -200 -130
rect -180 -150 -160 -130
rect -140 -150 -120 -130
rect -100 -150 -80 -130
rect -60 -150 -40 -130
rect -20 -150 0 -130
rect -865 -165 0 -150
<< nsubdiff >>
rect -865 850 0 865
rect -865 830 -845 850
rect -825 830 -805 850
rect -785 830 -765 850
rect -745 830 -725 850
rect -705 830 -685 850
rect -665 830 -645 850
rect -625 830 -605 850
rect -585 830 -565 850
rect -545 830 -525 850
rect -505 830 -485 850
rect -465 830 -445 850
rect -425 830 -405 850
rect -385 830 -365 850
rect -345 830 -325 850
rect -305 830 -285 850
rect -265 830 -245 850
rect -225 830 -205 850
rect -185 830 -160 850
rect -140 830 -120 850
rect -100 830 -80 850
rect -60 830 -40 850
rect -20 830 0 850
rect -865 815 0 830
<< psubdiffcont >>
rect -845 -150 -825 -130
rect -805 -150 -785 -130
rect -765 -150 -745 -130
rect -725 -150 -705 -130
rect -685 -150 -665 -130
rect -645 -150 -625 -130
rect -605 -150 -585 -130
rect -565 -150 -545 -130
rect -525 -150 -505 -130
rect -485 -150 -465 -130
rect -445 -150 -425 -130
rect -405 -150 -385 -130
rect -365 -150 -345 -130
rect -325 -150 -305 -130
rect -285 -150 -265 -130
rect -245 -150 -225 -130
rect -200 -150 -180 -130
rect -160 -150 -140 -130
rect -120 -150 -100 -130
rect -80 -150 -60 -130
rect -40 -150 -20 -130
<< nsubdiffcont >>
rect -845 830 -825 850
rect -805 830 -785 850
rect -765 830 -745 850
rect -725 830 -705 850
rect -685 830 -665 850
rect -645 830 -625 850
rect -605 830 -585 850
rect -565 830 -545 850
rect -525 830 -505 850
rect -485 830 -465 850
rect -445 830 -425 850
rect -405 830 -385 850
rect -365 830 -345 850
rect -325 830 -305 850
rect -285 830 -265 850
rect -245 830 -225 850
rect -205 830 -185 850
rect -160 830 -140 850
rect -120 830 -100 850
rect -80 830 -60 850
rect -40 830 -20 850
<< poly >>
rect -480 755 -465 770
rect -405 755 -390 770
rect -480 380 -465 455
rect -405 440 -390 455
rect -430 430 -390 440
rect -430 410 -420 430
rect -400 410 -390 430
rect -430 400 -390 410
rect -480 370 -440 380
rect -480 350 -470 370
rect -450 350 -440 370
rect -480 340 -440 350
rect -795 325 -780 340
rect -720 325 -705 340
rect -555 325 -540 340
rect -480 325 -465 340
rect -405 325 -390 400
rect -330 325 -315 340
rect -165 325 -150 340
rect -90 325 -75 340
rect -795 110 -780 175
rect -795 100 -755 110
rect -795 80 -785 100
rect -765 80 -755 100
rect -795 70 -755 80
rect -720 60 -705 175
rect -555 160 -540 175
rect -480 160 -465 175
rect -405 160 -390 175
rect -330 160 -315 175
rect -555 150 -515 160
rect -555 130 -545 150
rect -525 130 -515 150
rect -555 120 -515 130
rect -355 150 -315 160
rect -355 130 -345 150
rect -325 130 -315 150
rect -355 120 -315 130
rect -720 50 -680 60
rect -720 30 -710 50
rect -690 30 -680 50
rect -720 20 -680 30
rect -165 10 -150 175
rect -165 0 -125 10
rect -165 -20 -155 0
rect -135 -20 -125 0
rect -165 -30 -125 -20
rect -90 -50 -75 175
rect -90 -60 -50 -50
rect -90 -80 -80 -60
rect -60 -80 -50 -60
rect -90 -90 -50 -80
<< polycont >>
rect -420 410 -400 430
rect -470 350 -450 370
rect -785 80 -765 100
rect -545 130 -525 150
rect -345 130 -325 150
rect -710 30 -690 50
rect -155 -20 -135 0
rect -80 -80 -60 -60
<< locali >>
rect -865 850 0 860
rect -865 830 -845 850
rect -825 830 -805 850
rect -785 830 -765 850
rect -745 830 -725 850
rect -705 830 -685 850
rect -665 830 -645 850
rect -625 830 -605 850
rect -585 830 -565 850
rect -545 830 -525 850
rect -505 830 -485 850
rect -465 830 -445 850
rect -425 830 -405 850
rect -385 830 -365 850
rect -345 830 -325 850
rect -305 830 -285 850
rect -265 830 -245 850
rect -225 830 -205 850
rect -185 830 -160 850
rect -140 830 -120 850
rect -100 830 -80 850
rect -60 830 -40 850
rect -20 830 0 850
rect -865 820 0 830
rect -530 730 -490 740
rect -530 710 -520 730
rect -500 710 -490 730
rect -530 690 -490 710
rect -530 670 -520 690
rect -500 670 -490 690
rect -530 650 -490 670
rect -530 630 -520 650
rect -500 630 -490 650
rect -530 610 -490 630
rect -530 590 -520 610
rect -500 590 -490 610
rect -530 570 -490 590
rect -530 550 -520 570
rect -500 550 -490 570
rect -530 530 -490 550
rect -530 510 -520 530
rect -500 510 -490 530
rect -530 490 -490 510
rect -530 470 -520 490
rect -500 470 -490 490
rect -530 455 -490 470
rect -455 730 -415 740
rect -455 710 -445 730
rect -425 710 -415 730
rect -455 690 -415 710
rect -455 670 -445 690
rect -425 670 -415 690
rect -455 650 -415 670
rect -455 630 -445 650
rect -425 630 -415 650
rect -455 610 -415 630
rect -455 590 -445 610
rect -425 590 -415 610
rect -455 570 -415 590
rect -455 550 -445 570
rect -425 550 -415 570
rect -455 530 -415 550
rect -455 510 -445 530
rect -425 510 -415 530
rect -455 490 -415 510
rect -455 470 -445 490
rect -425 470 -415 490
rect -455 460 -415 470
rect -380 730 -340 740
rect -380 710 -370 730
rect -350 710 -340 730
rect -380 690 -340 710
rect -380 670 -370 690
rect -350 670 -340 690
rect -380 650 -340 670
rect -380 630 -370 650
rect -350 630 -340 650
rect -380 610 -340 630
rect -380 590 -370 610
rect -350 590 -340 610
rect -380 570 -340 590
rect -380 550 -370 570
rect -350 550 -340 570
rect -380 530 -340 550
rect -380 510 -370 530
rect -350 510 -340 530
rect -380 490 -340 510
rect -380 470 -370 490
rect -350 470 -340 490
rect -380 455 -340 470
rect -520 430 -500 455
rect -430 430 -390 440
rect -520 410 -420 430
rect -400 410 -390 430
rect -520 365 -500 410
rect -430 400 -390 410
rect -685 345 -500 365
rect -685 305 -665 345
rect -520 325 -500 345
rect -480 370 -440 380
rect -370 370 -350 455
rect -480 350 -470 370
rect -450 350 -35 370
rect -480 340 -440 350
rect -370 325 -350 350
rect -845 290 -805 305
rect -845 270 -835 290
rect -815 270 -805 290
rect -845 250 -805 270
rect -845 230 -835 250
rect -815 230 -805 250
rect -845 210 -805 230
rect -845 190 -835 210
rect -815 190 -805 210
rect -845 180 -805 190
rect -695 290 -655 305
rect -695 270 -685 290
rect -665 270 -655 290
rect -695 250 -655 270
rect -695 230 -685 250
rect -665 230 -655 250
rect -695 210 -655 230
rect -695 190 -685 210
rect -665 190 -655 210
rect -695 180 -655 190
rect -605 290 -565 305
rect -605 270 -595 290
rect -575 270 -565 290
rect -605 250 -565 270
rect -605 230 -595 250
rect -575 230 -565 250
rect -605 210 -565 230
rect -605 190 -595 210
rect -575 190 -565 210
rect -605 180 -565 190
rect -530 290 -490 325
rect -530 270 -520 290
rect -500 270 -490 290
rect -530 250 -490 270
rect -530 230 -520 250
rect -500 230 -490 250
rect -530 210 -490 230
rect -530 190 -520 210
rect -500 190 -490 210
rect -530 180 -490 190
rect -455 290 -415 305
rect -455 270 -445 290
rect -425 270 -415 290
rect -455 250 -415 270
rect -455 230 -445 250
rect -425 230 -415 250
rect -455 210 -415 230
rect -455 190 -445 210
rect -425 190 -415 210
rect -455 180 -415 190
rect -380 290 -340 325
rect -205 305 -185 350
rect -55 305 -35 350
rect -380 270 -370 290
rect -350 270 -340 290
rect -380 250 -340 270
rect -380 230 -370 250
rect -350 230 -340 250
rect -380 210 -340 230
rect -380 190 -370 210
rect -350 190 -340 210
rect -380 180 -340 190
rect -305 290 -265 305
rect -305 270 -295 290
rect -275 270 -265 290
rect -305 250 -265 270
rect -305 230 -295 250
rect -275 230 -265 250
rect -305 210 -265 230
rect -305 190 -295 210
rect -275 190 -265 210
rect -305 180 -265 190
rect -215 290 -175 305
rect -215 270 -205 290
rect -185 270 -175 290
rect -215 250 -175 270
rect -215 230 -205 250
rect -185 230 -175 250
rect -215 210 -175 230
rect -215 190 -205 210
rect -185 190 -175 210
rect -215 180 -175 190
rect -140 290 -100 305
rect -140 270 -130 290
rect -110 270 -100 290
rect -140 250 -100 270
rect -140 230 -130 250
rect -110 230 -100 250
rect -140 210 -100 230
rect -140 190 -130 210
rect -110 190 -100 210
rect -140 180 -100 190
rect -65 290 -25 305
rect -65 270 -55 290
rect -35 270 -25 290
rect -65 250 -25 270
rect -65 230 -55 250
rect -35 230 -25 250
rect -65 210 -25 230
rect -65 190 -55 210
rect -35 190 -25 210
rect -65 180 -25 190
rect -555 150 -515 160
rect -355 150 -315 160
rect -860 130 -545 150
rect -525 130 -345 150
rect -325 130 -315 150
rect -555 120 -515 130
rect -355 120 -315 130
rect -795 100 -755 110
rect -855 80 -785 100
rect -765 80 -755 100
rect -795 70 -755 80
rect -720 50 -680 60
rect -855 30 -710 50
rect -690 30 -680 50
rect -720 20 -680 30
rect -165 0 -125 10
rect -855 -20 -155 0
rect -135 -20 -125 0
rect -165 -30 -125 -20
rect -90 -60 -50 -50
rect -855 -80 -80 -60
rect -60 -80 -50 -60
rect -90 -90 -50 -80
rect -865 -130 0 -120
rect -865 -150 -845 -130
rect -825 -150 -805 -130
rect -785 -150 -765 -130
rect -745 -150 -725 -130
rect -705 -150 -685 -130
rect -665 -150 -645 -130
rect -625 -150 -605 -130
rect -585 -150 -565 -130
rect -545 -150 -525 -130
rect -505 -150 -485 -130
rect -465 -150 -445 -130
rect -425 -150 -405 -130
rect -385 -150 -365 -130
rect -345 -150 -325 -130
rect -305 -150 -285 -130
rect -265 -150 -245 -130
rect -225 -150 -200 -130
rect -180 -150 -160 -130
rect -140 -150 -120 -130
rect -100 -150 -80 -130
rect -60 -150 -40 -130
rect -20 -150 0 -130
rect -865 -160 0 -150
<< viali >>
rect -845 830 -825 850
rect -805 830 -785 850
rect -765 830 -745 850
rect -725 830 -705 850
rect -685 830 -665 850
rect -645 830 -625 850
rect -605 830 -585 850
rect -565 830 -545 850
rect -525 830 -505 850
rect -485 830 -465 850
rect -445 830 -425 850
rect -405 830 -385 850
rect -365 830 -345 850
rect -325 830 -305 850
rect -285 830 -265 850
rect -245 830 -225 850
rect -205 830 -185 850
rect -160 830 -140 850
rect -120 830 -100 850
rect -80 830 -60 850
rect -40 830 -20 850
rect -445 710 -425 730
rect -445 670 -425 690
rect -445 630 -425 650
rect -445 590 -425 610
rect -445 550 -425 570
rect -445 510 -425 530
rect -445 470 -425 490
rect -835 270 -815 290
rect -835 230 -815 250
rect -835 190 -815 210
rect -595 270 -575 290
rect -595 230 -575 250
rect -595 190 -575 210
rect -445 270 -425 290
rect -445 230 -425 250
rect -445 190 -425 210
rect -295 270 -275 290
rect -295 230 -275 250
rect -295 190 -275 210
rect -130 270 -110 290
rect -130 230 -110 250
rect -130 190 -110 210
rect -845 -150 -825 -130
rect -805 -150 -785 -130
rect -765 -150 -745 -130
rect -725 -150 -705 -130
rect -685 -150 -665 -130
rect -645 -150 -625 -130
rect -605 -150 -585 -130
rect -565 -150 -545 -130
rect -525 -150 -505 -130
rect -485 -150 -465 -130
rect -445 -150 -425 -130
rect -405 -150 -385 -130
rect -365 -150 -345 -130
rect -325 -150 -305 -130
rect -285 -150 -265 -130
rect -245 -150 -225 -130
rect -200 -150 -180 -130
rect -160 -150 -140 -130
rect -120 -150 -100 -130
rect -80 -150 -60 -130
rect -40 -150 -20 -130
<< metal1 >>
rect -865 850 0 865
rect -865 830 -845 850
rect -825 830 -805 850
rect -785 830 -765 850
rect -745 830 -725 850
rect -705 830 -685 850
rect -665 830 -645 850
rect -625 830 -605 850
rect -585 830 -565 850
rect -545 830 -525 850
rect -505 830 -485 850
rect -465 830 -445 850
rect -425 830 -405 850
rect -385 830 -365 850
rect -345 830 -325 850
rect -305 830 -285 850
rect -265 830 -245 850
rect -225 830 -205 850
rect -185 830 -160 850
rect -140 830 -120 850
rect -100 830 -80 850
rect -60 830 -40 850
rect -20 830 0 850
rect -865 815 0 830
rect -835 325 -815 815
rect -445 740 -425 815
rect -455 730 -415 740
rect -455 710 -445 730
rect -425 710 -415 730
rect -455 690 -415 710
rect -455 670 -445 690
rect -425 670 -415 690
rect -455 650 -415 670
rect -455 630 -445 650
rect -425 630 -415 650
rect -455 610 -415 630
rect -455 590 -445 610
rect -425 590 -415 610
rect -455 570 -415 590
rect -455 550 -445 570
rect -425 550 -415 570
rect -455 530 -415 550
rect -455 510 -445 530
rect -425 510 -415 530
rect -455 490 -415 510
rect -455 470 -445 490
rect -425 470 -415 490
rect -455 460 -415 470
rect -845 290 -805 325
rect -130 305 -110 815
rect -845 270 -835 290
rect -815 270 -805 290
rect -845 250 -805 270
rect -845 230 -835 250
rect -815 230 -805 250
rect -845 210 -805 230
rect -845 190 -835 210
rect -815 190 -805 210
rect -845 180 -805 190
rect -605 290 -565 305
rect -605 270 -595 290
rect -575 270 -565 290
rect -605 250 -565 270
rect -605 230 -595 250
rect -575 230 -565 250
rect -605 210 -565 230
rect -605 190 -595 210
rect -575 190 -565 210
rect -605 180 -565 190
rect -455 290 -415 305
rect -455 270 -445 290
rect -425 270 -415 290
rect -455 250 -415 270
rect -455 230 -445 250
rect -425 230 -415 250
rect -455 210 -415 230
rect -455 190 -445 210
rect -425 190 -415 210
rect -455 180 -415 190
rect -305 290 -265 305
rect -305 270 -295 290
rect -275 270 -265 290
rect -305 250 -265 270
rect -305 230 -295 250
rect -275 230 -265 250
rect -305 210 -265 230
rect -305 190 -295 210
rect -275 190 -265 210
rect -305 180 -265 190
rect -140 290 -100 305
rect -140 270 -130 290
rect -110 270 -100 290
rect -140 250 -100 270
rect -140 230 -130 250
rect -110 230 -100 250
rect -140 210 -100 230
rect -140 190 -130 210
rect -110 190 -100 210
rect -140 180 -100 190
rect -595 -115 -575 180
rect -445 -115 -425 180
rect -295 -115 -275 180
rect -865 -130 0 -115
rect -865 -150 -845 -130
rect -825 -150 -805 -130
rect -785 -150 -765 -130
rect -745 -150 -725 -130
rect -705 -150 -685 -130
rect -665 -150 -645 -130
rect -625 -150 -605 -130
rect -585 -150 -565 -130
rect -545 -150 -525 -130
rect -505 -150 -485 -130
rect -465 -150 -445 -130
rect -425 -150 -405 -130
rect -385 -150 -365 -130
rect -345 -150 -325 -130
rect -305 -150 -285 -130
rect -265 -150 -245 -130
rect -225 -150 -200 -130
rect -180 -150 -160 -130
rect -140 -150 -120 -130
rect -100 -150 -80 -130
rect -60 -150 -40 -130
rect -20 -150 0 -130
rect -865 -165 0 -150
<< labels >>
rlabel locali -640 135 -630 145 1 Dis
port 7 n
rlabel locali -240 355 -230 365 1 OUT
port 5 n
rlabel locali -625 350 -615 360 1 OUT_bar
port 6 n
rlabel locali -850 35 -840 45 1 B_bar
port 4 n
rlabel locali -850 85 -840 95 1 A_bar
port 2 n
rlabel locali -220 -15 -210 -5 1 A
port 1 n
rlabel locali -220 -75 -210 -65 1 B
port 3 n
rlabel metal1 -445 830 -425 850 1 CLK
port 8 n
rlabel metal1 -445 -150 -425 -130 5 GND!
port 9 s
<< end >>
