magic
tech sky130A
magscale 1 2
timestamp 1671307844
<< pwell >>
rect 35703 -2536 37555 -1492
rect 37607 -2536 39459 -1492
<< nmoslvt >>
rect 36029 -2518 36059 -1518
rect 36179 -2518 36209 -1518
rect 36329 -2518 36359 -1518
rect 36479 -2518 36509 -1518
rect 36629 -2518 36659 -1518
rect 36779 -2518 36809 -1518
rect 36929 -2518 36959 -1518
rect 37079 -2518 37109 -1518
rect 37229 -2518 37259 -1518
rect 37379 -2518 37409 -1518
rect 37933 -2510 37963 -1510
rect 38083 -2510 38113 -1510
rect 38233 -2510 38263 -1510
rect 38383 -2510 38413 -1510
rect 38533 -2510 38563 -1510
rect 38683 -2510 38713 -1510
rect 38833 -2510 38863 -1510
rect 38983 -2510 39013 -1510
rect 39133 -2510 39163 -1510
rect 39283 -2510 39313 -1510
<< ndiff >>
rect 35909 -1546 36029 -1518
rect 35909 -1580 35952 -1546
rect 35986 -1580 36029 -1546
rect 35909 -1614 36029 -1580
rect 35909 -1648 35952 -1614
rect 35986 -1648 36029 -1614
rect 35909 -1682 36029 -1648
rect 35909 -1716 35952 -1682
rect 35986 -1716 36029 -1682
rect 35909 -1750 36029 -1716
rect 35909 -1784 35952 -1750
rect 35986 -1784 36029 -1750
rect 35909 -1818 36029 -1784
rect 35909 -1852 35952 -1818
rect 35986 -1852 36029 -1818
rect 35909 -1886 36029 -1852
rect 35909 -1920 35952 -1886
rect 35986 -1920 36029 -1886
rect 35909 -1954 36029 -1920
rect 35909 -1988 35952 -1954
rect 35986 -1988 36029 -1954
rect 35909 -2022 36029 -1988
rect 35909 -2056 35952 -2022
rect 35986 -2056 36029 -2022
rect 35909 -2090 36029 -2056
rect 35909 -2124 35952 -2090
rect 35986 -2124 36029 -2090
rect 35909 -2158 36029 -2124
rect 35909 -2192 35952 -2158
rect 35986 -2192 36029 -2158
rect 35909 -2226 36029 -2192
rect 35909 -2260 35952 -2226
rect 35986 -2260 36029 -2226
rect 35909 -2294 36029 -2260
rect 35909 -2328 35952 -2294
rect 35986 -2328 36029 -2294
rect 35909 -2362 36029 -2328
rect 35909 -2396 35952 -2362
rect 35986 -2396 36029 -2362
rect 35909 -2430 36029 -2396
rect 35909 -2464 35952 -2430
rect 35986 -2464 36029 -2430
rect 35909 -2518 36029 -2464
rect 36059 -1546 36179 -1518
rect 36059 -1580 36102 -1546
rect 36136 -1580 36179 -1546
rect 36059 -1614 36179 -1580
rect 36059 -1648 36102 -1614
rect 36136 -1648 36179 -1614
rect 36059 -1682 36179 -1648
rect 36059 -1716 36102 -1682
rect 36136 -1716 36179 -1682
rect 36059 -1750 36179 -1716
rect 36059 -1784 36102 -1750
rect 36136 -1784 36179 -1750
rect 36059 -1818 36179 -1784
rect 36059 -1852 36102 -1818
rect 36136 -1852 36179 -1818
rect 36059 -1886 36179 -1852
rect 36059 -1920 36102 -1886
rect 36136 -1920 36179 -1886
rect 36059 -1954 36179 -1920
rect 36059 -1988 36102 -1954
rect 36136 -1988 36179 -1954
rect 36059 -2022 36179 -1988
rect 36059 -2056 36102 -2022
rect 36136 -2056 36179 -2022
rect 36059 -2090 36179 -2056
rect 36059 -2124 36102 -2090
rect 36136 -2124 36179 -2090
rect 36059 -2158 36179 -2124
rect 36059 -2192 36102 -2158
rect 36136 -2192 36179 -2158
rect 36059 -2226 36179 -2192
rect 36059 -2260 36102 -2226
rect 36136 -2260 36179 -2226
rect 36059 -2294 36179 -2260
rect 36059 -2328 36102 -2294
rect 36136 -2328 36179 -2294
rect 36059 -2362 36179 -2328
rect 36059 -2396 36102 -2362
rect 36136 -2396 36179 -2362
rect 36059 -2430 36179 -2396
rect 36059 -2464 36102 -2430
rect 36136 -2464 36179 -2430
rect 36059 -2518 36179 -2464
rect 36209 -1546 36329 -1518
rect 36209 -1580 36252 -1546
rect 36286 -1580 36329 -1546
rect 36209 -1614 36329 -1580
rect 36209 -1648 36252 -1614
rect 36286 -1648 36329 -1614
rect 36209 -1682 36329 -1648
rect 36209 -1716 36252 -1682
rect 36286 -1716 36329 -1682
rect 36209 -1750 36329 -1716
rect 36209 -1784 36252 -1750
rect 36286 -1784 36329 -1750
rect 36209 -1818 36329 -1784
rect 36209 -1852 36252 -1818
rect 36286 -1852 36329 -1818
rect 36209 -1886 36329 -1852
rect 36209 -1920 36252 -1886
rect 36286 -1920 36329 -1886
rect 36209 -1954 36329 -1920
rect 36209 -1988 36252 -1954
rect 36286 -1988 36329 -1954
rect 36209 -2022 36329 -1988
rect 36209 -2056 36252 -2022
rect 36286 -2056 36329 -2022
rect 36209 -2090 36329 -2056
rect 36209 -2124 36252 -2090
rect 36286 -2124 36329 -2090
rect 36209 -2158 36329 -2124
rect 36209 -2192 36252 -2158
rect 36286 -2192 36329 -2158
rect 36209 -2226 36329 -2192
rect 36209 -2260 36252 -2226
rect 36286 -2260 36329 -2226
rect 36209 -2294 36329 -2260
rect 36209 -2328 36252 -2294
rect 36286 -2328 36329 -2294
rect 36209 -2362 36329 -2328
rect 36209 -2396 36252 -2362
rect 36286 -2396 36329 -2362
rect 36209 -2430 36329 -2396
rect 36209 -2464 36252 -2430
rect 36286 -2464 36329 -2430
rect 36209 -2518 36329 -2464
rect 36359 -1546 36479 -1518
rect 36359 -1580 36402 -1546
rect 36436 -1580 36479 -1546
rect 36359 -1614 36479 -1580
rect 36359 -1648 36402 -1614
rect 36436 -1648 36479 -1614
rect 36359 -1682 36479 -1648
rect 36359 -1716 36402 -1682
rect 36436 -1716 36479 -1682
rect 36359 -1750 36479 -1716
rect 36359 -1784 36402 -1750
rect 36436 -1784 36479 -1750
rect 36359 -1818 36479 -1784
rect 36359 -1852 36402 -1818
rect 36436 -1852 36479 -1818
rect 36359 -1886 36479 -1852
rect 36359 -1920 36402 -1886
rect 36436 -1920 36479 -1886
rect 36359 -1954 36479 -1920
rect 36359 -1988 36402 -1954
rect 36436 -1988 36479 -1954
rect 36359 -2022 36479 -1988
rect 36359 -2056 36402 -2022
rect 36436 -2056 36479 -2022
rect 36359 -2090 36479 -2056
rect 36359 -2124 36402 -2090
rect 36436 -2124 36479 -2090
rect 36359 -2158 36479 -2124
rect 36359 -2192 36402 -2158
rect 36436 -2192 36479 -2158
rect 36359 -2226 36479 -2192
rect 36359 -2260 36402 -2226
rect 36436 -2260 36479 -2226
rect 36359 -2294 36479 -2260
rect 36359 -2328 36402 -2294
rect 36436 -2328 36479 -2294
rect 36359 -2362 36479 -2328
rect 36359 -2396 36402 -2362
rect 36436 -2396 36479 -2362
rect 36359 -2430 36479 -2396
rect 36359 -2464 36402 -2430
rect 36436 -2464 36479 -2430
rect 36359 -2518 36479 -2464
rect 36509 -1546 36629 -1518
rect 36509 -1580 36552 -1546
rect 36586 -1580 36629 -1546
rect 36509 -1614 36629 -1580
rect 36509 -1648 36552 -1614
rect 36586 -1648 36629 -1614
rect 36509 -1682 36629 -1648
rect 36509 -1716 36552 -1682
rect 36586 -1716 36629 -1682
rect 36509 -1750 36629 -1716
rect 36509 -1784 36552 -1750
rect 36586 -1784 36629 -1750
rect 36509 -1818 36629 -1784
rect 36509 -1852 36552 -1818
rect 36586 -1852 36629 -1818
rect 36509 -1886 36629 -1852
rect 36509 -1920 36552 -1886
rect 36586 -1920 36629 -1886
rect 36509 -1954 36629 -1920
rect 36509 -1988 36552 -1954
rect 36586 -1988 36629 -1954
rect 36509 -2022 36629 -1988
rect 36509 -2056 36552 -2022
rect 36586 -2056 36629 -2022
rect 36509 -2090 36629 -2056
rect 36509 -2124 36552 -2090
rect 36586 -2124 36629 -2090
rect 36509 -2158 36629 -2124
rect 36509 -2192 36552 -2158
rect 36586 -2192 36629 -2158
rect 36509 -2226 36629 -2192
rect 36509 -2260 36552 -2226
rect 36586 -2260 36629 -2226
rect 36509 -2294 36629 -2260
rect 36509 -2328 36552 -2294
rect 36586 -2328 36629 -2294
rect 36509 -2362 36629 -2328
rect 36509 -2396 36552 -2362
rect 36586 -2396 36629 -2362
rect 36509 -2430 36629 -2396
rect 36509 -2464 36552 -2430
rect 36586 -2464 36629 -2430
rect 36509 -2518 36629 -2464
rect 36659 -1546 36779 -1518
rect 36659 -1580 36702 -1546
rect 36736 -1580 36779 -1546
rect 36659 -1614 36779 -1580
rect 36659 -1648 36702 -1614
rect 36736 -1648 36779 -1614
rect 36659 -1682 36779 -1648
rect 36659 -1716 36702 -1682
rect 36736 -1716 36779 -1682
rect 36659 -1750 36779 -1716
rect 36659 -1784 36702 -1750
rect 36736 -1784 36779 -1750
rect 36659 -1818 36779 -1784
rect 36659 -1852 36702 -1818
rect 36736 -1852 36779 -1818
rect 36659 -1886 36779 -1852
rect 36659 -1920 36702 -1886
rect 36736 -1920 36779 -1886
rect 36659 -1954 36779 -1920
rect 36659 -1988 36702 -1954
rect 36736 -1988 36779 -1954
rect 36659 -2022 36779 -1988
rect 36659 -2056 36702 -2022
rect 36736 -2056 36779 -2022
rect 36659 -2090 36779 -2056
rect 36659 -2124 36702 -2090
rect 36736 -2124 36779 -2090
rect 36659 -2158 36779 -2124
rect 36659 -2192 36702 -2158
rect 36736 -2192 36779 -2158
rect 36659 -2226 36779 -2192
rect 36659 -2260 36702 -2226
rect 36736 -2260 36779 -2226
rect 36659 -2294 36779 -2260
rect 36659 -2328 36702 -2294
rect 36736 -2328 36779 -2294
rect 36659 -2362 36779 -2328
rect 36659 -2396 36702 -2362
rect 36736 -2396 36779 -2362
rect 36659 -2430 36779 -2396
rect 36659 -2464 36702 -2430
rect 36736 -2464 36779 -2430
rect 36659 -2518 36779 -2464
rect 36809 -1546 36929 -1518
rect 36809 -1580 36852 -1546
rect 36886 -1580 36929 -1546
rect 36809 -1614 36929 -1580
rect 36809 -1648 36852 -1614
rect 36886 -1648 36929 -1614
rect 36809 -1682 36929 -1648
rect 36809 -1716 36852 -1682
rect 36886 -1716 36929 -1682
rect 36809 -1750 36929 -1716
rect 36809 -1784 36852 -1750
rect 36886 -1784 36929 -1750
rect 36809 -1818 36929 -1784
rect 36809 -1852 36852 -1818
rect 36886 -1852 36929 -1818
rect 36809 -1886 36929 -1852
rect 36809 -1920 36852 -1886
rect 36886 -1920 36929 -1886
rect 36809 -1954 36929 -1920
rect 36809 -1988 36852 -1954
rect 36886 -1988 36929 -1954
rect 36809 -2022 36929 -1988
rect 36809 -2056 36852 -2022
rect 36886 -2056 36929 -2022
rect 36809 -2090 36929 -2056
rect 36809 -2124 36852 -2090
rect 36886 -2124 36929 -2090
rect 36809 -2158 36929 -2124
rect 36809 -2192 36852 -2158
rect 36886 -2192 36929 -2158
rect 36809 -2226 36929 -2192
rect 36809 -2260 36852 -2226
rect 36886 -2260 36929 -2226
rect 36809 -2294 36929 -2260
rect 36809 -2328 36852 -2294
rect 36886 -2328 36929 -2294
rect 36809 -2362 36929 -2328
rect 36809 -2396 36852 -2362
rect 36886 -2396 36929 -2362
rect 36809 -2430 36929 -2396
rect 36809 -2464 36852 -2430
rect 36886 -2464 36929 -2430
rect 36809 -2518 36929 -2464
rect 36959 -1546 37079 -1518
rect 36959 -1580 37002 -1546
rect 37036 -1580 37079 -1546
rect 36959 -1614 37079 -1580
rect 36959 -1648 37002 -1614
rect 37036 -1648 37079 -1614
rect 36959 -1682 37079 -1648
rect 36959 -1716 37002 -1682
rect 37036 -1716 37079 -1682
rect 36959 -1750 37079 -1716
rect 36959 -1784 37002 -1750
rect 37036 -1784 37079 -1750
rect 36959 -1818 37079 -1784
rect 36959 -1852 37002 -1818
rect 37036 -1852 37079 -1818
rect 36959 -1886 37079 -1852
rect 36959 -1920 37002 -1886
rect 37036 -1920 37079 -1886
rect 36959 -1954 37079 -1920
rect 36959 -1988 37002 -1954
rect 37036 -1988 37079 -1954
rect 36959 -2022 37079 -1988
rect 36959 -2056 37002 -2022
rect 37036 -2056 37079 -2022
rect 36959 -2090 37079 -2056
rect 36959 -2124 37002 -2090
rect 37036 -2124 37079 -2090
rect 36959 -2158 37079 -2124
rect 36959 -2192 37002 -2158
rect 37036 -2192 37079 -2158
rect 36959 -2226 37079 -2192
rect 36959 -2260 37002 -2226
rect 37036 -2260 37079 -2226
rect 36959 -2294 37079 -2260
rect 36959 -2328 37002 -2294
rect 37036 -2328 37079 -2294
rect 36959 -2362 37079 -2328
rect 36959 -2396 37002 -2362
rect 37036 -2396 37079 -2362
rect 36959 -2430 37079 -2396
rect 36959 -2464 37002 -2430
rect 37036 -2464 37079 -2430
rect 36959 -2518 37079 -2464
rect 37109 -1546 37229 -1518
rect 37109 -1580 37152 -1546
rect 37186 -1580 37229 -1546
rect 37109 -1614 37229 -1580
rect 37109 -1648 37152 -1614
rect 37186 -1648 37229 -1614
rect 37109 -1682 37229 -1648
rect 37109 -1716 37152 -1682
rect 37186 -1716 37229 -1682
rect 37109 -1750 37229 -1716
rect 37109 -1784 37152 -1750
rect 37186 -1784 37229 -1750
rect 37109 -1818 37229 -1784
rect 37109 -1852 37152 -1818
rect 37186 -1852 37229 -1818
rect 37109 -1886 37229 -1852
rect 37109 -1920 37152 -1886
rect 37186 -1920 37229 -1886
rect 37109 -1954 37229 -1920
rect 37109 -1988 37152 -1954
rect 37186 -1988 37229 -1954
rect 37109 -2022 37229 -1988
rect 37109 -2056 37152 -2022
rect 37186 -2056 37229 -2022
rect 37109 -2090 37229 -2056
rect 37109 -2124 37152 -2090
rect 37186 -2124 37229 -2090
rect 37109 -2158 37229 -2124
rect 37109 -2192 37152 -2158
rect 37186 -2192 37229 -2158
rect 37109 -2226 37229 -2192
rect 37109 -2260 37152 -2226
rect 37186 -2260 37229 -2226
rect 37109 -2294 37229 -2260
rect 37109 -2328 37152 -2294
rect 37186 -2328 37229 -2294
rect 37109 -2362 37229 -2328
rect 37109 -2396 37152 -2362
rect 37186 -2396 37229 -2362
rect 37109 -2430 37229 -2396
rect 37109 -2464 37152 -2430
rect 37186 -2464 37229 -2430
rect 37109 -2518 37229 -2464
rect 37259 -1546 37379 -1518
rect 37259 -1580 37302 -1546
rect 37336 -1580 37379 -1546
rect 37259 -1614 37379 -1580
rect 37259 -1648 37302 -1614
rect 37336 -1648 37379 -1614
rect 37259 -1682 37379 -1648
rect 37259 -1716 37302 -1682
rect 37336 -1716 37379 -1682
rect 37259 -1750 37379 -1716
rect 37259 -1784 37302 -1750
rect 37336 -1784 37379 -1750
rect 37259 -1818 37379 -1784
rect 37259 -1852 37302 -1818
rect 37336 -1852 37379 -1818
rect 37259 -1886 37379 -1852
rect 37259 -1920 37302 -1886
rect 37336 -1920 37379 -1886
rect 37259 -1954 37379 -1920
rect 37259 -1988 37302 -1954
rect 37336 -1988 37379 -1954
rect 37259 -2022 37379 -1988
rect 37259 -2056 37302 -2022
rect 37336 -2056 37379 -2022
rect 37259 -2090 37379 -2056
rect 37259 -2124 37302 -2090
rect 37336 -2124 37379 -2090
rect 37259 -2158 37379 -2124
rect 37259 -2192 37302 -2158
rect 37336 -2192 37379 -2158
rect 37259 -2226 37379 -2192
rect 37259 -2260 37302 -2226
rect 37336 -2260 37379 -2226
rect 37259 -2294 37379 -2260
rect 37259 -2328 37302 -2294
rect 37336 -2328 37379 -2294
rect 37259 -2362 37379 -2328
rect 37259 -2396 37302 -2362
rect 37336 -2396 37379 -2362
rect 37259 -2430 37379 -2396
rect 37259 -2464 37302 -2430
rect 37336 -2464 37379 -2430
rect 37259 -2518 37379 -2464
rect 37409 -1546 37529 -1518
rect 37409 -1580 37452 -1546
rect 37486 -1580 37529 -1546
rect 37409 -1614 37529 -1580
rect 37409 -1648 37452 -1614
rect 37486 -1648 37529 -1614
rect 37409 -1682 37529 -1648
rect 37409 -1716 37452 -1682
rect 37486 -1716 37529 -1682
rect 37409 -1750 37529 -1716
rect 37409 -1784 37452 -1750
rect 37486 -1784 37529 -1750
rect 37409 -1818 37529 -1784
rect 37409 -1852 37452 -1818
rect 37486 -1852 37529 -1818
rect 37409 -1886 37529 -1852
rect 37409 -1920 37452 -1886
rect 37486 -1920 37529 -1886
rect 37409 -1954 37529 -1920
rect 37409 -1988 37452 -1954
rect 37486 -1988 37529 -1954
rect 37409 -2022 37529 -1988
rect 37409 -2056 37452 -2022
rect 37486 -2056 37529 -2022
rect 37409 -2090 37529 -2056
rect 37409 -2124 37452 -2090
rect 37486 -2124 37529 -2090
rect 37409 -2158 37529 -2124
rect 37409 -2192 37452 -2158
rect 37486 -2192 37529 -2158
rect 37409 -2226 37529 -2192
rect 37409 -2260 37452 -2226
rect 37486 -2260 37529 -2226
rect 37409 -2294 37529 -2260
rect 37409 -2328 37452 -2294
rect 37486 -2328 37529 -2294
rect 37409 -2362 37529 -2328
rect 37409 -2396 37452 -2362
rect 37486 -2396 37529 -2362
rect 37409 -2430 37529 -2396
rect 37409 -2464 37452 -2430
rect 37486 -2464 37529 -2430
rect 37409 -2518 37529 -2464
rect 37813 -1546 37933 -1510
rect 37813 -1580 37856 -1546
rect 37890 -1580 37933 -1546
rect 37813 -1614 37933 -1580
rect 37813 -1648 37856 -1614
rect 37890 -1648 37933 -1614
rect 37813 -1682 37933 -1648
rect 37813 -1716 37856 -1682
rect 37890 -1716 37933 -1682
rect 37813 -1750 37933 -1716
rect 37813 -1784 37856 -1750
rect 37890 -1784 37933 -1750
rect 37813 -1818 37933 -1784
rect 37813 -1852 37856 -1818
rect 37890 -1852 37933 -1818
rect 37813 -1886 37933 -1852
rect 37813 -1920 37856 -1886
rect 37890 -1920 37933 -1886
rect 37813 -1954 37933 -1920
rect 37813 -1988 37856 -1954
rect 37890 -1988 37933 -1954
rect 37813 -2022 37933 -1988
rect 37813 -2056 37856 -2022
rect 37890 -2056 37933 -2022
rect 37813 -2090 37933 -2056
rect 37813 -2124 37856 -2090
rect 37890 -2124 37933 -2090
rect 37813 -2158 37933 -2124
rect 37813 -2192 37856 -2158
rect 37890 -2192 37933 -2158
rect 37813 -2226 37933 -2192
rect 37813 -2260 37856 -2226
rect 37890 -2260 37933 -2226
rect 37813 -2294 37933 -2260
rect 37813 -2328 37856 -2294
rect 37890 -2328 37933 -2294
rect 37813 -2362 37933 -2328
rect 37813 -2396 37856 -2362
rect 37890 -2396 37933 -2362
rect 37813 -2430 37933 -2396
rect 37813 -2464 37856 -2430
rect 37890 -2464 37933 -2430
rect 37813 -2510 37933 -2464
rect 37963 -1546 38083 -1510
rect 37963 -1580 38006 -1546
rect 38040 -1580 38083 -1546
rect 37963 -1614 38083 -1580
rect 37963 -1648 38006 -1614
rect 38040 -1648 38083 -1614
rect 37963 -1682 38083 -1648
rect 37963 -1716 38006 -1682
rect 38040 -1716 38083 -1682
rect 37963 -1750 38083 -1716
rect 37963 -1784 38006 -1750
rect 38040 -1784 38083 -1750
rect 37963 -1818 38083 -1784
rect 37963 -1852 38006 -1818
rect 38040 -1852 38083 -1818
rect 37963 -1886 38083 -1852
rect 37963 -1920 38006 -1886
rect 38040 -1920 38083 -1886
rect 37963 -1954 38083 -1920
rect 37963 -1988 38006 -1954
rect 38040 -1988 38083 -1954
rect 37963 -2022 38083 -1988
rect 37963 -2056 38006 -2022
rect 38040 -2056 38083 -2022
rect 37963 -2090 38083 -2056
rect 37963 -2124 38006 -2090
rect 38040 -2124 38083 -2090
rect 37963 -2158 38083 -2124
rect 37963 -2192 38006 -2158
rect 38040 -2192 38083 -2158
rect 37963 -2226 38083 -2192
rect 37963 -2260 38006 -2226
rect 38040 -2260 38083 -2226
rect 37963 -2294 38083 -2260
rect 37963 -2328 38006 -2294
rect 38040 -2328 38083 -2294
rect 37963 -2362 38083 -2328
rect 37963 -2396 38006 -2362
rect 38040 -2396 38083 -2362
rect 37963 -2430 38083 -2396
rect 37963 -2464 38006 -2430
rect 38040 -2464 38083 -2430
rect 37963 -2510 38083 -2464
rect 38113 -1546 38233 -1510
rect 38113 -1580 38156 -1546
rect 38190 -1580 38233 -1546
rect 38113 -1614 38233 -1580
rect 38113 -1648 38156 -1614
rect 38190 -1648 38233 -1614
rect 38113 -1682 38233 -1648
rect 38113 -1716 38156 -1682
rect 38190 -1716 38233 -1682
rect 38113 -1750 38233 -1716
rect 38113 -1784 38156 -1750
rect 38190 -1784 38233 -1750
rect 38113 -1818 38233 -1784
rect 38113 -1852 38156 -1818
rect 38190 -1852 38233 -1818
rect 38113 -1886 38233 -1852
rect 38113 -1920 38156 -1886
rect 38190 -1920 38233 -1886
rect 38113 -1954 38233 -1920
rect 38113 -1988 38156 -1954
rect 38190 -1988 38233 -1954
rect 38113 -2022 38233 -1988
rect 38113 -2056 38156 -2022
rect 38190 -2056 38233 -2022
rect 38113 -2090 38233 -2056
rect 38113 -2124 38156 -2090
rect 38190 -2124 38233 -2090
rect 38113 -2158 38233 -2124
rect 38113 -2192 38156 -2158
rect 38190 -2192 38233 -2158
rect 38113 -2226 38233 -2192
rect 38113 -2260 38156 -2226
rect 38190 -2260 38233 -2226
rect 38113 -2294 38233 -2260
rect 38113 -2328 38156 -2294
rect 38190 -2328 38233 -2294
rect 38113 -2362 38233 -2328
rect 38113 -2396 38156 -2362
rect 38190 -2396 38233 -2362
rect 38113 -2430 38233 -2396
rect 38113 -2464 38156 -2430
rect 38190 -2464 38233 -2430
rect 38113 -2510 38233 -2464
rect 38263 -1546 38383 -1510
rect 38263 -1580 38306 -1546
rect 38340 -1580 38383 -1546
rect 38263 -1614 38383 -1580
rect 38263 -1648 38306 -1614
rect 38340 -1648 38383 -1614
rect 38263 -1682 38383 -1648
rect 38263 -1716 38306 -1682
rect 38340 -1716 38383 -1682
rect 38263 -1750 38383 -1716
rect 38263 -1784 38306 -1750
rect 38340 -1784 38383 -1750
rect 38263 -1818 38383 -1784
rect 38263 -1852 38306 -1818
rect 38340 -1852 38383 -1818
rect 38263 -1886 38383 -1852
rect 38263 -1920 38306 -1886
rect 38340 -1920 38383 -1886
rect 38263 -1954 38383 -1920
rect 38263 -1988 38306 -1954
rect 38340 -1988 38383 -1954
rect 38263 -2022 38383 -1988
rect 38263 -2056 38306 -2022
rect 38340 -2056 38383 -2022
rect 38263 -2090 38383 -2056
rect 38263 -2124 38306 -2090
rect 38340 -2124 38383 -2090
rect 38263 -2158 38383 -2124
rect 38263 -2192 38306 -2158
rect 38340 -2192 38383 -2158
rect 38263 -2226 38383 -2192
rect 38263 -2260 38306 -2226
rect 38340 -2260 38383 -2226
rect 38263 -2294 38383 -2260
rect 38263 -2328 38306 -2294
rect 38340 -2328 38383 -2294
rect 38263 -2362 38383 -2328
rect 38263 -2396 38306 -2362
rect 38340 -2396 38383 -2362
rect 38263 -2430 38383 -2396
rect 38263 -2464 38306 -2430
rect 38340 -2464 38383 -2430
rect 38263 -2510 38383 -2464
rect 38413 -1546 38533 -1510
rect 38413 -1580 38456 -1546
rect 38490 -1580 38533 -1546
rect 38413 -1614 38533 -1580
rect 38413 -1648 38456 -1614
rect 38490 -1648 38533 -1614
rect 38413 -1682 38533 -1648
rect 38413 -1716 38456 -1682
rect 38490 -1716 38533 -1682
rect 38413 -1750 38533 -1716
rect 38413 -1784 38456 -1750
rect 38490 -1784 38533 -1750
rect 38413 -1818 38533 -1784
rect 38413 -1852 38456 -1818
rect 38490 -1852 38533 -1818
rect 38413 -1886 38533 -1852
rect 38413 -1920 38456 -1886
rect 38490 -1920 38533 -1886
rect 38413 -1954 38533 -1920
rect 38413 -1988 38456 -1954
rect 38490 -1988 38533 -1954
rect 38413 -2022 38533 -1988
rect 38413 -2056 38456 -2022
rect 38490 -2056 38533 -2022
rect 38413 -2090 38533 -2056
rect 38413 -2124 38456 -2090
rect 38490 -2124 38533 -2090
rect 38413 -2158 38533 -2124
rect 38413 -2192 38456 -2158
rect 38490 -2192 38533 -2158
rect 38413 -2226 38533 -2192
rect 38413 -2260 38456 -2226
rect 38490 -2260 38533 -2226
rect 38413 -2294 38533 -2260
rect 38413 -2328 38456 -2294
rect 38490 -2328 38533 -2294
rect 38413 -2362 38533 -2328
rect 38413 -2396 38456 -2362
rect 38490 -2396 38533 -2362
rect 38413 -2430 38533 -2396
rect 38413 -2464 38456 -2430
rect 38490 -2464 38533 -2430
rect 38413 -2510 38533 -2464
rect 38563 -1546 38683 -1510
rect 38563 -1580 38606 -1546
rect 38640 -1580 38683 -1546
rect 38563 -1614 38683 -1580
rect 38563 -1648 38606 -1614
rect 38640 -1648 38683 -1614
rect 38563 -1682 38683 -1648
rect 38563 -1716 38606 -1682
rect 38640 -1716 38683 -1682
rect 38563 -1750 38683 -1716
rect 38563 -1784 38606 -1750
rect 38640 -1784 38683 -1750
rect 38563 -1818 38683 -1784
rect 38563 -1852 38606 -1818
rect 38640 -1852 38683 -1818
rect 38563 -1886 38683 -1852
rect 38563 -1920 38606 -1886
rect 38640 -1920 38683 -1886
rect 38563 -1954 38683 -1920
rect 38563 -1988 38606 -1954
rect 38640 -1988 38683 -1954
rect 38563 -2022 38683 -1988
rect 38563 -2056 38606 -2022
rect 38640 -2056 38683 -2022
rect 38563 -2090 38683 -2056
rect 38563 -2124 38606 -2090
rect 38640 -2124 38683 -2090
rect 38563 -2158 38683 -2124
rect 38563 -2192 38606 -2158
rect 38640 -2192 38683 -2158
rect 38563 -2226 38683 -2192
rect 38563 -2260 38606 -2226
rect 38640 -2260 38683 -2226
rect 38563 -2294 38683 -2260
rect 38563 -2328 38606 -2294
rect 38640 -2328 38683 -2294
rect 38563 -2362 38683 -2328
rect 38563 -2396 38606 -2362
rect 38640 -2396 38683 -2362
rect 38563 -2430 38683 -2396
rect 38563 -2464 38606 -2430
rect 38640 -2464 38683 -2430
rect 38563 -2510 38683 -2464
rect 38713 -1546 38833 -1510
rect 38713 -1580 38756 -1546
rect 38790 -1580 38833 -1546
rect 38713 -1614 38833 -1580
rect 38713 -1648 38756 -1614
rect 38790 -1648 38833 -1614
rect 38713 -1682 38833 -1648
rect 38713 -1716 38756 -1682
rect 38790 -1716 38833 -1682
rect 38713 -1750 38833 -1716
rect 38713 -1784 38756 -1750
rect 38790 -1784 38833 -1750
rect 38713 -1818 38833 -1784
rect 38713 -1852 38756 -1818
rect 38790 -1852 38833 -1818
rect 38713 -1886 38833 -1852
rect 38713 -1920 38756 -1886
rect 38790 -1920 38833 -1886
rect 38713 -1954 38833 -1920
rect 38713 -1988 38756 -1954
rect 38790 -1988 38833 -1954
rect 38713 -2022 38833 -1988
rect 38713 -2056 38756 -2022
rect 38790 -2056 38833 -2022
rect 38713 -2090 38833 -2056
rect 38713 -2124 38756 -2090
rect 38790 -2124 38833 -2090
rect 38713 -2158 38833 -2124
rect 38713 -2192 38756 -2158
rect 38790 -2192 38833 -2158
rect 38713 -2226 38833 -2192
rect 38713 -2260 38756 -2226
rect 38790 -2260 38833 -2226
rect 38713 -2294 38833 -2260
rect 38713 -2328 38756 -2294
rect 38790 -2328 38833 -2294
rect 38713 -2362 38833 -2328
rect 38713 -2396 38756 -2362
rect 38790 -2396 38833 -2362
rect 38713 -2430 38833 -2396
rect 38713 -2464 38756 -2430
rect 38790 -2464 38833 -2430
rect 38713 -2510 38833 -2464
rect 38863 -1546 38983 -1510
rect 38863 -1580 38906 -1546
rect 38940 -1580 38983 -1546
rect 38863 -1614 38983 -1580
rect 38863 -1648 38906 -1614
rect 38940 -1648 38983 -1614
rect 38863 -1682 38983 -1648
rect 38863 -1716 38906 -1682
rect 38940 -1716 38983 -1682
rect 38863 -1750 38983 -1716
rect 38863 -1784 38906 -1750
rect 38940 -1784 38983 -1750
rect 38863 -1818 38983 -1784
rect 38863 -1852 38906 -1818
rect 38940 -1852 38983 -1818
rect 38863 -1886 38983 -1852
rect 38863 -1920 38906 -1886
rect 38940 -1920 38983 -1886
rect 38863 -1954 38983 -1920
rect 38863 -1988 38906 -1954
rect 38940 -1988 38983 -1954
rect 38863 -2022 38983 -1988
rect 38863 -2056 38906 -2022
rect 38940 -2056 38983 -2022
rect 38863 -2090 38983 -2056
rect 38863 -2124 38906 -2090
rect 38940 -2124 38983 -2090
rect 38863 -2158 38983 -2124
rect 38863 -2192 38906 -2158
rect 38940 -2192 38983 -2158
rect 38863 -2226 38983 -2192
rect 38863 -2260 38906 -2226
rect 38940 -2260 38983 -2226
rect 38863 -2294 38983 -2260
rect 38863 -2328 38906 -2294
rect 38940 -2328 38983 -2294
rect 38863 -2362 38983 -2328
rect 38863 -2396 38906 -2362
rect 38940 -2396 38983 -2362
rect 38863 -2430 38983 -2396
rect 38863 -2464 38906 -2430
rect 38940 -2464 38983 -2430
rect 38863 -2510 38983 -2464
rect 39013 -1546 39133 -1510
rect 39013 -1580 39056 -1546
rect 39090 -1580 39133 -1546
rect 39013 -1614 39133 -1580
rect 39013 -1648 39056 -1614
rect 39090 -1648 39133 -1614
rect 39013 -1682 39133 -1648
rect 39013 -1716 39056 -1682
rect 39090 -1716 39133 -1682
rect 39013 -1750 39133 -1716
rect 39013 -1784 39056 -1750
rect 39090 -1784 39133 -1750
rect 39013 -1818 39133 -1784
rect 39013 -1852 39056 -1818
rect 39090 -1852 39133 -1818
rect 39013 -1886 39133 -1852
rect 39013 -1920 39056 -1886
rect 39090 -1920 39133 -1886
rect 39013 -1954 39133 -1920
rect 39013 -1988 39056 -1954
rect 39090 -1988 39133 -1954
rect 39013 -2022 39133 -1988
rect 39013 -2056 39056 -2022
rect 39090 -2056 39133 -2022
rect 39013 -2090 39133 -2056
rect 39013 -2124 39056 -2090
rect 39090 -2124 39133 -2090
rect 39013 -2158 39133 -2124
rect 39013 -2192 39056 -2158
rect 39090 -2192 39133 -2158
rect 39013 -2226 39133 -2192
rect 39013 -2260 39056 -2226
rect 39090 -2260 39133 -2226
rect 39013 -2294 39133 -2260
rect 39013 -2328 39056 -2294
rect 39090 -2328 39133 -2294
rect 39013 -2362 39133 -2328
rect 39013 -2396 39056 -2362
rect 39090 -2396 39133 -2362
rect 39013 -2430 39133 -2396
rect 39013 -2464 39056 -2430
rect 39090 -2464 39133 -2430
rect 39013 -2510 39133 -2464
rect 39163 -1546 39283 -1510
rect 39163 -1580 39206 -1546
rect 39240 -1580 39283 -1546
rect 39163 -1614 39283 -1580
rect 39163 -1648 39206 -1614
rect 39240 -1648 39283 -1614
rect 39163 -1682 39283 -1648
rect 39163 -1716 39206 -1682
rect 39240 -1716 39283 -1682
rect 39163 -1750 39283 -1716
rect 39163 -1784 39206 -1750
rect 39240 -1784 39283 -1750
rect 39163 -1818 39283 -1784
rect 39163 -1852 39206 -1818
rect 39240 -1852 39283 -1818
rect 39163 -1886 39283 -1852
rect 39163 -1920 39206 -1886
rect 39240 -1920 39283 -1886
rect 39163 -1954 39283 -1920
rect 39163 -1988 39206 -1954
rect 39240 -1988 39283 -1954
rect 39163 -2022 39283 -1988
rect 39163 -2056 39206 -2022
rect 39240 -2056 39283 -2022
rect 39163 -2090 39283 -2056
rect 39163 -2124 39206 -2090
rect 39240 -2124 39283 -2090
rect 39163 -2158 39283 -2124
rect 39163 -2192 39206 -2158
rect 39240 -2192 39283 -2158
rect 39163 -2226 39283 -2192
rect 39163 -2260 39206 -2226
rect 39240 -2260 39283 -2226
rect 39163 -2294 39283 -2260
rect 39163 -2328 39206 -2294
rect 39240 -2328 39283 -2294
rect 39163 -2362 39283 -2328
rect 39163 -2396 39206 -2362
rect 39240 -2396 39283 -2362
rect 39163 -2430 39283 -2396
rect 39163 -2464 39206 -2430
rect 39240 -2464 39283 -2430
rect 39163 -2510 39283 -2464
rect 39313 -1546 39433 -1510
rect 39313 -1580 39356 -1546
rect 39390 -1580 39433 -1546
rect 39313 -1614 39433 -1580
rect 39313 -1648 39356 -1614
rect 39390 -1648 39433 -1614
rect 39313 -1682 39433 -1648
rect 39313 -1716 39356 -1682
rect 39390 -1716 39433 -1682
rect 39313 -1750 39433 -1716
rect 39313 -1784 39356 -1750
rect 39390 -1784 39433 -1750
rect 39313 -1818 39433 -1784
rect 39313 -1852 39356 -1818
rect 39390 -1852 39433 -1818
rect 39313 -1886 39433 -1852
rect 39313 -1920 39356 -1886
rect 39390 -1920 39433 -1886
rect 39313 -1954 39433 -1920
rect 39313 -1988 39356 -1954
rect 39390 -1988 39433 -1954
rect 39313 -2022 39433 -1988
rect 39313 -2056 39356 -2022
rect 39390 -2056 39433 -2022
rect 39313 -2090 39433 -2056
rect 39313 -2124 39356 -2090
rect 39390 -2124 39433 -2090
rect 39313 -2158 39433 -2124
rect 39313 -2192 39356 -2158
rect 39390 -2192 39433 -2158
rect 39313 -2226 39433 -2192
rect 39313 -2260 39356 -2226
rect 39390 -2260 39433 -2226
rect 39313 -2294 39433 -2260
rect 39313 -2328 39356 -2294
rect 39390 -2328 39433 -2294
rect 39313 -2362 39433 -2328
rect 39313 -2396 39356 -2362
rect 39390 -2396 39433 -2362
rect 39313 -2430 39433 -2396
rect 39313 -2464 39356 -2430
rect 39390 -2464 39433 -2430
rect 39313 -2510 39433 -2464
<< ndiffc >>
rect 35952 -1580 35986 -1546
rect 35952 -1648 35986 -1614
rect 35952 -1716 35986 -1682
rect 35952 -1784 35986 -1750
rect 35952 -1852 35986 -1818
rect 35952 -1920 35986 -1886
rect 35952 -1988 35986 -1954
rect 35952 -2056 35986 -2022
rect 35952 -2124 35986 -2090
rect 35952 -2192 35986 -2158
rect 35952 -2260 35986 -2226
rect 35952 -2328 35986 -2294
rect 35952 -2396 35986 -2362
rect 35952 -2464 35986 -2430
rect 36102 -1580 36136 -1546
rect 36102 -1648 36136 -1614
rect 36102 -1716 36136 -1682
rect 36102 -1784 36136 -1750
rect 36102 -1852 36136 -1818
rect 36102 -1920 36136 -1886
rect 36102 -1988 36136 -1954
rect 36102 -2056 36136 -2022
rect 36102 -2124 36136 -2090
rect 36102 -2192 36136 -2158
rect 36102 -2260 36136 -2226
rect 36102 -2328 36136 -2294
rect 36102 -2396 36136 -2362
rect 36102 -2464 36136 -2430
rect 36252 -1580 36286 -1546
rect 36252 -1648 36286 -1614
rect 36252 -1716 36286 -1682
rect 36252 -1784 36286 -1750
rect 36252 -1852 36286 -1818
rect 36252 -1920 36286 -1886
rect 36252 -1988 36286 -1954
rect 36252 -2056 36286 -2022
rect 36252 -2124 36286 -2090
rect 36252 -2192 36286 -2158
rect 36252 -2260 36286 -2226
rect 36252 -2328 36286 -2294
rect 36252 -2396 36286 -2362
rect 36252 -2464 36286 -2430
rect 36402 -1580 36436 -1546
rect 36402 -1648 36436 -1614
rect 36402 -1716 36436 -1682
rect 36402 -1784 36436 -1750
rect 36402 -1852 36436 -1818
rect 36402 -1920 36436 -1886
rect 36402 -1988 36436 -1954
rect 36402 -2056 36436 -2022
rect 36402 -2124 36436 -2090
rect 36402 -2192 36436 -2158
rect 36402 -2260 36436 -2226
rect 36402 -2328 36436 -2294
rect 36402 -2396 36436 -2362
rect 36402 -2464 36436 -2430
rect 36552 -1580 36586 -1546
rect 36552 -1648 36586 -1614
rect 36552 -1716 36586 -1682
rect 36552 -1784 36586 -1750
rect 36552 -1852 36586 -1818
rect 36552 -1920 36586 -1886
rect 36552 -1988 36586 -1954
rect 36552 -2056 36586 -2022
rect 36552 -2124 36586 -2090
rect 36552 -2192 36586 -2158
rect 36552 -2260 36586 -2226
rect 36552 -2328 36586 -2294
rect 36552 -2396 36586 -2362
rect 36552 -2464 36586 -2430
rect 36702 -1580 36736 -1546
rect 36702 -1648 36736 -1614
rect 36702 -1716 36736 -1682
rect 36702 -1784 36736 -1750
rect 36702 -1852 36736 -1818
rect 36702 -1920 36736 -1886
rect 36702 -1988 36736 -1954
rect 36702 -2056 36736 -2022
rect 36702 -2124 36736 -2090
rect 36702 -2192 36736 -2158
rect 36702 -2260 36736 -2226
rect 36702 -2328 36736 -2294
rect 36702 -2396 36736 -2362
rect 36702 -2464 36736 -2430
rect 36852 -1580 36886 -1546
rect 36852 -1648 36886 -1614
rect 36852 -1716 36886 -1682
rect 36852 -1784 36886 -1750
rect 36852 -1852 36886 -1818
rect 36852 -1920 36886 -1886
rect 36852 -1988 36886 -1954
rect 36852 -2056 36886 -2022
rect 36852 -2124 36886 -2090
rect 36852 -2192 36886 -2158
rect 36852 -2260 36886 -2226
rect 36852 -2328 36886 -2294
rect 36852 -2396 36886 -2362
rect 36852 -2464 36886 -2430
rect 37002 -1580 37036 -1546
rect 37002 -1648 37036 -1614
rect 37002 -1716 37036 -1682
rect 37002 -1784 37036 -1750
rect 37002 -1852 37036 -1818
rect 37002 -1920 37036 -1886
rect 37002 -1988 37036 -1954
rect 37002 -2056 37036 -2022
rect 37002 -2124 37036 -2090
rect 37002 -2192 37036 -2158
rect 37002 -2260 37036 -2226
rect 37002 -2328 37036 -2294
rect 37002 -2396 37036 -2362
rect 37002 -2464 37036 -2430
rect 37152 -1580 37186 -1546
rect 37152 -1648 37186 -1614
rect 37152 -1716 37186 -1682
rect 37152 -1784 37186 -1750
rect 37152 -1852 37186 -1818
rect 37152 -1920 37186 -1886
rect 37152 -1988 37186 -1954
rect 37152 -2056 37186 -2022
rect 37152 -2124 37186 -2090
rect 37152 -2192 37186 -2158
rect 37152 -2260 37186 -2226
rect 37152 -2328 37186 -2294
rect 37152 -2396 37186 -2362
rect 37152 -2464 37186 -2430
rect 37302 -1580 37336 -1546
rect 37302 -1648 37336 -1614
rect 37302 -1716 37336 -1682
rect 37302 -1784 37336 -1750
rect 37302 -1852 37336 -1818
rect 37302 -1920 37336 -1886
rect 37302 -1988 37336 -1954
rect 37302 -2056 37336 -2022
rect 37302 -2124 37336 -2090
rect 37302 -2192 37336 -2158
rect 37302 -2260 37336 -2226
rect 37302 -2328 37336 -2294
rect 37302 -2396 37336 -2362
rect 37302 -2464 37336 -2430
rect 37452 -1580 37486 -1546
rect 37452 -1648 37486 -1614
rect 37452 -1716 37486 -1682
rect 37452 -1784 37486 -1750
rect 37452 -1852 37486 -1818
rect 37452 -1920 37486 -1886
rect 37452 -1988 37486 -1954
rect 37452 -2056 37486 -2022
rect 37452 -2124 37486 -2090
rect 37452 -2192 37486 -2158
rect 37452 -2260 37486 -2226
rect 37452 -2328 37486 -2294
rect 37452 -2396 37486 -2362
rect 37452 -2464 37486 -2430
rect 37856 -1580 37890 -1546
rect 37856 -1648 37890 -1614
rect 37856 -1716 37890 -1682
rect 37856 -1784 37890 -1750
rect 37856 -1852 37890 -1818
rect 37856 -1920 37890 -1886
rect 37856 -1988 37890 -1954
rect 37856 -2056 37890 -2022
rect 37856 -2124 37890 -2090
rect 37856 -2192 37890 -2158
rect 37856 -2260 37890 -2226
rect 37856 -2328 37890 -2294
rect 37856 -2396 37890 -2362
rect 37856 -2464 37890 -2430
rect 38006 -1580 38040 -1546
rect 38006 -1648 38040 -1614
rect 38006 -1716 38040 -1682
rect 38006 -1784 38040 -1750
rect 38006 -1852 38040 -1818
rect 38006 -1920 38040 -1886
rect 38006 -1988 38040 -1954
rect 38006 -2056 38040 -2022
rect 38006 -2124 38040 -2090
rect 38006 -2192 38040 -2158
rect 38006 -2260 38040 -2226
rect 38006 -2328 38040 -2294
rect 38006 -2396 38040 -2362
rect 38006 -2464 38040 -2430
rect 38156 -1580 38190 -1546
rect 38156 -1648 38190 -1614
rect 38156 -1716 38190 -1682
rect 38156 -1784 38190 -1750
rect 38156 -1852 38190 -1818
rect 38156 -1920 38190 -1886
rect 38156 -1988 38190 -1954
rect 38156 -2056 38190 -2022
rect 38156 -2124 38190 -2090
rect 38156 -2192 38190 -2158
rect 38156 -2260 38190 -2226
rect 38156 -2328 38190 -2294
rect 38156 -2396 38190 -2362
rect 38156 -2464 38190 -2430
rect 38306 -1580 38340 -1546
rect 38306 -1648 38340 -1614
rect 38306 -1716 38340 -1682
rect 38306 -1784 38340 -1750
rect 38306 -1852 38340 -1818
rect 38306 -1920 38340 -1886
rect 38306 -1988 38340 -1954
rect 38306 -2056 38340 -2022
rect 38306 -2124 38340 -2090
rect 38306 -2192 38340 -2158
rect 38306 -2260 38340 -2226
rect 38306 -2328 38340 -2294
rect 38306 -2396 38340 -2362
rect 38306 -2464 38340 -2430
rect 38456 -1580 38490 -1546
rect 38456 -1648 38490 -1614
rect 38456 -1716 38490 -1682
rect 38456 -1784 38490 -1750
rect 38456 -1852 38490 -1818
rect 38456 -1920 38490 -1886
rect 38456 -1988 38490 -1954
rect 38456 -2056 38490 -2022
rect 38456 -2124 38490 -2090
rect 38456 -2192 38490 -2158
rect 38456 -2260 38490 -2226
rect 38456 -2328 38490 -2294
rect 38456 -2396 38490 -2362
rect 38456 -2464 38490 -2430
rect 38606 -1580 38640 -1546
rect 38606 -1648 38640 -1614
rect 38606 -1716 38640 -1682
rect 38606 -1784 38640 -1750
rect 38606 -1852 38640 -1818
rect 38606 -1920 38640 -1886
rect 38606 -1988 38640 -1954
rect 38606 -2056 38640 -2022
rect 38606 -2124 38640 -2090
rect 38606 -2192 38640 -2158
rect 38606 -2260 38640 -2226
rect 38606 -2328 38640 -2294
rect 38606 -2396 38640 -2362
rect 38606 -2464 38640 -2430
rect 38756 -1580 38790 -1546
rect 38756 -1648 38790 -1614
rect 38756 -1716 38790 -1682
rect 38756 -1784 38790 -1750
rect 38756 -1852 38790 -1818
rect 38756 -1920 38790 -1886
rect 38756 -1988 38790 -1954
rect 38756 -2056 38790 -2022
rect 38756 -2124 38790 -2090
rect 38756 -2192 38790 -2158
rect 38756 -2260 38790 -2226
rect 38756 -2328 38790 -2294
rect 38756 -2396 38790 -2362
rect 38756 -2464 38790 -2430
rect 38906 -1580 38940 -1546
rect 38906 -1648 38940 -1614
rect 38906 -1716 38940 -1682
rect 38906 -1784 38940 -1750
rect 38906 -1852 38940 -1818
rect 38906 -1920 38940 -1886
rect 38906 -1988 38940 -1954
rect 38906 -2056 38940 -2022
rect 38906 -2124 38940 -2090
rect 38906 -2192 38940 -2158
rect 38906 -2260 38940 -2226
rect 38906 -2328 38940 -2294
rect 38906 -2396 38940 -2362
rect 38906 -2464 38940 -2430
rect 39056 -1580 39090 -1546
rect 39056 -1648 39090 -1614
rect 39056 -1716 39090 -1682
rect 39056 -1784 39090 -1750
rect 39056 -1852 39090 -1818
rect 39056 -1920 39090 -1886
rect 39056 -1988 39090 -1954
rect 39056 -2056 39090 -2022
rect 39056 -2124 39090 -2090
rect 39056 -2192 39090 -2158
rect 39056 -2260 39090 -2226
rect 39056 -2328 39090 -2294
rect 39056 -2396 39090 -2362
rect 39056 -2464 39090 -2430
rect 39206 -1580 39240 -1546
rect 39206 -1648 39240 -1614
rect 39206 -1716 39240 -1682
rect 39206 -1784 39240 -1750
rect 39206 -1852 39240 -1818
rect 39206 -1920 39240 -1886
rect 39206 -1988 39240 -1954
rect 39206 -2056 39240 -2022
rect 39206 -2124 39240 -2090
rect 39206 -2192 39240 -2158
rect 39206 -2260 39240 -2226
rect 39206 -2328 39240 -2294
rect 39206 -2396 39240 -2362
rect 39206 -2464 39240 -2430
rect 39356 -1580 39390 -1546
rect 39356 -1648 39390 -1614
rect 39356 -1716 39390 -1682
rect 39356 -1784 39390 -1750
rect 39356 -1852 39390 -1818
rect 39356 -1920 39390 -1886
rect 39356 -1988 39390 -1954
rect 39356 -2056 39390 -2022
rect 39356 -2124 39390 -2090
rect 39356 -2192 39390 -2158
rect 39356 -2260 39390 -2226
rect 39356 -2328 39390 -2294
rect 39356 -2396 39390 -2362
rect 39356 -2464 39390 -2430
<< psubdiff >>
rect 35729 -1546 35849 -1518
rect 35729 -1580 35772 -1546
rect 35806 -1580 35849 -1546
rect 35729 -1614 35849 -1580
rect 35729 -1648 35772 -1614
rect 35806 -1648 35849 -1614
rect 35729 -1682 35849 -1648
rect 35729 -1716 35772 -1682
rect 35806 -1716 35849 -1682
rect 35729 -1750 35849 -1716
rect 35729 -1784 35772 -1750
rect 35806 -1784 35849 -1750
rect 35729 -1818 35849 -1784
rect 35729 -1852 35772 -1818
rect 35806 -1852 35849 -1818
rect 35729 -1886 35849 -1852
rect 35729 -1920 35772 -1886
rect 35806 -1920 35849 -1886
rect 35729 -1954 35849 -1920
rect 35729 -1988 35772 -1954
rect 35806 -1988 35849 -1954
rect 35729 -2022 35849 -1988
rect 35729 -2056 35772 -2022
rect 35806 -2056 35849 -2022
rect 35729 -2090 35849 -2056
rect 35729 -2124 35772 -2090
rect 35806 -2124 35849 -2090
rect 35729 -2158 35849 -2124
rect 35729 -2192 35772 -2158
rect 35806 -2192 35849 -2158
rect 35729 -2226 35849 -2192
rect 35729 -2260 35772 -2226
rect 35806 -2260 35849 -2226
rect 35729 -2294 35849 -2260
rect 35729 -2328 35772 -2294
rect 35806 -2328 35849 -2294
rect 35729 -2362 35849 -2328
rect 35729 -2396 35772 -2362
rect 35806 -2396 35849 -2362
rect 35729 -2430 35849 -2396
rect 35729 -2464 35772 -2430
rect 35806 -2464 35849 -2430
rect 35729 -2510 35849 -2464
rect 37633 -1546 37753 -1518
rect 37633 -1580 37676 -1546
rect 37710 -1580 37753 -1546
rect 37633 -1614 37753 -1580
rect 37633 -1648 37676 -1614
rect 37710 -1648 37753 -1614
rect 37633 -1682 37753 -1648
rect 37633 -1716 37676 -1682
rect 37710 -1716 37753 -1682
rect 37633 -1750 37753 -1716
rect 37633 -1784 37676 -1750
rect 37710 -1784 37753 -1750
rect 37633 -1818 37753 -1784
rect 37633 -1852 37676 -1818
rect 37710 -1852 37753 -1818
rect 37633 -1886 37753 -1852
rect 37633 -1920 37676 -1886
rect 37710 -1920 37753 -1886
rect 37633 -1954 37753 -1920
rect 37633 -1988 37676 -1954
rect 37710 -1988 37753 -1954
rect 37633 -2022 37753 -1988
rect 37633 -2056 37676 -2022
rect 37710 -2056 37753 -2022
rect 37633 -2090 37753 -2056
rect 37633 -2124 37676 -2090
rect 37710 -2124 37753 -2090
rect 37633 -2158 37753 -2124
rect 37633 -2192 37676 -2158
rect 37710 -2192 37753 -2158
rect 37633 -2226 37753 -2192
rect 37633 -2260 37676 -2226
rect 37710 -2260 37753 -2226
rect 37633 -2294 37753 -2260
rect 37633 -2328 37676 -2294
rect 37710 -2328 37753 -2294
rect 37633 -2362 37753 -2328
rect 37633 -2396 37676 -2362
rect 37710 -2396 37753 -2362
rect 37633 -2430 37753 -2396
rect 37633 -2464 37676 -2430
rect 37710 -2464 37753 -2430
rect 37633 -2510 37753 -2464
<< psubdiffcont >>
rect 35772 -1580 35806 -1546
rect 35772 -1648 35806 -1614
rect 35772 -1716 35806 -1682
rect 35772 -1784 35806 -1750
rect 35772 -1852 35806 -1818
rect 35772 -1920 35806 -1886
rect 35772 -1988 35806 -1954
rect 35772 -2056 35806 -2022
rect 35772 -2124 35806 -2090
rect 35772 -2192 35806 -2158
rect 35772 -2260 35806 -2226
rect 35772 -2328 35806 -2294
rect 35772 -2396 35806 -2362
rect 35772 -2464 35806 -2430
rect 37676 -1580 37710 -1546
rect 37676 -1648 37710 -1614
rect 37676 -1716 37710 -1682
rect 37676 -1784 37710 -1750
rect 37676 -1852 37710 -1818
rect 37676 -1920 37710 -1886
rect 37676 -1988 37710 -1954
rect 37676 -2056 37710 -2022
rect 37676 -2124 37710 -2090
rect 37676 -2192 37710 -2158
rect 37676 -2260 37710 -2226
rect 37676 -2328 37710 -2294
rect 37676 -2396 37710 -2362
rect 37676 -2464 37710 -2430
<< poly >>
rect 35541 -1436 35621 -1413
rect 35541 -1470 35564 -1436
rect 35598 -1438 35621 -1436
rect 35598 -1468 37409 -1438
rect 35598 -1470 35621 -1468
rect 35541 -1493 35621 -1470
rect 36029 -1518 36059 -1468
rect 36179 -1518 36209 -1468
rect 36329 -1518 36359 -1468
rect 36479 -1518 36509 -1468
rect 36629 -1518 36659 -1468
rect 36779 -1518 36809 -1468
rect 36929 -1518 36959 -1468
rect 37079 -1518 37109 -1468
rect 37229 -1518 37259 -1468
rect 37379 -1518 37409 -1468
rect 37933 -1510 37963 -1482
rect 38083 -1510 38113 -1482
rect 38233 -1510 38263 -1482
rect 38383 -1510 38413 -1482
rect 38533 -1510 38563 -1482
rect 38683 -1510 38713 -1482
rect 38833 -1510 38863 -1482
rect 38983 -1510 39013 -1483
rect 39133 -1510 39163 -1483
rect 39283 -1510 39313 -1483
rect 44121 -1849 44441 -1833
rect 44121 -1883 44162 -1849
rect 44196 -1883 44230 -1849
rect 44264 -1883 44298 -1849
rect 44332 -1883 44366 -1849
rect 44400 -1883 44441 -1849
rect 44121 -1906 44441 -1883
rect 44121 -2261 44441 -2238
rect 44121 -2295 44162 -2261
rect 44196 -2295 44230 -2261
rect 44264 -2295 44298 -2261
rect 44332 -2295 44366 -2261
rect 44400 -2295 44441 -2261
rect 44121 -2311 44441 -2295
rect 36029 -2544 36059 -2518
rect 36179 -2544 36209 -2518
rect 36329 -2544 36359 -2518
rect 36479 -2544 36509 -2518
rect 36629 -2545 36659 -2518
rect 36779 -2545 36809 -2518
rect 36929 -2545 36959 -2518
rect 37079 -2544 37109 -2518
rect 37229 -2545 37259 -2518
rect 37379 -2562 37409 -2518
rect 37933 -2560 37963 -2510
rect 38083 -2560 38113 -2510
rect 38233 -2560 38263 -2510
rect 38383 -2560 38413 -2510
rect 38533 -2560 38563 -2510
rect 38683 -2560 38713 -2510
rect 38833 -2560 38863 -2510
rect 38983 -2560 39013 -2510
rect 39133 -2560 39163 -2510
rect 39283 -2560 39313 -2510
rect 37933 -2562 39313 -2560
rect 37379 -2592 39313 -2562
<< polycont >>
rect 35564 -1470 35598 -1436
rect 44162 -1883 44196 -1849
rect 44230 -1883 44264 -1849
rect 44298 -1883 44332 -1849
rect 44366 -1883 44400 -1849
rect 44162 -2295 44196 -2261
rect 44230 -2295 44264 -2261
rect 44298 -2295 44332 -2261
rect 44366 -2295 44400 -2261
<< npolyres >>
rect 44121 -2238 44441 -1906
<< locali >>
rect 39432 9738 39512 9761
rect 39432 9704 39455 9738
rect 39489 9704 39512 9738
rect 39432 9681 39512 9704
rect 39552 9738 39632 9761
rect 39552 9704 39575 9738
rect 39609 9704 39632 9738
rect 39552 9681 39632 9704
rect 39432 9618 39512 9641
rect 39432 9584 39455 9618
rect 39489 9584 39512 9618
rect 39432 9561 39512 9584
rect 39552 9618 39632 9641
rect 39552 9584 39575 9618
rect 39609 9584 39632 9618
rect 39552 9561 39632 9584
rect 27940 2674 43396 2696
rect 27940 2640 27949 2674
rect 27983 2640 28029 2674
rect 28063 2640 28109 2674
rect 28143 2640 28189 2674
rect 28223 2640 28269 2674
rect 28303 2640 28349 2674
rect 28383 2640 28429 2674
rect 28463 2640 28509 2674
rect 28543 2640 28589 2674
rect 28623 2640 28669 2674
rect 28703 2640 28749 2674
rect 28783 2640 28829 2674
rect 28863 2640 28909 2674
rect 28943 2640 28989 2674
rect 29023 2640 29069 2674
rect 29103 2640 29149 2674
rect 29183 2640 29229 2674
rect 29263 2640 29309 2674
rect 29343 2640 29389 2674
rect 29423 2640 29469 2674
rect 29503 2640 29549 2674
rect 29583 2640 29629 2674
rect 29663 2640 29709 2674
rect 29743 2640 29789 2674
rect 29823 2640 29869 2674
rect 29903 2640 29949 2674
rect 29983 2640 30029 2674
rect 30063 2640 30109 2674
rect 30143 2640 30189 2674
rect 30223 2640 30269 2674
rect 30303 2640 30349 2674
rect 30383 2640 30429 2674
rect 30463 2640 30509 2674
rect 30543 2640 30589 2674
rect 30623 2640 30669 2674
rect 30703 2640 30749 2674
rect 30783 2640 30829 2674
rect 30863 2640 30910 2674
rect 30944 2640 30990 2674
rect 31024 2640 31070 2674
rect 31104 2640 31150 2674
rect 31184 2640 31230 2674
rect 31264 2640 31310 2674
rect 31344 2640 31390 2674
rect 31424 2640 31470 2674
rect 31504 2640 31550 2674
rect 31584 2640 31630 2674
rect 31664 2640 31710 2674
rect 31744 2640 31790 2674
rect 31824 2640 31870 2674
rect 31904 2640 31950 2674
rect 31984 2640 32030 2674
rect 32064 2640 32110 2674
rect 32144 2640 32190 2674
rect 32224 2640 32270 2674
rect 32304 2640 32350 2674
rect 32384 2640 32430 2674
rect 32464 2640 32510 2674
rect 32544 2640 32590 2674
rect 32624 2640 32670 2674
rect 32704 2640 32750 2674
rect 32784 2640 32830 2674
rect 32864 2640 32910 2674
rect 32944 2640 32990 2674
rect 33024 2640 33070 2674
rect 33104 2640 33150 2674
rect 33184 2640 33230 2674
rect 33264 2640 33310 2674
rect 33344 2640 33390 2674
rect 33424 2640 33470 2674
rect 33504 2640 33550 2674
rect 33584 2640 33630 2674
rect 33664 2640 33710 2674
rect 33744 2640 33790 2674
rect 33824 2640 33870 2674
rect 33904 2640 33950 2674
rect 33984 2640 34030 2674
rect 34064 2640 34110 2674
rect 34144 2640 34190 2674
rect 34224 2640 34270 2674
rect 34304 2640 34350 2674
rect 34384 2640 34430 2674
rect 34464 2640 34510 2674
rect 34544 2640 34590 2674
rect 34624 2640 34670 2674
rect 34704 2640 34750 2674
rect 34784 2640 34830 2674
rect 34864 2640 34910 2674
rect 34944 2640 34990 2674
rect 35024 2640 35070 2674
rect 35104 2640 35150 2674
rect 35184 2640 35242 2674
rect 35276 2640 35322 2674
rect 35356 2640 35402 2674
rect 35436 2640 35482 2674
rect 35516 2640 35562 2674
rect 35596 2640 35642 2674
rect 35676 2640 35722 2674
rect 35756 2640 35802 2674
rect 35836 2640 35882 2674
rect 35916 2640 35962 2674
rect 35996 2640 36042 2674
rect 36076 2640 36122 2674
rect 36156 2640 36202 2674
rect 36236 2640 36282 2674
rect 36316 2640 36362 2674
rect 36396 2640 36442 2674
rect 36476 2640 36522 2674
rect 36556 2640 36602 2674
rect 36636 2640 36682 2674
rect 36716 2640 36762 2674
rect 36796 2640 36842 2674
rect 36876 2640 36922 2674
rect 36956 2640 37002 2674
rect 37036 2640 37082 2674
rect 37116 2640 37162 2674
rect 37196 2640 37242 2674
rect 37276 2640 37322 2674
rect 37356 2640 37402 2674
rect 37436 2640 37482 2674
rect 37516 2640 37562 2674
rect 37596 2640 37642 2674
rect 37676 2640 37722 2674
rect 37756 2640 37802 2674
rect 37836 2640 37882 2674
rect 37916 2640 37962 2674
rect 37996 2640 38042 2674
rect 38076 2640 38122 2674
rect 38156 2640 38202 2674
rect 38236 2640 38282 2674
rect 38316 2640 38362 2674
rect 38396 2640 38442 2674
rect 38476 2640 38522 2674
rect 38556 2640 38602 2674
rect 38636 2640 38682 2674
rect 38716 2640 38762 2674
rect 38796 2640 38842 2674
rect 38876 2640 38922 2674
rect 38956 2640 39002 2674
rect 39036 2640 39083 2674
rect 39117 2640 39163 2674
rect 39197 2640 39243 2674
rect 39277 2640 39323 2674
rect 39357 2640 39403 2674
rect 39437 2640 39483 2674
rect 39517 2640 39563 2674
rect 39597 2640 39643 2674
rect 39677 2640 39723 2674
rect 39757 2640 39803 2674
rect 39837 2640 39883 2674
rect 39917 2640 39963 2674
rect 39997 2640 40043 2674
rect 40077 2640 40123 2674
rect 40157 2640 40203 2674
rect 40237 2640 40283 2674
rect 40317 2640 40363 2674
rect 40397 2640 40443 2674
rect 40477 2640 40523 2674
rect 40557 2640 40603 2674
rect 40637 2640 40683 2674
rect 40717 2640 40763 2674
rect 40797 2640 40843 2674
rect 40877 2640 40923 2674
rect 40957 2640 41003 2674
rect 41037 2640 41083 2674
rect 41117 2640 41163 2674
rect 41197 2640 41243 2674
rect 41277 2640 41323 2674
rect 41357 2640 41403 2674
rect 41437 2640 41483 2674
rect 41517 2640 41563 2674
rect 41597 2640 41643 2674
rect 41677 2640 41723 2674
rect 41757 2640 41803 2674
rect 41837 2640 41883 2674
rect 41917 2640 41963 2674
rect 41997 2640 42043 2674
rect 42077 2640 42123 2674
rect 42157 2640 42203 2674
rect 42237 2640 42283 2674
rect 42317 2640 42363 2674
rect 42397 2640 42443 2674
rect 42477 2640 42523 2674
rect 42557 2640 42603 2674
rect 42637 2640 42683 2674
rect 42717 2640 42763 2674
rect 42797 2640 42843 2674
rect 42877 2640 42923 2674
rect 42957 2640 43003 2674
rect 43037 2640 43083 2674
rect 43117 2640 43163 2674
rect 43197 2640 43243 2674
rect 43277 2640 43323 2674
rect 43357 2640 43396 2674
rect 27940 2584 43396 2640
rect 27940 2550 27949 2584
rect 27983 2550 28029 2584
rect 28063 2550 28109 2584
rect 28143 2550 28189 2584
rect 28223 2550 28269 2584
rect 28303 2550 28349 2584
rect 28383 2550 28429 2584
rect 28463 2550 28509 2584
rect 28543 2550 28589 2584
rect 28623 2550 28669 2584
rect 28703 2550 28749 2584
rect 28783 2550 28829 2584
rect 28863 2550 28909 2584
rect 28943 2550 28989 2584
rect 29023 2550 29069 2584
rect 29103 2550 29149 2584
rect 29183 2550 29229 2584
rect 29263 2550 29309 2584
rect 29343 2550 29389 2584
rect 29423 2550 29469 2584
rect 29503 2550 29549 2584
rect 29583 2550 29629 2584
rect 29663 2550 29709 2584
rect 29743 2550 29789 2584
rect 29823 2550 29869 2584
rect 29903 2550 29949 2584
rect 29983 2550 30029 2584
rect 30063 2550 30109 2584
rect 30143 2550 30189 2584
rect 30223 2550 30269 2584
rect 30303 2550 30349 2584
rect 30383 2550 30429 2584
rect 30463 2550 30509 2584
rect 30543 2550 30589 2584
rect 30623 2550 30669 2584
rect 30703 2550 30749 2584
rect 30783 2550 30829 2584
rect 30863 2550 30910 2584
rect 30944 2550 30990 2584
rect 31024 2550 31070 2584
rect 31104 2550 31150 2584
rect 31184 2550 31230 2584
rect 31264 2550 31310 2584
rect 31344 2550 31390 2584
rect 31424 2550 31470 2584
rect 31504 2550 31550 2584
rect 31584 2550 31630 2584
rect 31664 2550 31710 2584
rect 31744 2550 31790 2584
rect 31824 2550 31870 2584
rect 31904 2550 31950 2584
rect 31984 2550 32030 2584
rect 32064 2550 32110 2584
rect 32144 2550 32190 2584
rect 32224 2550 32270 2584
rect 32304 2550 32350 2584
rect 32384 2550 32430 2584
rect 32464 2550 32510 2584
rect 32544 2550 32590 2584
rect 32624 2550 32670 2584
rect 32704 2550 32750 2584
rect 32784 2550 32830 2584
rect 32864 2550 32910 2584
rect 32944 2550 32990 2584
rect 33024 2550 33070 2584
rect 33104 2550 33150 2584
rect 33184 2550 33230 2584
rect 33264 2550 33310 2584
rect 33344 2550 33390 2584
rect 33424 2550 33470 2584
rect 33504 2550 33550 2584
rect 33584 2550 33630 2584
rect 33664 2550 33710 2584
rect 33744 2550 33790 2584
rect 33824 2550 33870 2584
rect 33904 2550 33950 2584
rect 33984 2550 34030 2584
rect 34064 2550 34110 2584
rect 34144 2550 34190 2584
rect 34224 2550 34270 2584
rect 34304 2550 34350 2584
rect 34384 2550 34430 2584
rect 34464 2550 34510 2584
rect 34544 2550 34590 2584
rect 34624 2550 34670 2584
rect 34704 2550 34750 2584
rect 34784 2550 34830 2584
rect 34864 2550 34910 2584
rect 34944 2550 34990 2584
rect 35024 2550 35070 2584
rect 35104 2550 35150 2584
rect 35184 2550 35242 2584
rect 35276 2550 35322 2584
rect 35356 2550 35402 2584
rect 35436 2550 35482 2584
rect 35516 2550 35562 2584
rect 35596 2550 35642 2584
rect 35676 2550 35722 2584
rect 35756 2550 35802 2584
rect 35836 2550 35882 2584
rect 35916 2550 35962 2584
rect 35996 2550 36042 2584
rect 36076 2550 36122 2584
rect 36156 2550 36202 2584
rect 36236 2550 36282 2584
rect 36316 2550 36362 2584
rect 36396 2550 36442 2584
rect 36476 2550 36522 2584
rect 36556 2550 36602 2584
rect 36636 2550 36682 2584
rect 36716 2550 36762 2584
rect 36796 2550 36842 2584
rect 36876 2550 36922 2584
rect 36956 2550 37002 2584
rect 37036 2550 37082 2584
rect 37116 2550 37162 2584
rect 37196 2550 37242 2584
rect 37276 2550 37322 2584
rect 37356 2550 37402 2584
rect 37436 2550 37482 2584
rect 37516 2550 37562 2584
rect 37596 2550 37642 2584
rect 37676 2550 37722 2584
rect 37756 2550 37802 2584
rect 37836 2550 37882 2584
rect 37916 2550 37962 2584
rect 37996 2550 38042 2584
rect 38076 2550 38122 2584
rect 38156 2550 38202 2584
rect 38236 2550 38282 2584
rect 38316 2550 38362 2584
rect 38396 2550 38442 2584
rect 38476 2550 38522 2584
rect 38556 2550 38602 2584
rect 38636 2550 38682 2584
rect 38716 2550 38762 2584
rect 38796 2550 38842 2584
rect 38876 2550 38922 2584
rect 38956 2550 39002 2584
rect 39036 2550 39083 2584
rect 39117 2550 39163 2584
rect 39197 2550 39243 2584
rect 39277 2550 39323 2584
rect 39357 2550 39403 2584
rect 39437 2550 39483 2584
rect 39517 2550 39563 2584
rect 39597 2550 39643 2584
rect 39677 2550 39723 2584
rect 39757 2550 39803 2584
rect 39837 2550 39883 2584
rect 39917 2550 39963 2584
rect 39997 2550 40043 2584
rect 40077 2550 40123 2584
rect 40157 2550 40203 2584
rect 40237 2550 40283 2584
rect 40317 2550 40363 2584
rect 40397 2550 40443 2584
rect 40477 2550 40523 2584
rect 40557 2550 40603 2584
rect 40637 2550 40683 2584
rect 40717 2550 40763 2584
rect 40797 2550 40843 2584
rect 40877 2550 40923 2584
rect 40957 2550 41003 2584
rect 41037 2550 41083 2584
rect 41117 2550 41163 2584
rect 41197 2550 41243 2584
rect 41277 2550 41323 2584
rect 41357 2550 41403 2584
rect 41437 2550 41483 2584
rect 41517 2550 41563 2584
rect 41597 2550 41643 2584
rect 41677 2550 41723 2584
rect 41757 2550 41803 2584
rect 41837 2550 41883 2584
rect 41917 2550 41963 2584
rect 41997 2550 42043 2584
rect 42077 2550 42123 2584
rect 42157 2550 42203 2584
rect 42237 2550 42283 2584
rect 42317 2550 42363 2584
rect 42397 2550 42443 2584
rect 42477 2550 42523 2584
rect 42557 2550 42603 2584
rect 42637 2550 42683 2584
rect 42717 2550 42763 2584
rect 42797 2550 42843 2584
rect 42877 2550 42923 2584
rect 42957 2550 43003 2584
rect 43037 2550 43083 2584
rect 43117 2550 43163 2584
rect 43197 2550 43243 2584
rect 43277 2550 43323 2584
rect 43357 2550 43396 2584
rect 27940 2526 43396 2550
rect 32663 1600 33063 2526
rect 32523 1598 33201 1600
rect 32522 1560 33202 1598
rect 32522 1500 32560 1560
rect 32620 1500 32680 1560
rect 32740 1500 32980 1560
rect 33040 1550 33202 1560
rect 33040 1510 33110 1550
rect 33150 1510 33202 1550
rect 33040 1500 33202 1510
rect 32522 1440 33202 1500
rect 32522 1380 32560 1440
rect 32620 1380 32680 1440
rect 32740 1380 32980 1440
rect 33040 1380 33100 1440
rect 33160 1380 33202 1440
rect 32522 1338 33202 1380
rect 34256 1545 34516 1598
rect 34256 1511 34309 1545
rect 34343 1511 34429 1545
rect 34463 1511 34516 1545
rect 34256 1425 34516 1511
rect 34256 1391 34309 1425
rect 34343 1391 34429 1425
rect 34463 1391 34516 1425
rect 34256 1338 34516 1391
rect 34676 1545 34936 1598
rect 34676 1511 34729 1545
rect 34763 1511 34849 1545
rect 34883 1511 34936 1545
rect 34676 1425 34936 1511
rect 34676 1391 34729 1425
rect 34763 1391 34849 1425
rect 34883 1391 34936 1425
rect 34676 1338 34936 1391
rect 32523 1178 33201 1338
rect 32522 1140 33202 1178
rect 32522 1080 32560 1140
rect 32620 1125 32980 1140
rect 32620 1091 32695 1125
rect 32729 1091 32980 1125
rect 32620 1080 32980 1091
rect 33040 1080 33100 1140
rect 33160 1080 33202 1140
rect 32522 1020 33202 1080
rect 32522 960 32560 1020
rect 32620 960 32680 1020
rect 32740 960 32980 1020
rect 33040 960 33100 1020
rect 33160 960 33202 1020
rect 32522 919 33202 960
rect 32522 918 32782 919
rect 32942 918 33202 919
rect 34256 1125 34516 1178
rect 34256 1091 34309 1125
rect 34343 1091 34429 1125
rect 34463 1091 34516 1125
rect 34256 1005 34516 1091
rect 34256 971 34309 1005
rect 34343 971 34429 1005
rect 34463 971 34516 1005
rect 34256 918 34516 971
rect 34676 1125 34936 1178
rect 34676 1091 34729 1125
rect 34763 1091 34849 1125
rect 34883 1091 34936 1125
rect 34676 1005 34936 1091
rect 34676 971 34729 1005
rect 34763 971 34849 1005
rect 34883 971 34936 1005
rect 34676 918 34936 971
rect 44202 -28 44282 -27
rect 44322 -28 44402 -27
rect 44202 -32 44403 -28
rect 44202 -84 44218 -32
rect 44270 -84 44338 -32
rect 44390 -84 44403 -32
rect 44202 -85 44226 -84
rect 44260 -85 44346 -84
rect 44380 -85 44403 -84
rect 44202 -94 44403 -85
rect 44202 -107 44433 -94
rect 44203 -147 44433 -107
rect 44202 -152 44433 -147
rect 44202 -204 44218 -152
rect 44270 -204 44338 -152
rect 44390 -174 44433 -152
rect 44390 -204 44403 -174
rect 44202 -205 44226 -204
rect 44260 -205 44346 -204
rect 44380 -205 44403 -204
rect 44202 -227 44403 -205
rect 44203 -228 44403 -227
rect 35795 -487 35995 -464
rect 35795 -521 35818 -487
rect 35852 -521 35938 -487
rect 35972 -521 35995 -487
rect 35795 -530 35995 -521
rect 35795 -607 36445 -530
rect 35795 -641 35818 -607
rect 35852 -641 35938 -607
rect 35972 -610 36445 -607
rect 35972 -641 35995 -610
rect 35795 -664 35995 -641
rect 36365 -1109 36445 -610
rect 36365 -1154 36833 -1109
rect 36365 -1189 36834 -1154
rect 36634 -1405 36834 -1189
rect 35541 -1436 35621 -1413
rect 35541 -1470 35564 -1436
rect 35598 -1470 35621 -1436
rect 35541 -1493 35621 -1470
rect 36079 -1485 39460 -1405
rect 35749 -1546 36009 -1540
rect 35749 -1580 35772 -1546
rect 35806 -1580 35952 -1546
rect 35986 -1580 36009 -1546
rect 35749 -1614 36009 -1580
rect 35749 -1648 35772 -1614
rect 35806 -1648 35952 -1614
rect 35986 -1648 36009 -1614
rect 35749 -1682 36009 -1648
rect 35749 -1716 35772 -1682
rect 35806 -1716 35952 -1682
rect 35986 -1716 36009 -1682
rect 35749 -1750 36009 -1716
rect 35749 -1784 35772 -1750
rect 35806 -1784 35952 -1750
rect 35986 -1784 36009 -1750
rect 35749 -1818 36009 -1784
rect 35749 -1852 35772 -1818
rect 35806 -1852 35952 -1818
rect 35986 -1852 36009 -1818
rect 35749 -1886 36009 -1852
rect 35749 -1920 35772 -1886
rect 35806 -1920 35952 -1886
rect 35986 -1920 36009 -1886
rect 35749 -1954 36009 -1920
rect 35749 -1988 35772 -1954
rect 35806 -1988 35952 -1954
rect 35986 -1988 36009 -1954
rect 35749 -2022 36009 -1988
rect 35749 -2056 35772 -2022
rect 35806 -2056 35952 -2022
rect 35986 -2056 36009 -2022
rect 35749 -2090 36009 -2056
rect 35749 -2124 35772 -2090
rect 35806 -2124 35952 -2090
rect 35986 -2124 36009 -2090
rect 35749 -2158 36009 -2124
rect 35749 -2192 35772 -2158
rect 35806 -2192 35952 -2158
rect 35986 -2192 36009 -2158
rect 35749 -2226 36009 -2192
rect 35749 -2260 35772 -2226
rect 35806 -2260 35952 -2226
rect 35986 -2260 36009 -2226
rect 35749 -2294 36009 -2260
rect 35749 -2328 35772 -2294
rect 35806 -2328 35952 -2294
rect 35986 -2328 36009 -2294
rect 35749 -2362 36009 -2328
rect 35749 -2396 35772 -2362
rect 35806 -2396 35952 -2362
rect 35986 -2396 36009 -2362
rect 35749 -2430 36009 -2396
rect 35749 -2464 35772 -2430
rect 35806 -2464 35952 -2430
rect 35986 -2464 36009 -2430
rect 35749 -2490 36009 -2464
rect 36079 -1546 36159 -1485
rect 36079 -1580 36102 -1546
rect 36136 -1580 36159 -1546
rect 36079 -1614 36159 -1580
rect 36079 -1648 36102 -1614
rect 36136 -1648 36159 -1614
rect 36079 -1682 36159 -1648
rect 36079 -1716 36102 -1682
rect 36136 -1716 36159 -1682
rect 36079 -1750 36159 -1716
rect 36079 -1784 36102 -1750
rect 36136 -1784 36159 -1750
rect 36079 -1818 36159 -1784
rect 36079 -1852 36102 -1818
rect 36136 -1852 36159 -1818
rect 36079 -1886 36159 -1852
rect 36079 -1920 36102 -1886
rect 36136 -1920 36159 -1886
rect 36079 -1954 36159 -1920
rect 36079 -1988 36102 -1954
rect 36136 -1988 36159 -1954
rect 36079 -2022 36159 -1988
rect 36079 -2056 36102 -2022
rect 36136 -2056 36159 -2022
rect 36079 -2090 36159 -2056
rect 36079 -2124 36102 -2090
rect 36136 -2124 36159 -2090
rect 36079 -2158 36159 -2124
rect 36079 -2192 36102 -2158
rect 36136 -2192 36159 -2158
rect 36079 -2226 36159 -2192
rect 36079 -2260 36102 -2226
rect 36136 -2260 36159 -2226
rect 36079 -2294 36159 -2260
rect 36079 -2328 36102 -2294
rect 36136 -2328 36159 -2294
rect 36079 -2362 36159 -2328
rect 36079 -2396 36102 -2362
rect 36136 -2396 36159 -2362
rect 36079 -2430 36159 -2396
rect 36079 -2464 36102 -2430
rect 36136 -2464 36159 -2430
rect 36079 -2490 36159 -2464
rect 36229 -1546 36309 -1540
rect 36229 -1580 36252 -1546
rect 36286 -1580 36309 -1546
rect 36229 -1614 36309 -1580
rect 36229 -1648 36252 -1614
rect 36286 -1648 36309 -1614
rect 36229 -1682 36309 -1648
rect 36229 -1716 36252 -1682
rect 36286 -1716 36309 -1682
rect 36229 -1750 36309 -1716
rect 36229 -1784 36252 -1750
rect 36286 -1784 36309 -1750
rect 36229 -1818 36309 -1784
rect 36229 -1852 36252 -1818
rect 36286 -1852 36309 -1818
rect 36229 -1886 36309 -1852
rect 36229 -1920 36252 -1886
rect 36286 -1920 36309 -1886
rect 36229 -1954 36309 -1920
rect 36229 -1988 36252 -1954
rect 36286 -1988 36309 -1954
rect 36229 -2022 36309 -1988
rect 36229 -2056 36252 -2022
rect 36286 -2056 36309 -2022
rect 36229 -2090 36309 -2056
rect 36229 -2124 36252 -2090
rect 36286 -2124 36309 -2090
rect 36229 -2158 36309 -2124
rect 36229 -2192 36252 -2158
rect 36286 -2192 36309 -2158
rect 36229 -2226 36309 -2192
rect 36229 -2260 36252 -2226
rect 36286 -2260 36309 -2226
rect 36229 -2294 36309 -2260
rect 36229 -2328 36252 -2294
rect 36286 -2328 36309 -2294
rect 36229 -2362 36309 -2328
rect 36229 -2396 36252 -2362
rect 36286 -2396 36309 -2362
rect 36229 -2430 36309 -2396
rect 36229 -2464 36252 -2430
rect 36286 -2464 36309 -2430
rect 35929 -2545 36009 -2490
rect 36229 -2545 36309 -2464
rect 36379 -1546 36459 -1485
rect 36379 -1580 36402 -1546
rect 36436 -1580 36459 -1546
rect 36379 -1614 36459 -1580
rect 36379 -1648 36402 -1614
rect 36436 -1648 36459 -1614
rect 36379 -1682 36459 -1648
rect 36379 -1716 36402 -1682
rect 36436 -1716 36459 -1682
rect 36379 -1750 36459 -1716
rect 36379 -1784 36402 -1750
rect 36436 -1784 36459 -1750
rect 36379 -1818 36459 -1784
rect 36379 -1852 36402 -1818
rect 36436 -1852 36459 -1818
rect 36379 -1886 36459 -1852
rect 36379 -1920 36402 -1886
rect 36436 -1920 36459 -1886
rect 36379 -1954 36459 -1920
rect 36379 -1988 36402 -1954
rect 36436 -1988 36459 -1954
rect 36379 -2022 36459 -1988
rect 36379 -2056 36402 -2022
rect 36436 -2056 36459 -2022
rect 36379 -2090 36459 -2056
rect 36379 -2124 36402 -2090
rect 36436 -2124 36459 -2090
rect 36379 -2158 36459 -2124
rect 36379 -2192 36402 -2158
rect 36436 -2192 36459 -2158
rect 36379 -2226 36459 -2192
rect 36379 -2260 36402 -2226
rect 36436 -2260 36459 -2226
rect 36379 -2294 36459 -2260
rect 36379 -2328 36402 -2294
rect 36436 -2328 36459 -2294
rect 36379 -2362 36459 -2328
rect 36379 -2396 36402 -2362
rect 36436 -2396 36459 -2362
rect 36379 -2430 36459 -2396
rect 36379 -2464 36402 -2430
rect 36436 -2464 36459 -2430
rect 36379 -2490 36459 -2464
rect 36529 -1546 36609 -1540
rect 36529 -1580 36552 -1546
rect 36586 -1580 36609 -1546
rect 36529 -1614 36609 -1580
rect 36529 -1648 36552 -1614
rect 36586 -1648 36609 -1614
rect 36529 -1682 36609 -1648
rect 36529 -1716 36552 -1682
rect 36586 -1716 36609 -1682
rect 36529 -1750 36609 -1716
rect 36529 -1784 36552 -1750
rect 36586 -1784 36609 -1750
rect 36529 -1818 36609 -1784
rect 36529 -1852 36552 -1818
rect 36586 -1852 36609 -1818
rect 36529 -1886 36609 -1852
rect 36529 -1920 36552 -1886
rect 36586 -1920 36609 -1886
rect 36529 -1954 36609 -1920
rect 36529 -1988 36552 -1954
rect 36586 -1988 36609 -1954
rect 36529 -2022 36609 -1988
rect 36529 -2056 36552 -2022
rect 36586 -2056 36609 -2022
rect 36529 -2090 36609 -2056
rect 36529 -2124 36552 -2090
rect 36586 -2124 36609 -2090
rect 36529 -2158 36609 -2124
rect 36529 -2192 36552 -2158
rect 36586 -2192 36609 -2158
rect 36529 -2226 36609 -2192
rect 36529 -2260 36552 -2226
rect 36586 -2260 36609 -2226
rect 36529 -2294 36609 -2260
rect 36529 -2328 36552 -2294
rect 36586 -2328 36609 -2294
rect 36529 -2362 36609 -2328
rect 36529 -2396 36552 -2362
rect 36586 -2396 36609 -2362
rect 36529 -2430 36609 -2396
rect 36529 -2464 36552 -2430
rect 36586 -2464 36609 -2430
rect 36529 -2545 36609 -2464
rect 36679 -1546 36759 -1485
rect 36679 -1580 36702 -1546
rect 36736 -1580 36759 -1546
rect 36679 -1614 36759 -1580
rect 36679 -1648 36702 -1614
rect 36736 -1648 36759 -1614
rect 36679 -1682 36759 -1648
rect 36679 -1716 36702 -1682
rect 36736 -1716 36759 -1682
rect 36679 -1750 36759 -1716
rect 36679 -1784 36702 -1750
rect 36736 -1784 36759 -1750
rect 36679 -1818 36759 -1784
rect 36679 -1852 36702 -1818
rect 36736 -1852 36759 -1818
rect 36679 -1886 36759 -1852
rect 36679 -1920 36702 -1886
rect 36736 -1920 36759 -1886
rect 36679 -1954 36759 -1920
rect 36679 -1988 36702 -1954
rect 36736 -1988 36759 -1954
rect 36679 -2022 36759 -1988
rect 36679 -2056 36702 -2022
rect 36736 -2056 36759 -2022
rect 36679 -2090 36759 -2056
rect 36679 -2124 36702 -2090
rect 36736 -2124 36759 -2090
rect 36679 -2158 36759 -2124
rect 36679 -2192 36702 -2158
rect 36736 -2192 36759 -2158
rect 36679 -2226 36759 -2192
rect 36679 -2260 36702 -2226
rect 36736 -2260 36759 -2226
rect 36679 -2294 36759 -2260
rect 36679 -2328 36702 -2294
rect 36736 -2328 36759 -2294
rect 36679 -2362 36759 -2328
rect 36679 -2396 36702 -2362
rect 36736 -2396 36759 -2362
rect 36679 -2430 36759 -2396
rect 36679 -2464 36702 -2430
rect 36736 -2464 36759 -2430
rect 36679 -2490 36759 -2464
rect 36829 -1546 36909 -1540
rect 36829 -1580 36852 -1546
rect 36886 -1580 36909 -1546
rect 36829 -1614 36909 -1580
rect 36829 -1648 36852 -1614
rect 36886 -1648 36909 -1614
rect 36829 -1682 36909 -1648
rect 36829 -1716 36852 -1682
rect 36886 -1716 36909 -1682
rect 36829 -1750 36909 -1716
rect 36829 -1784 36852 -1750
rect 36886 -1784 36909 -1750
rect 36829 -1818 36909 -1784
rect 36829 -1852 36852 -1818
rect 36886 -1852 36909 -1818
rect 36829 -1886 36909 -1852
rect 36829 -1920 36852 -1886
rect 36886 -1920 36909 -1886
rect 36829 -1954 36909 -1920
rect 36829 -1988 36852 -1954
rect 36886 -1988 36909 -1954
rect 36829 -2022 36909 -1988
rect 36829 -2056 36852 -2022
rect 36886 -2056 36909 -2022
rect 36829 -2090 36909 -2056
rect 36829 -2124 36852 -2090
rect 36886 -2124 36909 -2090
rect 36829 -2158 36909 -2124
rect 36829 -2192 36852 -2158
rect 36886 -2192 36909 -2158
rect 36829 -2226 36909 -2192
rect 36829 -2260 36852 -2226
rect 36886 -2260 36909 -2226
rect 36829 -2294 36909 -2260
rect 36829 -2328 36852 -2294
rect 36886 -2328 36909 -2294
rect 36829 -2362 36909 -2328
rect 36829 -2396 36852 -2362
rect 36886 -2396 36909 -2362
rect 36829 -2430 36909 -2396
rect 36829 -2464 36852 -2430
rect 36886 -2464 36909 -2430
rect 36829 -2545 36909 -2464
rect 36979 -1546 37059 -1485
rect 36979 -1580 37002 -1546
rect 37036 -1580 37059 -1546
rect 36979 -1614 37059 -1580
rect 36979 -1648 37002 -1614
rect 37036 -1648 37059 -1614
rect 36979 -1682 37059 -1648
rect 36979 -1716 37002 -1682
rect 37036 -1716 37059 -1682
rect 36979 -1750 37059 -1716
rect 36979 -1784 37002 -1750
rect 37036 -1784 37059 -1750
rect 36979 -1818 37059 -1784
rect 36979 -1852 37002 -1818
rect 37036 -1852 37059 -1818
rect 36979 -1886 37059 -1852
rect 36979 -1920 37002 -1886
rect 37036 -1920 37059 -1886
rect 36979 -1954 37059 -1920
rect 36979 -1988 37002 -1954
rect 37036 -1988 37059 -1954
rect 36979 -2022 37059 -1988
rect 36979 -2056 37002 -2022
rect 37036 -2056 37059 -2022
rect 36979 -2090 37059 -2056
rect 36979 -2124 37002 -2090
rect 37036 -2124 37059 -2090
rect 36979 -2158 37059 -2124
rect 36979 -2192 37002 -2158
rect 37036 -2192 37059 -2158
rect 36979 -2226 37059 -2192
rect 36979 -2260 37002 -2226
rect 37036 -2260 37059 -2226
rect 36979 -2294 37059 -2260
rect 36979 -2328 37002 -2294
rect 37036 -2328 37059 -2294
rect 36979 -2362 37059 -2328
rect 36979 -2396 37002 -2362
rect 37036 -2396 37059 -2362
rect 36979 -2430 37059 -2396
rect 36979 -2464 37002 -2430
rect 37036 -2464 37059 -2430
rect 36979 -2490 37059 -2464
rect 37129 -1546 37209 -1540
rect 37129 -1580 37152 -1546
rect 37186 -1580 37209 -1546
rect 37129 -1614 37209 -1580
rect 37129 -1648 37152 -1614
rect 37186 -1648 37209 -1614
rect 37129 -1682 37209 -1648
rect 37129 -1716 37152 -1682
rect 37186 -1716 37209 -1682
rect 37129 -1750 37209 -1716
rect 37129 -1784 37152 -1750
rect 37186 -1784 37209 -1750
rect 37129 -1818 37209 -1784
rect 37129 -1852 37152 -1818
rect 37186 -1852 37209 -1818
rect 37129 -1886 37209 -1852
rect 37129 -1920 37152 -1886
rect 37186 -1920 37209 -1886
rect 37129 -1954 37209 -1920
rect 37129 -1988 37152 -1954
rect 37186 -1988 37209 -1954
rect 37129 -2022 37209 -1988
rect 37129 -2056 37152 -2022
rect 37186 -2056 37209 -2022
rect 37129 -2090 37209 -2056
rect 37129 -2124 37152 -2090
rect 37186 -2124 37209 -2090
rect 37129 -2158 37209 -2124
rect 37129 -2192 37152 -2158
rect 37186 -2192 37209 -2158
rect 37129 -2226 37209 -2192
rect 37129 -2260 37152 -2226
rect 37186 -2260 37209 -2226
rect 37129 -2294 37209 -2260
rect 37129 -2328 37152 -2294
rect 37186 -2328 37209 -2294
rect 37129 -2362 37209 -2328
rect 37129 -2396 37152 -2362
rect 37186 -2396 37209 -2362
rect 37129 -2430 37209 -2396
rect 37129 -2464 37152 -2430
rect 37186 -2464 37209 -2430
rect 37129 -2545 37209 -2464
rect 37279 -1546 37359 -1485
rect 37279 -1580 37302 -1546
rect 37336 -1580 37359 -1546
rect 37279 -1614 37359 -1580
rect 37279 -1648 37302 -1614
rect 37336 -1648 37359 -1614
rect 37279 -1682 37359 -1648
rect 37279 -1716 37302 -1682
rect 37336 -1716 37359 -1682
rect 37279 -1750 37359 -1716
rect 37279 -1784 37302 -1750
rect 37336 -1784 37359 -1750
rect 37279 -1818 37359 -1784
rect 37279 -1852 37302 -1818
rect 37336 -1852 37359 -1818
rect 37279 -1886 37359 -1852
rect 37279 -1920 37302 -1886
rect 37336 -1920 37359 -1886
rect 37279 -1954 37359 -1920
rect 37279 -1988 37302 -1954
rect 37336 -1988 37359 -1954
rect 37279 -2022 37359 -1988
rect 37279 -2056 37302 -2022
rect 37336 -2056 37359 -2022
rect 37279 -2090 37359 -2056
rect 37279 -2124 37302 -2090
rect 37336 -2124 37359 -2090
rect 37279 -2158 37359 -2124
rect 37279 -2192 37302 -2158
rect 37336 -2192 37359 -2158
rect 37279 -2226 37359 -2192
rect 37279 -2260 37302 -2226
rect 37336 -2260 37359 -2226
rect 37279 -2294 37359 -2260
rect 37279 -2328 37302 -2294
rect 37336 -2328 37359 -2294
rect 37279 -2362 37359 -2328
rect 37279 -2396 37302 -2362
rect 37336 -2396 37359 -2362
rect 37279 -2430 37359 -2396
rect 37279 -2464 37302 -2430
rect 37336 -2464 37359 -2430
rect 37279 -2490 37359 -2464
rect 37429 -1546 37509 -1540
rect 37429 -1580 37452 -1546
rect 37486 -1580 37509 -1546
rect 37429 -1614 37509 -1580
rect 37429 -1648 37452 -1614
rect 37486 -1648 37509 -1614
rect 37429 -1682 37509 -1648
rect 37429 -1716 37452 -1682
rect 37486 -1716 37509 -1682
rect 37429 -1750 37509 -1716
rect 37429 -1784 37452 -1750
rect 37486 -1784 37509 -1750
rect 37429 -1818 37509 -1784
rect 37429 -1852 37452 -1818
rect 37486 -1852 37509 -1818
rect 37429 -1886 37509 -1852
rect 37429 -1920 37452 -1886
rect 37486 -1920 37509 -1886
rect 37429 -1954 37509 -1920
rect 37429 -1988 37452 -1954
rect 37486 -1988 37509 -1954
rect 37429 -2022 37509 -1988
rect 37429 -2056 37452 -2022
rect 37486 -2056 37509 -2022
rect 37429 -2090 37509 -2056
rect 37429 -2124 37452 -2090
rect 37486 -2124 37509 -2090
rect 37429 -2158 37509 -2124
rect 37429 -2192 37452 -2158
rect 37486 -2192 37509 -2158
rect 37429 -2226 37509 -2192
rect 37429 -2260 37452 -2226
rect 37486 -2260 37509 -2226
rect 37429 -2294 37509 -2260
rect 37429 -2328 37452 -2294
rect 37486 -2328 37509 -2294
rect 37429 -2362 37509 -2328
rect 37429 -2396 37452 -2362
rect 37486 -2396 37509 -2362
rect 37429 -2430 37509 -2396
rect 37429 -2464 37452 -2430
rect 37486 -2464 37509 -2430
rect 37429 -2545 37509 -2464
rect 37653 -1542 37733 -1540
rect 37833 -1542 37913 -1540
rect 37653 -1546 37913 -1542
rect 37653 -1580 37676 -1546
rect 37710 -1580 37856 -1546
rect 37890 -1580 37913 -1546
rect 37653 -1614 37913 -1580
rect 37653 -1648 37676 -1614
rect 37710 -1648 37856 -1614
rect 37890 -1648 37913 -1614
rect 37653 -1682 37913 -1648
rect 37653 -1716 37676 -1682
rect 37710 -1716 37856 -1682
rect 37890 -1716 37913 -1682
rect 37653 -1750 37913 -1716
rect 37653 -1784 37676 -1750
rect 37710 -1784 37856 -1750
rect 37890 -1784 37913 -1750
rect 37653 -1818 37913 -1784
rect 37653 -1852 37676 -1818
rect 37710 -1852 37856 -1818
rect 37890 -1852 37913 -1818
rect 37653 -1886 37913 -1852
rect 37653 -1920 37676 -1886
rect 37710 -1920 37856 -1886
rect 37890 -1920 37913 -1886
rect 37653 -1954 37913 -1920
rect 37653 -1988 37676 -1954
rect 37710 -1988 37856 -1954
rect 37890 -1988 37913 -1954
rect 37653 -2022 37913 -1988
rect 37653 -2056 37676 -2022
rect 37710 -2056 37856 -2022
rect 37890 -2056 37913 -2022
rect 37653 -2090 37913 -2056
rect 37653 -2124 37676 -2090
rect 37710 -2124 37856 -2090
rect 37890 -2124 37913 -2090
rect 37653 -2158 37913 -2124
rect 37653 -2192 37676 -2158
rect 37710 -2192 37856 -2158
rect 37890 -2192 37913 -2158
rect 37653 -2226 37913 -2192
rect 37653 -2260 37676 -2226
rect 37710 -2260 37856 -2226
rect 37890 -2260 37913 -2226
rect 37653 -2294 37913 -2260
rect 37653 -2328 37676 -2294
rect 37710 -2328 37856 -2294
rect 37890 -2328 37913 -2294
rect 37653 -2362 37913 -2328
rect 37653 -2396 37676 -2362
rect 37710 -2396 37856 -2362
rect 37890 -2396 37913 -2362
rect 37653 -2430 37913 -2396
rect 37653 -2464 37676 -2430
rect 37710 -2464 37856 -2430
rect 37890 -2464 37913 -2430
rect 37653 -2490 37913 -2464
rect 37983 -1546 38063 -1485
rect 37983 -1580 38006 -1546
rect 38040 -1580 38063 -1546
rect 37983 -1614 38063 -1580
rect 37983 -1648 38006 -1614
rect 38040 -1648 38063 -1614
rect 37983 -1682 38063 -1648
rect 37983 -1716 38006 -1682
rect 38040 -1716 38063 -1682
rect 37983 -1750 38063 -1716
rect 37983 -1784 38006 -1750
rect 38040 -1784 38063 -1750
rect 37983 -1818 38063 -1784
rect 37983 -1852 38006 -1818
rect 38040 -1852 38063 -1818
rect 37983 -1886 38063 -1852
rect 37983 -1920 38006 -1886
rect 38040 -1920 38063 -1886
rect 37983 -1954 38063 -1920
rect 37983 -1988 38006 -1954
rect 38040 -1988 38063 -1954
rect 37983 -2022 38063 -1988
rect 37983 -2056 38006 -2022
rect 38040 -2056 38063 -2022
rect 37983 -2090 38063 -2056
rect 37983 -2124 38006 -2090
rect 38040 -2124 38063 -2090
rect 37983 -2158 38063 -2124
rect 37983 -2192 38006 -2158
rect 38040 -2192 38063 -2158
rect 37983 -2226 38063 -2192
rect 37983 -2260 38006 -2226
rect 38040 -2260 38063 -2226
rect 37983 -2294 38063 -2260
rect 37983 -2328 38006 -2294
rect 38040 -2328 38063 -2294
rect 37983 -2362 38063 -2328
rect 37983 -2396 38006 -2362
rect 38040 -2396 38063 -2362
rect 37983 -2430 38063 -2396
rect 37983 -2464 38006 -2430
rect 38040 -2464 38063 -2430
rect 37983 -2490 38063 -2464
rect 38133 -1546 38213 -1540
rect 38133 -1580 38156 -1546
rect 38190 -1580 38213 -1546
rect 38133 -1614 38213 -1580
rect 38133 -1648 38156 -1614
rect 38190 -1648 38213 -1614
rect 38133 -1682 38213 -1648
rect 38133 -1716 38156 -1682
rect 38190 -1716 38213 -1682
rect 38133 -1750 38213 -1716
rect 38133 -1784 38156 -1750
rect 38190 -1784 38213 -1750
rect 38133 -1818 38213 -1784
rect 38133 -1852 38156 -1818
rect 38190 -1852 38213 -1818
rect 38133 -1886 38213 -1852
rect 38133 -1920 38156 -1886
rect 38190 -1920 38213 -1886
rect 38133 -1954 38213 -1920
rect 38133 -1988 38156 -1954
rect 38190 -1988 38213 -1954
rect 38133 -2022 38213 -1988
rect 38133 -2056 38156 -2022
rect 38190 -2056 38213 -2022
rect 38133 -2090 38213 -2056
rect 38133 -2124 38156 -2090
rect 38190 -2124 38213 -2090
rect 38133 -2158 38213 -2124
rect 38133 -2192 38156 -2158
rect 38190 -2192 38213 -2158
rect 38133 -2226 38213 -2192
rect 38133 -2260 38156 -2226
rect 38190 -2260 38213 -2226
rect 38133 -2294 38213 -2260
rect 38133 -2328 38156 -2294
rect 38190 -2328 38213 -2294
rect 38133 -2362 38213 -2328
rect 38133 -2396 38156 -2362
rect 38190 -2396 38213 -2362
rect 38133 -2430 38213 -2396
rect 38133 -2464 38156 -2430
rect 38190 -2464 38213 -2430
rect 37833 -2545 37913 -2490
rect 38133 -2545 38213 -2464
rect 38283 -1546 38363 -1485
rect 38283 -1580 38306 -1546
rect 38340 -1580 38363 -1546
rect 38283 -1614 38363 -1580
rect 38283 -1648 38306 -1614
rect 38340 -1648 38363 -1614
rect 38283 -1682 38363 -1648
rect 38283 -1716 38306 -1682
rect 38340 -1716 38363 -1682
rect 38283 -1750 38363 -1716
rect 38283 -1784 38306 -1750
rect 38340 -1784 38363 -1750
rect 38283 -1818 38363 -1784
rect 38283 -1852 38306 -1818
rect 38340 -1852 38363 -1818
rect 38283 -1886 38363 -1852
rect 38283 -1920 38306 -1886
rect 38340 -1920 38363 -1886
rect 38283 -1954 38363 -1920
rect 38283 -1988 38306 -1954
rect 38340 -1988 38363 -1954
rect 38283 -2022 38363 -1988
rect 38283 -2056 38306 -2022
rect 38340 -2056 38363 -2022
rect 38283 -2090 38363 -2056
rect 38283 -2124 38306 -2090
rect 38340 -2124 38363 -2090
rect 38283 -2158 38363 -2124
rect 38283 -2192 38306 -2158
rect 38340 -2192 38363 -2158
rect 38283 -2226 38363 -2192
rect 38283 -2260 38306 -2226
rect 38340 -2260 38363 -2226
rect 38283 -2294 38363 -2260
rect 38283 -2328 38306 -2294
rect 38340 -2328 38363 -2294
rect 38283 -2362 38363 -2328
rect 38283 -2396 38306 -2362
rect 38340 -2396 38363 -2362
rect 38283 -2430 38363 -2396
rect 38283 -2464 38306 -2430
rect 38340 -2464 38363 -2430
rect 38283 -2490 38363 -2464
rect 38433 -1546 38513 -1540
rect 38433 -1580 38456 -1546
rect 38490 -1580 38513 -1546
rect 38433 -1614 38513 -1580
rect 38433 -1648 38456 -1614
rect 38490 -1648 38513 -1614
rect 38433 -1682 38513 -1648
rect 38433 -1716 38456 -1682
rect 38490 -1716 38513 -1682
rect 38433 -1750 38513 -1716
rect 38433 -1784 38456 -1750
rect 38490 -1784 38513 -1750
rect 38433 -1818 38513 -1784
rect 38433 -1852 38456 -1818
rect 38490 -1852 38513 -1818
rect 38433 -1886 38513 -1852
rect 38433 -1920 38456 -1886
rect 38490 -1920 38513 -1886
rect 38433 -1954 38513 -1920
rect 38433 -1988 38456 -1954
rect 38490 -1988 38513 -1954
rect 38433 -2022 38513 -1988
rect 38433 -2056 38456 -2022
rect 38490 -2056 38513 -2022
rect 38433 -2090 38513 -2056
rect 38433 -2124 38456 -2090
rect 38490 -2124 38513 -2090
rect 38433 -2158 38513 -2124
rect 38433 -2192 38456 -2158
rect 38490 -2192 38513 -2158
rect 38433 -2226 38513 -2192
rect 38433 -2260 38456 -2226
rect 38490 -2260 38513 -2226
rect 38433 -2294 38513 -2260
rect 38433 -2328 38456 -2294
rect 38490 -2328 38513 -2294
rect 38433 -2362 38513 -2328
rect 38433 -2396 38456 -2362
rect 38490 -2396 38513 -2362
rect 38433 -2430 38513 -2396
rect 38433 -2464 38456 -2430
rect 38490 -2464 38513 -2430
rect 38433 -2545 38513 -2464
rect 38583 -1546 38663 -1485
rect 38583 -1580 38606 -1546
rect 38640 -1580 38663 -1546
rect 38583 -1614 38663 -1580
rect 38583 -1648 38606 -1614
rect 38640 -1648 38663 -1614
rect 38583 -1682 38663 -1648
rect 38583 -1716 38606 -1682
rect 38640 -1716 38663 -1682
rect 38583 -1750 38663 -1716
rect 38583 -1784 38606 -1750
rect 38640 -1784 38663 -1750
rect 38583 -1818 38663 -1784
rect 38583 -1852 38606 -1818
rect 38640 -1852 38663 -1818
rect 38583 -1886 38663 -1852
rect 38583 -1920 38606 -1886
rect 38640 -1920 38663 -1886
rect 38583 -1954 38663 -1920
rect 38583 -1988 38606 -1954
rect 38640 -1988 38663 -1954
rect 38583 -2022 38663 -1988
rect 38583 -2056 38606 -2022
rect 38640 -2056 38663 -2022
rect 38583 -2090 38663 -2056
rect 38583 -2124 38606 -2090
rect 38640 -2124 38663 -2090
rect 38583 -2158 38663 -2124
rect 38583 -2192 38606 -2158
rect 38640 -2192 38663 -2158
rect 38583 -2226 38663 -2192
rect 38583 -2260 38606 -2226
rect 38640 -2260 38663 -2226
rect 38583 -2294 38663 -2260
rect 38583 -2328 38606 -2294
rect 38640 -2328 38663 -2294
rect 38583 -2362 38663 -2328
rect 38583 -2396 38606 -2362
rect 38640 -2396 38663 -2362
rect 38583 -2430 38663 -2396
rect 38583 -2464 38606 -2430
rect 38640 -2464 38663 -2430
rect 38583 -2490 38663 -2464
rect 38733 -1546 38813 -1540
rect 38733 -1580 38756 -1546
rect 38790 -1580 38813 -1546
rect 38733 -1614 38813 -1580
rect 38733 -1648 38756 -1614
rect 38790 -1648 38813 -1614
rect 38733 -1682 38813 -1648
rect 38733 -1716 38756 -1682
rect 38790 -1716 38813 -1682
rect 38733 -1750 38813 -1716
rect 38733 -1784 38756 -1750
rect 38790 -1784 38813 -1750
rect 38733 -1818 38813 -1784
rect 38733 -1852 38756 -1818
rect 38790 -1852 38813 -1818
rect 38733 -1886 38813 -1852
rect 38733 -1920 38756 -1886
rect 38790 -1920 38813 -1886
rect 38733 -1954 38813 -1920
rect 38733 -1988 38756 -1954
rect 38790 -1988 38813 -1954
rect 38733 -2022 38813 -1988
rect 38733 -2056 38756 -2022
rect 38790 -2056 38813 -2022
rect 38733 -2090 38813 -2056
rect 38733 -2124 38756 -2090
rect 38790 -2124 38813 -2090
rect 38733 -2158 38813 -2124
rect 38733 -2192 38756 -2158
rect 38790 -2192 38813 -2158
rect 38733 -2226 38813 -2192
rect 38733 -2260 38756 -2226
rect 38790 -2260 38813 -2226
rect 38733 -2294 38813 -2260
rect 38733 -2328 38756 -2294
rect 38790 -2328 38813 -2294
rect 38733 -2362 38813 -2328
rect 38733 -2396 38756 -2362
rect 38790 -2396 38813 -2362
rect 38733 -2430 38813 -2396
rect 38733 -2464 38756 -2430
rect 38790 -2464 38813 -2430
rect 38733 -2545 38813 -2464
rect 38883 -1546 38963 -1485
rect 38883 -1580 38906 -1546
rect 38940 -1580 38963 -1546
rect 38883 -1614 38963 -1580
rect 38883 -1648 38906 -1614
rect 38940 -1648 38963 -1614
rect 38883 -1682 38963 -1648
rect 38883 -1716 38906 -1682
rect 38940 -1716 38963 -1682
rect 38883 -1750 38963 -1716
rect 38883 -1784 38906 -1750
rect 38940 -1784 38963 -1750
rect 38883 -1818 38963 -1784
rect 38883 -1852 38906 -1818
rect 38940 -1852 38963 -1818
rect 38883 -1886 38963 -1852
rect 38883 -1920 38906 -1886
rect 38940 -1920 38963 -1886
rect 38883 -1954 38963 -1920
rect 38883 -1988 38906 -1954
rect 38940 -1988 38963 -1954
rect 38883 -2022 38963 -1988
rect 38883 -2056 38906 -2022
rect 38940 -2056 38963 -2022
rect 38883 -2090 38963 -2056
rect 38883 -2124 38906 -2090
rect 38940 -2124 38963 -2090
rect 38883 -2158 38963 -2124
rect 38883 -2192 38906 -2158
rect 38940 -2192 38963 -2158
rect 38883 -2226 38963 -2192
rect 38883 -2260 38906 -2226
rect 38940 -2260 38963 -2226
rect 38883 -2294 38963 -2260
rect 38883 -2328 38906 -2294
rect 38940 -2328 38963 -2294
rect 38883 -2362 38963 -2328
rect 38883 -2396 38906 -2362
rect 38940 -2396 38963 -2362
rect 38883 -2430 38963 -2396
rect 38883 -2464 38906 -2430
rect 38940 -2464 38963 -2430
rect 38883 -2490 38963 -2464
rect 39033 -1546 39113 -1540
rect 39033 -1580 39056 -1546
rect 39090 -1580 39113 -1546
rect 39033 -1614 39113 -1580
rect 39033 -1648 39056 -1614
rect 39090 -1648 39113 -1614
rect 39033 -1682 39113 -1648
rect 39033 -1716 39056 -1682
rect 39090 -1716 39113 -1682
rect 39033 -1750 39113 -1716
rect 39033 -1784 39056 -1750
rect 39090 -1784 39113 -1750
rect 39033 -1818 39113 -1784
rect 39033 -1852 39056 -1818
rect 39090 -1852 39113 -1818
rect 39033 -1886 39113 -1852
rect 39033 -1920 39056 -1886
rect 39090 -1920 39113 -1886
rect 39033 -1954 39113 -1920
rect 39033 -1988 39056 -1954
rect 39090 -1988 39113 -1954
rect 39033 -2022 39113 -1988
rect 39033 -2056 39056 -2022
rect 39090 -2056 39113 -2022
rect 39033 -2090 39113 -2056
rect 39033 -2124 39056 -2090
rect 39090 -2124 39113 -2090
rect 39033 -2158 39113 -2124
rect 39033 -2192 39056 -2158
rect 39090 -2192 39113 -2158
rect 39033 -2226 39113 -2192
rect 39033 -2260 39056 -2226
rect 39090 -2260 39113 -2226
rect 39033 -2294 39113 -2260
rect 39033 -2328 39056 -2294
rect 39090 -2328 39113 -2294
rect 39033 -2362 39113 -2328
rect 39033 -2396 39056 -2362
rect 39090 -2396 39113 -2362
rect 39033 -2430 39113 -2396
rect 39033 -2464 39056 -2430
rect 39090 -2464 39113 -2430
rect 39033 -2545 39113 -2464
rect 39183 -1546 39263 -1485
rect 39183 -1580 39206 -1546
rect 39240 -1580 39263 -1546
rect 39183 -1614 39263 -1580
rect 39183 -1648 39206 -1614
rect 39240 -1648 39263 -1614
rect 39183 -1682 39263 -1648
rect 39183 -1716 39206 -1682
rect 39240 -1716 39263 -1682
rect 39183 -1750 39263 -1716
rect 39183 -1784 39206 -1750
rect 39240 -1784 39263 -1750
rect 39183 -1818 39263 -1784
rect 39183 -1852 39206 -1818
rect 39240 -1852 39263 -1818
rect 39183 -1886 39263 -1852
rect 39183 -1920 39206 -1886
rect 39240 -1920 39263 -1886
rect 39183 -1954 39263 -1920
rect 39183 -1988 39206 -1954
rect 39240 -1988 39263 -1954
rect 39183 -2022 39263 -1988
rect 39183 -2056 39206 -2022
rect 39240 -2056 39263 -2022
rect 39183 -2090 39263 -2056
rect 39183 -2124 39206 -2090
rect 39240 -2124 39263 -2090
rect 39183 -2158 39263 -2124
rect 39183 -2192 39206 -2158
rect 39240 -2192 39263 -2158
rect 39183 -2226 39263 -2192
rect 39183 -2260 39206 -2226
rect 39240 -2260 39263 -2226
rect 39183 -2294 39263 -2260
rect 39183 -2328 39206 -2294
rect 39240 -2328 39263 -2294
rect 39183 -2362 39263 -2328
rect 39183 -2396 39206 -2362
rect 39240 -2396 39263 -2362
rect 39183 -2430 39263 -2396
rect 39183 -2464 39206 -2430
rect 39240 -2464 39263 -2430
rect 39183 -2490 39263 -2464
rect 39333 -1546 39413 -1540
rect 39333 -1580 39356 -1546
rect 39390 -1580 39413 -1546
rect 39333 -1614 39413 -1580
rect 39333 -1648 39356 -1614
rect 39390 -1648 39413 -1614
rect 39333 -1682 39413 -1648
rect 39333 -1716 39356 -1682
rect 39390 -1716 39413 -1682
rect 39333 -1750 39413 -1716
rect 39333 -1784 39356 -1750
rect 39390 -1784 39413 -1750
rect 39333 -1818 39413 -1784
rect 39333 -1852 39356 -1818
rect 39390 -1852 39413 -1818
rect 39333 -1886 39413 -1852
rect 44121 -1852 44162 -1849
rect 44196 -1852 44230 -1849
rect 44121 -1883 44156 -1852
rect 44196 -1883 44228 -1852
rect 44264 -1883 44298 -1849
rect 44332 -1852 44366 -1849
rect 44400 -1852 44441 -1849
rect 44334 -1883 44366 -1852
rect 44406 -1883 44441 -1852
rect 39333 -1920 39356 -1886
rect 39390 -1920 39413 -1886
rect 44137 -1886 44156 -1883
rect 44190 -1886 44228 -1883
rect 44262 -1886 44300 -1883
rect 44334 -1886 44372 -1883
rect 44406 -1886 44425 -1883
rect 44137 -1889 44425 -1886
rect 39333 -1954 39413 -1920
rect 39333 -1988 39356 -1954
rect 39390 -1988 39413 -1954
rect 39333 -2022 39413 -1988
rect 39333 -2056 39356 -2022
rect 39390 -2056 39413 -2022
rect 39333 -2090 39413 -2056
rect 39333 -2124 39356 -2090
rect 39390 -2124 39413 -2090
rect 39333 -2158 39413 -2124
rect 39333 -2192 39356 -2158
rect 39390 -2192 39413 -2158
rect 39333 -2226 39413 -2192
rect 39333 -2260 39356 -2226
rect 39390 -2260 39413 -2226
rect 39333 -2294 39413 -2260
rect 44137 -2258 44425 -2255
rect 44137 -2261 44156 -2258
rect 44190 -2261 44228 -2258
rect 44262 -2261 44300 -2258
rect 44334 -2261 44372 -2258
rect 44406 -2261 44425 -2258
rect 39333 -2328 39356 -2294
rect 39390 -2328 39413 -2294
rect 44121 -2292 44156 -2261
rect 44196 -2292 44228 -2261
rect 44121 -2295 44162 -2292
rect 44196 -2295 44230 -2292
rect 44264 -2295 44298 -2261
rect 44334 -2292 44366 -2261
rect 44406 -2292 44441 -2261
rect 44332 -2295 44366 -2292
rect 44400 -2295 44441 -2292
rect 39333 -2362 39413 -2328
rect 39333 -2396 39356 -2362
rect 39390 -2396 39413 -2362
rect 39333 -2430 39413 -2396
rect 39333 -2464 39356 -2430
rect 39390 -2464 39413 -2430
rect 39333 -2545 39413 -2464
rect 35929 -2625 39414 -2545
rect 35930 -2840 37300 -2625
rect 35312 -2862 51662 -2840
rect 35312 -2896 35347 -2862
rect 35381 -2896 35427 -2862
rect 35461 -2896 35507 -2862
rect 35541 -2896 35587 -2862
rect 35621 -2896 35667 -2862
rect 35701 -2896 35747 -2862
rect 35781 -2896 35827 -2862
rect 35861 -2896 35907 -2862
rect 35941 -2896 35987 -2862
rect 36021 -2896 36067 -2862
rect 36101 -2896 36147 -2862
rect 36181 -2896 36227 -2862
rect 36261 -2896 36307 -2862
rect 36341 -2896 36387 -2862
rect 36421 -2896 36467 -2862
rect 36501 -2896 36547 -2862
rect 36581 -2896 36627 -2862
rect 36661 -2896 36707 -2862
rect 36741 -2896 36787 -2862
rect 36821 -2896 36867 -2862
rect 36901 -2896 36947 -2862
rect 36981 -2896 37027 -2862
rect 37061 -2896 37107 -2862
rect 37141 -2896 37187 -2862
rect 37221 -2896 37267 -2862
rect 37301 -2896 37347 -2862
rect 37381 -2896 37427 -2862
rect 37461 -2896 37507 -2862
rect 37541 -2896 37587 -2862
rect 37621 -2896 37667 -2862
rect 37701 -2896 37747 -2862
rect 37781 -2896 37827 -2862
rect 37861 -2896 37907 -2862
rect 37941 -2896 37987 -2862
rect 38021 -2896 38067 -2862
rect 38101 -2896 38147 -2862
rect 38181 -2896 38227 -2862
rect 38261 -2896 38307 -2862
rect 38341 -2896 38387 -2862
rect 38421 -2896 38467 -2862
rect 38501 -2896 38547 -2862
rect 38581 -2896 38627 -2862
rect 38661 -2896 38707 -2862
rect 38741 -2896 38787 -2862
rect 38821 -2896 38867 -2862
rect 38901 -2896 38947 -2862
rect 38981 -2896 39027 -2862
rect 39061 -2896 39107 -2862
rect 39141 -2896 39188 -2862
rect 39222 -2896 39268 -2862
rect 39302 -2896 39348 -2862
rect 39382 -2896 39428 -2862
rect 39462 -2896 39508 -2862
rect 39542 -2896 39588 -2862
rect 39622 -2896 39668 -2862
rect 39702 -2896 39748 -2862
rect 39782 -2896 39828 -2862
rect 39862 -2896 39908 -2862
rect 39942 -2896 39988 -2862
rect 40022 -2896 40068 -2862
rect 40102 -2896 40148 -2862
rect 40182 -2896 40228 -2862
rect 40262 -2896 40308 -2862
rect 40342 -2896 40388 -2862
rect 40422 -2896 40468 -2862
rect 40502 -2896 40548 -2862
rect 40582 -2896 40628 -2862
rect 40662 -2896 40708 -2862
rect 40742 -2896 40788 -2862
rect 40822 -2896 40868 -2862
rect 40902 -2896 40948 -2862
rect 40982 -2896 41028 -2862
rect 41062 -2896 41108 -2862
rect 41142 -2896 41188 -2862
rect 41222 -2896 41268 -2862
rect 41302 -2896 41348 -2862
rect 41382 -2896 41428 -2862
rect 41462 -2896 41508 -2862
rect 41542 -2896 41588 -2862
rect 41622 -2896 41668 -2862
rect 41702 -2896 41748 -2862
rect 41782 -2896 41828 -2862
rect 41862 -2896 41908 -2862
rect 41942 -2896 41988 -2862
rect 42022 -2896 42068 -2862
rect 42102 -2896 42148 -2862
rect 42182 -2896 42228 -2862
rect 42262 -2896 42308 -2862
rect 42342 -2896 42388 -2862
rect 42422 -2896 42468 -2862
rect 42502 -2896 42548 -2862
rect 42582 -2896 42628 -2862
rect 42662 -2896 42708 -2862
rect 42742 -2896 42788 -2862
rect 42822 -2896 42868 -2862
rect 42902 -2896 42948 -2862
rect 42982 -2896 43028 -2862
rect 43062 -2896 43108 -2862
rect 43142 -2896 43188 -2862
rect 43222 -2896 43268 -2862
rect 43302 -2896 43348 -2862
rect 43382 -2896 43428 -2862
rect 43462 -2896 43508 -2862
rect 43542 -2896 43588 -2862
rect 43622 -2896 43668 -2862
rect 43702 -2896 43748 -2862
rect 43782 -2896 43828 -2862
rect 43862 -2896 43908 -2862
rect 43942 -2896 43988 -2862
rect 44022 -2896 44068 -2862
rect 44102 -2896 44148 -2862
rect 44182 -2896 44228 -2862
rect 44262 -2896 44308 -2862
rect 44342 -2896 44388 -2862
rect 44422 -2896 44468 -2862
rect 44502 -2896 44548 -2862
rect 44582 -2896 44628 -2862
rect 44662 -2896 44708 -2862
rect 44742 -2896 44788 -2862
rect 44822 -2896 44868 -2862
rect 44902 -2896 44948 -2862
rect 44982 -2896 45028 -2862
rect 45062 -2896 45108 -2862
rect 45142 -2896 45188 -2862
rect 45222 -2896 45268 -2862
rect 45302 -2896 45348 -2862
rect 45382 -2896 45428 -2862
rect 45462 -2896 45508 -2862
rect 45542 -2896 45588 -2862
rect 45622 -2896 45668 -2862
rect 45702 -2896 45748 -2862
rect 45782 -2896 45828 -2862
rect 45862 -2896 45908 -2862
rect 45942 -2896 45988 -2862
rect 46022 -2896 46068 -2862
rect 46102 -2896 46148 -2862
rect 46182 -2896 46228 -2862
rect 46262 -2896 46308 -2862
rect 46342 -2896 46388 -2862
rect 46422 -2896 46468 -2862
rect 46502 -2896 46548 -2862
rect 46582 -2896 46628 -2862
rect 46662 -2896 46708 -2862
rect 46742 -2896 46788 -2862
rect 46822 -2896 46868 -2862
rect 46902 -2896 46948 -2862
rect 46982 -2896 47028 -2862
rect 47062 -2896 47108 -2862
rect 47142 -2896 47188 -2862
rect 47222 -2896 47268 -2862
rect 47302 -2896 47349 -2862
rect 47383 -2896 47429 -2862
rect 47463 -2896 47509 -2862
rect 47543 -2896 47589 -2862
rect 47623 -2896 47669 -2862
rect 47703 -2896 47749 -2862
rect 47783 -2896 47829 -2862
rect 47863 -2896 47909 -2862
rect 47943 -2896 47989 -2862
rect 48023 -2896 48069 -2862
rect 48103 -2896 48149 -2862
rect 48183 -2896 48229 -2862
rect 48263 -2896 48309 -2862
rect 48343 -2896 48389 -2862
rect 48423 -2896 48469 -2862
rect 48503 -2896 48549 -2862
rect 48583 -2896 48629 -2862
rect 48663 -2896 48709 -2862
rect 48743 -2896 48789 -2862
rect 48823 -2896 48869 -2862
rect 48903 -2896 48949 -2862
rect 48983 -2896 49029 -2862
rect 49063 -2896 49109 -2862
rect 49143 -2896 49189 -2862
rect 49223 -2896 49269 -2862
rect 49303 -2896 49349 -2862
rect 49383 -2896 49429 -2862
rect 49463 -2896 49509 -2862
rect 49543 -2896 49589 -2862
rect 49623 -2896 49669 -2862
rect 49703 -2896 49749 -2862
rect 49783 -2896 49829 -2862
rect 49863 -2896 49909 -2862
rect 49943 -2896 49989 -2862
rect 50023 -2896 50069 -2862
rect 50103 -2896 50149 -2862
rect 50183 -2896 50229 -2862
rect 50263 -2896 50309 -2862
rect 50343 -2896 50389 -2862
rect 50423 -2896 50469 -2862
rect 50503 -2896 50549 -2862
rect 50583 -2896 50629 -2862
rect 50663 -2896 50709 -2862
rect 50743 -2896 50789 -2862
rect 50823 -2896 50869 -2862
rect 50903 -2896 50949 -2862
rect 50983 -2896 51029 -2862
rect 51063 -2896 51109 -2862
rect 51143 -2896 51189 -2862
rect 51223 -2896 51269 -2862
rect 51303 -2896 51349 -2862
rect 51383 -2896 51429 -2862
rect 51463 -2896 51509 -2862
rect 51543 -2896 51589 -2862
rect 51623 -2896 51662 -2862
rect 35312 -2952 51662 -2896
rect 35312 -2986 35347 -2952
rect 35381 -2986 35427 -2952
rect 35461 -2986 35507 -2952
rect 35541 -2986 35587 -2952
rect 35621 -2986 35667 -2952
rect 35701 -2986 35747 -2952
rect 35781 -2986 35827 -2952
rect 35861 -2986 35907 -2952
rect 35941 -2986 35987 -2952
rect 36021 -2986 36067 -2952
rect 36101 -2986 36147 -2952
rect 36181 -2986 36227 -2952
rect 36261 -2986 36307 -2952
rect 36341 -2986 36387 -2952
rect 36421 -2986 36467 -2952
rect 36501 -2986 36547 -2952
rect 36581 -2986 36627 -2952
rect 36661 -2986 36707 -2952
rect 36741 -2986 36787 -2952
rect 36821 -2986 36867 -2952
rect 36901 -2986 36947 -2952
rect 36981 -2986 37027 -2952
rect 37061 -2986 37107 -2952
rect 37141 -2986 37187 -2952
rect 37221 -2986 37267 -2952
rect 37301 -2986 37347 -2952
rect 37381 -2986 37427 -2952
rect 37461 -2986 37507 -2952
rect 37541 -2986 37587 -2952
rect 37621 -2986 37667 -2952
rect 37701 -2986 37747 -2952
rect 37781 -2986 37827 -2952
rect 37861 -2986 37907 -2952
rect 37941 -2986 37987 -2952
rect 38021 -2986 38067 -2952
rect 38101 -2986 38147 -2952
rect 38181 -2986 38227 -2952
rect 38261 -2986 38307 -2952
rect 38341 -2986 38387 -2952
rect 38421 -2986 38467 -2952
rect 38501 -2986 38547 -2952
rect 38581 -2986 38627 -2952
rect 38661 -2986 38707 -2952
rect 38741 -2986 38787 -2952
rect 38821 -2986 38867 -2952
rect 38901 -2986 38947 -2952
rect 38981 -2986 39027 -2952
rect 39061 -2986 39107 -2952
rect 39141 -2986 39188 -2952
rect 39222 -2986 39268 -2952
rect 39302 -2986 39348 -2952
rect 39382 -2986 39428 -2952
rect 39462 -2986 39508 -2952
rect 39542 -2986 39588 -2952
rect 39622 -2986 39668 -2952
rect 39702 -2986 39748 -2952
rect 39782 -2986 39828 -2952
rect 39862 -2986 39908 -2952
rect 39942 -2986 39988 -2952
rect 40022 -2986 40068 -2952
rect 40102 -2986 40148 -2952
rect 40182 -2986 40228 -2952
rect 40262 -2986 40308 -2952
rect 40342 -2986 40388 -2952
rect 40422 -2986 40468 -2952
rect 40502 -2986 40548 -2952
rect 40582 -2986 40628 -2952
rect 40662 -2986 40708 -2952
rect 40742 -2986 40788 -2952
rect 40822 -2986 40868 -2952
rect 40902 -2986 40948 -2952
rect 40982 -2986 41028 -2952
rect 41062 -2986 41108 -2952
rect 41142 -2986 41188 -2952
rect 41222 -2986 41268 -2952
rect 41302 -2986 41348 -2952
rect 41382 -2986 41428 -2952
rect 41462 -2986 41508 -2952
rect 41542 -2986 41588 -2952
rect 41622 -2986 41668 -2952
rect 41702 -2986 41748 -2952
rect 41782 -2986 41828 -2952
rect 41862 -2986 41908 -2952
rect 41942 -2986 41988 -2952
rect 42022 -2986 42068 -2952
rect 42102 -2986 42148 -2952
rect 42182 -2986 42228 -2952
rect 42262 -2986 42308 -2952
rect 42342 -2986 42388 -2952
rect 42422 -2986 42468 -2952
rect 42502 -2986 42548 -2952
rect 42582 -2986 42628 -2952
rect 42662 -2986 42708 -2952
rect 42742 -2986 42788 -2952
rect 42822 -2986 42868 -2952
rect 42902 -2986 42948 -2952
rect 42982 -2986 43028 -2952
rect 43062 -2986 43108 -2952
rect 43142 -2986 43188 -2952
rect 43222 -2986 43268 -2952
rect 43302 -2986 43348 -2952
rect 43382 -2986 43428 -2952
rect 43462 -2986 43508 -2952
rect 43542 -2986 43588 -2952
rect 43622 -2986 43668 -2952
rect 43702 -2986 43748 -2952
rect 43782 -2986 43828 -2952
rect 43862 -2986 43908 -2952
rect 43942 -2986 43988 -2952
rect 44022 -2986 44068 -2952
rect 44102 -2986 44148 -2952
rect 44182 -2986 44228 -2952
rect 44262 -2986 44308 -2952
rect 44342 -2986 44388 -2952
rect 44422 -2986 44468 -2952
rect 44502 -2986 44548 -2952
rect 44582 -2986 44628 -2952
rect 44662 -2986 44708 -2952
rect 44742 -2986 44788 -2952
rect 44822 -2986 44868 -2952
rect 44902 -2986 44948 -2952
rect 44982 -2986 45028 -2952
rect 45062 -2986 45108 -2952
rect 45142 -2986 45188 -2952
rect 45222 -2986 45268 -2952
rect 45302 -2986 45348 -2952
rect 45382 -2986 45428 -2952
rect 45462 -2986 45508 -2952
rect 45542 -2986 45588 -2952
rect 45622 -2986 45668 -2952
rect 45702 -2986 45748 -2952
rect 45782 -2986 45828 -2952
rect 45862 -2986 45908 -2952
rect 45942 -2986 45988 -2952
rect 46022 -2986 46068 -2952
rect 46102 -2986 46148 -2952
rect 46182 -2986 46228 -2952
rect 46262 -2986 46308 -2952
rect 46342 -2986 46388 -2952
rect 46422 -2986 46468 -2952
rect 46502 -2986 46548 -2952
rect 46582 -2986 46628 -2952
rect 46662 -2986 46708 -2952
rect 46742 -2986 46788 -2952
rect 46822 -2986 46868 -2952
rect 46902 -2986 46948 -2952
rect 46982 -2986 47028 -2952
rect 47062 -2986 47108 -2952
rect 47142 -2986 47188 -2952
rect 47222 -2986 47268 -2952
rect 47302 -2986 47349 -2952
rect 47383 -2986 47429 -2952
rect 47463 -2986 47509 -2952
rect 47543 -2986 47589 -2952
rect 47623 -2986 47669 -2952
rect 47703 -2986 47749 -2952
rect 47783 -2986 47829 -2952
rect 47863 -2986 47909 -2952
rect 47943 -2986 47989 -2952
rect 48023 -2986 48069 -2952
rect 48103 -2986 48149 -2952
rect 48183 -2986 48229 -2952
rect 48263 -2986 48309 -2952
rect 48343 -2986 48389 -2952
rect 48423 -2986 48469 -2952
rect 48503 -2986 48549 -2952
rect 48583 -2986 48629 -2952
rect 48663 -2986 48709 -2952
rect 48743 -2986 48789 -2952
rect 48823 -2986 48869 -2952
rect 48903 -2986 48949 -2952
rect 48983 -2986 49029 -2952
rect 49063 -2986 49109 -2952
rect 49143 -2986 49189 -2952
rect 49223 -2986 49269 -2952
rect 49303 -2986 49349 -2952
rect 49383 -2986 49429 -2952
rect 49463 -2986 49509 -2952
rect 49543 -2986 49589 -2952
rect 49623 -2986 49669 -2952
rect 49703 -2986 49749 -2952
rect 49783 -2986 49829 -2952
rect 49863 -2986 49909 -2952
rect 49943 -2986 49989 -2952
rect 50023 -2986 50069 -2952
rect 50103 -2986 50149 -2952
rect 50183 -2986 50229 -2952
rect 50263 -2986 50309 -2952
rect 50343 -2986 50389 -2952
rect 50423 -2986 50469 -2952
rect 50503 -2986 50549 -2952
rect 50583 -2986 50629 -2952
rect 50663 -2986 50709 -2952
rect 50743 -2986 50789 -2952
rect 50823 -2986 50869 -2952
rect 50903 -2986 50949 -2952
rect 50983 -2986 51029 -2952
rect 51063 -2986 51109 -2952
rect 51143 -2986 51189 -2952
rect 51223 -2986 51269 -2952
rect 51303 -2986 51349 -2952
rect 51383 -2986 51429 -2952
rect 51463 -2986 51509 -2952
rect 51543 -2986 51589 -2952
rect 51623 -2986 51662 -2952
rect 35312 -3010 51662 -2986
rect 39460 -3073 39540 -3050
rect 39460 -3107 39483 -3073
rect 39517 -3107 39540 -3073
rect 39460 -3130 39540 -3107
rect 39580 -3073 39660 -3050
rect 39580 -3107 39603 -3073
rect 39637 -3107 39660 -3073
rect 39580 -3130 39660 -3107
rect 39460 -3193 39540 -3170
rect 39460 -3227 39483 -3193
rect 39517 -3227 39540 -3193
rect 39460 -3250 39540 -3227
rect 39580 -3193 39660 -3170
rect 39580 -3227 39603 -3193
rect 39637 -3227 39660 -3193
rect 39580 -3250 39660 -3227
<< viali >>
rect 39455 9704 39489 9738
rect 39575 9704 39609 9738
rect 39455 9584 39489 9618
rect 39575 9584 39609 9618
rect 27949 2640 27983 2674
rect 28029 2640 28063 2674
rect 28109 2640 28143 2674
rect 28189 2640 28223 2674
rect 28269 2640 28303 2674
rect 28349 2640 28383 2674
rect 28429 2640 28463 2674
rect 28509 2640 28543 2674
rect 28589 2640 28623 2674
rect 28669 2640 28703 2674
rect 28749 2640 28783 2674
rect 28829 2640 28863 2674
rect 28909 2640 28943 2674
rect 28989 2640 29023 2674
rect 29069 2640 29103 2674
rect 29149 2640 29183 2674
rect 29229 2640 29263 2674
rect 29309 2640 29343 2674
rect 29389 2640 29423 2674
rect 29469 2640 29503 2674
rect 29549 2640 29583 2674
rect 29629 2640 29663 2674
rect 29709 2640 29743 2674
rect 29789 2640 29823 2674
rect 29869 2640 29903 2674
rect 29949 2640 29983 2674
rect 30029 2640 30063 2674
rect 30109 2640 30143 2674
rect 30189 2640 30223 2674
rect 30269 2640 30303 2674
rect 30349 2640 30383 2674
rect 30429 2640 30463 2674
rect 30509 2640 30543 2674
rect 30589 2640 30623 2674
rect 30669 2640 30703 2674
rect 30749 2640 30783 2674
rect 30829 2640 30863 2674
rect 30910 2640 30944 2674
rect 30990 2640 31024 2674
rect 31070 2640 31104 2674
rect 31150 2640 31184 2674
rect 31230 2640 31264 2674
rect 31310 2640 31344 2674
rect 31390 2640 31424 2674
rect 31470 2640 31504 2674
rect 31550 2640 31584 2674
rect 31630 2640 31664 2674
rect 31710 2640 31744 2674
rect 31790 2640 31824 2674
rect 31870 2640 31904 2674
rect 31950 2640 31984 2674
rect 32030 2640 32064 2674
rect 32110 2640 32144 2674
rect 32190 2640 32224 2674
rect 32270 2640 32304 2674
rect 32350 2640 32384 2674
rect 32430 2640 32464 2674
rect 32510 2640 32544 2674
rect 32590 2640 32624 2674
rect 32670 2640 32704 2674
rect 32750 2640 32784 2674
rect 32830 2640 32864 2674
rect 32910 2640 32944 2674
rect 32990 2640 33024 2674
rect 33070 2640 33104 2674
rect 33150 2640 33184 2674
rect 33230 2640 33264 2674
rect 33310 2640 33344 2674
rect 33390 2640 33424 2674
rect 33470 2640 33504 2674
rect 33550 2640 33584 2674
rect 33630 2640 33664 2674
rect 33710 2640 33744 2674
rect 33790 2640 33824 2674
rect 33870 2640 33904 2674
rect 33950 2640 33984 2674
rect 34030 2640 34064 2674
rect 34110 2640 34144 2674
rect 34190 2640 34224 2674
rect 34270 2640 34304 2674
rect 34350 2640 34384 2674
rect 34430 2640 34464 2674
rect 34510 2640 34544 2674
rect 34590 2640 34624 2674
rect 34670 2640 34704 2674
rect 34750 2640 34784 2674
rect 34830 2640 34864 2674
rect 34910 2640 34944 2674
rect 34990 2640 35024 2674
rect 35070 2640 35104 2674
rect 35150 2640 35184 2674
rect 35242 2640 35276 2674
rect 35322 2640 35356 2674
rect 35402 2640 35436 2674
rect 35482 2640 35516 2674
rect 35562 2640 35596 2674
rect 35642 2640 35676 2674
rect 35722 2640 35756 2674
rect 35802 2640 35836 2674
rect 35882 2640 35916 2674
rect 35962 2640 35996 2674
rect 36042 2640 36076 2674
rect 36122 2640 36156 2674
rect 36202 2640 36236 2674
rect 36282 2640 36316 2674
rect 36362 2640 36396 2674
rect 36442 2640 36476 2674
rect 36522 2640 36556 2674
rect 36602 2640 36636 2674
rect 36682 2640 36716 2674
rect 36762 2640 36796 2674
rect 36842 2640 36876 2674
rect 36922 2640 36956 2674
rect 37002 2640 37036 2674
rect 37082 2640 37116 2674
rect 37162 2640 37196 2674
rect 37242 2640 37276 2674
rect 37322 2640 37356 2674
rect 37402 2640 37436 2674
rect 37482 2640 37516 2674
rect 37562 2640 37596 2674
rect 37642 2640 37676 2674
rect 37722 2640 37756 2674
rect 37802 2640 37836 2674
rect 37882 2640 37916 2674
rect 37962 2640 37996 2674
rect 38042 2640 38076 2674
rect 38122 2640 38156 2674
rect 38202 2640 38236 2674
rect 38282 2640 38316 2674
rect 38362 2640 38396 2674
rect 38442 2640 38476 2674
rect 38522 2640 38556 2674
rect 38602 2640 38636 2674
rect 38682 2640 38716 2674
rect 38762 2640 38796 2674
rect 38842 2640 38876 2674
rect 38922 2640 38956 2674
rect 39002 2640 39036 2674
rect 39083 2640 39117 2674
rect 39163 2640 39197 2674
rect 39243 2640 39277 2674
rect 39323 2640 39357 2674
rect 39403 2640 39437 2674
rect 39483 2640 39517 2674
rect 39563 2640 39597 2674
rect 39643 2640 39677 2674
rect 39723 2640 39757 2674
rect 39803 2640 39837 2674
rect 39883 2640 39917 2674
rect 39963 2640 39997 2674
rect 40043 2640 40077 2674
rect 40123 2640 40157 2674
rect 40203 2640 40237 2674
rect 40283 2640 40317 2674
rect 40363 2640 40397 2674
rect 40443 2640 40477 2674
rect 40523 2640 40557 2674
rect 40603 2640 40637 2674
rect 40683 2640 40717 2674
rect 40763 2640 40797 2674
rect 40843 2640 40877 2674
rect 40923 2640 40957 2674
rect 41003 2640 41037 2674
rect 41083 2640 41117 2674
rect 41163 2640 41197 2674
rect 41243 2640 41277 2674
rect 41323 2640 41357 2674
rect 41403 2640 41437 2674
rect 41483 2640 41517 2674
rect 41563 2640 41597 2674
rect 41643 2640 41677 2674
rect 41723 2640 41757 2674
rect 41803 2640 41837 2674
rect 41883 2640 41917 2674
rect 41963 2640 41997 2674
rect 42043 2640 42077 2674
rect 42123 2640 42157 2674
rect 42203 2640 42237 2674
rect 42283 2640 42317 2674
rect 42363 2640 42397 2674
rect 42443 2640 42477 2674
rect 42523 2640 42557 2674
rect 42603 2640 42637 2674
rect 42683 2640 42717 2674
rect 42763 2640 42797 2674
rect 42843 2640 42877 2674
rect 42923 2640 42957 2674
rect 43003 2640 43037 2674
rect 43083 2640 43117 2674
rect 43163 2640 43197 2674
rect 43243 2640 43277 2674
rect 43323 2640 43357 2674
rect 27949 2550 27983 2584
rect 28029 2550 28063 2584
rect 28109 2550 28143 2584
rect 28189 2550 28223 2584
rect 28269 2550 28303 2584
rect 28349 2550 28383 2584
rect 28429 2550 28463 2584
rect 28509 2550 28543 2584
rect 28589 2550 28623 2584
rect 28669 2550 28703 2584
rect 28749 2550 28783 2584
rect 28829 2550 28863 2584
rect 28909 2550 28943 2584
rect 28989 2550 29023 2584
rect 29069 2550 29103 2584
rect 29149 2550 29183 2584
rect 29229 2550 29263 2584
rect 29309 2550 29343 2584
rect 29389 2550 29423 2584
rect 29469 2550 29503 2584
rect 29549 2550 29583 2584
rect 29629 2550 29663 2584
rect 29709 2550 29743 2584
rect 29789 2550 29823 2584
rect 29869 2550 29903 2584
rect 29949 2550 29983 2584
rect 30029 2550 30063 2584
rect 30109 2550 30143 2584
rect 30189 2550 30223 2584
rect 30269 2550 30303 2584
rect 30349 2550 30383 2584
rect 30429 2550 30463 2584
rect 30509 2550 30543 2584
rect 30589 2550 30623 2584
rect 30669 2550 30703 2584
rect 30749 2550 30783 2584
rect 30829 2550 30863 2584
rect 30910 2550 30944 2584
rect 30990 2550 31024 2584
rect 31070 2550 31104 2584
rect 31150 2550 31184 2584
rect 31230 2550 31264 2584
rect 31310 2550 31344 2584
rect 31390 2550 31424 2584
rect 31470 2550 31504 2584
rect 31550 2550 31584 2584
rect 31630 2550 31664 2584
rect 31710 2550 31744 2584
rect 31790 2550 31824 2584
rect 31870 2550 31904 2584
rect 31950 2550 31984 2584
rect 32030 2550 32064 2584
rect 32110 2550 32144 2584
rect 32190 2550 32224 2584
rect 32270 2550 32304 2584
rect 32350 2550 32384 2584
rect 32430 2550 32464 2584
rect 32510 2550 32544 2584
rect 32590 2550 32624 2584
rect 32670 2550 32704 2584
rect 32750 2550 32784 2584
rect 32830 2550 32864 2584
rect 32910 2550 32944 2584
rect 32990 2550 33024 2584
rect 33070 2550 33104 2584
rect 33150 2550 33184 2584
rect 33230 2550 33264 2584
rect 33310 2550 33344 2584
rect 33390 2550 33424 2584
rect 33470 2550 33504 2584
rect 33550 2550 33584 2584
rect 33630 2550 33664 2584
rect 33710 2550 33744 2584
rect 33790 2550 33824 2584
rect 33870 2550 33904 2584
rect 33950 2550 33984 2584
rect 34030 2550 34064 2584
rect 34110 2550 34144 2584
rect 34190 2550 34224 2584
rect 34270 2550 34304 2584
rect 34350 2550 34384 2584
rect 34430 2550 34464 2584
rect 34510 2550 34544 2584
rect 34590 2550 34624 2584
rect 34670 2550 34704 2584
rect 34750 2550 34784 2584
rect 34830 2550 34864 2584
rect 34910 2550 34944 2584
rect 34990 2550 35024 2584
rect 35070 2550 35104 2584
rect 35150 2550 35184 2584
rect 35242 2550 35276 2584
rect 35322 2550 35356 2584
rect 35402 2550 35436 2584
rect 35482 2550 35516 2584
rect 35562 2550 35596 2584
rect 35642 2550 35676 2584
rect 35722 2550 35756 2584
rect 35802 2550 35836 2584
rect 35882 2550 35916 2584
rect 35962 2550 35996 2584
rect 36042 2550 36076 2584
rect 36122 2550 36156 2584
rect 36202 2550 36236 2584
rect 36282 2550 36316 2584
rect 36362 2550 36396 2584
rect 36442 2550 36476 2584
rect 36522 2550 36556 2584
rect 36602 2550 36636 2584
rect 36682 2550 36716 2584
rect 36762 2550 36796 2584
rect 36842 2550 36876 2584
rect 36922 2550 36956 2584
rect 37002 2550 37036 2584
rect 37082 2550 37116 2584
rect 37162 2550 37196 2584
rect 37242 2550 37276 2584
rect 37322 2550 37356 2584
rect 37402 2550 37436 2584
rect 37482 2550 37516 2584
rect 37562 2550 37596 2584
rect 37642 2550 37676 2584
rect 37722 2550 37756 2584
rect 37802 2550 37836 2584
rect 37882 2550 37916 2584
rect 37962 2550 37996 2584
rect 38042 2550 38076 2584
rect 38122 2550 38156 2584
rect 38202 2550 38236 2584
rect 38282 2550 38316 2584
rect 38362 2550 38396 2584
rect 38442 2550 38476 2584
rect 38522 2550 38556 2584
rect 38602 2550 38636 2584
rect 38682 2550 38716 2584
rect 38762 2550 38796 2584
rect 38842 2550 38876 2584
rect 38922 2550 38956 2584
rect 39002 2550 39036 2584
rect 39083 2550 39117 2584
rect 39163 2550 39197 2584
rect 39243 2550 39277 2584
rect 39323 2550 39357 2584
rect 39403 2550 39437 2584
rect 39483 2550 39517 2584
rect 39563 2550 39597 2584
rect 39643 2550 39677 2584
rect 39723 2550 39757 2584
rect 39803 2550 39837 2584
rect 39883 2550 39917 2584
rect 39963 2550 39997 2584
rect 40043 2550 40077 2584
rect 40123 2550 40157 2584
rect 40203 2550 40237 2584
rect 40283 2550 40317 2584
rect 40363 2550 40397 2584
rect 40443 2550 40477 2584
rect 40523 2550 40557 2584
rect 40603 2550 40637 2584
rect 40683 2550 40717 2584
rect 40763 2550 40797 2584
rect 40843 2550 40877 2584
rect 40923 2550 40957 2584
rect 41003 2550 41037 2584
rect 41083 2550 41117 2584
rect 41163 2550 41197 2584
rect 41243 2550 41277 2584
rect 41323 2550 41357 2584
rect 41403 2550 41437 2584
rect 41483 2550 41517 2584
rect 41563 2550 41597 2584
rect 41643 2550 41677 2584
rect 41723 2550 41757 2584
rect 41803 2550 41837 2584
rect 41883 2550 41917 2584
rect 41963 2550 41997 2584
rect 42043 2550 42077 2584
rect 42123 2550 42157 2584
rect 42203 2550 42237 2584
rect 42283 2550 42317 2584
rect 42363 2550 42397 2584
rect 42443 2550 42477 2584
rect 42523 2550 42557 2584
rect 42603 2550 42637 2584
rect 42683 2550 42717 2584
rect 42763 2550 42797 2584
rect 42843 2550 42877 2584
rect 42923 2550 42957 2584
rect 43003 2550 43037 2584
rect 43083 2550 43117 2584
rect 43163 2550 43197 2584
rect 43243 2550 43277 2584
rect 43323 2550 43357 2584
rect 32560 1500 32620 1560
rect 32680 1500 32740 1560
rect 32980 1500 33040 1560
rect 33110 1510 33150 1550
rect 32560 1380 32620 1440
rect 32680 1380 32740 1440
rect 32980 1380 33040 1440
rect 33100 1380 33160 1440
rect 34309 1511 34343 1545
rect 34429 1511 34463 1545
rect 34309 1391 34343 1425
rect 34429 1391 34463 1425
rect 34729 1511 34763 1545
rect 34849 1511 34883 1545
rect 34729 1391 34763 1425
rect 34849 1391 34883 1425
rect 32560 1080 32620 1140
rect 32695 1091 32729 1125
rect 32980 1080 33040 1140
rect 33100 1080 33160 1140
rect 32560 960 32620 1020
rect 32680 960 32740 1020
rect 32980 960 33040 1020
rect 33100 960 33160 1020
rect 34309 1091 34343 1125
rect 34429 1091 34463 1125
rect 34309 971 34343 1005
rect 34429 971 34463 1005
rect 34729 1091 34763 1125
rect 34849 1091 34883 1125
rect 34729 971 34763 1005
rect 34849 971 34883 1005
rect 44218 -84 44270 -32
rect 44338 -84 44390 -32
rect 44226 -85 44260 -84
rect 44346 -85 44380 -84
rect 44218 -204 44270 -152
rect 44338 -204 44390 -152
rect 44226 -205 44260 -204
rect 44346 -205 44380 -204
rect 35818 -521 35852 -487
rect 35938 -521 35972 -487
rect 35818 -641 35852 -607
rect 35938 -641 35972 -607
rect 35564 -1470 35598 -1436
rect 44156 -1883 44162 -1852
rect 44162 -1883 44190 -1852
rect 44228 -1883 44230 -1852
rect 44230 -1883 44262 -1852
rect 44300 -1883 44332 -1852
rect 44332 -1883 44334 -1852
rect 44372 -1883 44400 -1852
rect 44400 -1883 44406 -1852
rect 44156 -1886 44190 -1883
rect 44228 -1886 44262 -1883
rect 44300 -1886 44334 -1883
rect 44372 -1886 44406 -1883
rect 44156 -2261 44190 -2258
rect 44228 -2261 44262 -2258
rect 44300 -2261 44334 -2258
rect 44372 -2261 44406 -2258
rect 44156 -2292 44162 -2261
rect 44162 -2292 44190 -2261
rect 44228 -2292 44230 -2261
rect 44230 -2292 44262 -2261
rect 44300 -2292 44332 -2261
rect 44332 -2292 44334 -2261
rect 44372 -2292 44400 -2261
rect 44400 -2292 44406 -2261
rect 35347 -2896 35381 -2862
rect 35427 -2896 35461 -2862
rect 35507 -2896 35541 -2862
rect 35587 -2896 35621 -2862
rect 35667 -2896 35701 -2862
rect 35747 -2896 35781 -2862
rect 35827 -2896 35861 -2862
rect 35907 -2896 35941 -2862
rect 35987 -2896 36021 -2862
rect 36067 -2896 36101 -2862
rect 36147 -2896 36181 -2862
rect 36227 -2896 36261 -2862
rect 36307 -2896 36341 -2862
rect 36387 -2896 36421 -2862
rect 36467 -2896 36501 -2862
rect 36547 -2896 36581 -2862
rect 36627 -2896 36661 -2862
rect 36707 -2896 36741 -2862
rect 36787 -2896 36821 -2862
rect 36867 -2896 36901 -2862
rect 36947 -2896 36981 -2862
rect 37027 -2896 37061 -2862
rect 37107 -2896 37141 -2862
rect 37187 -2896 37221 -2862
rect 37267 -2896 37301 -2862
rect 37347 -2896 37381 -2862
rect 37427 -2896 37461 -2862
rect 37507 -2896 37541 -2862
rect 37587 -2896 37621 -2862
rect 37667 -2896 37701 -2862
rect 37747 -2896 37781 -2862
rect 37827 -2896 37861 -2862
rect 37907 -2896 37941 -2862
rect 37987 -2896 38021 -2862
rect 38067 -2896 38101 -2862
rect 38147 -2896 38181 -2862
rect 38227 -2896 38261 -2862
rect 38307 -2896 38341 -2862
rect 38387 -2896 38421 -2862
rect 38467 -2896 38501 -2862
rect 38547 -2896 38581 -2862
rect 38627 -2896 38661 -2862
rect 38707 -2896 38741 -2862
rect 38787 -2896 38821 -2862
rect 38867 -2896 38901 -2862
rect 38947 -2896 38981 -2862
rect 39027 -2896 39061 -2862
rect 39107 -2896 39141 -2862
rect 39188 -2896 39222 -2862
rect 39268 -2896 39302 -2862
rect 39348 -2896 39382 -2862
rect 39428 -2896 39462 -2862
rect 39508 -2896 39542 -2862
rect 39588 -2896 39622 -2862
rect 39668 -2896 39702 -2862
rect 39748 -2896 39782 -2862
rect 39828 -2896 39862 -2862
rect 39908 -2896 39942 -2862
rect 39988 -2896 40022 -2862
rect 40068 -2896 40102 -2862
rect 40148 -2896 40182 -2862
rect 40228 -2896 40262 -2862
rect 40308 -2896 40342 -2862
rect 40388 -2896 40422 -2862
rect 40468 -2896 40502 -2862
rect 40548 -2896 40582 -2862
rect 40628 -2896 40662 -2862
rect 40708 -2896 40742 -2862
rect 40788 -2896 40822 -2862
rect 40868 -2896 40902 -2862
rect 40948 -2896 40982 -2862
rect 41028 -2896 41062 -2862
rect 41108 -2896 41142 -2862
rect 41188 -2896 41222 -2862
rect 41268 -2896 41302 -2862
rect 41348 -2896 41382 -2862
rect 41428 -2896 41462 -2862
rect 41508 -2896 41542 -2862
rect 41588 -2896 41622 -2862
rect 41668 -2896 41702 -2862
rect 41748 -2896 41782 -2862
rect 41828 -2896 41862 -2862
rect 41908 -2896 41942 -2862
rect 41988 -2896 42022 -2862
rect 42068 -2896 42102 -2862
rect 42148 -2896 42182 -2862
rect 42228 -2896 42262 -2862
rect 42308 -2896 42342 -2862
rect 42388 -2896 42422 -2862
rect 42468 -2896 42502 -2862
rect 42548 -2896 42582 -2862
rect 42628 -2896 42662 -2862
rect 42708 -2896 42742 -2862
rect 42788 -2896 42822 -2862
rect 42868 -2896 42902 -2862
rect 42948 -2896 42982 -2862
rect 43028 -2896 43062 -2862
rect 43108 -2896 43142 -2862
rect 43188 -2896 43222 -2862
rect 43268 -2896 43302 -2862
rect 43348 -2896 43382 -2862
rect 43428 -2896 43462 -2862
rect 43508 -2896 43542 -2862
rect 43588 -2896 43622 -2862
rect 43668 -2896 43702 -2862
rect 43748 -2896 43782 -2862
rect 43828 -2896 43862 -2862
rect 43908 -2896 43942 -2862
rect 43988 -2896 44022 -2862
rect 44068 -2896 44102 -2862
rect 44148 -2896 44182 -2862
rect 44228 -2896 44262 -2862
rect 44308 -2896 44342 -2862
rect 44388 -2896 44422 -2862
rect 44468 -2896 44502 -2862
rect 44548 -2896 44582 -2862
rect 44628 -2896 44662 -2862
rect 44708 -2896 44742 -2862
rect 44788 -2896 44822 -2862
rect 44868 -2896 44902 -2862
rect 44948 -2896 44982 -2862
rect 45028 -2896 45062 -2862
rect 45108 -2896 45142 -2862
rect 45188 -2896 45222 -2862
rect 45268 -2896 45302 -2862
rect 45348 -2896 45382 -2862
rect 45428 -2896 45462 -2862
rect 45508 -2896 45542 -2862
rect 45588 -2896 45622 -2862
rect 45668 -2896 45702 -2862
rect 45748 -2896 45782 -2862
rect 45828 -2896 45862 -2862
rect 45908 -2896 45942 -2862
rect 45988 -2896 46022 -2862
rect 46068 -2896 46102 -2862
rect 46148 -2896 46182 -2862
rect 46228 -2896 46262 -2862
rect 46308 -2896 46342 -2862
rect 46388 -2896 46422 -2862
rect 46468 -2896 46502 -2862
rect 46548 -2896 46582 -2862
rect 46628 -2896 46662 -2862
rect 46708 -2896 46742 -2862
rect 46788 -2896 46822 -2862
rect 46868 -2896 46902 -2862
rect 46948 -2896 46982 -2862
rect 47028 -2896 47062 -2862
rect 47108 -2896 47142 -2862
rect 47188 -2896 47222 -2862
rect 47268 -2896 47302 -2862
rect 47349 -2896 47383 -2862
rect 47429 -2896 47463 -2862
rect 47509 -2896 47543 -2862
rect 47589 -2896 47623 -2862
rect 47669 -2896 47703 -2862
rect 47749 -2896 47783 -2862
rect 47829 -2896 47863 -2862
rect 47909 -2896 47943 -2862
rect 47989 -2896 48023 -2862
rect 48069 -2896 48103 -2862
rect 48149 -2896 48183 -2862
rect 48229 -2896 48263 -2862
rect 48309 -2896 48343 -2862
rect 48389 -2896 48423 -2862
rect 48469 -2896 48503 -2862
rect 48549 -2896 48583 -2862
rect 48629 -2896 48663 -2862
rect 48709 -2896 48743 -2862
rect 48789 -2896 48823 -2862
rect 48869 -2896 48903 -2862
rect 48949 -2896 48983 -2862
rect 49029 -2896 49063 -2862
rect 49109 -2896 49143 -2862
rect 49189 -2896 49223 -2862
rect 49269 -2896 49303 -2862
rect 49349 -2896 49383 -2862
rect 49429 -2896 49463 -2862
rect 49509 -2896 49543 -2862
rect 49589 -2896 49623 -2862
rect 49669 -2896 49703 -2862
rect 49749 -2896 49783 -2862
rect 49829 -2896 49863 -2862
rect 49909 -2896 49943 -2862
rect 49989 -2896 50023 -2862
rect 50069 -2896 50103 -2862
rect 50149 -2896 50183 -2862
rect 50229 -2896 50263 -2862
rect 50309 -2896 50343 -2862
rect 50389 -2896 50423 -2862
rect 50469 -2896 50503 -2862
rect 50549 -2896 50583 -2862
rect 50629 -2896 50663 -2862
rect 50709 -2896 50743 -2862
rect 50789 -2896 50823 -2862
rect 50869 -2896 50903 -2862
rect 50949 -2896 50983 -2862
rect 51029 -2896 51063 -2862
rect 51109 -2896 51143 -2862
rect 51189 -2896 51223 -2862
rect 51269 -2896 51303 -2862
rect 51349 -2896 51383 -2862
rect 51429 -2896 51463 -2862
rect 51509 -2896 51543 -2862
rect 51589 -2896 51623 -2862
rect 35347 -2986 35381 -2952
rect 35427 -2986 35461 -2952
rect 35507 -2986 35541 -2952
rect 35587 -2986 35621 -2952
rect 35667 -2986 35701 -2952
rect 35747 -2986 35781 -2952
rect 35827 -2986 35861 -2952
rect 35907 -2986 35941 -2952
rect 35987 -2986 36021 -2952
rect 36067 -2986 36101 -2952
rect 36147 -2986 36181 -2952
rect 36227 -2986 36261 -2952
rect 36307 -2986 36341 -2952
rect 36387 -2986 36421 -2952
rect 36467 -2986 36501 -2952
rect 36547 -2986 36581 -2952
rect 36627 -2986 36661 -2952
rect 36707 -2986 36741 -2952
rect 36787 -2986 36821 -2952
rect 36867 -2986 36901 -2952
rect 36947 -2986 36981 -2952
rect 37027 -2986 37061 -2952
rect 37107 -2986 37141 -2952
rect 37187 -2986 37221 -2952
rect 37267 -2986 37301 -2952
rect 37347 -2986 37381 -2952
rect 37427 -2986 37461 -2952
rect 37507 -2986 37541 -2952
rect 37587 -2986 37621 -2952
rect 37667 -2986 37701 -2952
rect 37747 -2986 37781 -2952
rect 37827 -2986 37861 -2952
rect 37907 -2986 37941 -2952
rect 37987 -2986 38021 -2952
rect 38067 -2986 38101 -2952
rect 38147 -2986 38181 -2952
rect 38227 -2986 38261 -2952
rect 38307 -2986 38341 -2952
rect 38387 -2986 38421 -2952
rect 38467 -2986 38501 -2952
rect 38547 -2986 38581 -2952
rect 38627 -2986 38661 -2952
rect 38707 -2986 38741 -2952
rect 38787 -2986 38821 -2952
rect 38867 -2986 38901 -2952
rect 38947 -2986 38981 -2952
rect 39027 -2986 39061 -2952
rect 39107 -2986 39141 -2952
rect 39188 -2986 39222 -2952
rect 39268 -2986 39302 -2952
rect 39348 -2986 39382 -2952
rect 39428 -2986 39462 -2952
rect 39508 -2986 39542 -2952
rect 39588 -2986 39622 -2952
rect 39668 -2986 39702 -2952
rect 39748 -2986 39782 -2952
rect 39828 -2986 39862 -2952
rect 39908 -2986 39942 -2952
rect 39988 -2986 40022 -2952
rect 40068 -2986 40102 -2952
rect 40148 -2986 40182 -2952
rect 40228 -2986 40262 -2952
rect 40308 -2986 40342 -2952
rect 40388 -2986 40422 -2952
rect 40468 -2986 40502 -2952
rect 40548 -2986 40582 -2952
rect 40628 -2986 40662 -2952
rect 40708 -2986 40742 -2952
rect 40788 -2986 40822 -2952
rect 40868 -2986 40902 -2952
rect 40948 -2986 40982 -2952
rect 41028 -2986 41062 -2952
rect 41108 -2986 41142 -2952
rect 41188 -2986 41222 -2952
rect 41268 -2986 41302 -2952
rect 41348 -2986 41382 -2952
rect 41428 -2986 41462 -2952
rect 41508 -2986 41542 -2952
rect 41588 -2986 41622 -2952
rect 41668 -2986 41702 -2952
rect 41748 -2986 41782 -2952
rect 41828 -2986 41862 -2952
rect 41908 -2986 41942 -2952
rect 41988 -2986 42022 -2952
rect 42068 -2986 42102 -2952
rect 42148 -2986 42182 -2952
rect 42228 -2986 42262 -2952
rect 42308 -2986 42342 -2952
rect 42388 -2986 42422 -2952
rect 42468 -2986 42502 -2952
rect 42548 -2986 42582 -2952
rect 42628 -2986 42662 -2952
rect 42708 -2986 42742 -2952
rect 42788 -2986 42822 -2952
rect 42868 -2986 42902 -2952
rect 42948 -2986 42982 -2952
rect 43028 -2986 43062 -2952
rect 43108 -2986 43142 -2952
rect 43188 -2986 43222 -2952
rect 43268 -2986 43302 -2952
rect 43348 -2986 43382 -2952
rect 43428 -2986 43462 -2952
rect 43508 -2986 43542 -2952
rect 43588 -2986 43622 -2952
rect 43668 -2986 43702 -2952
rect 43748 -2986 43782 -2952
rect 43828 -2986 43862 -2952
rect 43908 -2986 43942 -2952
rect 43988 -2986 44022 -2952
rect 44068 -2986 44102 -2952
rect 44148 -2986 44182 -2952
rect 44228 -2986 44262 -2952
rect 44308 -2986 44342 -2952
rect 44388 -2986 44422 -2952
rect 44468 -2986 44502 -2952
rect 44548 -2986 44582 -2952
rect 44628 -2986 44662 -2952
rect 44708 -2986 44742 -2952
rect 44788 -2986 44822 -2952
rect 44868 -2986 44902 -2952
rect 44948 -2986 44982 -2952
rect 45028 -2986 45062 -2952
rect 45108 -2986 45142 -2952
rect 45188 -2986 45222 -2952
rect 45268 -2986 45302 -2952
rect 45348 -2986 45382 -2952
rect 45428 -2986 45462 -2952
rect 45508 -2986 45542 -2952
rect 45588 -2986 45622 -2952
rect 45668 -2986 45702 -2952
rect 45748 -2986 45782 -2952
rect 45828 -2986 45862 -2952
rect 45908 -2986 45942 -2952
rect 45988 -2986 46022 -2952
rect 46068 -2986 46102 -2952
rect 46148 -2986 46182 -2952
rect 46228 -2986 46262 -2952
rect 46308 -2986 46342 -2952
rect 46388 -2986 46422 -2952
rect 46468 -2986 46502 -2952
rect 46548 -2986 46582 -2952
rect 46628 -2986 46662 -2952
rect 46708 -2986 46742 -2952
rect 46788 -2986 46822 -2952
rect 46868 -2986 46902 -2952
rect 46948 -2986 46982 -2952
rect 47028 -2986 47062 -2952
rect 47108 -2986 47142 -2952
rect 47188 -2986 47222 -2952
rect 47268 -2986 47302 -2952
rect 47349 -2986 47383 -2952
rect 47429 -2986 47463 -2952
rect 47509 -2986 47543 -2952
rect 47589 -2986 47623 -2952
rect 47669 -2986 47703 -2952
rect 47749 -2986 47783 -2952
rect 47829 -2986 47863 -2952
rect 47909 -2986 47943 -2952
rect 47989 -2986 48023 -2952
rect 48069 -2986 48103 -2952
rect 48149 -2986 48183 -2952
rect 48229 -2986 48263 -2952
rect 48309 -2986 48343 -2952
rect 48389 -2986 48423 -2952
rect 48469 -2986 48503 -2952
rect 48549 -2986 48583 -2952
rect 48629 -2986 48663 -2952
rect 48709 -2986 48743 -2952
rect 48789 -2986 48823 -2952
rect 48869 -2986 48903 -2952
rect 48949 -2986 48983 -2952
rect 49029 -2986 49063 -2952
rect 49109 -2986 49143 -2952
rect 49189 -2986 49223 -2952
rect 49269 -2986 49303 -2952
rect 49349 -2986 49383 -2952
rect 49429 -2986 49463 -2952
rect 49509 -2986 49543 -2952
rect 49589 -2986 49623 -2952
rect 49669 -2986 49703 -2952
rect 49749 -2986 49783 -2952
rect 49829 -2986 49863 -2952
rect 49909 -2986 49943 -2952
rect 49989 -2986 50023 -2952
rect 50069 -2986 50103 -2952
rect 50149 -2986 50183 -2952
rect 50229 -2986 50263 -2952
rect 50309 -2986 50343 -2952
rect 50389 -2986 50423 -2952
rect 50469 -2986 50503 -2952
rect 50549 -2986 50583 -2952
rect 50629 -2986 50663 -2952
rect 50709 -2986 50743 -2952
rect 50789 -2986 50823 -2952
rect 50869 -2986 50903 -2952
rect 50949 -2986 50983 -2952
rect 51029 -2986 51063 -2952
rect 51109 -2986 51143 -2952
rect 51189 -2986 51223 -2952
rect 51269 -2986 51303 -2952
rect 51349 -2986 51383 -2952
rect 51429 -2986 51463 -2952
rect 51509 -2986 51543 -2952
rect 51589 -2986 51623 -2952
rect 39483 -3107 39517 -3073
rect 39603 -3107 39637 -3073
rect 39483 -3227 39517 -3193
rect 39603 -3227 39637 -3193
<< metal1 >>
rect 39402 9747 39662 9791
rect 39402 9695 39446 9747
rect 39498 9695 39566 9747
rect 39618 9695 39662 9747
rect 39402 9627 39662 9695
rect 39402 9575 39446 9627
rect 39498 9575 39566 9627
rect 39618 9575 39662 9627
rect 39402 9531 39662 9575
rect 27940 2674 43396 2706
rect 27940 2640 27949 2674
rect 27983 2640 28029 2674
rect 28063 2640 28109 2674
rect 28143 2640 28189 2674
rect 28223 2640 28269 2674
rect 28303 2640 28349 2674
rect 28383 2640 28429 2674
rect 28463 2640 28509 2674
rect 28543 2640 28589 2674
rect 28623 2640 28669 2674
rect 28703 2640 28749 2674
rect 28783 2640 28829 2674
rect 28863 2640 28909 2674
rect 28943 2640 28989 2674
rect 29023 2640 29069 2674
rect 29103 2640 29149 2674
rect 29183 2640 29229 2674
rect 29263 2640 29309 2674
rect 29343 2640 29389 2674
rect 29423 2640 29469 2674
rect 29503 2640 29549 2674
rect 29583 2640 29629 2674
rect 29663 2640 29709 2674
rect 29743 2640 29789 2674
rect 29823 2640 29869 2674
rect 29903 2640 29949 2674
rect 29983 2640 30029 2674
rect 30063 2640 30109 2674
rect 30143 2640 30189 2674
rect 30223 2640 30269 2674
rect 30303 2640 30349 2674
rect 30383 2640 30429 2674
rect 30463 2640 30509 2674
rect 30543 2640 30589 2674
rect 30623 2640 30669 2674
rect 30703 2640 30749 2674
rect 30783 2640 30829 2674
rect 30863 2640 30910 2674
rect 30944 2640 30990 2674
rect 31024 2640 31070 2674
rect 31104 2640 31150 2674
rect 31184 2640 31230 2674
rect 31264 2640 31310 2674
rect 31344 2640 31390 2674
rect 31424 2640 31470 2674
rect 31504 2640 31550 2674
rect 31584 2640 31630 2674
rect 31664 2640 31710 2674
rect 31744 2640 31790 2674
rect 31824 2640 31870 2674
rect 31904 2640 31950 2674
rect 31984 2640 32030 2674
rect 32064 2640 32110 2674
rect 32144 2640 32190 2674
rect 32224 2640 32270 2674
rect 32304 2640 32350 2674
rect 32384 2640 32430 2674
rect 32464 2640 32510 2674
rect 32544 2640 32590 2674
rect 32624 2640 32670 2674
rect 32704 2640 32750 2674
rect 32784 2640 32830 2674
rect 32864 2640 32910 2674
rect 32944 2640 32990 2674
rect 33024 2640 33070 2674
rect 33104 2640 33150 2674
rect 33184 2640 33230 2674
rect 33264 2640 33310 2674
rect 33344 2640 33390 2674
rect 33424 2640 33470 2674
rect 33504 2640 33550 2674
rect 33584 2640 33630 2674
rect 33664 2640 33710 2674
rect 33744 2640 33790 2674
rect 33824 2640 33870 2674
rect 33904 2640 33950 2674
rect 33984 2640 34030 2674
rect 34064 2640 34110 2674
rect 34144 2640 34190 2674
rect 34224 2640 34270 2674
rect 34304 2640 34350 2674
rect 34384 2640 34430 2674
rect 34464 2640 34510 2674
rect 34544 2640 34590 2674
rect 34624 2640 34670 2674
rect 34704 2640 34750 2674
rect 34784 2640 34830 2674
rect 34864 2640 34910 2674
rect 34944 2640 34990 2674
rect 35024 2640 35070 2674
rect 35104 2640 35150 2674
rect 35184 2640 35242 2674
rect 35276 2640 35322 2674
rect 35356 2640 35402 2674
rect 35436 2640 35482 2674
rect 35516 2640 35562 2674
rect 35596 2640 35642 2674
rect 35676 2640 35722 2674
rect 35756 2640 35802 2674
rect 35836 2640 35882 2674
rect 35916 2640 35962 2674
rect 35996 2640 36042 2674
rect 36076 2640 36122 2674
rect 36156 2640 36202 2674
rect 36236 2640 36282 2674
rect 36316 2640 36362 2674
rect 36396 2640 36442 2674
rect 36476 2640 36522 2674
rect 36556 2640 36602 2674
rect 36636 2640 36682 2674
rect 36716 2640 36762 2674
rect 36796 2640 36842 2674
rect 36876 2640 36922 2674
rect 36956 2640 37002 2674
rect 37036 2640 37082 2674
rect 37116 2640 37162 2674
rect 37196 2640 37242 2674
rect 37276 2640 37322 2674
rect 37356 2640 37402 2674
rect 37436 2640 37482 2674
rect 37516 2640 37562 2674
rect 37596 2640 37642 2674
rect 37676 2640 37722 2674
rect 37756 2640 37802 2674
rect 37836 2640 37882 2674
rect 37916 2640 37962 2674
rect 37996 2640 38042 2674
rect 38076 2640 38122 2674
rect 38156 2640 38202 2674
rect 38236 2640 38282 2674
rect 38316 2640 38362 2674
rect 38396 2640 38442 2674
rect 38476 2640 38522 2674
rect 38556 2640 38602 2674
rect 38636 2640 38682 2674
rect 38716 2640 38762 2674
rect 38796 2640 38842 2674
rect 38876 2640 38922 2674
rect 38956 2640 39002 2674
rect 39036 2640 39083 2674
rect 39117 2640 39163 2674
rect 39197 2640 39243 2674
rect 39277 2640 39323 2674
rect 39357 2640 39403 2674
rect 39437 2640 39483 2674
rect 39517 2640 39563 2674
rect 39597 2640 39643 2674
rect 39677 2640 39723 2674
rect 39757 2640 39803 2674
rect 39837 2640 39883 2674
rect 39917 2640 39963 2674
rect 39997 2640 40043 2674
rect 40077 2640 40123 2674
rect 40157 2640 40203 2674
rect 40237 2640 40283 2674
rect 40317 2640 40363 2674
rect 40397 2640 40443 2674
rect 40477 2640 40523 2674
rect 40557 2640 40603 2674
rect 40637 2640 40683 2674
rect 40717 2640 40763 2674
rect 40797 2640 40843 2674
rect 40877 2640 40923 2674
rect 40957 2640 41003 2674
rect 41037 2640 41083 2674
rect 41117 2640 41163 2674
rect 41197 2640 41243 2674
rect 41277 2640 41323 2674
rect 41357 2640 41403 2674
rect 41437 2640 41483 2674
rect 41517 2640 41563 2674
rect 41597 2640 41643 2674
rect 41677 2640 41723 2674
rect 41757 2640 41803 2674
rect 41837 2640 41883 2674
rect 41917 2640 41963 2674
rect 41997 2640 42043 2674
rect 42077 2640 42123 2674
rect 42157 2640 42203 2674
rect 42237 2640 42283 2674
rect 42317 2640 42363 2674
rect 42397 2640 42443 2674
rect 42477 2640 42523 2674
rect 42557 2640 42603 2674
rect 42637 2640 42683 2674
rect 42717 2640 42763 2674
rect 42797 2640 42843 2674
rect 42877 2640 42923 2674
rect 42957 2640 43003 2674
rect 43037 2640 43083 2674
rect 43117 2640 43163 2674
rect 43197 2640 43243 2674
rect 43277 2640 43323 2674
rect 43357 2640 43396 2674
rect 27940 2584 43396 2640
rect 27940 2550 27949 2584
rect 27983 2550 28029 2584
rect 28063 2550 28109 2584
rect 28143 2550 28189 2584
rect 28223 2550 28269 2584
rect 28303 2550 28349 2584
rect 28383 2550 28429 2584
rect 28463 2550 28509 2584
rect 28543 2550 28589 2584
rect 28623 2550 28669 2584
rect 28703 2550 28749 2584
rect 28783 2550 28829 2584
rect 28863 2550 28909 2584
rect 28943 2550 28989 2584
rect 29023 2550 29069 2584
rect 29103 2550 29149 2584
rect 29183 2550 29229 2584
rect 29263 2550 29309 2584
rect 29343 2550 29389 2584
rect 29423 2550 29469 2584
rect 29503 2550 29549 2584
rect 29583 2550 29629 2584
rect 29663 2550 29709 2584
rect 29743 2550 29789 2584
rect 29823 2550 29869 2584
rect 29903 2550 29949 2584
rect 29983 2550 30029 2584
rect 30063 2550 30109 2584
rect 30143 2550 30189 2584
rect 30223 2550 30269 2584
rect 30303 2550 30349 2584
rect 30383 2550 30429 2584
rect 30463 2550 30509 2584
rect 30543 2550 30589 2584
rect 30623 2550 30669 2584
rect 30703 2550 30749 2584
rect 30783 2550 30829 2584
rect 30863 2550 30910 2584
rect 30944 2550 30990 2584
rect 31024 2550 31070 2584
rect 31104 2550 31150 2584
rect 31184 2550 31230 2584
rect 31264 2550 31310 2584
rect 31344 2550 31390 2584
rect 31424 2550 31470 2584
rect 31504 2550 31550 2584
rect 31584 2550 31630 2584
rect 31664 2550 31710 2584
rect 31744 2550 31790 2584
rect 31824 2550 31870 2584
rect 31904 2550 31950 2584
rect 31984 2550 32030 2584
rect 32064 2550 32110 2584
rect 32144 2550 32190 2584
rect 32224 2550 32270 2584
rect 32304 2550 32350 2584
rect 32384 2550 32430 2584
rect 32464 2550 32510 2584
rect 32544 2550 32590 2584
rect 32624 2550 32670 2584
rect 32704 2550 32750 2584
rect 32784 2550 32830 2584
rect 32864 2550 32910 2584
rect 32944 2550 32990 2584
rect 33024 2550 33070 2584
rect 33104 2550 33150 2584
rect 33184 2550 33230 2584
rect 33264 2550 33310 2584
rect 33344 2550 33390 2584
rect 33424 2550 33470 2584
rect 33504 2550 33550 2584
rect 33584 2550 33630 2584
rect 33664 2550 33710 2584
rect 33744 2550 33790 2584
rect 33824 2550 33870 2584
rect 33904 2550 33950 2584
rect 33984 2550 34030 2584
rect 34064 2550 34110 2584
rect 34144 2550 34190 2584
rect 34224 2550 34270 2584
rect 34304 2550 34350 2584
rect 34384 2550 34430 2584
rect 34464 2550 34510 2584
rect 34544 2550 34590 2584
rect 34624 2550 34670 2584
rect 34704 2550 34750 2584
rect 34784 2550 34830 2584
rect 34864 2550 34910 2584
rect 34944 2550 34990 2584
rect 35024 2550 35070 2584
rect 35104 2550 35150 2584
rect 35184 2550 35242 2584
rect 35276 2550 35322 2584
rect 35356 2550 35402 2584
rect 35436 2550 35482 2584
rect 35516 2550 35562 2584
rect 35596 2550 35642 2584
rect 35676 2550 35722 2584
rect 35756 2550 35802 2584
rect 35836 2550 35882 2584
rect 35916 2550 35962 2584
rect 35996 2550 36042 2584
rect 36076 2550 36122 2584
rect 36156 2550 36202 2584
rect 36236 2550 36282 2584
rect 36316 2550 36362 2584
rect 36396 2550 36442 2584
rect 36476 2550 36522 2584
rect 36556 2550 36602 2584
rect 36636 2550 36682 2584
rect 36716 2550 36762 2584
rect 36796 2550 36842 2584
rect 36876 2550 36922 2584
rect 36956 2550 37002 2584
rect 37036 2550 37082 2584
rect 37116 2550 37162 2584
rect 37196 2550 37242 2584
rect 37276 2550 37322 2584
rect 37356 2550 37402 2584
rect 37436 2550 37482 2584
rect 37516 2550 37562 2584
rect 37596 2550 37642 2584
rect 37676 2550 37722 2584
rect 37756 2550 37802 2584
rect 37836 2550 37882 2584
rect 37916 2550 37962 2584
rect 37996 2550 38042 2584
rect 38076 2550 38122 2584
rect 38156 2550 38202 2584
rect 38236 2550 38282 2584
rect 38316 2550 38362 2584
rect 38396 2550 38442 2584
rect 38476 2550 38522 2584
rect 38556 2550 38602 2584
rect 38636 2550 38682 2584
rect 38716 2550 38762 2584
rect 38796 2550 38842 2584
rect 38876 2550 38922 2584
rect 38956 2550 39002 2584
rect 39036 2550 39083 2584
rect 39117 2550 39163 2584
rect 39197 2550 39243 2584
rect 39277 2550 39323 2584
rect 39357 2550 39403 2584
rect 39437 2550 39483 2584
rect 39517 2550 39563 2584
rect 39597 2550 39643 2584
rect 39677 2550 39723 2584
rect 39757 2550 39803 2584
rect 39837 2550 39883 2584
rect 39917 2550 39963 2584
rect 39997 2550 40043 2584
rect 40077 2550 40123 2584
rect 40157 2550 40203 2584
rect 40237 2550 40283 2584
rect 40317 2550 40363 2584
rect 40397 2550 40443 2584
rect 40477 2550 40523 2584
rect 40557 2550 40603 2584
rect 40637 2550 40683 2584
rect 40717 2550 40763 2584
rect 40797 2550 40843 2584
rect 40877 2550 40923 2584
rect 40957 2550 41003 2584
rect 41037 2550 41083 2584
rect 41117 2550 41163 2584
rect 41197 2550 41243 2584
rect 41277 2550 41323 2584
rect 41357 2550 41403 2584
rect 41437 2550 41483 2584
rect 41517 2550 41563 2584
rect 41597 2550 41643 2584
rect 41677 2550 41723 2584
rect 41757 2550 41803 2584
rect 41837 2550 41883 2584
rect 41917 2550 41963 2584
rect 41997 2550 42043 2584
rect 42077 2550 42123 2584
rect 42157 2550 42203 2584
rect 42237 2550 42283 2584
rect 42317 2550 42363 2584
rect 42397 2550 42443 2584
rect 42477 2550 42523 2584
rect 42557 2550 42603 2584
rect 42637 2550 42683 2584
rect 42717 2550 42763 2584
rect 42797 2550 42843 2584
rect 42877 2550 42923 2584
rect 42957 2550 43003 2584
rect 43037 2550 43083 2584
rect 43117 2550 43163 2584
rect 43197 2550 43243 2584
rect 43277 2550 43323 2584
rect 43357 2550 43396 2584
rect 27940 2516 43396 2550
rect 32522 1560 32782 1598
rect 32522 1500 32560 1560
rect 32620 1500 32680 1560
rect 32740 1500 32782 1560
rect 32522 1440 32782 1500
rect 32522 1380 32560 1440
rect 32620 1380 32680 1440
rect 32740 1380 32782 1440
rect 32522 1338 32782 1380
rect 32942 1560 33202 1598
rect 32942 1500 32980 1560
rect 33040 1554 33202 1560
rect 33040 1502 33106 1554
rect 33158 1502 33202 1554
rect 33040 1500 33202 1502
rect 32942 1440 33202 1500
rect 32942 1380 32980 1440
rect 33040 1380 33100 1440
rect 33160 1380 33202 1440
rect 32942 1338 33202 1380
rect 34256 1554 34516 1598
rect 34256 1502 34300 1554
rect 34352 1502 34420 1554
rect 34472 1502 34516 1554
rect 34256 1434 34516 1502
rect 34256 1382 34300 1434
rect 34352 1382 34420 1434
rect 34472 1382 34516 1434
rect 34256 1338 34516 1382
rect 34676 1554 34936 1598
rect 34676 1502 34720 1554
rect 34772 1502 34840 1554
rect 34892 1502 34936 1554
rect 34676 1434 34936 1502
rect 34676 1382 34720 1434
rect 34772 1382 34840 1434
rect 34892 1382 34936 1434
rect 34676 1338 34936 1382
rect 32522 1140 32782 1178
rect 32522 1080 32560 1140
rect 32620 1134 32782 1140
rect 32620 1082 32686 1134
rect 32738 1082 32782 1134
rect 32620 1080 32782 1082
rect 32522 1020 32782 1080
rect 32522 960 32560 1020
rect 32620 960 32680 1020
rect 32740 960 32782 1020
rect 32522 918 32782 960
rect 32942 1140 33202 1178
rect 32942 1080 32980 1140
rect 33040 1080 33100 1140
rect 33160 1080 33202 1140
rect 32942 1020 33202 1080
rect 32942 960 32980 1020
rect 33040 960 33100 1020
rect 33160 960 33202 1020
rect 32942 918 33202 960
rect 34256 1134 34516 1178
rect 34256 1082 34300 1134
rect 34352 1082 34420 1134
rect 34472 1082 34516 1134
rect 34256 1014 34516 1082
rect 34256 962 34300 1014
rect 34352 962 34420 1014
rect 34472 962 34516 1014
rect 34256 918 34516 962
rect 34676 1134 34936 1178
rect 34676 1082 34720 1134
rect 34772 1082 34840 1134
rect 34892 1082 34936 1134
rect 34676 1014 34936 1082
rect 34676 962 34720 1014
rect 34772 962 34840 1014
rect 34892 962 34936 1014
rect 34676 918 34936 962
rect 44172 2 44432 3
rect 44172 -32 44433 2
rect 44172 -35 44218 -32
rect 44172 -87 44214 -35
rect 44270 -35 44338 -32
rect 44270 -84 44334 -35
rect 44390 -84 44433 -32
rect 44269 -87 44334 -84
rect 44172 -94 44217 -87
rect 44269 -94 44337 -87
rect 44389 -94 44433 -84
rect 44172 -152 44433 -94
rect 44172 -155 44218 -152
rect 44172 -207 44214 -155
rect 44270 -155 44338 -152
rect 44270 -204 44334 -155
rect 44390 -204 44433 -152
rect 44269 -207 44334 -204
rect 44172 -214 44217 -207
rect 44269 -214 44337 -207
rect 44389 -214 44433 -204
rect 44172 -257 44433 -214
rect 44173 -258 44433 -257
rect 35765 -478 36025 -434
rect 35765 -530 35809 -478
rect 35861 -530 35929 -478
rect 35981 -530 36025 -478
rect 35765 -598 36025 -530
rect 35765 -650 35809 -598
rect 35861 -650 35929 -598
rect 35981 -650 36025 -598
rect 35765 -694 36025 -650
rect 35541 -1436 35621 -1413
rect 35541 -1470 35564 -1436
rect 35598 -1470 35621 -1436
rect 35541 -1493 35621 -1470
rect 44196 -1752 44396 -258
rect 44149 -1843 44409 -1752
rect 44125 -1852 44437 -1843
rect 44125 -1886 44156 -1852
rect 44190 -1886 44228 -1852
rect 44262 -1886 44300 -1852
rect 44334 -1886 44372 -1852
rect 44406 -1886 44437 -1852
rect 44125 -1895 44437 -1886
rect 44125 -2258 44437 -2249
rect 44125 -2292 44156 -2258
rect 44190 -2292 44228 -2258
rect 44262 -2292 44300 -2258
rect 44334 -2292 44372 -2258
rect 44406 -2292 44437 -2258
rect 44125 -2301 44437 -2292
rect 44152 -2830 44412 -2301
rect 35312 -2862 51662 -2830
rect 35312 -2896 35347 -2862
rect 35381 -2896 35427 -2862
rect 35461 -2896 35507 -2862
rect 35541 -2896 35587 -2862
rect 35621 -2896 35667 -2862
rect 35701 -2896 35747 -2862
rect 35781 -2896 35827 -2862
rect 35861 -2896 35907 -2862
rect 35941 -2896 35987 -2862
rect 36021 -2896 36067 -2862
rect 36101 -2896 36147 -2862
rect 36181 -2896 36227 -2862
rect 36261 -2896 36307 -2862
rect 36341 -2896 36387 -2862
rect 36421 -2896 36467 -2862
rect 36501 -2896 36547 -2862
rect 36581 -2896 36627 -2862
rect 36661 -2896 36707 -2862
rect 36741 -2896 36787 -2862
rect 36821 -2896 36867 -2862
rect 36901 -2896 36947 -2862
rect 36981 -2896 37027 -2862
rect 37061 -2896 37107 -2862
rect 37141 -2896 37187 -2862
rect 37221 -2896 37267 -2862
rect 37301 -2896 37347 -2862
rect 37381 -2896 37427 -2862
rect 37461 -2896 37507 -2862
rect 37541 -2896 37587 -2862
rect 37621 -2896 37667 -2862
rect 37701 -2896 37747 -2862
rect 37781 -2896 37827 -2862
rect 37861 -2896 37907 -2862
rect 37941 -2896 37987 -2862
rect 38021 -2896 38067 -2862
rect 38101 -2896 38147 -2862
rect 38181 -2896 38227 -2862
rect 38261 -2896 38307 -2862
rect 38341 -2896 38387 -2862
rect 38421 -2896 38467 -2862
rect 38501 -2896 38547 -2862
rect 38581 -2896 38627 -2862
rect 38661 -2896 38707 -2862
rect 38741 -2896 38787 -2862
rect 38821 -2896 38867 -2862
rect 38901 -2896 38947 -2862
rect 38981 -2896 39027 -2862
rect 39061 -2896 39107 -2862
rect 39141 -2896 39188 -2862
rect 39222 -2896 39268 -2862
rect 39302 -2896 39348 -2862
rect 39382 -2896 39428 -2862
rect 39462 -2896 39508 -2862
rect 39542 -2896 39588 -2862
rect 39622 -2896 39668 -2862
rect 39702 -2896 39748 -2862
rect 39782 -2896 39828 -2862
rect 39862 -2896 39908 -2862
rect 39942 -2896 39988 -2862
rect 40022 -2896 40068 -2862
rect 40102 -2896 40148 -2862
rect 40182 -2896 40228 -2862
rect 40262 -2896 40308 -2862
rect 40342 -2896 40388 -2862
rect 40422 -2896 40468 -2862
rect 40502 -2896 40548 -2862
rect 40582 -2896 40628 -2862
rect 40662 -2896 40708 -2862
rect 40742 -2896 40788 -2862
rect 40822 -2896 40868 -2862
rect 40902 -2896 40948 -2862
rect 40982 -2896 41028 -2862
rect 41062 -2896 41108 -2862
rect 41142 -2896 41188 -2862
rect 41222 -2896 41268 -2862
rect 41302 -2896 41348 -2862
rect 41382 -2896 41428 -2862
rect 41462 -2896 41508 -2862
rect 41542 -2896 41588 -2862
rect 41622 -2896 41668 -2862
rect 41702 -2896 41748 -2862
rect 41782 -2896 41828 -2862
rect 41862 -2896 41908 -2862
rect 41942 -2896 41988 -2862
rect 42022 -2896 42068 -2862
rect 42102 -2896 42148 -2862
rect 42182 -2896 42228 -2862
rect 42262 -2896 42308 -2862
rect 42342 -2896 42388 -2862
rect 42422 -2896 42468 -2862
rect 42502 -2896 42548 -2862
rect 42582 -2896 42628 -2862
rect 42662 -2896 42708 -2862
rect 42742 -2896 42788 -2862
rect 42822 -2896 42868 -2862
rect 42902 -2896 42948 -2862
rect 42982 -2896 43028 -2862
rect 43062 -2896 43108 -2862
rect 43142 -2896 43188 -2862
rect 43222 -2896 43268 -2862
rect 43302 -2896 43348 -2862
rect 43382 -2896 43428 -2862
rect 43462 -2896 43508 -2862
rect 43542 -2896 43588 -2862
rect 43622 -2896 43668 -2862
rect 43702 -2896 43748 -2862
rect 43782 -2896 43828 -2862
rect 43862 -2896 43908 -2862
rect 43942 -2896 43988 -2862
rect 44022 -2896 44068 -2862
rect 44102 -2896 44148 -2862
rect 44182 -2896 44228 -2862
rect 44262 -2896 44308 -2862
rect 44342 -2896 44388 -2862
rect 44422 -2896 44468 -2862
rect 44502 -2896 44548 -2862
rect 44582 -2896 44628 -2862
rect 44662 -2896 44708 -2862
rect 44742 -2896 44788 -2862
rect 44822 -2896 44868 -2862
rect 44902 -2896 44948 -2862
rect 44982 -2896 45028 -2862
rect 45062 -2896 45108 -2862
rect 45142 -2896 45188 -2862
rect 45222 -2896 45268 -2862
rect 45302 -2896 45348 -2862
rect 45382 -2896 45428 -2862
rect 45462 -2896 45508 -2862
rect 45542 -2896 45588 -2862
rect 45622 -2896 45668 -2862
rect 45702 -2896 45748 -2862
rect 45782 -2896 45828 -2862
rect 45862 -2896 45908 -2862
rect 45942 -2896 45988 -2862
rect 46022 -2896 46068 -2862
rect 46102 -2896 46148 -2862
rect 46182 -2896 46228 -2862
rect 46262 -2896 46308 -2862
rect 46342 -2896 46388 -2862
rect 46422 -2896 46468 -2862
rect 46502 -2896 46548 -2862
rect 46582 -2896 46628 -2862
rect 46662 -2896 46708 -2862
rect 46742 -2896 46788 -2862
rect 46822 -2896 46868 -2862
rect 46902 -2896 46948 -2862
rect 46982 -2896 47028 -2862
rect 47062 -2896 47108 -2862
rect 47142 -2896 47188 -2862
rect 47222 -2896 47268 -2862
rect 47302 -2896 47349 -2862
rect 47383 -2896 47429 -2862
rect 47463 -2896 47509 -2862
rect 47543 -2896 47589 -2862
rect 47623 -2896 47669 -2862
rect 47703 -2896 47749 -2862
rect 47783 -2896 47829 -2862
rect 47863 -2896 47909 -2862
rect 47943 -2896 47989 -2862
rect 48023 -2896 48069 -2862
rect 48103 -2896 48149 -2862
rect 48183 -2896 48229 -2862
rect 48263 -2896 48309 -2862
rect 48343 -2896 48389 -2862
rect 48423 -2896 48469 -2862
rect 48503 -2896 48549 -2862
rect 48583 -2896 48629 -2862
rect 48663 -2896 48709 -2862
rect 48743 -2896 48789 -2862
rect 48823 -2896 48869 -2862
rect 48903 -2896 48949 -2862
rect 48983 -2896 49029 -2862
rect 49063 -2896 49109 -2862
rect 49143 -2896 49189 -2862
rect 49223 -2896 49269 -2862
rect 49303 -2896 49349 -2862
rect 49383 -2896 49429 -2862
rect 49463 -2896 49509 -2862
rect 49543 -2896 49589 -2862
rect 49623 -2896 49669 -2862
rect 49703 -2896 49749 -2862
rect 49783 -2896 49829 -2862
rect 49863 -2896 49909 -2862
rect 49943 -2896 49989 -2862
rect 50023 -2896 50069 -2862
rect 50103 -2896 50149 -2862
rect 50183 -2896 50229 -2862
rect 50263 -2896 50309 -2862
rect 50343 -2896 50389 -2862
rect 50423 -2896 50469 -2862
rect 50503 -2896 50549 -2862
rect 50583 -2896 50629 -2862
rect 50663 -2896 50709 -2862
rect 50743 -2896 50789 -2862
rect 50823 -2896 50869 -2862
rect 50903 -2896 50949 -2862
rect 50983 -2896 51029 -2862
rect 51063 -2896 51109 -2862
rect 51143 -2896 51189 -2862
rect 51223 -2896 51269 -2862
rect 51303 -2896 51349 -2862
rect 51383 -2896 51429 -2862
rect 51463 -2896 51509 -2862
rect 51543 -2896 51589 -2862
rect 51623 -2896 51662 -2862
rect 35312 -2952 51662 -2896
rect 35312 -2986 35347 -2952
rect 35381 -2986 35427 -2952
rect 35461 -2986 35507 -2952
rect 35541 -2986 35587 -2952
rect 35621 -2986 35667 -2952
rect 35701 -2986 35747 -2952
rect 35781 -2986 35827 -2952
rect 35861 -2986 35907 -2952
rect 35941 -2986 35987 -2952
rect 36021 -2986 36067 -2952
rect 36101 -2986 36147 -2952
rect 36181 -2986 36227 -2952
rect 36261 -2986 36307 -2952
rect 36341 -2986 36387 -2952
rect 36421 -2986 36467 -2952
rect 36501 -2986 36547 -2952
rect 36581 -2986 36627 -2952
rect 36661 -2986 36707 -2952
rect 36741 -2986 36787 -2952
rect 36821 -2986 36867 -2952
rect 36901 -2986 36947 -2952
rect 36981 -2986 37027 -2952
rect 37061 -2986 37107 -2952
rect 37141 -2986 37187 -2952
rect 37221 -2986 37267 -2952
rect 37301 -2986 37347 -2952
rect 37381 -2986 37427 -2952
rect 37461 -2986 37507 -2952
rect 37541 -2986 37587 -2952
rect 37621 -2986 37667 -2952
rect 37701 -2986 37747 -2952
rect 37781 -2986 37827 -2952
rect 37861 -2986 37907 -2952
rect 37941 -2986 37987 -2952
rect 38021 -2986 38067 -2952
rect 38101 -2986 38147 -2952
rect 38181 -2986 38227 -2952
rect 38261 -2986 38307 -2952
rect 38341 -2986 38387 -2952
rect 38421 -2986 38467 -2952
rect 38501 -2986 38547 -2952
rect 38581 -2986 38627 -2952
rect 38661 -2986 38707 -2952
rect 38741 -2986 38787 -2952
rect 38821 -2986 38867 -2952
rect 38901 -2986 38947 -2952
rect 38981 -2986 39027 -2952
rect 39061 -2986 39107 -2952
rect 39141 -2986 39188 -2952
rect 39222 -2986 39268 -2952
rect 39302 -2986 39348 -2952
rect 39382 -2986 39428 -2952
rect 39462 -2986 39508 -2952
rect 39542 -2986 39588 -2952
rect 39622 -2986 39668 -2952
rect 39702 -2986 39748 -2952
rect 39782 -2986 39828 -2952
rect 39862 -2986 39908 -2952
rect 39942 -2986 39988 -2952
rect 40022 -2986 40068 -2952
rect 40102 -2986 40148 -2952
rect 40182 -2986 40228 -2952
rect 40262 -2986 40308 -2952
rect 40342 -2986 40388 -2952
rect 40422 -2986 40468 -2952
rect 40502 -2986 40548 -2952
rect 40582 -2986 40628 -2952
rect 40662 -2986 40708 -2952
rect 40742 -2986 40788 -2952
rect 40822 -2986 40868 -2952
rect 40902 -2986 40948 -2952
rect 40982 -2986 41028 -2952
rect 41062 -2986 41108 -2952
rect 41142 -2986 41188 -2952
rect 41222 -2986 41268 -2952
rect 41302 -2986 41348 -2952
rect 41382 -2986 41428 -2952
rect 41462 -2986 41508 -2952
rect 41542 -2986 41588 -2952
rect 41622 -2986 41668 -2952
rect 41702 -2986 41748 -2952
rect 41782 -2986 41828 -2952
rect 41862 -2986 41908 -2952
rect 41942 -2986 41988 -2952
rect 42022 -2986 42068 -2952
rect 42102 -2986 42148 -2952
rect 42182 -2986 42228 -2952
rect 42262 -2986 42308 -2952
rect 42342 -2986 42388 -2952
rect 42422 -2986 42468 -2952
rect 42502 -2986 42548 -2952
rect 42582 -2986 42628 -2952
rect 42662 -2986 42708 -2952
rect 42742 -2986 42788 -2952
rect 42822 -2986 42868 -2952
rect 42902 -2986 42948 -2952
rect 42982 -2986 43028 -2952
rect 43062 -2986 43108 -2952
rect 43142 -2986 43188 -2952
rect 43222 -2986 43268 -2952
rect 43302 -2986 43348 -2952
rect 43382 -2986 43428 -2952
rect 43462 -2986 43508 -2952
rect 43542 -2986 43588 -2952
rect 43622 -2986 43668 -2952
rect 43702 -2986 43748 -2952
rect 43782 -2986 43828 -2952
rect 43862 -2986 43908 -2952
rect 43942 -2986 43988 -2952
rect 44022 -2986 44068 -2952
rect 44102 -2986 44148 -2952
rect 44182 -2986 44228 -2952
rect 44262 -2986 44308 -2952
rect 44342 -2986 44388 -2952
rect 44422 -2986 44468 -2952
rect 44502 -2986 44548 -2952
rect 44582 -2986 44628 -2952
rect 44662 -2986 44708 -2952
rect 44742 -2986 44788 -2952
rect 44822 -2986 44868 -2952
rect 44902 -2986 44948 -2952
rect 44982 -2986 45028 -2952
rect 45062 -2986 45108 -2952
rect 45142 -2986 45188 -2952
rect 45222 -2986 45268 -2952
rect 45302 -2986 45348 -2952
rect 45382 -2986 45428 -2952
rect 45462 -2986 45508 -2952
rect 45542 -2986 45588 -2952
rect 45622 -2986 45668 -2952
rect 45702 -2986 45748 -2952
rect 45782 -2986 45828 -2952
rect 45862 -2986 45908 -2952
rect 45942 -2986 45988 -2952
rect 46022 -2986 46068 -2952
rect 46102 -2986 46148 -2952
rect 46182 -2986 46228 -2952
rect 46262 -2986 46308 -2952
rect 46342 -2986 46388 -2952
rect 46422 -2986 46468 -2952
rect 46502 -2986 46548 -2952
rect 46582 -2986 46628 -2952
rect 46662 -2986 46708 -2952
rect 46742 -2986 46788 -2952
rect 46822 -2986 46868 -2952
rect 46902 -2986 46948 -2952
rect 46982 -2986 47028 -2952
rect 47062 -2986 47108 -2952
rect 47142 -2986 47188 -2952
rect 47222 -2986 47268 -2952
rect 47302 -2986 47349 -2952
rect 47383 -2986 47429 -2952
rect 47463 -2986 47509 -2952
rect 47543 -2986 47589 -2952
rect 47623 -2986 47669 -2952
rect 47703 -2986 47749 -2952
rect 47783 -2986 47829 -2952
rect 47863 -2986 47909 -2952
rect 47943 -2986 47989 -2952
rect 48023 -2986 48069 -2952
rect 48103 -2986 48149 -2952
rect 48183 -2986 48229 -2952
rect 48263 -2986 48309 -2952
rect 48343 -2986 48389 -2952
rect 48423 -2986 48469 -2952
rect 48503 -2986 48549 -2952
rect 48583 -2986 48629 -2952
rect 48663 -2986 48709 -2952
rect 48743 -2986 48789 -2952
rect 48823 -2986 48869 -2952
rect 48903 -2986 48949 -2952
rect 48983 -2986 49029 -2952
rect 49063 -2986 49109 -2952
rect 49143 -2986 49189 -2952
rect 49223 -2986 49269 -2952
rect 49303 -2986 49349 -2952
rect 49383 -2986 49429 -2952
rect 49463 -2986 49509 -2952
rect 49543 -2986 49589 -2952
rect 49623 -2986 49669 -2952
rect 49703 -2986 49749 -2952
rect 49783 -2986 49829 -2952
rect 49863 -2986 49909 -2952
rect 49943 -2986 49989 -2952
rect 50023 -2986 50069 -2952
rect 50103 -2986 50149 -2952
rect 50183 -2986 50229 -2952
rect 50263 -2986 50309 -2952
rect 50343 -2986 50389 -2952
rect 50423 -2986 50469 -2952
rect 50503 -2986 50549 -2952
rect 50583 -2986 50629 -2952
rect 50663 -2986 50709 -2952
rect 50743 -2986 50789 -2952
rect 50823 -2986 50869 -2952
rect 50903 -2986 50949 -2952
rect 50983 -2986 51029 -2952
rect 51063 -2986 51109 -2952
rect 51143 -2986 51189 -2952
rect 51223 -2986 51269 -2952
rect 51303 -2986 51349 -2952
rect 51383 -2986 51429 -2952
rect 51463 -2986 51509 -2952
rect 51543 -2986 51589 -2952
rect 51623 -2986 51662 -2952
rect 35312 -3020 51662 -2986
rect 39430 -3064 39690 -3020
rect 39430 -3116 39474 -3064
rect 39526 -3116 39594 -3064
rect 39646 -3116 39690 -3064
rect 39430 -3184 39690 -3116
rect 39430 -3236 39474 -3184
rect 39526 -3236 39594 -3184
rect 39646 -3236 39690 -3184
rect 39430 -3280 39690 -3236
<< via1 >>
rect 39446 9738 39498 9747
rect 39446 9704 39455 9738
rect 39455 9704 39489 9738
rect 39489 9704 39498 9738
rect 39446 9695 39498 9704
rect 39566 9738 39618 9747
rect 39566 9704 39575 9738
rect 39575 9704 39609 9738
rect 39609 9704 39618 9738
rect 39566 9695 39618 9704
rect 39446 9618 39498 9627
rect 39446 9584 39455 9618
rect 39455 9584 39489 9618
rect 39489 9584 39498 9618
rect 39446 9575 39498 9584
rect 39566 9618 39618 9627
rect 39566 9584 39575 9618
rect 39575 9584 39609 9618
rect 39609 9584 39618 9618
rect 39566 9575 39618 9584
rect 32566 1502 32618 1554
rect 32686 1502 32738 1554
rect 32566 1382 32618 1434
rect 32686 1382 32738 1434
rect 32980 1500 33040 1560
rect 33106 1550 33158 1554
rect 33106 1510 33110 1550
rect 33110 1510 33150 1550
rect 33150 1510 33158 1550
rect 33106 1502 33158 1510
rect 32980 1380 33040 1440
rect 33100 1380 33160 1440
rect 34300 1545 34352 1554
rect 34300 1511 34309 1545
rect 34309 1511 34343 1545
rect 34343 1511 34352 1545
rect 34300 1502 34352 1511
rect 34420 1545 34472 1554
rect 34420 1511 34429 1545
rect 34429 1511 34463 1545
rect 34463 1511 34472 1545
rect 34420 1502 34472 1511
rect 34300 1425 34352 1434
rect 34300 1391 34309 1425
rect 34309 1391 34343 1425
rect 34343 1391 34352 1425
rect 34300 1382 34352 1391
rect 34420 1425 34472 1434
rect 34420 1391 34429 1425
rect 34429 1391 34463 1425
rect 34463 1391 34472 1425
rect 34420 1382 34472 1391
rect 34720 1545 34772 1554
rect 34720 1511 34729 1545
rect 34729 1511 34763 1545
rect 34763 1511 34772 1545
rect 34720 1502 34772 1511
rect 34840 1545 34892 1554
rect 34840 1511 34849 1545
rect 34849 1511 34883 1545
rect 34883 1511 34892 1545
rect 34840 1502 34892 1511
rect 34720 1425 34772 1434
rect 34720 1391 34729 1425
rect 34729 1391 34763 1425
rect 34763 1391 34772 1425
rect 34720 1382 34772 1391
rect 34840 1425 34892 1434
rect 34840 1391 34849 1425
rect 34849 1391 34883 1425
rect 34883 1391 34892 1425
rect 34840 1382 34892 1391
rect 32560 1080 32620 1140
rect 32686 1125 32738 1134
rect 32686 1091 32695 1125
rect 32695 1091 32729 1125
rect 32729 1091 32738 1125
rect 32686 1082 32738 1091
rect 32560 960 32620 1020
rect 32680 960 32740 1020
rect 32980 1080 33040 1140
rect 33100 1080 33160 1140
rect 32980 960 33040 1020
rect 33100 960 33160 1020
rect 34300 1125 34352 1134
rect 34300 1091 34309 1125
rect 34309 1091 34343 1125
rect 34343 1091 34352 1125
rect 34300 1082 34352 1091
rect 34420 1125 34472 1134
rect 34420 1091 34429 1125
rect 34429 1091 34463 1125
rect 34463 1091 34472 1125
rect 34420 1082 34472 1091
rect 34300 1005 34352 1014
rect 34300 971 34309 1005
rect 34309 971 34343 1005
rect 34343 971 34352 1005
rect 34300 962 34352 971
rect 34420 1005 34472 1014
rect 34420 971 34429 1005
rect 34429 971 34463 1005
rect 34463 971 34472 1005
rect 34420 962 34472 971
rect 34720 1125 34772 1134
rect 34720 1091 34729 1125
rect 34729 1091 34763 1125
rect 34763 1091 34772 1125
rect 34720 1082 34772 1091
rect 34840 1125 34892 1134
rect 34840 1091 34849 1125
rect 34849 1091 34883 1125
rect 34883 1091 34892 1125
rect 34840 1082 34892 1091
rect 34720 1005 34772 1014
rect 34720 971 34729 1005
rect 34729 971 34763 1005
rect 34763 971 34772 1005
rect 34720 962 34772 971
rect 34840 1005 34892 1014
rect 34840 971 34849 1005
rect 34849 971 34883 1005
rect 34883 971 34892 1005
rect 34840 962 34892 971
rect 44214 -84 44218 -35
rect 44218 -84 44270 -32
rect 44334 -84 44338 -35
rect 44338 -84 44390 -32
rect 44214 -85 44226 -84
rect 44226 -85 44260 -84
rect 44260 -85 44269 -84
rect 44214 -87 44269 -85
rect 44334 -85 44346 -84
rect 44346 -85 44380 -84
rect 44380 -85 44389 -84
rect 44334 -87 44389 -85
rect 44217 -94 44269 -87
rect 44337 -94 44389 -87
rect 44214 -204 44218 -155
rect 44218 -204 44270 -152
rect 44334 -204 44338 -155
rect 44338 -204 44390 -152
rect 44214 -205 44226 -204
rect 44226 -205 44260 -204
rect 44260 -205 44269 -204
rect 44214 -207 44269 -205
rect 44334 -205 44346 -204
rect 44346 -205 44380 -204
rect 44380 -205 44389 -204
rect 44334 -207 44389 -205
rect 44217 -214 44269 -207
rect 44337 -214 44389 -207
rect 35809 -487 35861 -478
rect 35809 -521 35818 -487
rect 35818 -521 35852 -487
rect 35852 -521 35861 -487
rect 35809 -530 35861 -521
rect 35929 -487 35981 -478
rect 35929 -521 35938 -487
rect 35938 -521 35972 -487
rect 35972 -521 35981 -487
rect 35929 -530 35981 -521
rect 35809 -607 35861 -598
rect 35809 -641 35818 -607
rect 35818 -641 35852 -607
rect 35852 -641 35861 -607
rect 35809 -650 35861 -641
rect 35929 -607 35981 -598
rect 35929 -641 35938 -607
rect 35938 -641 35972 -607
rect 35972 -641 35981 -607
rect 35929 -650 35981 -641
rect 39474 -3073 39526 -3064
rect 39474 -3107 39483 -3073
rect 39483 -3107 39517 -3073
rect 39517 -3107 39526 -3073
rect 39474 -3116 39526 -3107
rect 39594 -3073 39646 -3064
rect 39594 -3107 39603 -3073
rect 39603 -3107 39637 -3073
rect 39637 -3107 39646 -3073
rect 39594 -3116 39646 -3107
rect 39474 -3193 39526 -3184
rect 39474 -3227 39483 -3193
rect 39483 -3227 39517 -3193
rect 39517 -3227 39526 -3193
rect 39474 -3236 39526 -3227
rect 39594 -3193 39646 -3184
rect 39594 -3227 39603 -3193
rect 39603 -3227 39637 -3193
rect 39637 -3227 39646 -3193
rect 39594 -3236 39646 -3227
<< metal2 >>
rect 39402 9749 39662 9791
rect 39402 9693 39444 9749
rect 39500 9693 39564 9749
rect 39620 9693 39662 9749
rect 39402 9629 39662 9693
rect 39402 9573 39444 9629
rect 39500 9573 39564 9629
rect 39620 9573 39662 9629
rect 39402 9531 39662 9573
rect 32522 1560 32782 1598
rect 32522 1500 32560 1560
rect 32620 1500 32680 1560
rect 32740 1500 32782 1560
rect 32522 1440 32782 1500
rect 32522 1380 32560 1440
rect 32620 1380 32680 1440
rect 32740 1380 32782 1440
rect 32522 1338 32782 1380
rect 32942 1560 33202 1598
rect 32942 1500 32980 1560
rect 33040 1500 33100 1560
rect 33160 1500 33202 1560
rect 32942 1440 33202 1500
rect 32942 1380 32980 1440
rect 33040 1380 33100 1440
rect 33160 1380 33202 1440
rect 32942 1338 33202 1380
rect 34256 1554 34516 1598
rect 34256 1502 34300 1554
rect 34352 1502 34420 1554
rect 34472 1502 34516 1554
rect 34256 1434 34516 1502
rect 34256 1382 34300 1434
rect 34352 1382 34420 1434
rect 34472 1382 34516 1434
rect 34256 1338 34516 1382
rect 34676 1554 34936 1598
rect 34676 1502 34720 1554
rect 34772 1502 34840 1554
rect 34892 1502 34936 1554
rect 34676 1434 34936 1502
rect 34676 1382 34720 1434
rect 34772 1382 34840 1434
rect 34892 1382 34936 1434
rect 34676 1338 34936 1382
rect 32522 1140 32782 1178
rect 32522 1080 32560 1140
rect 32620 1134 32782 1140
rect 32620 1082 32686 1134
rect 32738 1082 32782 1134
rect 32620 1080 32782 1082
rect 32522 1020 32782 1080
rect 32522 960 32560 1020
rect 32620 960 32680 1020
rect 32740 960 32782 1020
rect 32522 918 32782 960
rect 32942 1140 33202 1178
rect 32942 1080 32980 1140
rect 33040 1080 33100 1140
rect 33160 1080 33202 1140
rect 32942 1020 33202 1080
rect 32942 960 32980 1020
rect 33040 960 33100 1020
rect 33160 960 33202 1020
rect 32942 918 33202 960
rect 34256 1134 34516 1178
rect 34256 1082 34300 1134
rect 34352 1082 34420 1134
rect 34472 1082 34516 1134
rect 34256 1014 34516 1082
rect 34256 962 34300 1014
rect 34352 962 34420 1014
rect 34472 962 34516 1014
rect 34256 918 34516 962
rect 34676 1134 34936 1178
rect 34676 1082 34720 1134
rect 34772 1082 34840 1134
rect 34892 1082 34936 1134
rect 34676 1014 34936 1082
rect 34676 962 34720 1014
rect 34772 962 34840 1014
rect 34892 962 34936 1014
rect 34676 918 34936 962
rect 44172 2 44432 3
rect 44172 -32 44433 2
rect 44172 -33 44218 -32
rect 44270 -33 44338 -32
rect 44172 -89 44212 -33
rect 44270 -40 44332 -33
rect 44172 -96 44215 -89
rect 44271 -89 44332 -40
rect 44390 -40 44433 -32
rect 44271 -96 44335 -89
rect 44391 -96 44433 -40
rect 44172 -152 44433 -96
rect 44172 -153 44218 -152
rect 44270 -153 44338 -152
rect 44172 -209 44212 -153
rect 44270 -160 44332 -153
rect 44172 -216 44215 -209
rect 44271 -209 44332 -160
rect 44390 -160 44433 -152
rect 44271 -216 44335 -209
rect 44391 -216 44433 -160
rect 44172 -257 44433 -216
rect 44173 -258 44433 -257
rect 35765 -476 36025 -434
rect 35765 -532 35807 -476
rect 35863 -532 35927 -476
rect 35983 -532 36025 -476
rect 35765 -596 36025 -532
rect 35765 -652 35807 -596
rect 35863 -652 35927 -596
rect 35983 -652 36025 -596
rect 35765 -694 36025 -652
rect 39430 -3062 39690 -3020
rect 39430 -3118 39472 -3062
rect 39528 -3118 39592 -3062
rect 39648 -3118 39690 -3062
rect 39430 -3182 39690 -3118
rect 39430 -3238 39472 -3182
rect 39528 -3238 39592 -3182
rect 39648 -3238 39690 -3182
rect 39430 -3280 39690 -3238
<< via2 >>
rect 39444 9747 39500 9749
rect 39444 9695 39446 9747
rect 39446 9695 39498 9747
rect 39498 9695 39500 9747
rect 39444 9693 39500 9695
rect 39564 9747 39620 9749
rect 39564 9695 39566 9747
rect 39566 9695 39618 9747
rect 39618 9695 39620 9747
rect 39564 9693 39620 9695
rect 39444 9627 39500 9629
rect 39444 9575 39446 9627
rect 39446 9575 39498 9627
rect 39498 9575 39500 9627
rect 39444 9573 39500 9575
rect 39564 9627 39620 9629
rect 39564 9575 39566 9627
rect 39566 9575 39618 9627
rect 39618 9575 39620 9627
rect 39564 9573 39620 9575
rect 32560 1554 32620 1560
rect 32560 1502 32566 1554
rect 32566 1502 32618 1554
rect 32618 1502 32620 1554
rect 32560 1500 32620 1502
rect 32680 1554 32740 1560
rect 32680 1502 32686 1554
rect 32686 1502 32738 1554
rect 32738 1502 32740 1554
rect 32680 1500 32740 1502
rect 32560 1434 32620 1440
rect 32560 1382 32566 1434
rect 32566 1382 32618 1434
rect 32618 1382 32620 1434
rect 32560 1380 32620 1382
rect 32680 1434 32740 1440
rect 32680 1382 32686 1434
rect 32686 1382 32738 1434
rect 32738 1382 32740 1434
rect 32680 1380 32740 1382
rect 32980 1500 33040 1560
rect 33100 1554 33160 1560
rect 33100 1502 33106 1554
rect 33106 1502 33158 1554
rect 33158 1502 33160 1554
rect 33100 1500 33160 1502
rect 32980 1380 33040 1440
rect 33100 1380 33160 1440
rect 32560 1080 32620 1140
rect 32560 960 32620 1020
rect 32680 960 32740 1020
rect 32980 1080 33040 1140
rect 33100 1080 33160 1140
rect 32980 960 33040 1020
rect 33100 960 33160 1020
rect 44212 -35 44218 -33
rect 44218 -35 44268 -33
rect 44212 -87 44214 -35
rect 44214 -40 44268 -35
rect 44332 -35 44338 -33
rect 44338 -35 44388 -33
rect 44214 -84 44270 -40
rect 44270 -84 44271 -40
rect 44214 -87 44269 -84
rect 44212 -89 44217 -87
rect 44215 -94 44217 -89
rect 44217 -94 44269 -87
rect 44269 -94 44271 -84
rect 44332 -87 44334 -35
rect 44334 -40 44388 -35
rect 44334 -84 44390 -40
rect 44390 -84 44391 -40
rect 44334 -87 44389 -84
rect 44332 -89 44337 -87
rect 44215 -96 44271 -94
rect 44335 -94 44337 -89
rect 44337 -94 44389 -87
rect 44389 -94 44391 -84
rect 44335 -96 44391 -94
rect 44212 -155 44218 -153
rect 44218 -155 44268 -153
rect 44212 -207 44214 -155
rect 44214 -160 44268 -155
rect 44332 -155 44338 -153
rect 44338 -155 44388 -153
rect 44214 -204 44270 -160
rect 44270 -204 44271 -160
rect 44214 -207 44269 -204
rect 44212 -209 44217 -207
rect 44215 -214 44217 -209
rect 44217 -214 44269 -207
rect 44269 -214 44271 -204
rect 44332 -207 44334 -155
rect 44334 -160 44388 -155
rect 44334 -204 44390 -160
rect 44390 -204 44391 -160
rect 44334 -207 44389 -204
rect 44332 -209 44337 -207
rect 44215 -216 44271 -214
rect 44335 -214 44337 -209
rect 44337 -214 44389 -207
rect 44389 -214 44391 -204
rect 44335 -216 44391 -214
rect 35807 -478 35863 -476
rect 35807 -530 35809 -478
rect 35809 -530 35861 -478
rect 35861 -530 35863 -478
rect 35807 -532 35863 -530
rect 35927 -478 35983 -476
rect 35927 -530 35929 -478
rect 35929 -530 35981 -478
rect 35981 -530 35983 -478
rect 35927 -532 35983 -530
rect 35807 -598 35863 -596
rect 35807 -650 35809 -598
rect 35809 -650 35861 -598
rect 35861 -650 35863 -598
rect 35807 -652 35863 -650
rect 35927 -598 35983 -596
rect 35927 -650 35929 -598
rect 35929 -650 35981 -598
rect 35981 -650 35983 -598
rect 35927 -652 35983 -650
rect 39472 -3064 39528 -3062
rect 39472 -3116 39474 -3064
rect 39474 -3116 39526 -3064
rect 39526 -3116 39528 -3064
rect 39472 -3118 39528 -3116
rect 39592 -3064 39648 -3062
rect 39592 -3116 39594 -3064
rect 39594 -3116 39646 -3064
rect 39646 -3116 39648 -3064
rect 39592 -3118 39648 -3116
rect 39472 -3184 39528 -3182
rect 39472 -3236 39474 -3184
rect 39474 -3236 39526 -3184
rect 39526 -3236 39528 -3184
rect 39472 -3238 39528 -3236
rect 39592 -3184 39648 -3182
rect 39592 -3236 39594 -3184
rect 39594 -3236 39646 -3184
rect 39646 -3236 39648 -3184
rect 39592 -3238 39648 -3236
<< metal3 >>
rect 35700 9791 39650 9878
rect 35700 9753 39662 9791
rect 35700 9689 39440 9753
rect 39504 9689 39560 9753
rect 39624 9689 39662 9753
rect 35700 9633 39662 9689
rect 35700 9569 39440 9633
rect 39504 9569 39560 9633
rect 39624 9569 39662 9633
rect 35700 9531 39662 9569
rect 35700 9478 39650 9531
rect 32522 1560 32782 1598
rect 32522 1496 32560 1560
rect 32624 1496 32680 1560
rect 32744 1496 32782 1560
rect 32522 1440 32782 1496
rect 32522 1376 32560 1440
rect 32624 1376 32680 1440
rect 32744 1376 32782 1440
rect 32522 1338 32782 1376
rect 32942 1560 33202 1598
rect 32942 1496 32980 1560
rect 33044 1496 33100 1560
rect 33164 1496 33202 1560
rect 32942 1440 33202 1496
rect 32942 1376 32980 1440
rect 33044 1376 33100 1440
rect 33164 1376 33202 1440
rect 32942 1338 33202 1376
rect 34256 1560 34516 1598
rect 34256 1496 34294 1560
rect 34358 1496 34414 1560
rect 34478 1496 34516 1560
rect 34256 1440 34516 1496
rect 34256 1376 34294 1440
rect 34358 1376 34414 1440
rect 34478 1376 34516 1440
rect 34256 1338 34516 1376
rect 34676 1560 34936 1598
rect 34676 1496 34714 1560
rect 34778 1496 34834 1560
rect 34898 1496 34936 1560
rect 34676 1440 34936 1496
rect 34676 1376 34714 1440
rect 34778 1376 34834 1440
rect 34898 1376 34936 1440
rect 34676 1338 34936 1376
rect 32522 1140 32782 1178
rect 32522 1076 32560 1140
rect 32624 1076 32680 1140
rect 32744 1076 32782 1140
rect 32522 1020 32782 1076
rect 32522 956 32560 1020
rect 32624 956 32680 1020
rect 32744 956 32782 1020
rect 32522 918 32782 956
rect 32942 1140 33202 1178
rect 32942 1076 32980 1140
rect 33044 1076 33100 1140
rect 33164 1076 33202 1140
rect 32942 1020 33202 1076
rect 32942 956 32980 1020
rect 33044 956 33100 1020
rect 33164 956 33202 1020
rect 32942 918 33202 956
rect 34256 1140 34516 1178
rect 34256 1076 34294 1140
rect 34358 1076 34414 1140
rect 34478 1076 34516 1140
rect 34256 1020 34516 1076
rect 34256 956 34294 1020
rect 34358 956 34414 1020
rect 34478 956 34516 1020
rect 34256 918 34516 956
rect 34676 1140 34936 1178
rect 34676 1076 34714 1140
rect 34778 1076 34834 1140
rect 34898 1076 34936 1140
rect 34676 1020 34936 1076
rect 34676 956 34714 1020
rect 34778 956 34834 1020
rect 34898 956 34936 1020
rect 34676 918 34936 956
rect 35700 -472 36100 9478
rect 35700 -536 35803 -472
rect 35867 -536 35923 -472
rect 35987 -536 36100 -472
rect 35700 -592 36100 -536
rect 35700 -656 35803 -592
rect 35867 -656 35923 -592
rect 35987 -656 36100 -592
rect 35700 -775 36100 -656
rect 36725 1784 39434 1817
rect 36725 1720 39350 1784
rect 39414 1720 39434 1784
rect 36725 1704 39434 1720
rect 36725 1640 39350 1704
rect 39414 1640 39434 1704
rect 36725 1624 39434 1640
rect 36725 1560 39350 1624
rect 39414 1560 39434 1624
rect 36725 1544 39434 1560
rect 36725 1480 39350 1544
rect 39414 1480 39434 1544
rect 36725 1464 39434 1480
rect 36725 1400 39350 1464
rect 39414 1400 39434 1464
rect 36725 1384 39434 1400
rect 36725 1320 39350 1384
rect 39414 1320 39434 1384
rect 36725 1304 39434 1320
rect 36725 1240 39350 1304
rect 39414 1240 39434 1304
rect 36725 1224 39434 1240
rect 36725 1160 39350 1224
rect 39414 1160 39434 1224
rect 36725 1144 39434 1160
rect 36725 1080 39350 1144
rect 39414 1080 39434 1144
rect 36725 1064 39434 1080
rect 36725 1000 39350 1064
rect 39414 1000 39434 1064
rect 36725 984 39434 1000
rect 36725 920 39350 984
rect 39414 920 39434 984
rect 36725 904 39434 920
rect 36725 840 39350 904
rect 39414 840 39434 904
rect 36725 824 39434 840
rect 36725 760 39350 824
rect 39414 760 39434 824
rect 36725 744 39434 760
rect 36725 680 39350 744
rect 39414 680 39434 744
rect 36725 664 39434 680
rect 36725 600 39350 664
rect 39414 600 39434 664
rect 36725 584 39434 600
rect 36725 520 39350 584
rect 39414 520 39434 584
rect 36725 504 39434 520
rect 36725 440 39350 504
rect 39414 440 39434 504
rect 36725 424 39434 440
rect 36725 360 39350 424
rect 39414 360 39434 424
rect 36725 344 39434 360
rect 36725 280 39350 344
rect 39414 280 39434 344
rect 36725 264 39434 280
rect 36725 200 39350 264
rect 39414 200 39434 264
rect 36725 184 39434 200
rect 36725 120 39350 184
rect 39414 120 39434 184
rect 36725 104 39434 120
rect 36725 40 39350 104
rect 39414 40 39434 104
rect 36725 24 39434 40
rect 36725 -40 39350 24
rect 39414 -40 39434 24
rect 44552 1620 46611 1668
rect 44552 1556 44572 1620
rect 44636 1556 46611 1620
rect 44552 1540 46611 1556
rect 44552 1476 44572 1540
rect 44636 1476 46611 1540
rect 44552 1460 46611 1476
rect 44552 1396 44572 1460
rect 44636 1396 46611 1460
rect 44552 1380 46611 1396
rect 44552 1316 44572 1380
rect 44636 1316 46611 1380
rect 44552 1300 46611 1316
rect 44552 1236 44572 1300
rect 44636 1236 46611 1300
rect 44552 1220 46611 1236
rect 44552 1156 44572 1220
rect 44636 1156 46611 1220
rect 44552 1140 46611 1156
rect 44552 1076 44572 1140
rect 44636 1076 46611 1140
rect 44552 1060 46611 1076
rect 44552 996 44572 1060
rect 44636 996 46611 1060
rect 44552 980 46611 996
rect 44552 916 44572 980
rect 44636 916 46611 980
rect 44552 900 46611 916
rect 44552 836 44572 900
rect 44636 836 46611 900
rect 44552 820 46611 836
rect 44552 756 44572 820
rect 44636 756 46611 820
rect 44552 740 46611 756
rect 44552 676 44572 740
rect 44636 676 46611 740
rect 44552 660 46611 676
rect 44552 596 44572 660
rect 44636 596 46611 660
rect 44552 580 46611 596
rect 44552 516 44572 580
rect 44636 516 46611 580
rect 44552 500 46611 516
rect 44552 436 44572 500
rect 44636 470 46611 500
rect 44636 436 46610 470
rect 44552 420 46610 436
rect 44552 356 44572 420
rect 44636 356 46610 420
rect 44552 340 46610 356
rect 44552 276 44572 340
rect 44636 276 46610 340
rect 44552 260 46610 276
rect 44552 196 44572 260
rect 44636 196 46610 260
rect 44552 180 46610 196
rect 44552 116 44572 180
rect 44636 116 46610 180
rect 44552 100 46610 116
rect 44552 36 44572 100
rect 44636 36 46610 100
rect 44552 20 46610 36
rect 36725 -56 39434 -40
rect 36725 -120 39350 -56
rect 39414 -120 39434 -56
rect 36725 -136 39434 -120
rect 36725 -200 39350 -136
rect 39414 -200 39434 -136
rect 36725 -216 39434 -200
rect 36725 -280 39350 -216
rect 39414 -280 39434 -216
rect 44172 -33 44433 3
rect 44172 -36 44212 -33
rect 44268 -36 44332 -33
rect 44388 -36 44433 -33
rect 44172 -100 44211 -36
rect 44275 -100 44331 -36
rect 44395 -100 44433 -36
rect 44172 -153 44433 -100
rect 44172 -156 44212 -153
rect 44268 -156 44332 -153
rect 44388 -156 44433 -153
rect 44172 -220 44211 -156
rect 44275 -220 44331 -156
rect 44395 -220 44433 -156
rect 44172 -258 44433 -220
rect 44552 -44 44572 20
rect 44636 -44 46610 20
rect 44552 -60 46610 -44
rect 44552 -124 44572 -60
rect 44636 -124 46610 -60
rect 44552 -140 46610 -124
rect 44552 -204 44572 -140
rect 44636 -199 46610 -140
rect 44636 -204 46611 -199
rect 44552 -220 46611 -204
rect 36725 -296 39434 -280
rect 36725 -360 39350 -296
rect 39414 -360 39434 -296
rect 44552 -284 44572 -220
rect 44636 -284 46611 -220
rect 44552 -332 46611 -284
rect 36725 -376 39434 -360
rect 36725 -440 39350 -376
rect 39414 -440 39434 -376
rect 36725 -456 39434 -440
rect 36725 -520 39350 -456
rect 39414 -520 39434 -456
rect 36725 -536 39434 -520
rect 36725 -600 39350 -536
rect 39414 -600 39434 -536
rect 36725 -616 39434 -600
rect 36725 -680 39350 -616
rect 39414 -680 39434 -616
rect 36725 -696 39434 -680
rect 36725 -760 39350 -696
rect 39414 -760 39434 -696
rect 36725 -793 39434 -760
rect 39430 -3058 39690 -3020
rect 39430 -3122 39468 -3058
rect 39532 -3122 39588 -3058
rect 39652 -3122 39690 -3058
rect 39430 -3178 39690 -3122
rect 39430 -3242 39468 -3178
rect 39532 -3242 39588 -3178
rect 39652 -3242 39690 -3178
rect 39430 -3280 39690 -3242
<< via3 >>
rect 39440 9749 39504 9753
rect 39440 9693 39444 9749
rect 39444 9693 39500 9749
rect 39500 9693 39504 9749
rect 39440 9689 39504 9693
rect 39560 9749 39624 9753
rect 39560 9693 39564 9749
rect 39564 9693 39620 9749
rect 39620 9693 39624 9749
rect 39560 9689 39624 9693
rect 39440 9629 39504 9633
rect 39440 9573 39444 9629
rect 39444 9573 39500 9629
rect 39500 9573 39504 9629
rect 39440 9569 39504 9573
rect 39560 9629 39624 9633
rect 39560 9573 39564 9629
rect 39564 9573 39620 9629
rect 39620 9573 39624 9629
rect 39560 9569 39624 9573
rect 32560 1500 32620 1560
rect 32620 1500 32624 1560
rect 32560 1496 32624 1500
rect 32680 1500 32740 1560
rect 32740 1500 32744 1560
rect 32680 1496 32744 1500
rect 32560 1380 32620 1440
rect 32620 1380 32624 1440
rect 32560 1376 32624 1380
rect 32680 1380 32740 1440
rect 32740 1380 32744 1440
rect 32680 1376 32744 1380
rect 32980 1500 33040 1560
rect 33040 1500 33044 1560
rect 32980 1496 33044 1500
rect 33100 1500 33160 1560
rect 33160 1500 33164 1560
rect 33100 1496 33164 1500
rect 32980 1380 33040 1440
rect 33040 1380 33044 1440
rect 32980 1376 33044 1380
rect 33100 1380 33160 1440
rect 33160 1380 33164 1440
rect 33100 1376 33164 1380
rect 34294 1496 34358 1560
rect 34414 1496 34478 1560
rect 34294 1376 34358 1440
rect 34414 1376 34478 1440
rect 34714 1496 34778 1560
rect 34834 1496 34898 1560
rect 34714 1376 34778 1440
rect 34834 1376 34898 1440
rect 32560 1080 32620 1140
rect 32620 1080 32624 1140
rect 32560 1076 32624 1080
rect 32680 1076 32744 1140
rect 32560 960 32620 1020
rect 32620 960 32624 1020
rect 32560 956 32624 960
rect 32680 960 32740 1020
rect 32740 960 32744 1020
rect 32680 956 32744 960
rect 32980 1080 33040 1140
rect 33040 1080 33044 1140
rect 32980 1076 33044 1080
rect 33100 1080 33160 1140
rect 33160 1080 33164 1140
rect 33100 1076 33164 1080
rect 32980 960 33040 1020
rect 33040 960 33044 1020
rect 32980 956 33044 960
rect 33100 960 33160 1020
rect 33160 960 33164 1020
rect 33100 956 33164 960
rect 34294 1076 34358 1140
rect 34414 1076 34478 1140
rect 34294 956 34358 1020
rect 34414 956 34478 1020
rect 34714 1076 34778 1140
rect 34834 1076 34898 1140
rect 34714 956 34778 1020
rect 34834 956 34898 1020
rect 35803 -476 35867 -472
rect 35803 -532 35807 -476
rect 35807 -532 35863 -476
rect 35863 -532 35867 -476
rect 35803 -536 35867 -532
rect 35923 -476 35987 -472
rect 35923 -532 35927 -476
rect 35927 -532 35983 -476
rect 35983 -532 35987 -476
rect 35923 -536 35987 -532
rect 35803 -596 35867 -592
rect 35803 -652 35807 -596
rect 35807 -652 35863 -596
rect 35863 -652 35867 -596
rect 35803 -656 35867 -652
rect 35923 -596 35987 -592
rect 35923 -652 35927 -596
rect 35927 -652 35983 -596
rect 35983 -652 35987 -596
rect 35923 -656 35987 -652
rect 39350 1720 39414 1784
rect 39350 1640 39414 1704
rect 39350 1560 39414 1624
rect 39350 1480 39414 1544
rect 39350 1400 39414 1464
rect 39350 1320 39414 1384
rect 39350 1240 39414 1304
rect 39350 1160 39414 1224
rect 39350 1080 39414 1144
rect 39350 1000 39414 1064
rect 39350 920 39414 984
rect 39350 840 39414 904
rect 39350 760 39414 824
rect 39350 680 39414 744
rect 39350 600 39414 664
rect 39350 520 39414 584
rect 39350 440 39414 504
rect 39350 360 39414 424
rect 39350 280 39414 344
rect 39350 200 39414 264
rect 39350 120 39414 184
rect 39350 40 39414 104
rect 39350 -40 39414 24
rect 44572 1556 44636 1620
rect 44572 1476 44636 1540
rect 44572 1396 44636 1460
rect 44572 1316 44636 1380
rect 44572 1236 44636 1300
rect 44572 1156 44636 1220
rect 44572 1076 44636 1140
rect 44572 996 44636 1060
rect 44572 916 44636 980
rect 44572 836 44636 900
rect 44572 756 44636 820
rect 44572 676 44636 740
rect 44572 596 44636 660
rect 44572 516 44636 580
rect 44572 436 44636 500
rect 44572 356 44636 420
rect 44572 276 44636 340
rect 44572 196 44636 260
rect 44572 116 44636 180
rect 44572 36 44636 100
rect 39350 -120 39414 -56
rect 39350 -200 39414 -136
rect 39350 -280 39414 -216
rect 44211 -89 44212 -36
rect 44212 -40 44268 -36
rect 44268 -40 44275 -36
rect 44212 -89 44271 -40
rect 44211 -96 44215 -89
rect 44215 -96 44271 -89
rect 44271 -96 44275 -40
rect 44211 -100 44275 -96
rect 44331 -89 44332 -36
rect 44332 -40 44388 -36
rect 44388 -40 44395 -36
rect 44332 -89 44391 -40
rect 44331 -96 44335 -89
rect 44335 -96 44391 -89
rect 44391 -96 44395 -40
rect 44331 -100 44395 -96
rect 44211 -209 44212 -156
rect 44212 -160 44268 -156
rect 44268 -160 44275 -156
rect 44212 -209 44271 -160
rect 44211 -216 44215 -209
rect 44215 -216 44271 -209
rect 44271 -216 44275 -160
rect 44211 -220 44275 -216
rect 44331 -209 44332 -156
rect 44332 -160 44388 -156
rect 44388 -160 44395 -156
rect 44332 -209 44391 -160
rect 44331 -216 44335 -209
rect 44335 -216 44391 -209
rect 44391 -216 44395 -160
rect 44331 -220 44395 -216
rect 44572 -44 44636 20
rect 44572 -124 44636 -60
rect 44572 -204 44636 -140
rect 39350 -360 39414 -296
rect 44572 -284 44636 -220
rect 39350 -440 39414 -376
rect 39350 -520 39414 -456
rect 39350 -600 39414 -536
rect 39350 -680 39414 -616
rect 39350 -760 39414 -696
rect 39468 -3062 39532 -3058
rect 39468 -3118 39472 -3062
rect 39472 -3118 39528 -3062
rect 39528 -3118 39532 -3062
rect 39468 -3122 39532 -3118
rect 39588 -3062 39652 -3058
rect 39588 -3118 39592 -3062
rect 39592 -3118 39648 -3062
rect 39648 -3118 39652 -3062
rect 39588 -3122 39652 -3118
rect 39468 -3182 39532 -3178
rect 39468 -3238 39472 -3182
rect 39472 -3238 39528 -3182
rect 39528 -3238 39532 -3182
rect 39468 -3242 39532 -3238
rect 39588 -3182 39652 -3178
rect 39588 -3238 39592 -3182
rect 39592 -3238 39648 -3182
rect 39648 -3238 39652 -3182
rect 39588 -3242 39652 -3238
<< mimcap >>
rect 36825 1664 39235 1717
rect 36825 -640 36878 1664
rect 39182 -640 39235 1664
rect 44751 1500 46511 1568
rect 44751 -164 44799 1500
rect 46463 -164 46511 1500
rect 44751 -232 46511 -164
rect 36825 -693 39235 -640
<< mimcapcontact >>
rect 36878 -640 39182 1664
rect 44799 -164 46463 1500
<< metal4 >>
rect 29031 39132 64231 39332
rect 29031 4332 29231 39132
rect 29631 38532 63631 38732
rect 29631 4932 29831 38532
rect 30231 37932 63031 38132
rect 30231 5532 30431 37932
rect 30831 37332 62431 37532
rect 30831 6132 31031 37332
rect 31431 36732 61831 36932
rect 31431 6732 31631 36732
rect 32031 36132 61231 36332
rect 32031 7332 32231 36132
rect 32631 35532 60631 35732
rect 32631 7932 32831 35532
rect 33231 34932 60031 35132
rect 33231 8532 33431 34932
rect 33831 34332 59431 34532
rect 33831 9132 34031 34332
rect 39402 9753 39662 9791
rect 39402 9689 39440 9753
rect 39504 9689 39560 9753
rect 39624 9732 39662 9753
rect 59231 9732 59431 34332
rect 39624 9689 59431 9732
rect 39402 9633 59431 9689
rect 39402 9569 39440 9633
rect 39504 9569 39560 9633
rect 39624 9569 59431 9633
rect 39402 9532 59431 9569
rect 39402 9531 39662 9532
rect 59831 9132 60031 34932
rect 33831 8932 60031 9132
rect 60431 8532 60631 35532
rect 33231 8332 60631 8532
rect 61031 7932 61231 36132
rect 32631 7732 61231 7932
rect 61631 7332 61831 36732
rect 32031 7132 61831 7332
rect 62231 6732 62431 37332
rect 31431 6532 62431 6732
rect 62831 6132 63031 37932
rect 30831 5932 63031 6132
rect 63431 5532 63631 38532
rect 30231 5332 63631 5532
rect 64031 4932 64231 39132
rect 29631 4732 64231 4932
rect 29031 4132 47085 4332
rect 39334 1784 39430 1805
rect 39334 1720 39350 1784
rect 39414 1720 39430 1784
rect 39334 1704 39430 1720
rect 35431 1664 39196 1678
rect 35431 1663 36878 1664
rect 32522 1586 32782 1598
rect 32522 1350 32534 1586
rect 32770 1350 32782 1586
rect 32522 1338 32782 1350
rect 32942 1586 33202 1598
rect 32942 1350 32954 1586
rect 33190 1350 33202 1586
rect 32942 1338 33202 1350
rect 34229 1586 36878 1663
rect 34229 1350 34268 1586
rect 34504 1350 34688 1586
rect 34924 1350 36878 1586
rect 32522 1166 32782 1178
rect 32522 930 32534 1166
rect 32770 930 32782 1166
rect 32522 918 32782 930
rect 32942 1166 33202 1178
rect 32942 930 32954 1166
rect 33190 930 33202 1166
rect 32942 918 33202 930
rect 34229 1166 36878 1350
rect 34229 930 34268 1166
rect 34504 930 34688 1166
rect 34924 930 36878 1166
rect 34229 863 36878 930
rect 35431 -472 36878 863
rect 35431 -536 35803 -472
rect 35867 -536 35923 -472
rect 35987 -536 36878 -472
rect 35431 -592 36878 -536
rect 35431 -656 35803 -592
rect 35867 -656 35923 -592
rect 35987 -640 36878 -592
rect 39182 -640 39196 1664
rect 35987 -654 39196 -640
rect 39334 1640 39350 1704
rect 39414 1640 39430 1704
rect 39334 1624 39430 1640
rect 39334 1560 39350 1624
rect 39414 1560 39430 1624
rect 39334 1544 39430 1560
rect 39334 1480 39350 1544
rect 39414 1480 39430 1544
rect 39334 1464 39430 1480
rect 39334 1400 39350 1464
rect 39414 1400 39430 1464
rect 39334 1384 39430 1400
rect 39334 1320 39350 1384
rect 39414 1320 39430 1384
rect 39334 1304 39430 1320
rect 39334 1240 39350 1304
rect 39414 1240 39430 1304
rect 39334 1224 39430 1240
rect 39334 1160 39350 1224
rect 39414 1160 39430 1224
rect 39334 1144 39430 1160
rect 39334 1080 39350 1144
rect 39414 1080 39430 1144
rect 39334 1064 39430 1080
rect 39334 1000 39350 1064
rect 39414 1000 39430 1064
rect 39334 984 39430 1000
rect 39334 920 39350 984
rect 39414 920 39430 984
rect 39334 904 39430 920
rect 39334 840 39350 904
rect 39414 840 39430 904
rect 39334 824 39430 840
rect 39334 760 39350 824
rect 39414 760 39430 824
rect 39334 744 39430 760
rect 39334 680 39350 744
rect 39414 680 39430 744
rect 39334 664 39430 680
rect 39334 600 39350 664
rect 39414 600 39430 664
rect 39334 584 39430 600
rect 39334 520 39350 584
rect 39414 520 39430 584
rect 39334 504 39430 520
rect 39334 440 39350 504
rect 39414 440 39430 504
rect 39334 424 39430 440
rect 39334 360 39350 424
rect 39414 360 39430 424
rect 39334 344 39430 360
rect 39334 280 39350 344
rect 39414 280 39430 344
rect 44556 1620 44652 1656
rect 44556 1556 44572 1620
rect 44636 1556 44652 1620
rect 44556 1540 44652 1556
rect 44556 1476 44572 1540
rect 44636 1476 44652 1540
rect 46825 1529 47085 4132
rect 44556 1460 44652 1476
rect 44556 1396 44572 1460
rect 44636 1396 44652 1460
rect 44556 1380 44652 1396
rect 44556 1316 44572 1380
rect 44636 1316 44652 1380
rect 44556 1300 44652 1316
rect 44556 1236 44572 1300
rect 44636 1236 44652 1300
rect 44556 1220 44652 1236
rect 44556 1156 44572 1220
rect 44636 1156 44652 1220
rect 44556 1140 44652 1156
rect 44556 1076 44572 1140
rect 44636 1076 44652 1140
rect 44556 1060 44652 1076
rect 44556 996 44572 1060
rect 44636 996 44652 1060
rect 44556 980 44652 996
rect 44556 916 44572 980
rect 44636 916 44652 980
rect 44556 900 44652 916
rect 44556 836 44572 900
rect 44636 836 44652 900
rect 44556 820 44652 836
rect 44556 756 44572 820
rect 44636 756 44652 820
rect 44556 740 44652 756
rect 44556 676 44572 740
rect 44636 676 44652 740
rect 44556 660 44652 676
rect 44556 596 44572 660
rect 44636 596 44652 660
rect 44556 580 44652 596
rect 44556 516 44572 580
rect 44636 516 44652 580
rect 44556 500 44652 516
rect 44556 436 44572 500
rect 44636 436 44652 500
rect 44556 420 44652 436
rect 44556 356 44572 420
rect 44636 356 44652 420
rect 44556 343 44652 356
rect 39334 264 39430 280
rect 39334 200 39350 264
rect 39414 200 39430 264
rect 39334 184 39430 200
rect 39334 120 39350 184
rect 39414 120 39430 184
rect 39334 104 39430 120
rect 39334 40 39350 104
rect 39414 40 39430 104
rect 39334 24 39430 40
rect 39334 -40 39350 24
rect 39414 -40 39430 24
rect 39334 -56 39430 -40
rect 39334 -120 39350 -56
rect 39414 -120 39430 -56
rect 39334 -136 39430 -120
rect 39334 -200 39350 -136
rect 39414 -200 39430 -136
rect 39334 -216 39430 -200
rect 39334 -280 39350 -216
rect 39414 -280 39430 -216
rect 39334 -296 39430 -280
rect 39334 -360 39350 -296
rect 39414 -324 39430 -296
rect 44011 340 44652 343
rect 44011 276 44572 340
rect 44636 276 44652 340
rect 44011 260 44652 276
rect 44011 196 44572 260
rect 44636 196 44652 260
rect 44011 180 44652 196
rect 44011 116 44572 180
rect 44636 116 44652 180
rect 44011 100 44652 116
rect 44011 36 44572 100
rect 44636 36 44652 100
rect 44011 20 44652 36
rect 44011 -36 44572 20
rect 44011 -100 44211 -36
rect 44275 -100 44331 -36
rect 44395 -44 44572 -36
rect 44636 -44 44652 20
rect 44395 -60 44652 -44
rect 44395 -100 44572 -60
rect 44011 -124 44572 -100
rect 44636 -124 44652 -60
rect 44011 -140 44652 -124
rect 44011 -156 44572 -140
rect 44011 -220 44211 -156
rect 44275 -220 44331 -156
rect 44395 -204 44572 -156
rect 44636 -204 44652 -140
rect 44790 1500 47085 1529
rect 44790 -164 44799 1500
rect 46463 1084 47085 1500
rect 46463 -164 46472 1084
rect 44790 -193 46472 -164
rect 44395 -220 44652 -204
rect 44011 -284 44572 -220
rect 44636 -284 44652 -220
rect 44011 -320 44652 -284
rect 39414 -360 39690 -324
rect 39334 -376 39690 -360
rect 39334 -440 39350 -376
rect 39414 -440 39690 -376
rect 39334 -456 39690 -440
rect 39334 -520 39350 -456
rect 39414 -520 39690 -456
rect 39334 -536 39690 -520
rect 39334 -600 39350 -536
rect 39414 -600 39690 -536
rect 39334 -616 39690 -600
rect 35987 -656 36864 -654
rect 35431 -924 36864 -656
rect 39334 -680 39350 -616
rect 39414 -680 39690 -616
rect 39334 -696 39690 -680
rect 39334 -760 39350 -696
rect 39414 -760 39690 -696
rect 39334 -781 39690 -760
rect 39430 -3058 39690 -781
rect 39430 -3122 39468 -3058
rect 39532 -3122 39588 -3058
rect 39652 -3122 39690 -3058
rect 39430 -3178 39690 -3122
rect 39430 -3242 39468 -3178
rect 39532 -3242 39588 -3178
rect 39652 -3242 39690 -3178
rect 39430 -3280 39690 -3242
<< via4 >>
rect 32534 1560 32770 1586
rect 32534 1496 32560 1560
rect 32560 1496 32624 1560
rect 32624 1496 32680 1560
rect 32680 1496 32744 1560
rect 32744 1496 32770 1560
rect 32534 1440 32770 1496
rect 32534 1376 32560 1440
rect 32560 1376 32624 1440
rect 32624 1376 32680 1440
rect 32680 1376 32744 1440
rect 32744 1376 32770 1440
rect 32534 1350 32770 1376
rect 32954 1560 33190 1586
rect 32954 1496 32980 1560
rect 32980 1496 33044 1560
rect 33044 1496 33100 1560
rect 33100 1496 33164 1560
rect 33164 1496 33190 1560
rect 32954 1440 33190 1496
rect 32954 1376 32980 1440
rect 32980 1376 33044 1440
rect 33044 1376 33100 1440
rect 33100 1376 33164 1440
rect 33164 1376 33190 1440
rect 32954 1350 33190 1376
rect 34268 1560 34504 1586
rect 34268 1496 34294 1560
rect 34294 1496 34358 1560
rect 34358 1496 34414 1560
rect 34414 1496 34478 1560
rect 34478 1496 34504 1560
rect 34268 1440 34504 1496
rect 34268 1376 34294 1440
rect 34294 1376 34358 1440
rect 34358 1376 34414 1440
rect 34414 1376 34478 1440
rect 34478 1376 34504 1440
rect 34268 1350 34504 1376
rect 34688 1560 34924 1586
rect 34688 1496 34714 1560
rect 34714 1496 34778 1560
rect 34778 1496 34834 1560
rect 34834 1496 34898 1560
rect 34898 1496 34924 1560
rect 34688 1440 34924 1496
rect 34688 1376 34714 1440
rect 34714 1376 34778 1440
rect 34778 1376 34834 1440
rect 34834 1376 34898 1440
rect 34898 1376 34924 1440
rect 34688 1350 34924 1376
rect 32534 1140 32770 1166
rect 32534 1076 32560 1140
rect 32560 1076 32624 1140
rect 32624 1076 32680 1140
rect 32680 1076 32744 1140
rect 32744 1076 32770 1140
rect 32534 1020 32770 1076
rect 32534 956 32560 1020
rect 32560 956 32624 1020
rect 32624 956 32680 1020
rect 32680 956 32744 1020
rect 32744 956 32770 1020
rect 32534 930 32770 956
rect 32954 1140 33190 1166
rect 32954 1076 32980 1140
rect 32980 1076 33044 1140
rect 33044 1076 33100 1140
rect 33100 1076 33164 1140
rect 33164 1076 33190 1140
rect 32954 1020 33190 1076
rect 32954 956 32980 1020
rect 32980 956 33044 1020
rect 33044 956 33100 1020
rect 33100 956 33164 1020
rect 33164 956 33190 1020
rect 32954 930 33190 956
rect 34268 1140 34504 1166
rect 34268 1076 34294 1140
rect 34294 1076 34358 1140
rect 34358 1076 34414 1140
rect 34414 1076 34478 1140
rect 34478 1076 34504 1140
rect 34268 1020 34504 1076
rect 34268 956 34294 1020
rect 34294 956 34358 1020
rect 34358 956 34414 1020
rect 34414 956 34478 1020
rect 34478 956 34504 1020
rect 34268 930 34504 956
rect 34688 1140 34924 1166
rect 34688 1076 34714 1140
rect 34714 1076 34778 1140
rect 34778 1076 34834 1140
rect 34834 1076 34898 1140
rect 34898 1076 34924 1140
rect 34688 1020 34924 1076
rect 34688 956 34714 1020
rect 34714 956 34778 1020
rect 34778 956 34834 1020
rect 34834 956 34898 1020
rect 34898 956 34924 1020
rect 34688 930 34924 956
<< metal5 >>
rect 32441 1665 33282 1678
rect 34175 1665 35016 1678
rect 32441 1586 35016 1665
rect 32441 1350 32534 1586
rect 32770 1350 32954 1586
rect 33190 1350 34268 1586
rect 34504 1350 34688 1586
rect 34924 1350 35016 1586
rect 32441 1166 35016 1350
rect 32441 930 32534 1166
rect 32770 930 32954 1166
rect 33190 930 34268 1166
rect 34504 930 34688 1166
rect 34924 930 35016 1166
rect 32441 865 35016 930
rect 32441 838 33282 865
rect 34175 838 35016 865
<< labels >>
flabel metal1 s 35558 -1479 35603 -1429 2 FreeSans 2000 0 0 0 Input
port 1 nsew
flabel metal1 s 39022 -2989 39234 -2862 2 FreeSans 2000 0 0 0 Ground
port 2 nsew
flabel metal1 s 34828 2547 35029 2675 2 FreeSans 2000 0 0 0 VDD
port 3 nsew
<< properties >>
string path -24.085 18.975 -16.135 18.975 -16.140 18.975 
<< end >>
