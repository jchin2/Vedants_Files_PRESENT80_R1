magic
tech sky130A
magscale 1 2
timestamp 1671041739
<< xpolycontact >>
rect -512 69 -442 501
rect -512 -501 -442 -69
<< xpolyres >>
rect -512 -69 -442 69
<< viali >>
rect -494 447 -460 481
rect -494 375 -460 409
rect -494 303 -460 337
rect -494 231 -460 265
rect -494 159 -460 193
rect -494 87 -460 121
rect -494 -122 -460 -88
rect -494 -194 -460 -160
rect -494 -266 -460 -232
rect -494 -338 -460 -304
rect -494 -410 -460 -376
rect -494 -482 -460 -448
<< metal1 >>
rect -502 481 -452 495
rect -502 447 -494 481
rect -460 447 -452 481
rect -502 409 -452 447
rect -502 375 -494 409
rect -460 375 -452 409
rect -502 337 -452 375
rect -502 303 -494 337
rect -460 303 -452 337
rect -502 265 -452 303
rect -502 231 -494 265
rect -460 231 -452 265
rect -502 193 -452 231
rect -502 159 -494 193
rect -460 159 -452 193
rect -502 121 -452 159
rect -502 87 -494 121
rect -460 87 -452 121
rect -502 74 -452 87
rect -502 -88 -452 -74
rect -502 -122 -494 -88
rect -460 -122 -452 -88
rect -502 -160 -452 -122
rect -502 -194 -494 -160
rect -460 -194 -452 -160
rect -502 -232 -452 -194
rect -502 -266 -494 -232
rect -460 -266 -452 -232
rect -502 -304 -452 -266
rect -502 -338 -494 -304
rect -460 -338 -452 -304
rect -502 -376 -452 -338
rect -502 -410 -494 -376
rect -460 -410 -452 -376
rect -502 -448 -452 -410
rect -502 -482 -494 -448
rect -460 -482 -452 -448
rect -502 -495 -452 -482
<< end >>
