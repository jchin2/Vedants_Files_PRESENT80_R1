magic
tech sky130A
magscale 1 2
timestamp 1671306811
<< poly >>
rect -160 223 160 239
rect -160 189 -119 223
rect -85 189 -51 223
rect -17 189 17 223
rect 51 189 85 223
rect 119 189 160 223
rect -160 166 160 189
rect -160 -189 160 -166
rect -160 -223 -119 -189
rect -85 -223 -51 -189
rect -17 -223 17 -189
rect 51 -223 85 -189
rect 119 -223 160 -189
rect -160 -239 160 -223
<< polycont >>
rect -119 189 -85 223
rect -51 189 -17 223
rect 17 189 51 223
rect 85 189 119 223
rect -119 -223 -85 -189
rect -51 -223 -17 -189
rect 17 -223 51 -189
rect 85 -223 119 -189
<< npolyres >>
rect -160 -166 160 166
<< locali >>
rect -160 220 -119 223
rect -85 220 -51 223
rect -160 189 -125 220
rect -85 189 -53 220
rect -17 189 17 223
rect 51 220 85 223
rect 119 220 160 223
rect 53 189 85 220
rect 125 189 160 220
rect -144 186 -125 189
rect -91 186 -53 189
rect -19 186 19 189
rect 53 186 91 189
rect 125 186 144 189
rect -144 183 144 186
rect -144 -186 144 -183
rect -144 -189 -125 -186
rect -91 -189 -53 -186
rect -19 -189 19 -186
rect 53 -189 91 -186
rect 125 -189 144 -186
rect -160 -220 -125 -189
rect -85 -220 -53 -189
rect -160 -223 -119 -220
rect -85 -223 -51 -220
rect -17 -223 17 -189
rect 53 -220 85 -189
rect 125 -220 160 -189
rect 51 -223 85 -220
rect 119 -223 160 -220
<< viali >>
rect -125 189 -119 220
rect -119 189 -91 220
rect -53 189 -51 220
rect -51 189 -19 220
rect 19 189 51 220
rect 51 189 53 220
rect 91 189 119 220
rect 119 189 125 220
rect -125 186 -91 189
rect -53 186 -19 189
rect 19 186 53 189
rect 91 186 125 189
rect -125 -189 -91 -186
rect -53 -189 -19 -186
rect 19 -189 53 -186
rect 91 -189 125 -186
rect -125 -220 -119 -189
rect -119 -220 -91 -189
rect -53 -220 -51 -189
rect -51 -220 -19 -189
rect 19 -220 51 -189
rect 51 -220 53 -189
rect 91 -220 119 -189
rect 119 -220 125 -189
<< metal1 >>
rect -156 220 156 229
rect -156 186 -125 220
rect -91 186 -53 220
rect -19 186 19 220
rect 53 186 91 220
rect 125 186 156 220
rect -156 177 156 186
rect -156 -186 156 -177
rect -156 -220 -125 -186
rect -91 -220 -53 -186
rect -19 -220 19 -186
rect 53 -220 91 -186
rect 125 -220 156 -186
rect -156 -229 156 -220
<< end >>
