magic
tech sky130A
magscale 1 2
timestamp 1672683112
<< nwell >>
rect -3390 1760 -1900 1950
rect -3050 1370 -2230 1760
<< pwell >>
rect -3356 594 -1924 1186
<< nmos >>
rect -3210 860 -3180 1160
rect -2880 860 -2850 1160
rect -2730 860 -2700 1160
rect -2580 860 -2550 1160
rect -2430 860 -2400 1160
rect -2100 860 -2070 1160
<< pmos >>
rect -2880 1420 -2850 1720
rect -2730 1420 -2700 1720
rect -2580 1420 -2550 1720
rect -2430 1420 -2400 1720
<< ndiff >>
rect -3330 1087 -3210 1160
rect -3330 1053 -3287 1087
rect -3253 1053 -3210 1087
rect -3330 1007 -3210 1053
rect -3330 973 -3287 1007
rect -3253 973 -3210 1007
rect -3330 927 -3210 973
rect -3330 893 -3287 927
rect -3253 893 -3210 927
rect -3330 860 -3210 893
rect -3180 1087 -3060 1160
rect -3180 1053 -3137 1087
rect -3103 1053 -3060 1087
rect -3180 1007 -3060 1053
rect -3180 973 -3137 1007
rect -3103 973 -3060 1007
rect -3180 927 -3060 973
rect -3180 893 -3137 927
rect -3103 893 -3060 927
rect -3180 860 -3060 893
rect -3000 1087 -2880 1160
rect -3000 1053 -2957 1087
rect -2923 1053 -2880 1087
rect -3000 1007 -2880 1053
rect -3000 973 -2957 1007
rect -2923 973 -2880 1007
rect -3000 927 -2880 973
rect -3000 893 -2957 927
rect -2923 893 -2880 927
rect -3000 860 -2880 893
rect -2850 1087 -2730 1160
rect -2850 1053 -2807 1087
rect -2773 1053 -2730 1087
rect -2850 1007 -2730 1053
rect -2850 973 -2807 1007
rect -2773 973 -2730 1007
rect -2850 927 -2730 973
rect -2850 893 -2807 927
rect -2773 893 -2730 927
rect -2850 860 -2730 893
rect -2700 1087 -2580 1160
rect -2700 1053 -2657 1087
rect -2623 1053 -2580 1087
rect -2700 1007 -2580 1053
rect -2700 973 -2657 1007
rect -2623 973 -2580 1007
rect -2700 927 -2580 973
rect -2700 893 -2657 927
rect -2623 893 -2580 927
rect -2700 860 -2580 893
rect -2550 1087 -2430 1160
rect -2550 1053 -2507 1087
rect -2473 1053 -2430 1087
rect -2550 1007 -2430 1053
rect -2550 973 -2507 1007
rect -2473 973 -2430 1007
rect -2550 927 -2430 973
rect -2550 893 -2507 927
rect -2473 893 -2430 927
rect -2550 860 -2430 893
rect -2400 1087 -2280 1160
rect -2400 1053 -2357 1087
rect -2323 1053 -2280 1087
rect -2400 1007 -2280 1053
rect -2400 973 -2357 1007
rect -2323 973 -2280 1007
rect -2400 927 -2280 973
rect -2400 893 -2357 927
rect -2323 893 -2280 927
rect -2400 860 -2280 893
rect -2220 1087 -2100 1160
rect -2220 1053 -2177 1087
rect -2143 1053 -2100 1087
rect -2220 1007 -2100 1053
rect -2220 973 -2177 1007
rect -2143 973 -2100 1007
rect -2220 927 -2100 973
rect -2220 893 -2177 927
rect -2143 893 -2100 927
rect -2220 860 -2100 893
rect -2070 1087 -1950 1160
rect -2070 1053 -2027 1087
rect -1993 1053 -1950 1087
rect -2070 1007 -1950 1053
rect -2070 973 -2027 1007
rect -1993 973 -1950 1007
rect -2070 927 -1950 973
rect -2070 893 -2027 927
rect -1993 893 -1950 927
rect -2070 860 -1950 893
<< pdiff >>
rect -3000 1647 -2880 1720
rect -3000 1613 -2957 1647
rect -2923 1613 -2880 1647
rect -3000 1567 -2880 1613
rect -3000 1533 -2957 1567
rect -2923 1533 -2880 1567
rect -3000 1487 -2880 1533
rect -3000 1453 -2957 1487
rect -2923 1453 -2880 1487
rect -3000 1420 -2880 1453
rect -2850 1647 -2730 1720
rect -2850 1613 -2807 1647
rect -2773 1613 -2730 1647
rect -2850 1567 -2730 1613
rect -2850 1533 -2807 1567
rect -2773 1533 -2730 1567
rect -2850 1487 -2730 1533
rect -2850 1453 -2807 1487
rect -2773 1453 -2730 1487
rect -2850 1420 -2730 1453
rect -2700 1647 -2580 1720
rect -2700 1613 -2657 1647
rect -2623 1613 -2580 1647
rect -2700 1567 -2580 1613
rect -2700 1533 -2657 1567
rect -2623 1533 -2580 1567
rect -2700 1487 -2580 1533
rect -2700 1453 -2657 1487
rect -2623 1453 -2580 1487
rect -2700 1420 -2580 1453
rect -2550 1647 -2430 1720
rect -2550 1613 -2507 1647
rect -2473 1613 -2430 1647
rect -2550 1567 -2430 1613
rect -2550 1533 -2507 1567
rect -2473 1533 -2430 1567
rect -2550 1487 -2430 1533
rect -2550 1453 -2507 1487
rect -2473 1453 -2430 1487
rect -2550 1420 -2430 1453
rect -2400 1647 -2280 1720
rect -2400 1613 -2357 1647
rect -2323 1613 -2280 1647
rect -2400 1567 -2280 1613
rect -2400 1533 -2357 1567
rect -2323 1533 -2280 1567
rect -2400 1487 -2280 1533
rect -2400 1453 -2357 1487
rect -2323 1453 -2280 1487
rect -2400 1420 -2280 1453
<< ndiffc >>
rect -3287 1053 -3253 1087
rect -3287 973 -3253 1007
rect -3287 893 -3253 927
rect -3137 1053 -3103 1087
rect -3137 973 -3103 1007
rect -3137 893 -3103 927
rect -2957 1053 -2923 1087
rect -2957 973 -2923 1007
rect -2957 893 -2923 927
rect -2807 1053 -2773 1087
rect -2807 973 -2773 1007
rect -2807 893 -2773 927
rect -2657 1053 -2623 1087
rect -2657 973 -2623 1007
rect -2657 893 -2623 927
rect -2507 1053 -2473 1087
rect -2507 973 -2473 1007
rect -2507 893 -2473 927
rect -2357 1053 -2323 1087
rect -2357 973 -2323 1007
rect -2357 893 -2323 927
rect -2177 1053 -2143 1087
rect -2177 973 -2143 1007
rect -2177 893 -2143 927
rect -2027 1053 -1993 1087
rect -2027 973 -1993 1007
rect -2027 893 -1993 927
<< pdiffc >>
rect -2957 1613 -2923 1647
rect -2957 1533 -2923 1567
rect -2957 1453 -2923 1487
rect -2807 1613 -2773 1647
rect -2807 1533 -2773 1567
rect -2807 1453 -2773 1487
rect -2657 1613 -2623 1647
rect -2657 1533 -2623 1567
rect -2657 1453 -2623 1487
rect -2507 1613 -2473 1647
rect -2507 1533 -2473 1567
rect -2507 1453 -2473 1487
rect -2357 1613 -2323 1647
rect -2357 1533 -2323 1567
rect -2357 1453 -2323 1487
<< psubdiff >>
rect -3330 687 -1950 720
rect -3330 653 -3297 687
rect -3263 653 -3217 687
rect -3183 653 -3137 687
rect -3103 653 -3057 687
rect -3023 653 -2977 687
rect -2943 653 -2897 687
rect -2863 653 -2817 687
rect -2783 653 -2737 687
rect -2703 653 -2657 687
rect -2623 653 -2577 687
rect -2543 653 -2497 687
rect -2463 653 -2417 687
rect -2383 653 -2337 687
rect -2303 653 -2257 687
rect -2223 653 -2177 687
rect -2143 653 -2097 687
rect -2063 653 -2017 687
rect -1983 653 -1950 687
rect -3330 620 -1950 653
<< nsubdiff >>
rect -3330 1867 -1950 1900
rect -3330 1833 -3297 1867
rect -3263 1833 -3217 1867
rect -3183 1833 -3137 1867
rect -3103 1833 -3057 1867
rect -3023 1833 -2977 1867
rect -2943 1833 -2897 1867
rect -2863 1833 -2817 1867
rect -2783 1833 -2737 1867
rect -2703 1833 -2657 1867
rect -2623 1833 -2577 1867
rect -2543 1833 -2497 1867
rect -2463 1833 -2417 1867
rect -2383 1833 -2337 1867
rect -2303 1833 -2257 1867
rect -2223 1833 -2177 1867
rect -2143 1833 -2097 1867
rect -2063 1833 -2017 1867
rect -1983 1833 -1950 1867
rect -3330 1800 -1950 1833
<< psubdiffcont >>
rect -3297 653 -3263 687
rect -3217 653 -3183 687
rect -3137 653 -3103 687
rect -3057 653 -3023 687
rect -2977 653 -2943 687
rect -2897 653 -2863 687
rect -2817 653 -2783 687
rect -2737 653 -2703 687
rect -2657 653 -2623 687
rect -2577 653 -2543 687
rect -2497 653 -2463 687
rect -2417 653 -2383 687
rect -2337 653 -2303 687
rect -2257 653 -2223 687
rect -2177 653 -2143 687
rect -2097 653 -2063 687
rect -2017 653 -1983 687
<< nsubdiffcont >>
rect -3297 1833 -3263 1867
rect -3217 1833 -3183 1867
rect -3137 1833 -3103 1867
rect -3057 1833 -3023 1867
rect -2977 1833 -2943 1867
rect -2897 1833 -2863 1867
rect -2817 1833 -2783 1867
rect -2737 1833 -2703 1867
rect -2657 1833 -2623 1867
rect -2577 1833 -2543 1867
rect -2497 1833 -2463 1867
rect -2417 1833 -2383 1867
rect -2337 1833 -2303 1867
rect -2257 1833 -2223 1867
rect -2177 1833 -2143 1867
rect -2097 1833 -2063 1867
rect -2017 1833 -1983 1867
<< poly >>
rect -2880 1750 -2700 1780
rect -2880 1720 -2850 1750
rect -2730 1720 -2700 1750
rect -2580 1750 -2400 1780
rect -2580 1720 -2550 1750
rect -2430 1720 -2400 1750
rect -2100 1487 -2020 1510
rect -2100 1453 -2077 1487
rect -2043 1453 -2020 1487
rect -2100 1430 -2020 1453
rect -2880 1390 -2850 1420
rect -3260 1247 -3180 1270
rect -3260 1213 -3237 1247
rect -3203 1213 -3180 1247
rect -3260 1190 -3180 1213
rect -2730 1265 -2700 1420
rect -2580 1390 -2550 1420
rect -2430 1390 -2400 1420
rect -2630 1367 -2550 1390
rect -2630 1333 -2607 1367
rect -2573 1333 -2550 1367
rect -2630 1310 -2550 1333
rect -2730 1242 -2650 1265
rect -2730 1208 -2707 1242
rect -2673 1208 -2650 1242
rect -3210 1160 -3180 1190
rect -2880 1160 -2850 1190
rect -2730 1185 -2650 1208
rect -2730 1160 -2700 1185
rect -2580 1160 -2550 1310
rect -2430 1160 -2400 1190
rect -2100 1160 -2070 1430
rect -3210 830 -3180 860
rect -2880 830 -2850 860
rect -2730 830 -2700 860
rect -2580 830 -2550 860
rect -2430 830 -2400 860
rect -2100 830 -2070 860
rect -2880 807 -2800 830
rect -2880 773 -2857 807
rect -2823 773 -2800 807
rect -2880 750 -2800 773
rect -2480 807 -2400 830
rect -2480 773 -2457 807
rect -2423 773 -2400 807
rect -2480 750 -2400 773
<< polycont >>
rect -2077 1453 -2043 1487
rect -3237 1213 -3203 1247
rect -2607 1333 -2573 1367
rect -2707 1208 -2673 1242
rect -2857 773 -2823 807
rect -2457 773 -2423 807
<< locali >>
rect -3330 1867 -1950 1890
rect -3330 1833 -3297 1867
rect -3263 1833 -3217 1867
rect -3183 1833 -3137 1867
rect -3103 1833 -3057 1867
rect -3023 1833 -2977 1867
rect -2943 1833 -2897 1867
rect -2863 1833 -2817 1867
rect -2783 1833 -2737 1867
rect -2703 1833 -2657 1867
rect -2623 1833 -2577 1867
rect -2543 1833 -2497 1867
rect -2463 1833 -2417 1867
rect -2383 1833 -2337 1867
rect -2303 1833 -2257 1867
rect -2223 1833 -2177 1867
rect -2143 1833 -2097 1867
rect -2063 1833 -2017 1867
rect -1983 1833 -1950 1867
rect -3330 1810 -1950 1833
rect -2980 1647 -2900 1680
rect -2980 1613 -2957 1647
rect -2923 1613 -2900 1647
rect -2980 1567 -2900 1613
rect -2980 1533 -2957 1567
rect -2923 1533 -2900 1567
rect -3130 1490 -3050 1510
rect -3330 1487 -3050 1490
rect -3330 1453 -3107 1487
rect -3073 1453 -3050 1487
rect -3330 1450 -3050 1453
rect -3130 1430 -3050 1450
rect -2980 1487 -2900 1533
rect -2980 1453 -2957 1487
rect -2923 1453 -2900 1487
rect -2980 1430 -2900 1453
rect -2830 1647 -2750 1680
rect -2830 1613 -2807 1647
rect -2773 1613 -2750 1647
rect -2830 1567 -2750 1613
rect -2830 1533 -2807 1567
rect -2773 1533 -2750 1567
rect -2830 1487 -2750 1533
rect -2830 1453 -2807 1487
rect -2773 1453 -2750 1487
rect -2830 1420 -2750 1453
rect -2680 1647 -2600 1680
rect -2680 1613 -2657 1647
rect -2623 1613 -2600 1647
rect -2680 1567 -2600 1613
rect -2680 1533 -2657 1567
rect -2623 1533 -2600 1567
rect -2680 1487 -2600 1533
rect -2680 1453 -2657 1487
rect -2623 1453 -2600 1487
rect -2680 1430 -2600 1453
rect -2530 1647 -2450 1680
rect -2530 1613 -2507 1647
rect -2473 1613 -2450 1647
rect -2530 1567 -2450 1613
rect -2530 1533 -2507 1567
rect -2473 1533 -2450 1567
rect -2530 1487 -2450 1533
rect -2530 1453 -2507 1487
rect -2473 1453 -2450 1487
rect -2530 1420 -2450 1453
rect -2380 1647 -2300 1680
rect -2380 1613 -2357 1647
rect -2323 1613 -2300 1647
rect -2380 1567 -2300 1613
rect -2380 1533 -2357 1567
rect -2323 1533 -2300 1567
rect -2380 1487 -2300 1533
rect -2380 1453 -2357 1487
rect -2323 1453 -2300 1487
rect -2380 1430 -2300 1453
rect -2230 1490 -2150 1510
rect -2100 1490 -2020 1510
rect -2230 1487 -2020 1490
rect -2230 1453 -2207 1487
rect -2173 1453 -2077 1487
rect -2043 1453 -2020 1487
rect -2230 1450 -2020 1453
rect -2230 1430 -2150 1450
rect -2100 1430 -2020 1450
rect -2810 1370 -2770 1420
rect -2630 1370 -2550 1390
rect -2810 1367 -2550 1370
rect -2810 1333 -2607 1367
rect -2573 1333 -2550 1367
rect -2810 1330 -2550 1333
rect -3260 1250 -3180 1270
rect -3330 1247 -3180 1250
rect -3330 1213 -3237 1247
rect -3203 1213 -3180 1247
rect -3330 1210 -3180 1213
rect -3260 1190 -3180 1210
rect -2810 1200 -2770 1330
rect -2630 1310 -2550 1330
rect -3140 1160 -2770 1200
rect -2730 1250 -2650 1265
rect -2510 1250 -2470 1420
rect -2230 1370 -2150 1390
rect -2230 1367 -1950 1370
rect -2230 1333 -2207 1367
rect -2173 1333 -1950 1367
rect -2230 1330 -1950 1333
rect -2230 1310 -2150 1330
rect -2730 1242 -2470 1250
rect -2730 1208 -2707 1242
rect -2673 1210 -2470 1242
rect -2673 1208 -2650 1210
rect -2730 1185 -2650 1208
rect -2510 1200 -2470 1210
rect -2510 1160 -1950 1200
rect -3140 1120 -3100 1160
rect -2810 1120 -2770 1160
rect -3310 1087 -3230 1120
rect -3310 1053 -3287 1087
rect -3253 1053 -3230 1087
rect -3310 1007 -3230 1053
rect -3310 973 -3287 1007
rect -3253 973 -3230 1007
rect -3310 927 -3230 973
rect -3310 893 -3287 927
rect -3253 893 -3230 927
rect -3310 870 -3230 893
rect -3160 1087 -3080 1120
rect -3160 1053 -3137 1087
rect -3103 1053 -3080 1087
rect -3160 1007 -3080 1053
rect -3160 973 -3137 1007
rect -3103 973 -3080 1007
rect -3160 927 -3080 973
rect -3160 893 -3137 927
rect -3103 893 -3080 927
rect -3160 870 -3080 893
rect -2980 1087 -2900 1120
rect -2980 1053 -2957 1087
rect -2923 1053 -2900 1087
rect -2980 1007 -2900 1053
rect -2980 973 -2957 1007
rect -2923 973 -2900 1007
rect -2980 927 -2900 973
rect -2980 893 -2957 927
rect -2923 893 -2900 927
rect -2980 870 -2900 893
rect -2830 1087 -2750 1120
rect -2830 1053 -2807 1087
rect -2773 1053 -2750 1087
rect -2830 1007 -2750 1053
rect -2830 973 -2807 1007
rect -2773 973 -2750 1007
rect -2830 927 -2750 973
rect -2830 893 -2807 927
rect -2773 893 -2750 927
rect -2830 870 -2750 893
rect -2680 1087 -2600 1120
rect -2680 1053 -2657 1087
rect -2623 1053 -2600 1087
rect -2680 1007 -2600 1053
rect -2680 973 -2657 1007
rect -2623 973 -2600 1007
rect -2680 927 -2600 973
rect -2680 893 -2657 927
rect -2623 893 -2600 927
rect -2680 870 -2600 893
rect -2530 1087 -2450 1160
rect -2180 1120 -2140 1160
rect -2530 1053 -2507 1087
rect -2473 1053 -2450 1087
rect -2530 1007 -2450 1053
rect -2530 973 -2507 1007
rect -2473 973 -2450 1007
rect -2530 927 -2450 973
rect -2530 893 -2507 927
rect -2473 893 -2450 927
rect -2530 870 -2450 893
rect -2380 1087 -2300 1120
rect -2380 1053 -2357 1087
rect -2323 1053 -2300 1087
rect -2380 1007 -2300 1053
rect -2380 973 -2357 1007
rect -2323 973 -2300 1007
rect -2380 927 -2300 973
rect -2380 893 -2357 927
rect -2323 893 -2300 927
rect -2380 870 -2300 893
rect -2200 1087 -2120 1120
rect -2200 1053 -2177 1087
rect -2143 1053 -2120 1087
rect -2200 1007 -2120 1053
rect -2200 973 -2177 1007
rect -2143 973 -2120 1007
rect -2200 927 -2120 973
rect -2200 893 -2177 927
rect -2143 893 -2120 927
rect -2200 870 -2120 893
rect -2050 1087 -1970 1120
rect -2050 1053 -2027 1087
rect -1993 1053 -1970 1087
rect -2050 1007 -1970 1053
rect -2050 973 -2027 1007
rect -1993 973 -1970 1007
rect -2050 927 -1970 973
rect -2050 893 -2027 927
rect -1993 893 -1970 927
rect -2050 870 -1970 893
rect -2880 810 -2800 830
rect -2480 810 -2400 830
rect -3330 807 -2400 810
rect -3330 773 -2857 807
rect -2823 773 -2457 807
rect -2423 773 -2400 807
rect -3330 770 -2400 773
rect -2880 750 -2800 770
rect -2480 750 -2400 770
rect -3330 687 -1950 710
rect -3330 653 -3297 687
rect -3263 653 -3217 687
rect -3183 653 -3137 687
rect -3103 653 -3057 687
rect -3023 653 -2977 687
rect -2943 653 -2897 687
rect -2863 653 -2817 687
rect -2783 653 -2737 687
rect -2703 653 -2657 687
rect -2623 653 -2577 687
rect -2543 653 -2497 687
rect -2463 653 -2417 687
rect -2383 653 -2337 687
rect -2303 653 -2257 687
rect -2223 653 -2177 687
rect -2143 653 -2097 687
rect -2063 653 -2017 687
rect -1983 653 -1950 687
rect -3330 630 -1950 653
<< viali >>
rect -3297 1833 -3263 1867
rect -3217 1833 -3183 1867
rect -3137 1833 -3103 1867
rect -3057 1833 -3023 1867
rect -2977 1833 -2943 1867
rect -2897 1833 -2863 1867
rect -2817 1833 -2783 1867
rect -2737 1833 -2703 1867
rect -2657 1833 -2623 1867
rect -2577 1833 -2543 1867
rect -2497 1833 -2463 1867
rect -2417 1833 -2383 1867
rect -2337 1833 -2303 1867
rect -2257 1833 -2223 1867
rect -2177 1833 -2143 1867
rect -2097 1833 -2063 1867
rect -2017 1833 -1983 1867
rect -2957 1613 -2923 1647
rect -2957 1533 -2923 1567
rect -3107 1453 -3073 1487
rect -2957 1453 -2923 1487
rect -2657 1613 -2623 1647
rect -2657 1533 -2623 1567
rect -2657 1453 -2623 1487
rect -2357 1613 -2323 1647
rect -2357 1533 -2323 1567
rect -2357 1453 -2323 1487
rect -2207 1453 -2173 1487
rect -2607 1333 -2573 1367
rect -2207 1333 -2173 1367
rect -3287 1053 -3253 1087
rect -3287 973 -3253 1007
rect -3287 893 -3253 927
rect -2957 1053 -2923 1087
rect -2957 973 -2923 1007
rect -2957 893 -2923 927
rect -2657 1053 -2623 1087
rect -2657 973 -2623 1007
rect -2657 893 -2623 927
rect -2357 1053 -2323 1087
rect -2357 973 -2323 1007
rect -2357 893 -2323 927
rect -2027 1053 -1993 1087
rect -2027 973 -1993 1007
rect -2027 893 -1993 927
rect -3297 653 -3263 687
rect -3217 653 -3183 687
rect -3137 653 -3103 687
rect -3057 653 -3023 687
rect -2977 653 -2943 687
rect -2897 653 -2863 687
rect -2817 653 -2783 687
rect -2737 653 -2703 687
rect -2657 653 -2623 687
rect -2577 653 -2543 687
rect -2497 653 -2463 687
rect -2417 653 -2383 687
rect -2337 653 -2303 687
rect -2257 653 -2223 687
rect -2177 653 -2143 687
rect -2097 653 -2063 687
rect -2017 653 -1983 687
<< metal1 >>
rect -3330 1867 -1950 1900
rect -3330 1833 -3297 1867
rect -3263 1833 -3217 1867
rect -3183 1833 -3137 1867
rect -3103 1833 -3057 1867
rect -3023 1833 -2977 1867
rect -2943 1833 -2897 1867
rect -2863 1833 -2817 1867
rect -2783 1833 -2737 1867
rect -2703 1833 -2657 1867
rect -2623 1833 -2577 1867
rect -2543 1833 -2497 1867
rect -2463 1833 -2417 1867
rect -2383 1833 -2337 1867
rect -2303 1833 -2257 1867
rect -2223 1833 -2177 1867
rect -2143 1833 -2097 1867
rect -2063 1833 -2017 1867
rect -1983 1833 -1950 1867
rect -3330 1800 -1950 1833
rect -3310 1087 -3230 1800
rect -2980 1647 -2900 1800
rect -2980 1613 -2957 1647
rect -2923 1613 -2900 1647
rect -2980 1567 -2900 1613
rect -2980 1533 -2957 1567
rect -2923 1533 -2900 1567
rect -3130 1496 -3050 1510
rect -3130 1444 -3116 1496
rect -3064 1444 -3050 1496
rect -3130 1430 -3050 1444
rect -2980 1487 -2900 1533
rect -2980 1453 -2957 1487
rect -2923 1453 -2900 1487
rect -2980 1430 -2900 1453
rect -2680 1647 -2600 1800
rect -2680 1613 -2657 1647
rect -2623 1613 -2600 1647
rect -2680 1567 -2600 1613
rect -2680 1533 -2657 1567
rect -2623 1533 -2600 1567
rect -2680 1487 -2600 1533
rect -2680 1453 -2657 1487
rect -2623 1453 -2600 1487
rect -2680 1430 -2600 1453
rect -2380 1647 -2300 1800
rect -2380 1613 -2357 1647
rect -2323 1613 -2300 1647
rect -2380 1567 -2300 1613
rect -2380 1533 -2357 1567
rect -2323 1533 -2300 1567
rect -2380 1487 -2300 1533
rect -2380 1453 -2357 1487
rect -2323 1453 -2300 1487
rect -2380 1430 -2300 1453
rect -2230 1496 -2150 1510
rect -2230 1444 -2216 1496
rect -2164 1444 -2150 1496
rect -2230 1430 -2150 1444
rect -2630 1370 -2550 1390
rect -2230 1370 -2150 1390
rect -2630 1367 -2150 1370
rect -2630 1333 -2607 1367
rect -2573 1333 -2207 1367
rect -2173 1333 -2150 1367
rect -2630 1330 -2150 1333
rect -2630 1310 -2550 1330
rect -2230 1310 -2150 1330
rect -3310 1053 -3287 1087
rect -3253 1053 -3230 1087
rect -3310 1007 -3230 1053
rect -3310 973 -3287 1007
rect -3253 973 -3230 1007
rect -3310 927 -3230 973
rect -3310 893 -3287 927
rect -3253 893 -3230 927
rect -3310 870 -3230 893
rect -2980 1087 -2900 1120
rect -2980 1053 -2957 1087
rect -2923 1053 -2900 1087
rect -2980 1007 -2900 1053
rect -2980 973 -2957 1007
rect -2923 973 -2900 1007
rect -2980 927 -2900 973
rect -2980 893 -2957 927
rect -2923 893 -2900 927
rect -2980 870 -2900 893
rect -2680 1087 -2600 1120
rect -2680 1053 -2657 1087
rect -2623 1053 -2600 1087
rect -2680 1007 -2600 1053
rect -2680 973 -2657 1007
rect -2623 973 -2600 1007
rect -2680 927 -2600 973
rect -2680 893 -2657 927
rect -2623 893 -2600 927
rect -2680 870 -2600 893
rect -2380 1087 -2300 1120
rect -2380 1053 -2357 1087
rect -2323 1053 -2300 1087
rect -2380 1007 -2300 1053
rect -2380 973 -2357 1007
rect -2323 973 -2300 1007
rect -2380 927 -2300 973
rect -2380 893 -2357 927
rect -2323 893 -2300 927
rect -2380 870 -2300 893
rect -2050 1087 -1970 1800
rect -2050 1053 -2027 1087
rect -1993 1053 -1970 1087
rect -2050 1007 -1970 1053
rect -2050 973 -2027 1007
rect -1993 973 -1970 1007
rect -2050 927 -1970 973
rect -2050 893 -2027 927
rect -1993 893 -1970 927
rect -2050 870 -1970 893
rect -2960 720 -2920 870
rect -2660 720 -2620 870
rect -2360 720 -2320 870
rect -3330 687 -1950 720
rect -3330 653 -3297 687
rect -3263 653 -3217 687
rect -3183 653 -3137 687
rect -3103 653 -3057 687
rect -3023 653 -2977 687
rect -2943 653 -2897 687
rect -2863 653 -2817 687
rect -2783 653 -2737 687
rect -2703 653 -2657 687
rect -2623 653 -2577 687
rect -2543 653 -2497 687
rect -2463 653 -2417 687
rect -2383 653 -2337 687
rect -2303 653 -2257 687
rect -2223 653 -2177 687
rect -2143 653 -2097 687
rect -2063 653 -2017 687
rect -1983 653 -1950 687
rect -3330 620 -1950 653
<< via1 >>
rect -3116 1487 -3064 1496
rect -3116 1453 -3107 1487
rect -3107 1453 -3073 1487
rect -3073 1453 -3064 1487
rect -3116 1444 -3064 1453
rect -2216 1487 -2164 1496
rect -2216 1453 -2207 1487
rect -2207 1453 -2173 1487
rect -2173 1453 -2164 1487
rect -2216 1444 -2164 1453
<< metal2 >>
rect -3130 1496 -3050 1510
rect -3130 1444 -3116 1496
rect -3064 1490 -3050 1496
rect -2230 1496 -2150 1510
rect -2230 1490 -2216 1496
rect -3064 1450 -2216 1490
rect -3064 1444 -3050 1450
rect -3130 1430 -3050 1444
rect -2230 1444 -2216 1450
rect -2164 1444 -2150 1496
rect -2230 1430 -2150 1444
<< labels >>
rlabel locali s -2710 1205 -2670 1245 4 OUT_bar
port 1 nsew
rlabel locali s -2080 1450 -2040 1490 4 A
port 2 nsew
rlabel locali s -3240 1210 -3200 1250 4 A_bar
port 3 nsew
rlabel locali s -2860 770 -2820 810 4 Dis
port 4 nsew
rlabel metal1 s -2610 1330 -2570 1370 4 OUT
port 5 nsew
rlabel metal1 s -2660 650 -2620 690 4 GND!
port 6 nsew
rlabel metal1 s -2660 1830 -2620 1870 4 CLK
port 7 nsew
<< end >>
