* NGSPICE file created from EESPFAL_4in_NAND_magic_checked.ext - technology: sky130A

.subckt EESPFAL_4in_NAND_magic_checked OUT A A_bar B B_bar C C_bar D D_bar Dis OUT_bar
+ GND CLK
X0 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=3.6e+12p pd=1.68e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X1 CLK B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=8.5e+12p pd=3.68e+07u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n1040_180# B a_n1190_180# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 OUT_bar OUT CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u M=2
X4 CLK D_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n1340_180# D OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT_bar A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar C_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X11 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK A a_n1040_180# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_n1190_180# C a_n1340_180# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

