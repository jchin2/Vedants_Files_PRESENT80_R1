magic
tech sky130A
timestamp 1666311795
<< nwell >>
rect -1385 905 -75 995
rect -870 540 -600 905
<< nmos >>
rect -1240 285 -1225 435
rect -1165 285 -1150 435
rect -1090 285 -1075 435
rect -1015 285 -1000 435
rect -850 285 -835 435
rect -775 285 -760 435
rect -700 285 -685 435
rect -625 285 -610 435
rect -460 285 -445 435
rect -385 285 -370 435
rect -310 285 -295 435
rect -235 285 -220 435
<< pmos >>
rect -775 565 -760 865
rect -700 565 -685 865
<< ndiff >>
rect -1300 400 -1240 435
rect -1300 380 -1280 400
rect -1260 380 -1240 400
rect -1300 360 -1240 380
rect -1300 340 -1280 360
rect -1260 340 -1240 360
rect -1300 320 -1240 340
rect -1300 300 -1280 320
rect -1260 300 -1240 320
rect -1300 285 -1240 300
rect -1225 285 -1165 435
rect -1150 400 -1090 435
rect -1150 380 -1130 400
rect -1110 380 -1090 400
rect -1150 360 -1090 380
rect -1150 340 -1130 360
rect -1110 340 -1090 360
rect -1150 320 -1090 340
rect -1150 300 -1130 320
rect -1110 300 -1090 320
rect -1150 285 -1090 300
rect -1075 285 -1015 435
rect -1000 400 -940 435
rect -1000 380 -980 400
rect -960 380 -940 400
rect -1000 360 -940 380
rect -1000 340 -980 360
rect -960 340 -940 360
rect -1000 320 -940 340
rect -1000 300 -980 320
rect -960 300 -940 320
rect -1000 285 -940 300
rect -910 400 -850 435
rect -910 380 -890 400
rect -870 380 -850 400
rect -910 360 -850 380
rect -910 340 -890 360
rect -870 340 -850 360
rect -910 320 -850 340
rect -910 300 -890 320
rect -870 300 -850 320
rect -910 285 -850 300
rect -835 400 -775 435
rect -835 380 -815 400
rect -795 380 -775 400
rect -835 360 -775 380
rect -835 340 -815 360
rect -795 340 -775 360
rect -835 320 -775 340
rect -835 300 -815 320
rect -795 300 -775 320
rect -835 285 -775 300
rect -760 400 -700 435
rect -760 380 -740 400
rect -720 380 -700 400
rect -760 360 -700 380
rect -760 340 -740 360
rect -720 340 -700 360
rect -760 320 -700 340
rect -760 300 -740 320
rect -720 300 -700 320
rect -760 285 -700 300
rect -685 400 -625 435
rect -685 380 -665 400
rect -645 380 -625 400
rect -685 360 -625 380
rect -685 340 -665 360
rect -645 340 -625 360
rect -685 320 -625 340
rect -685 300 -665 320
rect -645 300 -625 320
rect -685 285 -625 300
rect -610 400 -550 435
rect -610 380 -590 400
rect -570 380 -550 400
rect -610 360 -550 380
rect -610 340 -590 360
rect -570 340 -550 360
rect -610 320 -550 340
rect -610 300 -590 320
rect -570 300 -550 320
rect -610 285 -550 300
rect -520 400 -460 435
rect -520 380 -500 400
rect -480 380 -460 400
rect -520 360 -460 380
rect -520 340 -500 360
rect -480 340 -460 360
rect -520 320 -460 340
rect -520 300 -500 320
rect -480 300 -460 320
rect -520 285 -460 300
rect -445 285 -385 435
rect -370 400 -310 435
rect -370 380 -350 400
rect -330 380 -310 400
rect -370 360 -310 380
rect -370 340 -350 360
rect -330 340 -310 360
rect -370 320 -310 340
rect -370 300 -350 320
rect -330 300 -310 320
rect -370 285 -310 300
rect -295 285 -235 435
rect -220 400 -160 435
rect -220 380 -200 400
rect -180 380 -160 400
rect -220 360 -160 380
rect -220 340 -200 360
rect -180 340 -160 360
rect -220 320 -160 340
rect -220 300 -200 320
rect -180 300 -160 320
rect -220 285 -160 300
<< pdiff >>
rect -835 840 -775 865
rect -835 820 -815 840
rect -795 820 -775 840
rect -835 800 -775 820
rect -835 780 -815 800
rect -795 780 -775 800
rect -835 760 -775 780
rect -835 740 -815 760
rect -795 740 -775 760
rect -835 720 -775 740
rect -835 700 -815 720
rect -795 700 -775 720
rect -835 680 -775 700
rect -835 660 -815 680
rect -795 660 -775 680
rect -835 640 -775 660
rect -835 620 -815 640
rect -795 620 -775 640
rect -835 600 -775 620
rect -835 580 -815 600
rect -795 580 -775 600
rect -835 565 -775 580
rect -760 840 -700 865
rect -760 820 -740 840
rect -720 820 -700 840
rect -760 800 -700 820
rect -760 780 -740 800
rect -720 780 -700 800
rect -760 760 -700 780
rect -760 740 -740 760
rect -720 740 -700 760
rect -760 720 -700 740
rect -760 700 -740 720
rect -720 700 -700 720
rect -760 680 -700 700
rect -760 660 -740 680
rect -720 660 -700 680
rect -760 640 -700 660
rect -760 620 -740 640
rect -720 620 -700 640
rect -760 600 -700 620
rect -760 580 -740 600
rect -720 580 -700 600
rect -760 565 -700 580
rect -685 840 -625 865
rect -685 820 -665 840
rect -645 820 -625 840
rect -685 800 -625 820
rect -685 780 -665 800
rect -645 780 -625 800
rect -685 760 -625 780
rect -685 740 -665 760
rect -645 740 -625 760
rect -685 720 -625 740
rect -685 700 -665 720
rect -645 700 -625 720
rect -685 680 -625 700
rect -685 660 -665 680
rect -645 660 -625 680
rect -685 640 -625 660
rect -685 620 -665 640
rect -645 620 -625 640
rect -685 600 -625 620
rect -685 580 -665 600
rect -645 580 -625 600
rect -685 565 -625 580
<< ndiffc >>
rect -1280 380 -1260 400
rect -1280 340 -1260 360
rect -1280 300 -1260 320
rect -1130 380 -1110 400
rect -1130 340 -1110 360
rect -1130 300 -1110 320
rect -980 380 -960 400
rect -980 340 -960 360
rect -980 300 -960 320
rect -890 380 -870 400
rect -890 340 -870 360
rect -890 300 -870 320
rect -815 380 -795 400
rect -815 340 -795 360
rect -815 300 -795 320
rect -740 380 -720 400
rect -740 340 -720 360
rect -740 300 -720 320
rect -665 380 -645 400
rect -665 340 -645 360
rect -665 300 -645 320
rect -590 380 -570 400
rect -590 340 -570 360
rect -590 300 -570 320
rect -500 380 -480 400
rect -500 340 -480 360
rect -500 300 -480 320
rect -350 380 -330 400
rect -350 340 -330 360
rect -350 300 -330 320
rect -200 380 -180 400
rect -200 340 -180 360
rect -200 300 -180 320
<< pdiffc >>
rect -815 820 -795 840
rect -815 780 -795 800
rect -815 740 -795 760
rect -815 700 -795 720
rect -815 660 -795 680
rect -815 620 -795 640
rect -815 580 -795 600
rect -740 820 -720 840
rect -740 780 -720 800
rect -740 740 -720 760
rect -740 700 -720 720
rect -740 660 -720 680
rect -740 620 -720 640
rect -740 580 -720 600
rect -665 820 -645 840
rect -665 780 -645 800
rect -665 740 -645 760
rect -665 700 -645 720
rect -665 660 -645 680
rect -665 620 -645 640
rect -665 580 -645 600
<< psubdiff >>
rect -1360 400 -1300 435
rect -1360 380 -1340 400
rect -1320 380 -1300 400
rect -1360 360 -1300 380
rect -1360 340 -1340 360
rect -1320 340 -1300 360
rect -1360 320 -1300 340
rect -1360 300 -1340 320
rect -1320 300 -1300 320
rect -1360 285 -1300 300
rect -160 400 -100 435
rect -160 380 -140 400
rect -120 380 -100 400
rect -160 360 -100 380
rect -160 340 -140 360
rect -120 340 -100 360
rect -160 320 -100 340
rect -160 300 -140 320
rect -120 300 -100 320
rect -160 285 -100 300
rect -1380 -10 -75 5
rect -1380 -30 -1360 -10
rect -1340 -30 -1320 -10
rect -1300 -30 -1280 -10
rect -1260 -30 -1240 -10
rect -1220 -30 -1200 -10
rect -1180 -30 -1160 -10
rect -1140 -30 -1120 -10
rect -1100 -30 -1080 -10
rect -1060 -30 -1040 -10
rect -1020 -30 -1000 -10
rect -980 -30 -960 -10
rect -940 -30 -920 -10
rect -900 -30 -880 -10
rect -860 -30 -840 -10
rect -820 -30 -800 -10
rect -780 -30 -760 -10
rect -740 -30 -720 -10
rect -700 -30 -680 -10
rect -660 -30 -635 -10
rect -615 -30 -595 -10
rect -575 -30 -555 -10
rect -535 -30 -515 -10
rect -495 -30 -475 -10
rect -455 -30 -435 -10
rect -415 -30 -395 -10
rect -375 -30 -355 -10
rect -335 -30 -315 -10
rect -295 -30 -275 -10
rect -255 -30 -235 -10
rect -215 -30 -195 -10
rect -175 -30 -155 -10
rect -135 -30 -115 -10
rect -95 -30 -75 -10
rect -1380 -45 -75 -30
<< nsubdiff >>
rect -1365 960 -95 975
rect -1365 940 -1345 960
rect -1325 940 -1305 960
rect -1285 940 -1265 960
rect -1245 940 -1225 960
rect -1205 940 -1185 960
rect -1165 940 -1140 960
rect -1120 940 -1100 960
rect -1080 940 -1060 960
rect -1040 940 -1020 960
rect -1000 940 -980 960
rect -960 940 -940 960
rect -920 940 -900 960
rect -880 940 -860 960
rect -840 940 -820 960
rect -800 940 -780 960
rect -760 940 -740 960
rect -720 940 -700 960
rect -680 940 -660 960
rect -640 940 -620 960
rect -600 940 -580 960
rect -560 940 -540 960
rect -520 940 -500 960
rect -480 940 -455 960
rect -435 940 -415 960
rect -395 940 -375 960
rect -355 940 -335 960
rect -315 940 -295 960
rect -275 940 -255 960
rect -235 940 -215 960
rect -195 940 -175 960
rect -155 940 -135 960
rect -115 940 -95 960
rect -1365 925 -95 940
<< psubdiffcont >>
rect -1340 380 -1320 400
rect -1340 340 -1320 360
rect -1340 300 -1320 320
rect -140 380 -120 400
rect -140 340 -120 360
rect -140 300 -120 320
rect -1360 -30 -1340 -10
rect -1320 -30 -1300 -10
rect -1280 -30 -1260 -10
rect -1240 -30 -1220 -10
rect -1200 -30 -1180 -10
rect -1160 -30 -1140 -10
rect -1120 -30 -1100 -10
rect -1080 -30 -1060 -10
rect -1040 -30 -1020 -10
rect -1000 -30 -980 -10
rect -960 -30 -940 -10
rect -920 -30 -900 -10
rect -880 -30 -860 -10
rect -840 -30 -820 -10
rect -800 -30 -780 -10
rect -760 -30 -740 -10
rect -720 -30 -700 -10
rect -680 -30 -660 -10
rect -635 -30 -615 -10
rect -595 -30 -575 -10
rect -555 -30 -535 -10
rect -515 -30 -495 -10
rect -475 -30 -455 -10
rect -435 -30 -415 -10
rect -395 -30 -375 -10
rect -355 -30 -335 -10
rect -315 -30 -295 -10
rect -275 -30 -255 -10
rect -235 -30 -215 -10
rect -195 -30 -175 -10
rect -155 -30 -135 -10
rect -115 -30 -95 -10
<< nsubdiffcont >>
rect -1345 940 -1325 960
rect -1305 940 -1285 960
rect -1265 940 -1245 960
rect -1225 940 -1205 960
rect -1185 940 -1165 960
rect -1140 940 -1120 960
rect -1100 940 -1080 960
rect -1060 940 -1040 960
rect -1020 940 -1000 960
rect -980 940 -960 960
rect -940 940 -920 960
rect -900 940 -880 960
rect -860 940 -840 960
rect -820 940 -800 960
rect -780 940 -760 960
rect -740 940 -720 960
rect -700 940 -680 960
rect -660 940 -640 960
rect -620 940 -600 960
rect -580 940 -560 960
rect -540 940 -520 960
rect -500 940 -480 960
rect -455 940 -435 960
rect -415 940 -395 960
rect -375 940 -355 960
rect -335 940 -315 960
rect -295 940 -275 960
rect -255 940 -235 960
rect -215 940 -195 960
rect -175 940 -155 960
rect -135 940 -115 960
<< poly >>
rect -775 865 -760 880
rect -700 865 -685 880
rect -775 490 -760 565
rect -700 550 -685 565
rect -725 540 -685 550
rect -725 520 -715 540
rect -695 520 -685 540
rect -725 510 -685 520
rect -775 480 -735 490
rect -775 460 -765 480
rect -745 460 -735 480
rect -775 450 -735 460
rect -1240 435 -1225 450
rect -1165 435 -1150 450
rect -1090 435 -1075 450
rect -1015 435 -1000 450
rect -850 435 -835 450
rect -775 435 -760 450
rect -700 435 -685 510
rect -625 435 -610 450
rect -460 435 -445 450
rect -385 435 -370 450
rect -310 435 -295 450
rect -235 435 -220 450
rect -1240 60 -1225 285
rect -1165 165 -1150 285
rect -1090 220 -1075 285
rect -1090 210 -1050 220
rect -1090 190 -1080 210
rect -1060 190 -1050 210
rect -1090 180 -1050 190
rect -1165 155 -1125 165
rect -1165 135 -1155 155
rect -1135 135 -1125 155
rect -1165 125 -1125 135
rect -1015 115 -1000 285
rect -850 270 -835 285
rect -775 270 -760 285
rect -700 270 -685 285
rect -625 270 -610 285
rect -850 260 -810 270
rect -850 240 -840 260
rect -820 240 -810 260
rect -850 230 -810 240
rect -650 260 -610 270
rect -650 240 -640 260
rect -620 240 -610 260
rect -650 230 -610 240
rect -1015 105 -975 115
rect -1015 85 -1005 105
rect -985 85 -975 105
rect -1015 75 -975 85
rect -460 60 -445 285
rect -385 220 -370 285
rect -385 210 -345 220
rect -385 190 -375 210
rect -355 190 -345 210
rect -385 180 -345 190
rect -310 165 -295 285
rect -310 155 -270 165
rect -310 135 -300 155
rect -280 135 -270 155
rect -310 125 -270 135
rect -235 115 -220 285
rect -235 105 -195 115
rect -235 85 -225 105
rect -205 85 -195 105
rect -235 75 -195 85
rect -1240 50 -1200 60
rect -1240 30 -1230 50
rect -1210 30 -1200 50
rect -1240 20 -1200 30
rect -460 50 -420 60
rect -460 30 -450 50
rect -430 30 -420 50
rect -460 20 -420 30
<< polycont >>
rect -715 520 -695 540
rect -765 460 -745 480
rect -1080 190 -1060 210
rect -1155 135 -1135 155
rect -840 240 -820 260
rect -640 240 -620 260
rect -1005 85 -985 105
rect -375 190 -355 210
rect -300 135 -280 155
rect -225 85 -205 105
rect -1230 30 -1210 50
rect -450 30 -430 50
<< locali >>
rect -1365 960 -95 970
rect -1365 940 -1345 960
rect -1325 940 -1305 960
rect -1285 940 -1265 960
rect -1245 940 -1225 960
rect -1205 940 -1185 960
rect -1165 940 -1140 960
rect -1120 940 -1100 960
rect -1080 940 -1060 960
rect -1040 940 -1020 960
rect -1000 940 -980 960
rect -960 940 -940 960
rect -920 940 -900 960
rect -880 940 -860 960
rect -840 940 -820 960
rect -800 940 -780 960
rect -760 940 -740 960
rect -720 940 -700 960
rect -680 940 -660 960
rect -640 940 -620 960
rect -600 940 -580 960
rect -560 940 -540 960
rect -520 940 -500 960
rect -480 940 -455 960
rect -435 940 -415 960
rect -395 940 -375 960
rect -355 940 -335 960
rect -315 940 -295 960
rect -275 940 -255 960
rect -235 940 -215 960
rect -195 940 -175 960
rect -155 940 -135 960
rect -115 940 -95 960
rect -1365 930 -95 940
rect -825 840 -785 850
rect -825 820 -815 840
rect -795 820 -785 840
rect -825 800 -785 820
rect -825 780 -815 800
rect -795 780 -785 800
rect -825 760 -785 780
rect -825 740 -815 760
rect -795 740 -785 760
rect -825 720 -785 740
rect -825 700 -815 720
rect -795 700 -785 720
rect -825 680 -785 700
rect -825 660 -815 680
rect -795 660 -785 680
rect -825 640 -785 660
rect -825 620 -815 640
rect -795 620 -785 640
rect -825 600 -785 620
rect -825 580 -815 600
rect -795 580 -785 600
rect -825 565 -785 580
rect -750 840 -710 850
rect -750 820 -740 840
rect -720 820 -710 840
rect -750 800 -710 820
rect -750 780 -740 800
rect -720 780 -710 800
rect -750 760 -710 780
rect -750 740 -740 760
rect -720 740 -710 760
rect -750 720 -710 740
rect -750 700 -740 720
rect -720 700 -710 720
rect -750 680 -710 700
rect -750 660 -740 680
rect -720 660 -710 680
rect -750 640 -710 660
rect -750 620 -740 640
rect -720 620 -710 640
rect -750 600 -710 620
rect -750 580 -740 600
rect -720 580 -710 600
rect -750 570 -710 580
rect -675 840 -635 850
rect -675 820 -665 840
rect -645 820 -635 840
rect -675 800 -635 820
rect -675 780 -665 800
rect -645 780 -635 800
rect -675 760 -635 780
rect -675 740 -665 760
rect -645 740 -635 760
rect -675 720 -635 740
rect -675 700 -665 720
rect -645 700 -635 720
rect -675 680 -635 700
rect -675 660 -665 680
rect -645 660 -635 680
rect -675 640 -635 660
rect -675 620 -665 640
rect -645 620 -635 640
rect -675 600 -635 620
rect -675 580 -665 600
rect -645 580 -635 600
rect -675 565 -635 580
rect -815 540 -795 565
rect -725 540 -685 550
rect -815 520 -715 540
rect -695 520 -685 540
rect -815 475 -795 520
rect -725 510 -685 520
rect -1280 455 -795 475
rect -1280 415 -1260 455
rect -980 415 -960 455
rect -815 435 -795 455
rect -775 480 -735 490
rect -665 480 -645 565
rect -775 460 -765 480
rect -745 460 -180 480
rect -775 450 -735 460
rect -665 435 -645 460
rect -1350 400 -1310 415
rect -1350 380 -1340 400
rect -1320 380 -1310 400
rect -1350 360 -1310 380
rect -1350 340 -1340 360
rect -1320 340 -1310 360
rect -1350 320 -1310 340
rect -1350 300 -1340 320
rect -1320 300 -1310 320
rect -1350 290 -1310 300
rect -1290 400 -1250 415
rect -1290 380 -1280 400
rect -1260 380 -1250 400
rect -1290 360 -1250 380
rect -1290 340 -1280 360
rect -1260 340 -1250 360
rect -1290 320 -1250 340
rect -1290 300 -1280 320
rect -1260 300 -1250 320
rect -1290 290 -1250 300
rect -1140 400 -1100 415
rect -1140 380 -1130 400
rect -1110 380 -1100 400
rect -1140 360 -1100 380
rect -1140 340 -1130 360
rect -1110 340 -1100 360
rect -1140 320 -1100 340
rect -1140 300 -1130 320
rect -1110 300 -1100 320
rect -1140 290 -1100 300
rect -990 400 -950 415
rect -990 380 -980 400
rect -960 380 -950 400
rect -990 360 -950 380
rect -990 340 -980 360
rect -960 340 -950 360
rect -990 320 -950 340
rect -990 300 -980 320
rect -960 300 -950 320
rect -990 290 -950 300
rect -900 400 -860 415
rect -900 380 -890 400
rect -870 380 -860 400
rect -900 360 -860 380
rect -900 340 -890 360
rect -870 340 -860 360
rect -900 320 -860 340
rect -900 300 -890 320
rect -870 300 -860 320
rect -900 290 -860 300
rect -825 400 -785 435
rect -825 380 -815 400
rect -795 380 -785 400
rect -825 360 -785 380
rect -825 340 -815 360
rect -795 340 -785 360
rect -825 320 -785 340
rect -825 300 -815 320
rect -795 300 -785 320
rect -825 290 -785 300
rect -750 400 -710 415
rect -750 380 -740 400
rect -720 380 -710 400
rect -750 360 -710 380
rect -750 340 -740 360
rect -720 340 -710 360
rect -750 320 -710 340
rect -750 300 -740 320
rect -720 300 -710 320
rect -750 290 -710 300
rect -675 400 -635 435
rect -500 415 -480 460
rect -200 415 -180 460
rect -675 380 -665 400
rect -645 380 -635 400
rect -675 360 -635 380
rect -675 340 -665 360
rect -645 340 -635 360
rect -675 320 -635 340
rect -675 300 -665 320
rect -645 300 -635 320
rect -675 290 -635 300
rect -600 400 -560 415
rect -600 380 -590 400
rect -570 380 -560 400
rect -600 360 -560 380
rect -600 340 -590 360
rect -570 340 -560 360
rect -600 320 -560 340
rect -600 300 -590 320
rect -570 300 -560 320
rect -600 290 -560 300
rect -510 400 -470 415
rect -510 380 -500 400
rect -480 380 -470 400
rect -510 360 -470 380
rect -510 340 -500 360
rect -480 340 -470 360
rect -510 320 -470 340
rect -510 300 -500 320
rect -480 300 -470 320
rect -510 290 -470 300
rect -360 400 -320 415
rect -360 380 -350 400
rect -330 380 -320 400
rect -360 360 -320 380
rect -360 340 -350 360
rect -330 340 -320 360
rect -360 320 -320 340
rect -360 300 -350 320
rect -330 300 -320 320
rect -360 290 -320 300
rect -210 400 -170 415
rect -210 380 -200 400
rect -180 380 -170 400
rect -210 360 -170 380
rect -210 340 -200 360
rect -180 340 -170 360
rect -210 320 -170 340
rect -210 300 -200 320
rect -180 300 -170 320
rect -210 290 -170 300
rect -150 400 -110 415
rect -150 380 -140 400
rect -120 380 -110 400
rect -150 360 -110 380
rect -150 340 -140 360
rect -120 340 -110 360
rect -150 320 -110 340
rect -150 300 -140 320
rect -120 300 -110 320
rect -150 290 -110 300
rect -850 260 -810 270
rect -650 260 -610 270
rect -1300 240 -840 260
rect -820 240 -640 260
rect -620 240 -610 260
rect -850 230 -810 240
rect -650 230 -610 240
rect -1090 210 -1050 220
rect -385 210 -345 220
rect -1300 190 -1080 210
rect -1060 190 -375 210
rect -355 190 -345 210
rect -1090 180 -1050 190
rect -385 180 -345 190
rect -1165 155 -1125 165
rect -310 155 -270 165
rect -1300 135 -1155 155
rect -1135 135 -300 155
rect -280 135 -270 155
rect -1165 125 -1125 135
rect -310 125 -270 135
rect -1015 105 -975 115
rect -235 105 -195 115
rect -1300 85 -1005 105
rect -985 85 -225 105
rect -205 85 -195 105
rect -1015 75 -975 85
rect -235 75 -195 85
rect -1240 50 -1200 60
rect -460 50 -420 60
rect -1300 30 -1230 50
rect -1210 30 -450 50
rect -430 30 -420 50
rect -1240 20 -1200 30
rect -460 20 -420 30
rect -1380 -10 -75 0
rect -1380 -30 -1360 -10
rect -1340 -30 -1320 -10
rect -1300 -30 -1280 -10
rect -1260 -30 -1240 -10
rect -1220 -30 -1200 -10
rect -1180 -30 -1160 -10
rect -1140 -30 -1120 -10
rect -1100 -30 -1080 -10
rect -1060 -30 -1040 -10
rect -1020 -30 -1000 -10
rect -980 -30 -960 -10
rect -940 -30 -920 -10
rect -900 -30 -880 -10
rect -860 -30 -840 -10
rect -820 -30 -800 -10
rect -780 -30 -760 -10
rect -740 -30 -720 -10
rect -700 -30 -680 -10
rect -660 -30 -635 -10
rect -615 -30 -595 -10
rect -575 -30 -555 -10
rect -535 -30 -515 -10
rect -495 -30 -475 -10
rect -455 -30 -435 -10
rect -415 -30 -395 -10
rect -375 -30 -355 -10
rect -335 -30 -315 -10
rect -295 -30 -275 -10
rect -255 -30 -235 -10
rect -215 -30 -195 -10
rect -175 -30 -155 -10
rect -135 -30 -115 -10
rect -95 -30 -75 -10
rect -1380 -40 -75 -30
<< viali >>
rect -1345 940 -1325 960
rect -1305 940 -1285 960
rect -1265 940 -1245 960
rect -1225 940 -1205 960
rect -1185 940 -1165 960
rect -1140 940 -1120 960
rect -1100 940 -1080 960
rect -1060 940 -1040 960
rect -1020 940 -1000 960
rect -980 940 -960 960
rect -940 940 -920 960
rect -900 940 -880 960
rect -860 940 -840 960
rect -820 940 -800 960
rect -780 940 -760 960
rect -740 940 -720 960
rect -700 940 -680 960
rect -660 940 -640 960
rect -620 940 -600 960
rect -580 940 -560 960
rect -540 940 -520 960
rect -500 940 -480 960
rect -455 940 -435 960
rect -415 940 -395 960
rect -375 940 -355 960
rect -335 940 -315 960
rect -295 940 -275 960
rect -255 940 -235 960
rect -215 940 -195 960
rect -175 940 -155 960
rect -135 940 -115 960
rect -740 820 -720 840
rect -740 780 -720 800
rect -740 740 -720 760
rect -740 700 -720 720
rect -740 660 -720 680
rect -740 620 -720 640
rect -740 580 -720 600
rect -1340 380 -1320 400
rect -1340 340 -1320 360
rect -1340 300 -1320 320
rect -1130 380 -1110 400
rect -1130 340 -1110 360
rect -1130 300 -1110 320
rect -890 380 -870 400
rect -890 340 -870 360
rect -890 300 -870 320
rect -740 380 -720 400
rect -740 340 -720 360
rect -740 300 -720 320
rect -590 380 -570 400
rect -590 340 -570 360
rect -590 300 -570 320
rect -350 380 -330 400
rect -350 340 -330 360
rect -350 300 -330 320
rect -140 380 -120 400
rect -140 340 -120 360
rect -140 300 -120 320
rect -1360 -30 -1340 -10
rect -1320 -30 -1300 -10
rect -1280 -30 -1260 -10
rect -1240 -30 -1220 -10
rect -1200 -30 -1180 -10
rect -1160 -30 -1140 -10
rect -1120 -30 -1100 -10
rect -1080 -30 -1060 -10
rect -1040 -30 -1020 -10
rect -1000 -30 -980 -10
rect -960 -30 -940 -10
rect -920 -30 -900 -10
rect -880 -30 -860 -10
rect -840 -30 -820 -10
rect -800 -30 -780 -10
rect -760 -30 -740 -10
rect -720 -30 -700 -10
rect -680 -30 -660 -10
rect -635 -30 -615 -10
rect -595 -30 -575 -10
rect -555 -30 -535 -10
rect -515 -30 -495 -10
rect -475 -30 -455 -10
rect -435 -30 -415 -10
rect -395 -30 -375 -10
rect -355 -30 -335 -10
rect -315 -30 -295 -10
rect -275 -30 -255 -10
rect -235 -30 -215 -10
rect -195 -30 -175 -10
rect -155 -30 -135 -10
rect -115 -30 -95 -10
<< metal1 >>
rect -1365 960 -95 975
rect -1365 940 -1345 960
rect -1325 940 -1305 960
rect -1285 940 -1265 960
rect -1245 940 -1225 960
rect -1205 940 -1185 960
rect -1165 940 -1140 960
rect -1120 940 -1100 960
rect -1080 940 -1060 960
rect -1040 940 -1020 960
rect -1000 940 -980 960
rect -960 940 -940 960
rect -920 940 -900 960
rect -880 940 -860 960
rect -840 940 -820 960
rect -800 940 -780 960
rect -760 940 -740 960
rect -720 940 -700 960
rect -680 940 -660 960
rect -640 940 -620 960
rect -600 940 -580 960
rect -560 940 -540 960
rect -520 940 -500 960
rect -480 940 -455 960
rect -435 940 -415 960
rect -395 940 -375 960
rect -355 940 -335 960
rect -315 940 -295 960
rect -275 940 -255 960
rect -235 940 -215 960
rect -195 940 -175 960
rect -155 940 -135 960
rect -115 940 -95 960
rect -1365 925 -95 940
rect -1130 415 -1110 925
rect -740 850 -720 925
rect -750 840 -710 850
rect -750 820 -740 840
rect -720 820 -710 840
rect -750 800 -710 820
rect -750 780 -740 800
rect -720 780 -710 800
rect -750 760 -710 780
rect -750 740 -740 760
rect -720 740 -710 760
rect -750 720 -710 740
rect -750 700 -740 720
rect -720 700 -710 720
rect -750 680 -710 700
rect -750 660 -740 680
rect -720 660 -710 680
rect -750 640 -710 660
rect -750 620 -740 640
rect -720 620 -710 640
rect -750 600 -710 620
rect -750 580 -740 600
rect -720 580 -710 600
rect -750 570 -710 580
rect -350 415 -330 925
rect -1350 400 -1310 415
rect -1350 380 -1340 400
rect -1320 380 -1310 400
rect -1350 360 -1310 380
rect -1350 340 -1340 360
rect -1320 340 -1310 360
rect -1350 320 -1310 340
rect -1350 300 -1340 320
rect -1320 300 -1310 320
rect -1350 5 -1310 300
rect -1140 400 -1100 415
rect -1140 380 -1130 400
rect -1110 380 -1100 400
rect -1140 360 -1100 380
rect -1140 340 -1130 360
rect -1110 340 -1100 360
rect -1140 320 -1100 340
rect -1140 300 -1130 320
rect -1110 300 -1100 320
rect -1140 290 -1100 300
rect -900 400 -860 415
rect -900 380 -890 400
rect -870 380 -860 400
rect -900 360 -860 380
rect -900 340 -890 360
rect -870 340 -860 360
rect -900 320 -860 340
rect -900 300 -890 320
rect -870 300 -860 320
rect -900 290 -860 300
rect -750 400 -710 415
rect -750 380 -740 400
rect -720 380 -710 400
rect -750 360 -710 380
rect -750 340 -740 360
rect -720 340 -710 360
rect -750 320 -710 340
rect -750 300 -740 320
rect -720 300 -710 320
rect -750 290 -710 300
rect -600 400 -560 415
rect -600 380 -590 400
rect -570 380 -560 400
rect -600 360 -560 380
rect -600 340 -590 360
rect -570 340 -560 360
rect -600 320 -560 340
rect -600 300 -590 320
rect -570 300 -560 320
rect -600 290 -560 300
rect -360 400 -320 415
rect -360 380 -350 400
rect -330 380 -320 400
rect -360 360 -320 380
rect -360 340 -350 360
rect -330 340 -320 360
rect -360 320 -320 340
rect -360 300 -350 320
rect -330 300 -320 320
rect -360 290 -320 300
rect -150 400 -110 415
rect -150 380 -140 400
rect -120 380 -110 400
rect -150 360 -110 380
rect -150 340 -140 360
rect -120 340 -110 360
rect -150 320 -110 340
rect -150 300 -140 320
rect -120 300 -110 320
rect -890 5 -870 290
rect -740 5 -720 290
rect -590 5 -570 290
rect -150 5 -110 300
rect -1380 -10 -75 5
rect -1380 -30 -1360 -10
rect -1340 -30 -1320 -10
rect -1300 -30 -1280 -10
rect -1260 -30 -1240 -10
rect -1220 -30 -1200 -10
rect -1180 -30 -1160 -10
rect -1140 -30 -1120 -10
rect -1100 -30 -1080 -10
rect -1060 -30 -1040 -10
rect -1020 -30 -1000 -10
rect -980 -30 -960 -10
rect -940 -30 -920 -10
rect -900 -30 -880 -10
rect -860 -30 -840 -10
rect -820 -30 -800 -10
rect -780 -30 -760 -10
rect -740 -30 -720 -10
rect -700 -30 -680 -10
rect -660 -30 -635 -10
rect -615 -30 -595 -10
rect -575 -30 -555 -10
rect -535 -30 -515 -10
rect -495 -30 -475 -10
rect -455 -30 -435 -10
rect -415 -30 -395 -10
rect -375 -30 -355 -10
rect -335 -30 -315 -10
rect -295 -30 -275 -10
rect -255 -30 -235 -10
rect -215 -30 -195 -10
rect -175 -30 -155 -10
rect -135 -30 -115 -10
rect -95 -30 -75 -10
rect -1380 -45 -75 -30
<< labels >>
rlabel locali -1295 140 -1285 150 1 A_bar
port 2 n
rlabel locali -1295 90 -1285 100 1 B
port 3 n
rlabel locali -1295 35 -1285 45 1 B_bar
port 4 n
rlabel metal1 -740 940 -720 960 7 CLK
port 9 w
rlabel metal1 -880 -30 -860 -10 7 GND!
port 8 w
rlabel locali -1295 245 -1285 255 7 Dis
port 7 w
rlabel locali -1295 195 -1285 205 7 A
port 1 w
rlabel locali -575 465 -565 475 3 OUT
port 5 e
rlabel locali -900 460 -890 470 7 OUT_bar
port 6 w
<< end >>
