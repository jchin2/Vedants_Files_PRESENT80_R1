magic
tech sky130A
magscale 1 2
timestamp 1671076365
<< pwell >>
rect -9674 -44917 -6288 -43965
rect -5568 -44917 -2156 -43965
rect -6643 -48202 -5151 -47150
<< nmoslvt >>
rect -9408 -44891 -9378 -43991
rect -9258 -44891 -9228 -43991
rect -9108 -44891 -9078 -43991
rect -8958 -44891 -8928 -43991
rect -8808 -44891 -8778 -43991
rect -8658 -44891 -8628 -43991
rect -8508 -44891 -8478 -43991
rect -8358 -44891 -8328 -43991
rect -8208 -44891 -8178 -43991
rect -8058 -44891 -8028 -43991
rect -7908 -44891 -7878 -43991
rect -7758 -44891 -7728 -43991
rect -7608 -44891 -7578 -43991
rect -7458 -44891 -7428 -43991
rect -7308 -44891 -7278 -43991
rect -7158 -44891 -7128 -43991
rect -7008 -44891 -6978 -43991
rect -6858 -44891 -6828 -43991
rect -6708 -44891 -6678 -43991
rect -6558 -44891 -6528 -43991
rect -5302 -44891 -5272 -43991
rect -5152 -44891 -5122 -43991
rect -5002 -44891 -4972 -43991
rect -4852 -44891 -4822 -43991
rect -4702 -44891 -4672 -43991
rect -4552 -44891 -4522 -43991
rect -4402 -44891 -4372 -43991
rect -4252 -44891 -4222 -43991
rect -4102 -44891 -4072 -43991
rect -3952 -44891 -3922 -43991
rect -3802 -44891 -3772 -43991
rect -3652 -44891 -3622 -43991
rect -3502 -44891 -3472 -43991
rect -3352 -44891 -3322 -43991
rect -3202 -44891 -3172 -43991
rect -3052 -44891 -3022 -43991
rect -2902 -44891 -2872 -43991
rect -2752 -44891 -2722 -43991
rect -2602 -44891 -2572 -43991
rect -2452 -44891 -2422 -43991
rect -6377 -48176 -6347 -47176
rect -6227 -48176 -6197 -47176
rect -6077 -48176 -6047 -47176
rect -5927 -48176 -5897 -47176
rect -5777 -48176 -5747 -47176
rect -5627 -48176 -5597 -47176
rect -5477 -48176 -5447 -47176
rect -5327 -48176 -5297 -47176
<< ndiff >>
rect -9528 -44050 -9408 -43991
rect -9528 -44084 -9485 -44050
rect -9451 -44084 -9408 -44050
rect -9528 -44118 -9408 -44084
rect -9528 -44152 -9485 -44118
rect -9451 -44152 -9408 -44118
rect -9528 -44186 -9408 -44152
rect -9528 -44220 -9485 -44186
rect -9451 -44220 -9408 -44186
rect -9528 -44254 -9408 -44220
rect -9528 -44288 -9485 -44254
rect -9451 -44288 -9408 -44254
rect -9528 -44322 -9408 -44288
rect -9528 -44356 -9485 -44322
rect -9451 -44356 -9408 -44322
rect -9528 -44390 -9408 -44356
rect -9528 -44424 -9485 -44390
rect -9451 -44424 -9408 -44390
rect -9528 -44458 -9408 -44424
rect -9528 -44492 -9485 -44458
rect -9451 -44492 -9408 -44458
rect -9528 -44526 -9408 -44492
rect -9528 -44560 -9485 -44526
rect -9451 -44560 -9408 -44526
rect -9528 -44594 -9408 -44560
rect -9528 -44628 -9485 -44594
rect -9451 -44628 -9408 -44594
rect -9528 -44662 -9408 -44628
rect -9528 -44696 -9485 -44662
rect -9451 -44696 -9408 -44662
rect -9528 -44730 -9408 -44696
rect -9528 -44764 -9485 -44730
rect -9451 -44764 -9408 -44730
rect -9528 -44798 -9408 -44764
rect -9528 -44832 -9485 -44798
rect -9451 -44832 -9408 -44798
rect -9528 -44891 -9408 -44832
rect -9378 -44050 -9258 -43991
rect -9378 -44084 -9335 -44050
rect -9301 -44084 -9258 -44050
rect -9378 -44118 -9258 -44084
rect -9378 -44152 -9335 -44118
rect -9301 -44152 -9258 -44118
rect -9378 -44186 -9258 -44152
rect -9378 -44220 -9335 -44186
rect -9301 -44220 -9258 -44186
rect -9378 -44254 -9258 -44220
rect -9378 -44288 -9335 -44254
rect -9301 -44288 -9258 -44254
rect -9378 -44322 -9258 -44288
rect -9378 -44356 -9335 -44322
rect -9301 -44356 -9258 -44322
rect -9378 -44390 -9258 -44356
rect -9378 -44424 -9335 -44390
rect -9301 -44424 -9258 -44390
rect -9378 -44458 -9258 -44424
rect -9378 -44492 -9335 -44458
rect -9301 -44492 -9258 -44458
rect -9378 -44526 -9258 -44492
rect -9378 -44560 -9335 -44526
rect -9301 -44560 -9258 -44526
rect -9378 -44594 -9258 -44560
rect -9378 -44628 -9335 -44594
rect -9301 -44628 -9258 -44594
rect -9378 -44662 -9258 -44628
rect -9378 -44696 -9335 -44662
rect -9301 -44696 -9258 -44662
rect -9378 -44730 -9258 -44696
rect -9378 -44764 -9335 -44730
rect -9301 -44764 -9258 -44730
rect -9378 -44798 -9258 -44764
rect -9378 -44832 -9335 -44798
rect -9301 -44832 -9258 -44798
rect -9378 -44891 -9258 -44832
rect -9228 -44050 -9108 -43991
rect -9228 -44084 -9185 -44050
rect -9151 -44084 -9108 -44050
rect -9228 -44118 -9108 -44084
rect -9228 -44152 -9185 -44118
rect -9151 -44152 -9108 -44118
rect -9228 -44186 -9108 -44152
rect -9228 -44220 -9185 -44186
rect -9151 -44220 -9108 -44186
rect -9228 -44254 -9108 -44220
rect -9228 -44288 -9185 -44254
rect -9151 -44288 -9108 -44254
rect -9228 -44322 -9108 -44288
rect -9228 -44356 -9185 -44322
rect -9151 -44356 -9108 -44322
rect -9228 -44390 -9108 -44356
rect -9228 -44424 -9185 -44390
rect -9151 -44424 -9108 -44390
rect -9228 -44458 -9108 -44424
rect -9228 -44492 -9185 -44458
rect -9151 -44492 -9108 -44458
rect -9228 -44526 -9108 -44492
rect -9228 -44560 -9185 -44526
rect -9151 -44560 -9108 -44526
rect -9228 -44594 -9108 -44560
rect -9228 -44628 -9185 -44594
rect -9151 -44628 -9108 -44594
rect -9228 -44662 -9108 -44628
rect -9228 -44696 -9185 -44662
rect -9151 -44696 -9108 -44662
rect -9228 -44730 -9108 -44696
rect -9228 -44764 -9185 -44730
rect -9151 -44764 -9108 -44730
rect -9228 -44798 -9108 -44764
rect -9228 -44832 -9185 -44798
rect -9151 -44832 -9108 -44798
rect -9228 -44891 -9108 -44832
rect -9078 -44050 -8958 -43991
rect -9078 -44084 -9035 -44050
rect -9001 -44084 -8958 -44050
rect -9078 -44118 -8958 -44084
rect -9078 -44152 -9035 -44118
rect -9001 -44152 -8958 -44118
rect -9078 -44186 -8958 -44152
rect -9078 -44220 -9035 -44186
rect -9001 -44220 -8958 -44186
rect -9078 -44254 -8958 -44220
rect -9078 -44288 -9035 -44254
rect -9001 -44288 -8958 -44254
rect -9078 -44322 -8958 -44288
rect -9078 -44356 -9035 -44322
rect -9001 -44356 -8958 -44322
rect -9078 -44390 -8958 -44356
rect -9078 -44424 -9035 -44390
rect -9001 -44424 -8958 -44390
rect -9078 -44458 -8958 -44424
rect -9078 -44492 -9035 -44458
rect -9001 -44492 -8958 -44458
rect -9078 -44526 -8958 -44492
rect -9078 -44560 -9035 -44526
rect -9001 -44560 -8958 -44526
rect -9078 -44594 -8958 -44560
rect -9078 -44628 -9035 -44594
rect -9001 -44628 -8958 -44594
rect -9078 -44662 -8958 -44628
rect -9078 -44696 -9035 -44662
rect -9001 -44696 -8958 -44662
rect -9078 -44730 -8958 -44696
rect -9078 -44764 -9035 -44730
rect -9001 -44764 -8958 -44730
rect -9078 -44798 -8958 -44764
rect -9078 -44832 -9035 -44798
rect -9001 -44832 -8958 -44798
rect -9078 -44891 -8958 -44832
rect -8928 -44050 -8808 -43991
rect -8928 -44084 -8885 -44050
rect -8851 -44084 -8808 -44050
rect -8928 -44118 -8808 -44084
rect -8928 -44152 -8885 -44118
rect -8851 -44152 -8808 -44118
rect -8928 -44186 -8808 -44152
rect -8928 -44220 -8885 -44186
rect -8851 -44220 -8808 -44186
rect -8928 -44254 -8808 -44220
rect -8928 -44288 -8885 -44254
rect -8851 -44288 -8808 -44254
rect -8928 -44322 -8808 -44288
rect -8928 -44356 -8885 -44322
rect -8851 -44356 -8808 -44322
rect -8928 -44390 -8808 -44356
rect -8928 -44424 -8885 -44390
rect -8851 -44424 -8808 -44390
rect -8928 -44458 -8808 -44424
rect -8928 -44492 -8885 -44458
rect -8851 -44492 -8808 -44458
rect -8928 -44526 -8808 -44492
rect -8928 -44560 -8885 -44526
rect -8851 -44560 -8808 -44526
rect -8928 -44594 -8808 -44560
rect -8928 -44628 -8885 -44594
rect -8851 -44628 -8808 -44594
rect -8928 -44662 -8808 -44628
rect -8928 -44696 -8885 -44662
rect -8851 -44696 -8808 -44662
rect -8928 -44730 -8808 -44696
rect -8928 -44764 -8885 -44730
rect -8851 -44764 -8808 -44730
rect -8928 -44798 -8808 -44764
rect -8928 -44832 -8885 -44798
rect -8851 -44832 -8808 -44798
rect -8928 -44891 -8808 -44832
rect -8778 -44050 -8658 -43991
rect -8778 -44084 -8735 -44050
rect -8701 -44084 -8658 -44050
rect -8778 -44118 -8658 -44084
rect -8778 -44152 -8735 -44118
rect -8701 -44152 -8658 -44118
rect -8778 -44186 -8658 -44152
rect -8778 -44220 -8735 -44186
rect -8701 -44220 -8658 -44186
rect -8778 -44254 -8658 -44220
rect -8778 -44288 -8735 -44254
rect -8701 -44288 -8658 -44254
rect -8778 -44322 -8658 -44288
rect -8778 -44356 -8735 -44322
rect -8701 -44356 -8658 -44322
rect -8778 -44390 -8658 -44356
rect -8778 -44424 -8735 -44390
rect -8701 -44424 -8658 -44390
rect -8778 -44458 -8658 -44424
rect -8778 -44492 -8735 -44458
rect -8701 -44492 -8658 -44458
rect -8778 -44526 -8658 -44492
rect -8778 -44560 -8735 -44526
rect -8701 -44560 -8658 -44526
rect -8778 -44594 -8658 -44560
rect -8778 -44628 -8735 -44594
rect -8701 -44628 -8658 -44594
rect -8778 -44662 -8658 -44628
rect -8778 -44696 -8735 -44662
rect -8701 -44696 -8658 -44662
rect -8778 -44730 -8658 -44696
rect -8778 -44764 -8735 -44730
rect -8701 -44764 -8658 -44730
rect -8778 -44798 -8658 -44764
rect -8778 -44832 -8735 -44798
rect -8701 -44832 -8658 -44798
rect -8778 -44891 -8658 -44832
rect -8628 -44050 -8508 -43991
rect -8628 -44084 -8585 -44050
rect -8551 -44084 -8508 -44050
rect -8628 -44118 -8508 -44084
rect -8628 -44152 -8585 -44118
rect -8551 -44152 -8508 -44118
rect -8628 -44186 -8508 -44152
rect -8628 -44220 -8585 -44186
rect -8551 -44220 -8508 -44186
rect -8628 -44254 -8508 -44220
rect -8628 -44288 -8585 -44254
rect -8551 -44288 -8508 -44254
rect -8628 -44322 -8508 -44288
rect -8628 -44356 -8585 -44322
rect -8551 -44356 -8508 -44322
rect -8628 -44390 -8508 -44356
rect -8628 -44424 -8585 -44390
rect -8551 -44424 -8508 -44390
rect -8628 -44458 -8508 -44424
rect -8628 -44492 -8585 -44458
rect -8551 -44492 -8508 -44458
rect -8628 -44526 -8508 -44492
rect -8628 -44560 -8585 -44526
rect -8551 -44560 -8508 -44526
rect -8628 -44594 -8508 -44560
rect -8628 -44628 -8585 -44594
rect -8551 -44628 -8508 -44594
rect -8628 -44662 -8508 -44628
rect -8628 -44696 -8585 -44662
rect -8551 -44696 -8508 -44662
rect -8628 -44730 -8508 -44696
rect -8628 -44764 -8585 -44730
rect -8551 -44764 -8508 -44730
rect -8628 -44798 -8508 -44764
rect -8628 -44832 -8585 -44798
rect -8551 -44832 -8508 -44798
rect -8628 -44891 -8508 -44832
rect -8478 -44050 -8358 -43991
rect -8478 -44084 -8435 -44050
rect -8401 -44084 -8358 -44050
rect -8478 -44118 -8358 -44084
rect -8478 -44152 -8435 -44118
rect -8401 -44152 -8358 -44118
rect -8478 -44186 -8358 -44152
rect -8478 -44220 -8435 -44186
rect -8401 -44220 -8358 -44186
rect -8478 -44254 -8358 -44220
rect -8478 -44288 -8435 -44254
rect -8401 -44288 -8358 -44254
rect -8478 -44322 -8358 -44288
rect -8478 -44356 -8435 -44322
rect -8401 -44356 -8358 -44322
rect -8478 -44390 -8358 -44356
rect -8478 -44424 -8435 -44390
rect -8401 -44424 -8358 -44390
rect -8478 -44458 -8358 -44424
rect -8478 -44492 -8435 -44458
rect -8401 -44492 -8358 -44458
rect -8478 -44526 -8358 -44492
rect -8478 -44560 -8435 -44526
rect -8401 -44560 -8358 -44526
rect -8478 -44594 -8358 -44560
rect -8478 -44628 -8435 -44594
rect -8401 -44628 -8358 -44594
rect -8478 -44662 -8358 -44628
rect -8478 -44696 -8435 -44662
rect -8401 -44696 -8358 -44662
rect -8478 -44730 -8358 -44696
rect -8478 -44764 -8435 -44730
rect -8401 -44764 -8358 -44730
rect -8478 -44798 -8358 -44764
rect -8478 -44832 -8435 -44798
rect -8401 -44832 -8358 -44798
rect -8478 -44891 -8358 -44832
rect -8328 -44050 -8208 -43991
rect -8328 -44084 -8285 -44050
rect -8251 -44084 -8208 -44050
rect -8328 -44118 -8208 -44084
rect -8328 -44152 -8285 -44118
rect -8251 -44152 -8208 -44118
rect -8328 -44186 -8208 -44152
rect -8328 -44220 -8285 -44186
rect -8251 -44220 -8208 -44186
rect -8328 -44254 -8208 -44220
rect -8328 -44288 -8285 -44254
rect -8251 -44288 -8208 -44254
rect -8328 -44322 -8208 -44288
rect -8328 -44356 -8285 -44322
rect -8251 -44356 -8208 -44322
rect -8328 -44390 -8208 -44356
rect -8328 -44424 -8285 -44390
rect -8251 -44424 -8208 -44390
rect -8328 -44458 -8208 -44424
rect -8328 -44492 -8285 -44458
rect -8251 -44492 -8208 -44458
rect -8328 -44526 -8208 -44492
rect -8328 -44560 -8285 -44526
rect -8251 -44560 -8208 -44526
rect -8328 -44594 -8208 -44560
rect -8328 -44628 -8285 -44594
rect -8251 -44628 -8208 -44594
rect -8328 -44662 -8208 -44628
rect -8328 -44696 -8285 -44662
rect -8251 -44696 -8208 -44662
rect -8328 -44730 -8208 -44696
rect -8328 -44764 -8285 -44730
rect -8251 -44764 -8208 -44730
rect -8328 -44798 -8208 -44764
rect -8328 -44832 -8285 -44798
rect -8251 -44832 -8208 -44798
rect -8328 -44891 -8208 -44832
rect -8178 -44060 -8058 -43991
rect -8178 -44094 -8135 -44060
rect -8101 -44094 -8058 -44060
rect -8178 -44128 -8058 -44094
rect -8178 -44162 -8135 -44128
rect -8101 -44162 -8058 -44128
rect -8178 -44196 -8058 -44162
rect -8178 -44230 -8135 -44196
rect -8101 -44230 -8058 -44196
rect -8178 -44264 -8058 -44230
rect -8178 -44298 -8135 -44264
rect -8101 -44298 -8058 -44264
rect -8178 -44332 -8058 -44298
rect -8178 -44366 -8135 -44332
rect -8101 -44366 -8058 -44332
rect -8178 -44400 -8058 -44366
rect -8178 -44434 -8135 -44400
rect -8101 -44434 -8058 -44400
rect -8178 -44468 -8058 -44434
rect -8178 -44502 -8135 -44468
rect -8101 -44502 -8058 -44468
rect -8178 -44536 -8058 -44502
rect -8178 -44570 -8135 -44536
rect -8101 -44570 -8058 -44536
rect -8178 -44604 -8058 -44570
rect -8178 -44638 -8135 -44604
rect -8101 -44638 -8058 -44604
rect -8178 -44672 -8058 -44638
rect -8178 -44706 -8135 -44672
rect -8101 -44706 -8058 -44672
rect -8178 -44740 -8058 -44706
rect -8178 -44774 -8135 -44740
rect -8101 -44774 -8058 -44740
rect -8178 -44808 -8058 -44774
rect -8178 -44842 -8135 -44808
rect -8101 -44842 -8058 -44808
rect -8178 -44891 -8058 -44842
rect -8028 -44050 -7908 -43991
rect -8028 -44084 -7985 -44050
rect -7951 -44084 -7908 -44050
rect -8028 -44118 -7908 -44084
rect -8028 -44152 -7985 -44118
rect -7951 -44152 -7908 -44118
rect -8028 -44186 -7908 -44152
rect -8028 -44220 -7985 -44186
rect -7951 -44220 -7908 -44186
rect -8028 -44254 -7908 -44220
rect -8028 -44288 -7985 -44254
rect -7951 -44288 -7908 -44254
rect -8028 -44322 -7908 -44288
rect -8028 -44356 -7985 -44322
rect -7951 -44356 -7908 -44322
rect -8028 -44390 -7908 -44356
rect -8028 -44424 -7985 -44390
rect -7951 -44424 -7908 -44390
rect -8028 -44458 -7908 -44424
rect -8028 -44492 -7985 -44458
rect -7951 -44492 -7908 -44458
rect -8028 -44526 -7908 -44492
rect -8028 -44560 -7985 -44526
rect -7951 -44560 -7908 -44526
rect -8028 -44594 -7908 -44560
rect -8028 -44628 -7985 -44594
rect -7951 -44628 -7908 -44594
rect -8028 -44662 -7908 -44628
rect -8028 -44696 -7985 -44662
rect -7951 -44696 -7908 -44662
rect -8028 -44730 -7908 -44696
rect -8028 -44764 -7985 -44730
rect -7951 -44764 -7908 -44730
rect -8028 -44798 -7908 -44764
rect -8028 -44832 -7985 -44798
rect -7951 -44832 -7908 -44798
rect -8028 -44891 -7908 -44832
rect -7878 -44050 -7758 -43991
rect -7878 -44084 -7835 -44050
rect -7801 -44084 -7758 -44050
rect -7878 -44118 -7758 -44084
rect -7878 -44152 -7835 -44118
rect -7801 -44152 -7758 -44118
rect -7878 -44186 -7758 -44152
rect -7878 -44220 -7835 -44186
rect -7801 -44220 -7758 -44186
rect -7878 -44254 -7758 -44220
rect -7878 -44288 -7835 -44254
rect -7801 -44288 -7758 -44254
rect -7878 -44322 -7758 -44288
rect -7878 -44356 -7835 -44322
rect -7801 -44356 -7758 -44322
rect -7878 -44390 -7758 -44356
rect -7878 -44424 -7835 -44390
rect -7801 -44424 -7758 -44390
rect -7878 -44458 -7758 -44424
rect -7878 -44492 -7835 -44458
rect -7801 -44492 -7758 -44458
rect -7878 -44526 -7758 -44492
rect -7878 -44560 -7835 -44526
rect -7801 -44560 -7758 -44526
rect -7878 -44594 -7758 -44560
rect -7878 -44628 -7835 -44594
rect -7801 -44628 -7758 -44594
rect -7878 -44662 -7758 -44628
rect -7878 -44696 -7835 -44662
rect -7801 -44696 -7758 -44662
rect -7878 -44730 -7758 -44696
rect -7878 -44764 -7835 -44730
rect -7801 -44764 -7758 -44730
rect -7878 -44798 -7758 -44764
rect -7878 -44832 -7835 -44798
rect -7801 -44832 -7758 -44798
rect -7878 -44891 -7758 -44832
rect -7728 -44050 -7608 -43991
rect -7728 -44084 -7685 -44050
rect -7651 -44084 -7608 -44050
rect -7728 -44118 -7608 -44084
rect -7728 -44152 -7685 -44118
rect -7651 -44152 -7608 -44118
rect -7728 -44186 -7608 -44152
rect -7728 -44220 -7685 -44186
rect -7651 -44220 -7608 -44186
rect -7728 -44254 -7608 -44220
rect -7728 -44288 -7685 -44254
rect -7651 -44288 -7608 -44254
rect -7728 -44322 -7608 -44288
rect -7728 -44356 -7685 -44322
rect -7651 -44356 -7608 -44322
rect -7728 -44390 -7608 -44356
rect -7728 -44424 -7685 -44390
rect -7651 -44424 -7608 -44390
rect -7728 -44458 -7608 -44424
rect -7728 -44492 -7685 -44458
rect -7651 -44492 -7608 -44458
rect -7728 -44526 -7608 -44492
rect -7728 -44560 -7685 -44526
rect -7651 -44560 -7608 -44526
rect -7728 -44594 -7608 -44560
rect -7728 -44628 -7685 -44594
rect -7651 -44628 -7608 -44594
rect -7728 -44662 -7608 -44628
rect -7728 -44696 -7685 -44662
rect -7651 -44696 -7608 -44662
rect -7728 -44730 -7608 -44696
rect -7728 -44764 -7685 -44730
rect -7651 -44764 -7608 -44730
rect -7728 -44798 -7608 -44764
rect -7728 -44832 -7685 -44798
rect -7651 -44832 -7608 -44798
rect -7728 -44891 -7608 -44832
rect -7578 -44050 -7458 -43991
rect -7578 -44084 -7535 -44050
rect -7501 -44084 -7458 -44050
rect -7578 -44118 -7458 -44084
rect -7578 -44152 -7535 -44118
rect -7501 -44152 -7458 -44118
rect -7578 -44186 -7458 -44152
rect -7578 -44220 -7535 -44186
rect -7501 -44220 -7458 -44186
rect -7578 -44254 -7458 -44220
rect -7578 -44288 -7535 -44254
rect -7501 -44288 -7458 -44254
rect -7578 -44322 -7458 -44288
rect -7578 -44356 -7535 -44322
rect -7501 -44356 -7458 -44322
rect -7578 -44390 -7458 -44356
rect -7578 -44424 -7535 -44390
rect -7501 -44424 -7458 -44390
rect -7578 -44458 -7458 -44424
rect -7578 -44492 -7535 -44458
rect -7501 -44492 -7458 -44458
rect -7578 -44526 -7458 -44492
rect -7578 -44560 -7535 -44526
rect -7501 -44560 -7458 -44526
rect -7578 -44594 -7458 -44560
rect -7578 -44628 -7535 -44594
rect -7501 -44628 -7458 -44594
rect -7578 -44662 -7458 -44628
rect -7578 -44696 -7535 -44662
rect -7501 -44696 -7458 -44662
rect -7578 -44730 -7458 -44696
rect -7578 -44764 -7535 -44730
rect -7501 -44764 -7458 -44730
rect -7578 -44798 -7458 -44764
rect -7578 -44832 -7535 -44798
rect -7501 -44832 -7458 -44798
rect -7578 -44891 -7458 -44832
rect -7428 -44050 -7308 -43991
rect -7428 -44084 -7385 -44050
rect -7351 -44084 -7308 -44050
rect -7428 -44118 -7308 -44084
rect -7428 -44152 -7385 -44118
rect -7351 -44152 -7308 -44118
rect -7428 -44186 -7308 -44152
rect -7428 -44220 -7385 -44186
rect -7351 -44220 -7308 -44186
rect -7428 -44254 -7308 -44220
rect -7428 -44288 -7385 -44254
rect -7351 -44288 -7308 -44254
rect -7428 -44322 -7308 -44288
rect -7428 -44356 -7385 -44322
rect -7351 -44356 -7308 -44322
rect -7428 -44390 -7308 -44356
rect -7428 -44424 -7385 -44390
rect -7351 -44424 -7308 -44390
rect -7428 -44458 -7308 -44424
rect -7428 -44492 -7385 -44458
rect -7351 -44492 -7308 -44458
rect -7428 -44526 -7308 -44492
rect -7428 -44560 -7385 -44526
rect -7351 -44560 -7308 -44526
rect -7428 -44594 -7308 -44560
rect -7428 -44628 -7385 -44594
rect -7351 -44628 -7308 -44594
rect -7428 -44662 -7308 -44628
rect -7428 -44696 -7385 -44662
rect -7351 -44696 -7308 -44662
rect -7428 -44730 -7308 -44696
rect -7428 -44764 -7385 -44730
rect -7351 -44764 -7308 -44730
rect -7428 -44798 -7308 -44764
rect -7428 -44832 -7385 -44798
rect -7351 -44832 -7308 -44798
rect -7428 -44891 -7308 -44832
rect -7278 -44050 -7158 -43991
rect -7278 -44084 -7235 -44050
rect -7201 -44084 -7158 -44050
rect -7278 -44118 -7158 -44084
rect -7278 -44152 -7235 -44118
rect -7201 -44152 -7158 -44118
rect -7278 -44186 -7158 -44152
rect -7278 -44220 -7235 -44186
rect -7201 -44220 -7158 -44186
rect -7278 -44254 -7158 -44220
rect -7278 -44288 -7235 -44254
rect -7201 -44288 -7158 -44254
rect -7278 -44322 -7158 -44288
rect -7278 -44356 -7235 -44322
rect -7201 -44356 -7158 -44322
rect -7278 -44390 -7158 -44356
rect -7278 -44424 -7235 -44390
rect -7201 -44424 -7158 -44390
rect -7278 -44458 -7158 -44424
rect -7278 -44492 -7235 -44458
rect -7201 -44492 -7158 -44458
rect -7278 -44526 -7158 -44492
rect -7278 -44560 -7235 -44526
rect -7201 -44560 -7158 -44526
rect -7278 -44594 -7158 -44560
rect -7278 -44628 -7235 -44594
rect -7201 -44628 -7158 -44594
rect -7278 -44662 -7158 -44628
rect -7278 -44696 -7235 -44662
rect -7201 -44696 -7158 -44662
rect -7278 -44730 -7158 -44696
rect -7278 -44764 -7235 -44730
rect -7201 -44764 -7158 -44730
rect -7278 -44798 -7158 -44764
rect -7278 -44832 -7235 -44798
rect -7201 -44832 -7158 -44798
rect -7278 -44891 -7158 -44832
rect -7128 -44050 -7008 -43991
rect -7128 -44084 -7085 -44050
rect -7051 -44084 -7008 -44050
rect -7128 -44118 -7008 -44084
rect -7128 -44152 -7085 -44118
rect -7051 -44152 -7008 -44118
rect -7128 -44186 -7008 -44152
rect -7128 -44220 -7085 -44186
rect -7051 -44220 -7008 -44186
rect -7128 -44254 -7008 -44220
rect -7128 -44288 -7085 -44254
rect -7051 -44288 -7008 -44254
rect -7128 -44322 -7008 -44288
rect -7128 -44356 -7085 -44322
rect -7051 -44356 -7008 -44322
rect -7128 -44390 -7008 -44356
rect -7128 -44424 -7085 -44390
rect -7051 -44424 -7008 -44390
rect -7128 -44458 -7008 -44424
rect -7128 -44492 -7085 -44458
rect -7051 -44492 -7008 -44458
rect -7128 -44526 -7008 -44492
rect -7128 -44560 -7085 -44526
rect -7051 -44560 -7008 -44526
rect -7128 -44594 -7008 -44560
rect -7128 -44628 -7085 -44594
rect -7051 -44628 -7008 -44594
rect -7128 -44662 -7008 -44628
rect -7128 -44696 -7085 -44662
rect -7051 -44696 -7008 -44662
rect -7128 -44730 -7008 -44696
rect -7128 -44764 -7085 -44730
rect -7051 -44764 -7008 -44730
rect -7128 -44798 -7008 -44764
rect -7128 -44832 -7085 -44798
rect -7051 -44832 -7008 -44798
rect -7128 -44891 -7008 -44832
rect -6978 -44050 -6858 -43991
rect -6978 -44084 -6935 -44050
rect -6901 -44084 -6858 -44050
rect -6978 -44118 -6858 -44084
rect -6978 -44152 -6935 -44118
rect -6901 -44152 -6858 -44118
rect -6978 -44186 -6858 -44152
rect -6978 -44220 -6935 -44186
rect -6901 -44220 -6858 -44186
rect -6978 -44254 -6858 -44220
rect -6978 -44288 -6935 -44254
rect -6901 -44288 -6858 -44254
rect -6978 -44322 -6858 -44288
rect -6978 -44356 -6935 -44322
rect -6901 -44356 -6858 -44322
rect -6978 -44390 -6858 -44356
rect -6978 -44424 -6935 -44390
rect -6901 -44424 -6858 -44390
rect -6978 -44458 -6858 -44424
rect -6978 -44492 -6935 -44458
rect -6901 -44492 -6858 -44458
rect -6978 -44526 -6858 -44492
rect -6978 -44560 -6935 -44526
rect -6901 -44560 -6858 -44526
rect -6978 -44594 -6858 -44560
rect -6978 -44628 -6935 -44594
rect -6901 -44628 -6858 -44594
rect -6978 -44662 -6858 -44628
rect -6978 -44696 -6935 -44662
rect -6901 -44696 -6858 -44662
rect -6978 -44730 -6858 -44696
rect -6978 -44764 -6935 -44730
rect -6901 -44764 -6858 -44730
rect -6978 -44798 -6858 -44764
rect -6978 -44832 -6935 -44798
rect -6901 -44832 -6858 -44798
rect -6978 -44891 -6858 -44832
rect -6828 -44050 -6708 -43991
rect -6828 -44084 -6785 -44050
rect -6751 -44084 -6708 -44050
rect -6828 -44118 -6708 -44084
rect -6828 -44152 -6785 -44118
rect -6751 -44152 -6708 -44118
rect -6828 -44186 -6708 -44152
rect -6828 -44220 -6785 -44186
rect -6751 -44220 -6708 -44186
rect -6828 -44254 -6708 -44220
rect -6828 -44288 -6785 -44254
rect -6751 -44288 -6708 -44254
rect -6828 -44322 -6708 -44288
rect -6828 -44356 -6785 -44322
rect -6751 -44356 -6708 -44322
rect -6828 -44390 -6708 -44356
rect -6828 -44424 -6785 -44390
rect -6751 -44424 -6708 -44390
rect -6828 -44458 -6708 -44424
rect -6828 -44492 -6785 -44458
rect -6751 -44492 -6708 -44458
rect -6828 -44526 -6708 -44492
rect -6828 -44560 -6785 -44526
rect -6751 -44560 -6708 -44526
rect -6828 -44594 -6708 -44560
rect -6828 -44628 -6785 -44594
rect -6751 -44628 -6708 -44594
rect -6828 -44662 -6708 -44628
rect -6828 -44696 -6785 -44662
rect -6751 -44696 -6708 -44662
rect -6828 -44730 -6708 -44696
rect -6828 -44764 -6785 -44730
rect -6751 -44764 -6708 -44730
rect -6828 -44798 -6708 -44764
rect -6828 -44832 -6785 -44798
rect -6751 -44832 -6708 -44798
rect -6828 -44891 -6708 -44832
rect -6678 -44060 -6558 -43991
rect -6678 -44094 -6635 -44060
rect -6601 -44094 -6558 -44060
rect -6678 -44128 -6558 -44094
rect -6678 -44162 -6635 -44128
rect -6601 -44162 -6558 -44128
rect -6678 -44196 -6558 -44162
rect -6678 -44230 -6635 -44196
rect -6601 -44230 -6558 -44196
rect -6678 -44264 -6558 -44230
rect -6678 -44298 -6635 -44264
rect -6601 -44298 -6558 -44264
rect -6678 -44332 -6558 -44298
rect -6678 -44366 -6635 -44332
rect -6601 -44366 -6558 -44332
rect -6678 -44400 -6558 -44366
rect -6678 -44434 -6635 -44400
rect -6601 -44434 -6558 -44400
rect -6678 -44468 -6558 -44434
rect -6678 -44502 -6635 -44468
rect -6601 -44502 -6558 -44468
rect -6678 -44536 -6558 -44502
rect -6678 -44570 -6635 -44536
rect -6601 -44570 -6558 -44536
rect -6678 -44604 -6558 -44570
rect -6678 -44638 -6635 -44604
rect -6601 -44638 -6558 -44604
rect -6678 -44672 -6558 -44638
rect -6678 -44706 -6635 -44672
rect -6601 -44706 -6558 -44672
rect -6678 -44740 -6558 -44706
rect -6678 -44774 -6635 -44740
rect -6601 -44774 -6558 -44740
rect -6678 -44808 -6558 -44774
rect -6678 -44842 -6635 -44808
rect -6601 -44842 -6558 -44808
rect -6678 -44891 -6558 -44842
rect -6528 -44050 -6408 -43991
rect -6528 -44084 -6485 -44050
rect -6451 -44084 -6408 -44050
rect -6528 -44118 -6408 -44084
rect -6528 -44152 -6485 -44118
rect -6451 -44152 -6408 -44118
rect -6528 -44186 -6408 -44152
rect -6528 -44220 -6485 -44186
rect -6451 -44220 -6408 -44186
rect -6528 -44254 -6408 -44220
rect -6528 -44288 -6485 -44254
rect -6451 -44288 -6408 -44254
rect -6528 -44322 -6408 -44288
rect -6528 -44356 -6485 -44322
rect -6451 -44356 -6408 -44322
rect -6528 -44390 -6408 -44356
rect -6528 -44424 -6485 -44390
rect -6451 -44424 -6408 -44390
rect -6528 -44458 -6408 -44424
rect -6528 -44492 -6485 -44458
rect -6451 -44492 -6408 -44458
rect -6528 -44526 -6408 -44492
rect -6528 -44560 -6485 -44526
rect -6451 -44560 -6408 -44526
rect -6528 -44594 -6408 -44560
rect -6528 -44628 -6485 -44594
rect -6451 -44628 -6408 -44594
rect -6528 -44662 -6408 -44628
rect -6528 -44696 -6485 -44662
rect -6451 -44696 -6408 -44662
rect -6528 -44730 -6408 -44696
rect -6528 -44764 -6485 -44730
rect -6451 -44764 -6408 -44730
rect -6528 -44798 -6408 -44764
rect -6528 -44832 -6485 -44798
rect -6451 -44832 -6408 -44798
rect -6528 -44891 -6408 -44832
rect -5422 -44050 -5302 -43991
rect -5422 -44084 -5379 -44050
rect -5345 -44084 -5302 -44050
rect -5422 -44118 -5302 -44084
rect -5422 -44152 -5379 -44118
rect -5345 -44152 -5302 -44118
rect -5422 -44186 -5302 -44152
rect -5422 -44220 -5379 -44186
rect -5345 -44220 -5302 -44186
rect -5422 -44254 -5302 -44220
rect -5422 -44288 -5379 -44254
rect -5345 -44288 -5302 -44254
rect -5422 -44322 -5302 -44288
rect -5422 -44356 -5379 -44322
rect -5345 -44356 -5302 -44322
rect -5422 -44390 -5302 -44356
rect -5422 -44424 -5379 -44390
rect -5345 -44424 -5302 -44390
rect -5422 -44458 -5302 -44424
rect -5422 -44492 -5379 -44458
rect -5345 -44492 -5302 -44458
rect -5422 -44526 -5302 -44492
rect -5422 -44560 -5379 -44526
rect -5345 -44560 -5302 -44526
rect -5422 -44594 -5302 -44560
rect -5422 -44628 -5379 -44594
rect -5345 -44628 -5302 -44594
rect -5422 -44662 -5302 -44628
rect -5422 -44696 -5379 -44662
rect -5345 -44696 -5302 -44662
rect -5422 -44730 -5302 -44696
rect -5422 -44764 -5379 -44730
rect -5345 -44764 -5302 -44730
rect -5422 -44798 -5302 -44764
rect -5422 -44832 -5379 -44798
rect -5345 -44832 -5302 -44798
rect -5422 -44891 -5302 -44832
rect -5272 -44060 -5152 -43991
rect -5272 -44094 -5229 -44060
rect -5195 -44094 -5152 -44060
rect -5272 -44128 -5152 -44094
rect -5272 -44162 -5229 -44128
rect -5195 -44162 -5152 -44128
rect -5272 -44196 -5152 -44162
rect -5272 -44230 -5229 -44196
rect -5195 -44230 -5152 -44196
rect -5272 -44264 -5152 -44230
rect -5272 -44298 -5229 -44264
rect -5195 -44298 -5152 -44264
rect -5272 -44332 -5152 -44298
rect -5272 -44366 -5229 -44332
rect -5195 -44366 -5152 -44332
rect -5272 -44400 -5152 -44366
rect -5272 -44434 -5229 -44400
rect -5195 -44434 -5152 -44400
rect -5272 -44468 -5152 -44434
rect -5272 -44502 -5229 -44468
rect -5195 -44502 -5152 -44468
rect -5272 -44536 -5152 -44502
rect -5272 -44570 -5229 -44536
rect -5195 -44570 -5152 -44536
rect -5272 -44604 -5152 -44570
rect -5272 -44638 -5229 -44604
rect -5195 -44638 -5152 -44604
rect -5272 -44672 -5152 -44638
rect -5272 -44706 -5229 -44672
rect -5195 -44706 -5152 -44672
rect -5272 -44740 -5152 -44706
rect -5272 -44774 -5229 -44740
rect -5195 -44774 -5152 -44740
rect -5272 -44808 -5152 -44774
rect -5272 -44842 -5229 -44808
rect -5195 -44842 -5152 -44808
rect -5272 -44891 -5152 -44842
rect -5122 -44050 -5002 -43991
rect -5122 -44084 -5079 -44050
rect -5045 -44084 -5002 -44050
rect -5122 -44118 -5002 -44084
rect -5122 -44152 -5079 -44118
rect -5045 -44152 -5002 -44118
rect -5122 -44186 -5002 -44152
rect -5122 -44220 -5079 -44186
rect -5045 -44220 -5002 -44186
rect -5122 -44254 -5002 -44220
rect -5122 -44288 -5079 -44254
rect -5045 -44288 -5002 -44254
rect -5122 -44322 -5002 -44288
rect -5122 -44356 -5079 -44322
rect -5045 -44356 -5002 -44322
rect -5122 -44390 -5002 -44356
rect -5122 -44424 -5079 -44390
rect -5045 -44424 -5002 -44390
rect -5122 -44458 -5002 -44424
rect -5122 -44492 -5079 -44458
rect -5045 -44492 -5002 -44458
rect -5122 -44526 -5002 -44492
rect -5122 -44560 -5079 -44526
rect -5045 -44560 -5002 -44526
rect -5122 -44594 -5002 -44560
rect -5122 -44628 -5079 -44594
rect -5045 -44628 -5002 -44594
rect -5122 -44662 -5002 -44628
rect -5122 -44696 -5079 -44662
rect -5045 -44696 -5002 -44662
rect -5122 -44730 -5002 -44696
rect -5122 -44764 -5079 -44730
rect -5045 -44764 -5002 -44730
rect -5122 -44798 -5002 -44764
rect -5122 -44832 -5079 -44798
rect -5045 -44832 -5002 -44798
rect -5122 -44891 -5002 -44832
rect -4972 -44050 -4852 -43991
rect -4972 -44084 -4929 -44050
rect -4895 -44084 -4852 -44050
rect -4972 -44118 -4852 -44084
rect -4972 -44152 -4929 -44118
rect -4895 -44152 -4852 -44118
rect -4972 -44186 -4852 -44152
rect -4972 -44220 -4929 -44186
rect -4895 -44220 -4852 -44186
rect -4972 -44254 -4852 -44220
rect -4972 -44288 -4929 -44254
rect -4895 -44288 -4852 -44254
rect -4972 -44322 -4852 -44288
rect -4972 -44356 -4929 -44322
rect -4895 -44356 -4852 -44322
rect -4972 -44390 -4852 -44356
rect -4972 -44424 -4929 -44390
rect -4895 -44424 -4852 -44390
rect -4972 -44458 -4852 -44424
rect -4972 -44492 -4929 -44458
rect -4895 -44492 -4852 -44458
rect -4972 -44526 -4852 -44492
rect -4972 -44560 -4929 -44526
rect -4895 -44560 -4852 -44526
rect -4972 -44594 -4852 -44560
rect -4972 -44628 -4929 -44594
rect -4895 -44628 -4852 -44594
rect -4972 -44662 -4852 -44628
rect -4972 -44696 -4929 -44662
rect -4895 -44696 -4852 -44662
rect -4972 -44730 -4852 -44696
rect -4972 -44764 -4929 -44730
rect -4895 -44764 -4852 -44730
rect -4972 -44798 -4852 -44764
rect -4972 -44832 -4929 -44798
rect -4895 -44832 -4852 -44798
rect -4972 -44891 -4852 -44832
rect -4822 -44050 -4702 -43991
rect -4822 -44084 -4779 -44050
rect -4745 -44084 -4702 -44050
rect -4822 -44118 -4702 -44084
rect -4822 -44152 -4779 -44118
rect -4745 -44152 -4702 -44118
rect -4822 -44186 -4702 -44152
rect -4822 -44220 -4779 -44186
rect -4745 -44220 -4702 -44186
rect -4822 -44254 -4702 -44220
rect -4822 -44288 -4779 -44254
rect -4745 -44288 -4702 -44254
rect -4822 -44322 -4702 -44288
rect -4822 -44356 -4779 -44322
rect -4745 -44356 -4702 -44322
rect -4822 -44390 -4702 -44356
rect -4822 -44424 -4779 -44390
rect -4745 -44424 -4702 -44390
rect -4822 -44458 -4702 -44424
rect -4822 -44492 -4779 -44458
rect -4745 -44492 -4702 -44458
rect -4822 -44526 -4702 -44492
rect -4822 -44560 -4779 -44526
rect -4745 -44560 -4702 -44526
rect -4822 -44594 -4702 -44560
rect -4822 -44628 -4779 -44594
rect -4745 -44628 -4702 -44594
rect -4822 -44662 -4702 -44628
rect -4822 -44696 -4779 -44662
rect -4745 -44696 -4702 -44662
rect -4822 -44730 -4702 -44696
rect -4822 -44764 -4779 -44730
rect -4745 -44764 -4702 -44730
rect -4822 -44798 -4702 -44764
rect -4822 -44832 -4779 -44798
rect -4745 -44832 -4702 -44798
rect -4822 -44891 -4702 -44832
rect -4672 -44050 -4552 -43991
rect -4672 -44084 -4629 -44050
rect -4595 -44084 -4552 -44050
rect -4672 -44118 -4552 -44084
rect -4672 -44152 -4629 -44118
rect -4595 -44152 -4552 -44118
rect -4672 -44186 -4552 -44152
rect -4672 -44220 -4629 -44186
rect -4595 -44220 -4552 -44186
rect -4672 -44254 -4552 -44220
rect -4672 -44288 -4629 -44254
rect -4595 -44288 -4552 -44254
rect -4672 -44322 -4552 -44288
rect -4672 -44356 -4629 -44322
rect -4595 -44356 -4552 -44322
rect -4672 -44390 -4552 -44356
rect -4672 -44424 -4629 -44390
rect -4595 -44424 -4552 -44390
rect -4672 -44458 -4552 -44424
rect -4672 -44492 -4629 -44458
rect -4595 -44492 -4552 -44458
rect -4672 -44526 -4552 -44492
rect -4672 -44560 -4629 -44526
rect -4595 -44560 -4552 -44526
rect -4672 -44594 -4552 -44560
rect -4672 -44628 -4629 -44594
rect -4595 -44628 -4552 -44594
rect -4672 -44662 -4552 -44628
rect -4672 -44696 -4629 -44662
rect -4595 -44696 -4552 -44662
rect -4672 -44730 -4552 -44696
rect -4672 -44764 -4629 -44730
rect -4595 -44764 -4552 -44730
rect -4672 -44798 -4552 -44764
rect -4672 -44832 -4629 -44798
rect -4595 -44832 -4552 -44798
rect -4672 -44891 -4552 -44832
rect -4522 -44050 -4402 -43991
rect -4522 -44084 -4479 -44050
rect -4445 -44084 -4402 -44050
rect -4522 -44118 -4402 -44084
rect -4522 -44152 -4479 -44118
rect -4445 -44152 -4402 -44118
rect -4522 -44186 -4402 -44152
rect -4522 -44220 -4479 -44186
rect -4445 -44220 -4402 -44186
rect -4522 -44254 -4402 -44220
rect -4522 -44288 -4479 -44254
rect -4445 -44288 -4402 -44254
rect -4522 -44322 -4402 -44288
rect -4522 -44356 -4479 -44322
rect -4445 -44356 -4402 -44322
rect -4522 -44390 -4402 -44356
rect -4522 -44424 -4479 -44390
rect -4445 -44424 -4402 -44390
rect -4522 -44458 -4402 -44424
rect -4522 -44492 -4479 -44458
rect -4445 -44492 -4402 -44458
rect -4522 -44526 -4402 -44492
rect -4522 -44560 -4479 -44526
rect -4445 -44560 -4402 -44526
rect -4522 -44594 -4402 -44560
rect -4522 -44628 -4479 -44594
rect -4445 -44628 -4402 -44594
rect -4522 -44662 -4402 -44628
rect -4522 -44696 -4479 -44662
rect -4445 -44696 -4402 -44662
rect -4522 -44730 -4402 -44696
rect -4522 -44764 -4479 -44730
rect -4445 -44764 -4402 -44730
rect -4522 -44798 -4402 -44764
rect -4522 -44832 -4479 -44798
rect -4445 -44832 -4402 -44798
rect -4522 -44891 -4402 -44832
rect -4372 -44050 -4252 -43991
rect -4372 -44084 -4329 -44050
rect -4295 -44084 -4252 -44050
rect -4372 -44118 -4252 -44084
rect -4372 -44152 -4329 -44118
rect -4295 -44152 -4252 -44118
rect -4372 -44186 -4252 -44152
rect -4372 -44220 -4329 -44186
rect -4295 -44220 -4252 -44186
rect -4372 -44254 -4252 -44220
rect -4372 -44288 -4329 -44254
rect -4295 -44288 -4252 -44254
rect -4372 -44322 -4252 -44288
rect -4372 -44356 -4329 -44322
rect -4295 -44356 -4252 -44322
rect -4372 -44390 -4252 -44356
rect -4372 -44424 -4329 -44390
rect -4295 -44424 -4252 -44390
rect -4372 -44458 -4252 -44424
rect -4372 -44492 -4329 -44458
rect -4295 -44492 -4252 -44458
rect -4372 -44526 -4252 -44492
rect -4372 -44560 -4329 -44526
rect -4295 -44560 -4252 -44526
rect -4372 -44594 -4252 -44560
rect -4372 -44628 -4329 -44594
rect -4295 -44628 -4252 -44594
rect -4372 -44662 -4252 -44628
rect -4372 -44696 -4329 -44662
rect -4295 -44696 -4252 -44662
rect -4372 -44730 -4252 -44696
rect -4372 -44764 -4329 -44730
rect -4295 -44764 -4252 -44730
rect -4372 -44798 -4252 -44764
rect -4372 -44832 -4329 -44798
rect -4295 -44832 -4252 -44798
rect -4372 -44891 -4252 -44832
rect -4222 -44050 -4102 -43991
rect -4222 -44084 -4179 -44050
rect -4145 -44084 -4102 -44050
rect -4222 -44118 -4102 -44084
rect -4222 -44152 -4179 -44118
rect -4145 -44152 -4102 -44118
rect -4222 -44186 -4102 -44152
rect -4222 -44220 -4179 -44186
rect -4145 -44220 -4102 -44186
rect -4222 -44254 -4102 -44220
rect -4222 -44288 -4179 -44254
rect -4145 -44288 -4102 -44254
rect -4222 -44322 -4102 -44288
rect -4222 -44356 -4179 -44322
rect -4145 -44356 -4102 -44322
rect -4222 -44390 -4102 -44356
rect -4222 -44424 -4179 -44390
rect -4145 -44424 -4102 -44390
rect -4222 -44458 -4102 -44424
rect -4222 -44492 -4179 -44458
rect -4145 -44492 -4102 -44458
rect -4222 -44526 -4102 -44492
rect -4222 -44560 -4179 -44526
rect -4145 -44560 -4102 -44526
rect -4222 -44594 -4102 -44560
rect -4222 -44628 -4179 -44594
rect -4145 -44628 -4102 -44594
rect -4222 -44662 -4102 -44628
rect -4222 -44696 -4179 -44662
rect -4145 -44696 -4102 -44662
rect -4222 -44730 -4102 -44696
rect -4222 -44764 -4179 -44730
rect -4145 -44764 -4102 -44730
rect -4222 -44798 -4102 -44764
rect -4222 -44832 -4179 -44798
rect -4145 -44832 -4102 -44798
rect -4222 -44891 -4102 -44832
rect -4072 -44050 -3952 -43991
rect -4072 -44084 -4029 -44050
rect -3995 -44084 -3952 -44050
rect -4072 -44118 -3952 -44084
rect -4072 -44152 -4029 -44118
rect -3995 -44152 -3952 -44118
rect -4072 -44186 -3952 -44152
rect -4072 -44220 -4029 -44186
rect -3995 -44220 -3952 -44186
rect -4072 -44254 -3952 -44220
rect -4072 -44288 -4029 -44254
rect -3995 -44288 -3952 -44254
rect -4072 -44322 -3952 -44288
rect -4072 -44356 -4029 -44322
rect -3995 -44356 -3952 -44322
rect -4072 -44390 -3952 -44356
rect -4072 -44424 -4029 -44390
rect -3995 -44424 -3952 -44390
rect -4072 -44458 -3952 -44424
rect -4072 -44492 -4029 -44458
rect -3995 -44492 -3952 -44458
rect -4072 -44526 -3952 -44492
rect -4072 -44560 -4029 -44526
rect -3995 -44560 -3952 -44526
rect -4072 -44594 -3952 -44560
rect -4072 -44628 -4029 -44594
rect -3995 -44628 -3952 -44594
rect -4072 -44662 -3952 -44628
rect -4072 -44696 -4029 -44662
rect -3995 -44696 -3952 -44662
rect -4072 -44730 -3952 -44696
rect -4072 -44764 -4029 -44730
rect -3995 -44764 -3952 -44730
rect -4072 -44798 -3952 -44764
rect -4072 -44832 -4029 -44798
rect -3995 -44832 -3952 -44798
rect -4072 -44891 -3952 -44832
rect -3922 -44050 -3802 -43991
rect -3922 -44084 -3879 -44050
rect -3845 -44084 -3802 -44050
rect -3922 -44118 -3802 -44084
rect -3922 -44152 -3879 -44118
rect -3845 -44152 -3802 -44118
rect -3922 -44186 -3802 -44152
rect -3922 -44220 -3879 -44186
rect -3845 -44220 -3802 -44186
rect -3922 -44254 -3802 -44220
rect -3922 -44288 -3879 -44254
rect -3845 -44288 -3802 -44254
rect -3922 -44322 -3802 -44288
rect -3922 -44356 -3879 -44322
rect -3845 -44356 -3802 -44322
rect -3922 -44390 -3802 -44356
rect -3922 -44424 -3879 -44390
rect -3845 -44424 -3802 -44390
rect -3922 -44458 -3802 -44424
rect -3922 -44492 -3879 -44458
rect -3845 -44492 -3802 -44458
rect -3922 -44526 -3802 -44492
rect -3922 -44560 -3879 -44526
rect -3845 -44560 -3802 -44526
rect -3922 -44594 -3802 -44560
rect -3922 -44628 -3879 -44594
rect -3845 -44628 -3802 -44594
rect -3922 -44662 -3802 -44628
rect -3922 -44696 -3879 -44662
rect -3845 -44696 -3802 -44662
rect -3922 -44730 -3802 -44696
rect -3922 -44764 -3879 -44730
rect -3845 -44764 -3802 -44730
rect -3922 -44798 -3802 -44764
rect -3922 -44832 -3879 -44798
rect -3845 -44832 -3802 -44798
rect -3922 -44891 -3802 -44832
rect -3772 -44060 -3652 -43991
rect -3772 -44094 -3729 -44060
rect -3695 -44094 -3652 -44060
rect -3772 -44128 -3652 -44094
rect -3772 -44162 -3729 -44128
rect -3695 -44162 -3652 -44128
rect -3772 -44196 -3652 -44162
rect -3772 -44230 -3729 -44196
rect -3695 -44230 -3652 -44196
rect -3772 -44264 -3652 -44230
rect -3772 -44298 -3729 -44264
rect -3695 -44298 -3652 -44264
rect -3772 -44332 -3652 -44298
rect -3772 -44366 -3729 -44332
rect -3695 -44366 -3652 -44332
rect -3772 -44400 -3652 -44366
rect -3772 -44434 -3729 -44400
rect -3695 -44434 -3652 -44400
rect -3772 -44468 -3652 -44434
rect -3772 -44502 -3729 -44468
rect -3695 -44502 -3652 -44468
rect -3772 -44536 -3652 -44502
rect -3772 -44570 -3729 -44536
rect -3695 -44570 -3652 -44536
rect -3772 -44604 -3652 -44570
rect -3772 -44638 -3729 -44604
rect -3695 -44638 -3652 -44604
rect -3772 -44672 -3652 -44638
rect -3772 -44706 -3729 -44672
rect -3695 -44706 -3652 -44672
rect -3772 -44740 -3652 -44706
rect -3772 -44774 -3729 -44740
rect -3695 -44774 -3652 -44740
rect -3772 -44808 -3652 -44774
rect -3772 -44842 -3729 -44808
rect -3695 -44842 -3652 -44808
rect -3772 -44891 -3652 -44842
rect -3622 -44050 -3502 -43991
rect -3622 -44084 -3579 -44050
rect -3545 -44084 -3502 -44050
rect -3622 -44118 -3502 -44084
rect -3622 -44152 -3579 -44118
rect -3545 -44152 -3502 -44118
rect -3622 -44186 -3502 -44152
rect -3622 -44220 -3579 -44186
rect -3545 -44220 -3502 -44186
rect -3622 -44254 -3502 -44220
rect -3622 -44288 -3579 -44254
rect -3545 -44288 -3502 -44254
rect -3622 -44322 -3502 -44288
rect -3622 -44356 -3579 -44322
rect -3545 -44356 -3502 -44322
rect -3622 -44390 -3502 -44356
rect -3622 -44424 -3579 -44390
rect -3545 -44424 -3502 -44390
rect -3622 -44458 -3502 -44424
rect -3622 -44492 -3579 -44458
rect -3545 -44492 -3502 -44458
rect -3622 -44526 -3502 -44492
rect -3622 -44560 -3579 -44526
rect -3545 -44560 -3502 -44526
rect -3622 -44594 -3502 -44560
rect -3622 -44628 -3579 -44594
rect -3545 -44628 -3502 -44594
rect -3622 -44662 -3502 -44628
rect -3622 -44696 -3579 -44662
rect -3545 -44696 -3502 -44662
rect -3622 -44730 -3502 -44696
rect -3622 -44764 -3579 -44730
rect -3545 -44764 -3502 -44730
rect -3622 -44798 -3502 -44764
rect -3622 -44832 -3579 -44798
rect -3545 -44832 -3502 -44798
rect -3622 -44891 -3502 -44832
rect -3472 -44050 -3352 -43991
rect -3472 -44084 -3429 -44050
rect -3395 -44084 -3352 -44050
rect -3472 -44118 -3352 -44084
rect -3472 -44152 -3429 -44118
rect -3395 -44152 -3352 -44118
rect -3472 -44186 -3352 -44152
rect -3472 -44220 -3429 -44186
rect -3395 -44220 -3352 -44186
rect -3472 -44254 -3352 -44220
rect -3472 -44288 -3429 -44254
rect -3395 -44288 -3352 -44254
rect -3472 -44322 -3352 -44288
rect -3472 -44356 -3429 -44322
rect -3395 -44356 -3352 -44322
rect -3472 -44390 -3352 -44356
rect -3472 -44424 -3429 -44390
rect -3395 -44424 -3352 -44390
rect -3472 -44458 -3352 -44424
rect -3472 -44492 -3429 -44458
rect -3395 -44492 -3352 -44458
rect -3472 -44526 -3352 -44492
rect -3472 -44560 -3429 -44526
rect -3395 -44560 -3352 -44526
rect -3472 -44594 -3352 -44560
rect -3472 -44628 -3429 -44594
rect -3395 -44628 -3352 -44594
rect -3472 -44662 -3352 -44628
rect -3472 -44696 -3429 -44662
rect -3395 -44696 -3352 -44662
rect -3472 -44730 -3352 -44696
rect -3472 -44764 -3429 -44730
rect -3395 -44764 -3352 -44730
rect -3472 -44798 -3352 -44764
rect -3472 -44832 -3429 -44798
rect -3395 -44832 -3352 -44798
rect -3472 -44891 -3352 -44832
rect -3322 -44050 -3202 -43991
rect -3322 -44084 -3279 -44050
rect -3245 -44084 -3202 -44050
rect -3322 -44118 -3202 -44084
rect -3322 -44152 -3279 -44118
rect -3245 -44152 -3202 -44118
rect -3322 -44186 -3202 -44152
rect -3322 -44220 -3279 -44186
rect -3245 -44220 -3202 -44186
rect -3322 -44254 -3202 -44220
rect -3322 -44288 -3279 -44254
rect -3245 -44288 -3202 -44254
rect -3322 -44322 -3202 -44288
rect -3322 -44356 -3279 -44322
rect -3245 -44356 -3202 -44322
rect -3322 -44390 -3202 -44356
rect -3322 -44424 -3279 -44390
rect -3245 -44424 -3202 -44390
rect -3322 -44458 -3202 -44424
rect -3322 -44492 -3279 -44458
rect -3245 -44492 -3202 -44458
rect -3322 -44526 -3202 -44492
rect -3322 -44560 -3279 -44526
rect -3245 -44560 -3202 -44526
rect -3322 -44594 -3202 -44560
rect -3322 -44628 -3279 -44594
rect -3245 -44628 -3202 -44594
rect -3322 -44662 -3202 -44628
rect -3322 -44696 -3279 -44662
rect -3245 -44696 -3202 -44662
rect -3322 -44730 -3202 -44696
rect -3322 -44764 -3279 -44730
rect -3245 -44764 -3202 -44730
rect -3322 -44798 -3202 -44764
rect -3322 -44832 -3279 -44798
rect -3245 -44832 -3202 -44798
rect -3322 -44891 -3202 -44832
rect -3172 -44050 -3052 -43991
rect -3172 -44084 -3129 -44050
rect -3095 -44084 -3052 -44050
rect -3172 -44118 -3052 -44084
rect -3172 -44152 -3129 -44118
rect -3095 -44152 -3052 -44118
rect -3172 -44186 -3052 -44152
rect -3172 -44220 -3129 -44186
rect -3095 -44220 -3052 -44186
rect -3172 -44254 -3052 -44220
rect -3172 -44288 -3129 -44254
rect -3095 -44288 -3052 -44254
rect -3172 -44322 -3052 -44288
rect -3172 -44356 -3129 -44322
rect -3095 -44356 -3052 -44322
rect -3172 -44390 -3052 -44356
rect -3172 -44424 -3129 -44390
rect -3095 -44424 -3052 -44390
rect -3172 -44458 -3052 -44424
rect -3172 -44492 -3129 -44458
rect -3095 -44492 -3052 -44458
rect -3172 -44526 -3052 -44492
rect -3172 -44560 -3129 -44526
rect -3095 -44560 -3052 -44526
rect -3172 -44594 -3052 -44560
rect -3172 -44628 -3129 -44594
rect -3095 -44628 -3052 -44594
rect -3172 -44662 -3052 -44628
rect -3172 -44696 -3129 -44662
rect -3095 -44696 -3052 -44662
rect -3172 -44730 -3052 -44696
rect -3172 -44764 -3129 -44730
rect -3095 -44764 -3052 -44730
rect -3172 -44798 -3052 -44764
rect -3172 -44832 -3129 -44798
rect -3095 -44832 -3052 -44798
rect -3172 -44891 -3052 -44832
rect -3022 -44050 -2902 -43991
rect -3022 -44084 -2979 -44050
rect -2945 -44084 -2902 -44050
rect -3022 -44118 -2902 -44084
rect -3022 -44152 -2979 -44118
rect -2945 -44152 -2902 -44118
rect -3022 -44186 -2902 -44152
rect -3022 -44220 -2979 -44186
rect -2945 -44220 -2902 -44186
rect -3022 -44254 -2902 -44220
rect -3022 -44288 -2979 -44254
rect -2945 -44288 -2902 -44254
rect -3022 -44322 -2902 -44288
rect -3022 -44356 -2979 -44322
rect -2945 -44356 -2902 -44322
rect -3022 -44390 -2902 -44356
rect -3022 -44424 -2979 -44390
rect -2945 -44424 -2902 -44390
rect -3022 -44458 -2902 -44424
rect -3022 -44492 -2979 -44458
rect -2945 -44492 -2902 -44458
rect -3022 -44526 -2902 -44492
rect -3022 -44560 -2979 -44526
rect -2945 -44560 -2902 -44526
rect -3022 -44594 -2902 -44560
rect -3022 -44628 -2979 -44594
rect -2945 -44628 -2902 -44594
rect -3022 -44662 -2902 -44628
rect -3022 -44696 -2979 -44662
rect -2945 -44696 -2902 -44662
rect -3022 -44730 -2902 -44696
rect -3022 -44764 -2979 -44730
rect -2945 -44764 -2902 -44730
rect -3022 -44798 -2902 -44764
rect -3022 -44832 -2979 -44798
rect -2945 -44832 -2902 -44798
rect -3022 -44891 -2902 -44832
rect -2872 -44050 -2752 -43991
rect -2872 -44084 -2829 -44050
rect -2795 -44084 -2752 -44050
rect -2872 -44118 -2752 -44084
rect -2872 -44152 -2829 -44118
rect -2795 -44152 -2752 -44118
rect -2872 -44186 -2752 -44152
rect -2872 -44220 -2829 -44186
rect -2795 -44220 -2752 -44186
rect -2872 -44254 -2752 -44220
rect -2872 -44288 -2829 -44254
rect -2795 -44288 -2752 -44254
rect -2872 -44322 -2752 -44288
rect -2872 -44356 -2829 -44322
rect -2795 -44356 -2752 -44322
rect -2872 -44390 -2752 -44356
rect -2872 -44424 -2829 -44390
rect -2795 -44424 -2752 -44390
rect -2872 -44458 -2752 -44424
rect -2872 -44492 -2829 -44458
rect -2795 -44492 -2752 -44458
rect -2872 -44526 -2752 -44492
rect -2872 -44560 -2829 -44526
rect -2795 -44560 -2752 -44526
rect -2872 -44594 -2752 -44560
rect -2872 -44628 -2829 -44594
rect -2795 -44628 -2752 -44594
rect -2872 -44662 -2752 -44628
rect -2872 -44696 -2829 -44662
rect -2795 -44696 -2752 -44662
rect -2872 -44730 -2752 -44696
rect -2872 -44764 -2829 -44730
rect -2795 -44764 -2752 -44730
rect -2872 -44798 -2752 -44764
rect -2872 -44832 -2829 -44798
rect -2795 -44832 -2752 -44798
rect -2872 -44891 -2752 -44832
rect -2722 -44050 -2602 -43991
rect -2722 -44084 -2679 -44050
rect -2645 -44084 -2602 -44050
rect -2722 -44118 -2602 -44084
rect -2722 -44152 -2679 -44118
rect -2645 -44152 -2602 -44118
rect -2722 -44186 -2602 -44152
rect -2722 -44220 -2679 -44186
rect -2645 -44220 -2602 -44186
rect -2722 -44254 -2602 -44220
rect -2722 -44288 -2679 -44254
rect -2645 -44288 -2602 -44254
rect -2722 -44322 -2602 -44288
rect -2722 -44356 -2679 -44322
rect -2645 -44356 -2602 -44322
rect -2722 -44390 -2602 -44356
rect -2722 -44424 -2679 -44390
rect -2645 -44424 -2602 -44390
rect -2722 -44458 -2602 -44424
rect -2722 -44492 -2679 -44458
rect -2645 -44492 -2602 -44458
rect -2722 -44526 -2602 -44492
rect -2722 -44560 -2679 -44526
rect -2645 -44560 -2602 -44526
rect -2722 -44594 -2602 -44560
rect -2722 -44628 -2679 -44594
rect -2645 -44628 -2602 -44594
rect -2722 -44662 -2602 -44628
rect -2722 -44696 -2679 -44662
rect -2645 -44696 -2602 -44662
rect -2722 -44730 -2602 -44696
rect -2722 -44764 -2679 -44730
rect -2645 -44764 -2602 -44730
rect -2722 -44798 -2602 -44764
rect -2722 -44832 -2679 -44798
rect -2645 -44832 -2602 -44798
rect -2722 -44891 -2602 -44832
rect -2572 -44050 -2452 -43991
rect -2572 -44084 -2529 -44050
rect -2495 -44084 -2452 -44050
rect -2572 -44118 -2452 -44084
rect -2572 -44152 -2529 -44118
rect -2495 -44152 -2452 -44118
rect -2572 -44186 -2452 -44152
rect -2572 -44220 -2529 -44186
rect -2495 -44220 -2452 -44186
rect -2572 -44254 -2452 -44220
rect -2572 -44288 -2529 -44254
rect -2495 -44288 -2452 -44254
rect -2572 -44322 -2452 -44288
rect -2572 -44356 -2529 -44322
rect -2495 -44356 -2452 -44322
rect -2572 -44390 -2452 -44356
rect -2572 -44424 -2529 -44390
rect -2495 -44424 -2452 -44390
rect -2572 -44458 -2452 -44424
rect -2572 -44492 -2529 -44458
rect -2495 -44492 -2452 -44458
rect -2572 -44526 -2452 -44492
rect -2572 -44560 -2529 -44526
rect -2495 -44560 -2452 -44526
rect -2572 -44594 -2452 -44560
rect -2572 -44628 -2529 -44594
rect -2495 -44628 -2452 -44594
rect -2572 -44662 -2452 -44628
rect -2572 -44696 -2529 -44662
rect -2495 -44696 -2452 -44662
rect -2572 -44730 -2452 -44696
rect -2572 -44764 -2529 -44730
rect -2495 -44764 -2452 -44730
rect -2572 -44798 -2452 -44764
rect -2572 -44832 -2529 -44798
rect -2495 -44832 -2452 -44798
rect -2572 -44891 -2452 -44832
rect -2422 -44050 -2302 -43991
rect -2422 -44084 -2379 -44050
rect -2345 -44084 -2302 -44050
rect -2422 -44118 -2302 -44084
rect -2422 -44152 -2379 -44118
rect -2345 -44152 -2302 -44118
rect -2422 -44186 -2302 -44152
rect -2422 -44220 -2379 -44186
rect -2345 -44220 -2302 -44186
rect -2422 -44254 -2302 -44220
rect -2422 -44288 -2379 -44254
rect -2345 -44288 -2302 -44254
rect -2422 -44322 -2302 -44288
rect -2422 -44356 -2379 -44322
rect -2345 -44356 -2302 -44322
rect -2422 -44390 -2302 -44356
rect -2422 -44424 -2379 -44390
rect -2345 -44424 -2302 -44390
rect -2422 -44458 -2302 -44424
rect -2422 -44492 -2379 -44458
rect -2345 -44492 -2302 -44458
rect -2422 -44526 -2302 -44492
rect -2422 -44560 -2379 -44526
rect -2345 -44560 -2302 -44526
rect -2422 -44594 -2302 -44560
rect -2422 -44628 -2379 -44594
rect -2345 -44628 -2302 -44594
rect -2422 -44662 -2302 -44628
rect -2422 -44696 -2379 -44662
rect -2345 -44696 -2302 -44662
rect -2422 -44730 -2302 -44696
rect -2422 -44764 -2379 -44730
rect -2345 -44764 -2302 -44730
rect -2422 -44798 -2302 -44764
rect -2422 -44832 -2379 -44798
rect -2345 -44832 -2302 -44798
rect -2422 -44891 -2302 -44832
rect -6497 -47234 -6377 -47176
rect -6497 -47268 -6454 -47234
rect -6420 -47268 -6377 -47234
rect -6497 -47335 -6377 -47268
rect -6497 -47369 -6454 -47335
rect -6420 -47369 -6377 -47335
rect -6497 -47403 -6377 -47369
rect -6497 -47437 -6454 -47403
rect -6420 -47437 -6377 -47403
rect -6497 -47471 -6377 -47437
rect -6497 -47505 -6454 -47471
rect -6420 -47505 -6377 -47471
rect -6497 -47539 -6377 -47505
rect -6497 -47573 -6454 -47539
rect -6420 -47573 -6377 -47539
rect -6497 -47607 -6377 -47573
rect -6497 -47641 -6454 -47607
rect -6420 -47641 -6377 -47607
rect -6497 -47675 -6377 -47641
rect -6497 -47709 -6454 -47675
rect -6420 -47709 -6377 -47675
rect -6497 -47743 -6377 -47709
rect -6497 -47777 -6454 -47743
rect -6420 -47777 -6377 -47743
rect -6497 -47811 -6377 -47777
rect -6497 -47845 -6454 -47811
rect -6420 -47845 -6377 -47811
rect -6497 -47879 -6377 -47845
rect -6497 -47913 -6454 -47879
rect -6420 -47913 -6377 -47879
rect -6497 -47947 -6377 -47913
rect -6497 -47981 -6454 -47947
rect -6420 -47981 -6377 -47947
rect -6497 -48015 -6377 -47981
rect -6497 -48049 -6454 -48015
rect -6420 -48049 -6377 -48015
rect -6497 -48083 -6377 -48049
rect -6497 -48117 -6454 -48083
rect -6420 -48117 -6377 -48083
rect -6497 -48176 -6377 -48117
rect -6347 -47234 -6227 -47176
rect -6347 -47268 -6304 -47234
rect -6270 -47268 -6227 -47234
rect -6347 -47345 -6227 -47268
rect -6347 -47379 -6304 -47345
rect -6270 -47379 -6227 -47345
rect -6347 -47413 -6227 -47379
rect -6347 -47447 -6304 -47413
rect -6270 -47447 -6227 -47413
rect -6347 -47481 -6227 -47447
rect -6347 -47515 -6304 -47481
rect -6270 -47515 -6227 -47481
rect -6347 -47549 -6227 -47515
rect -6347 -47583 -6304 -47549
rect -6270 -47583 -6227 -47549
rect -6347 -47617 -6227 -47583
rect -6347 -47651 -6304 -47617
rect -6270 -47651 -6227 -47617
rect -6347 -47685 -6227 -47651
rect -6347 -47719 -6304 -47685
rect -6270 -47719 -6227 -47685
rect -6347 -47753 -6227 -47719
rect -6347 -47787 -6304 -47753
rect -6270 -47787 -6227 -47753
rect -6347 -47821 -6227 -47787
rect -6347 -47855 -6304 -47821
rect -6270 -47855 -6227 -47821
rect -6347 -47889 -6227 -47855
rect -6347 -47923 -6304 -47889
rect -6270 -47923 -6227 -47889
rect -6347 -47957 -6227 -47923
rect -6347 -47991 -6304 -47957
rect -6270 -47991 -6227 -47957
rect -6347 -48025 -6227 -47991
rect -6347 -48059 -6304 -48025
rect -6270 -48059 -6227 -48025
rect -6347 -48093 -6227 -48059
rect -6347 -48127 -6304 -48093
rect -6270 -48127 -6227 -48093
rect -6347 -48176 -6227 -48127
rect -6197 -47234 -6077 -47176
rect -6197 -47268 -6154 -47234
rect -6120 -47268 -6077 -47234
rect -6197 -47335 -6077 -47268
rect -6197 -47369 -6154 -47335
rect -6120 -47369 -6077 -47335
rect -6197 -47403 -6077 -47369
rect -6197 -47437 -6154 -47403
rect -6120 -47437 -6077 -47403
rect -6197 -47471 -6077 -47437
rect -6197 -47505 -6154 -47471
rect -6120 -47505 -6077 -47471
rect -6197 -47539 -6077 -47505
rect -6197 -47573 -6154 -47539
rect -6120 -47573 -6077 -47539
rect -6197 -47607 -6077 -47573
rect -6197 -47641 -6154 -47607
rect -6120 -47641 -6077 -47607
rect -6197 -47675 -6077 -47641
rect -6197 -47709 -6154 -47675
rect -6120 -47709 -6077 -47675
rect -6197 -47743 -6077 -47709
rect -6197 -47777 -6154 -47743
rect -6120 -47777 -6077 -47743
rect -6197 -47811 -6077 -47777
rect -6197 -47845 -6154 -47811
rect -6120 -47845 -6077 -47811
rect -6197 -47879 -6077 -47845
rect -6197 -47913 -6154 -47879
rect -6120 -47913 -6077 -47879
rect -6197 -47947 -6077 -47913
rect -6197 -47981 -6154 -47947
rect -6120 -47981 -6077 -47947
rect -6197 -48015 -6077 -47981
rect -6197 -48049 -6154 -48015
rect -6120 -48049 -6077 -48015
rect -6197 -48083 -6077 -48049
rect -6197 -48117 -6154 -48083
rect -6120 -48117 -6077 -48083
rect -6197 -48176 -6077 -48117
rect -6047 -47234 -5927 -47176
rect -6047 -47268 -6004 -47234
rect -5970 -47268 -5927 -47234
rect -6047 -47335 -5927 -47268
rect -6047 -47369 -6004 -47335
rect -5970 -47369 -5927 -47335
rect -6047 -47403 -5927 -47369
rect -6047 -47437 -6004 -47403
rect -5970 -47437 -5927 -47403
rect -6047 -47471 -5927 -47437
rect -6047 -47505 -6004 -47471
rect -5970 -47505 -5927 -47471
rect -6047 -47539 -5927 -47505
rect -6047 -47573 -6004 -47539
rect -5970 -47573 -5927 -47539
rect -6047 -47607 -5927 -47573
rect -6047 -47641 -6004 -47607
rect -5970 -47641 -5927 -47607
rect -6047 -47675 -5927 -47641
rect -6047 -47709 -6004 -47675
rect -5970 -47709 -5927 -47675
rect -6047 -47743 -5927 -47709
rect -6047 -47777 -6004 -47743
rect -5970 -47777 -5927 -47743
rect -6047 -47811 -5927 -47777
rect -6047 -47845 -6004 -47811
rect -5970 -47845 -5927 -47811
rect -6047 -47879 -5927 -47845
rect -6047 -47913 -6004 -47879
rect -5970 -47913 -5927 -47879
rect -6047 -47947 -5927 -47913
rect -6047 -47981 -6004 -47947
rect -5970 -47981 -5927 -47947
rect -6047 -48015 -5927 -47981
rect -6047 -48049 -6004 -48015
rect -5970 -48049 -5927 -48015
rect -6047 -48083 -5927 -48049
rect -6047 -48117 -6004 -48083
rect -5970 -48117 -5927 -48083
rect -6047 -48176 -5927 -48117
rect -5897 -47234 -5777 -47176
rect -5897 -47268 -5854 -47234
rect -5820 -47268 -5777 -47234
rect -5897 -47335 -5777 -47268
rect -5897 -47369 -5854 -47335
rect -5820 -47369 -5777 -47335
rect -5897 -47403 -5777 -47369
rect -5897 -47437 -5854 -47403
rect -5820 -47437 -5777 -47403
rect -5897 -47471 -5777 -47437
rect -5897 -47505 -5854 -47471
rect -5820 -47505 -5777 -47471
rect -5897 -47539 -5777 -47505
rect -5897 -47573 -5854 -47539
rect -5820 -47573 -5777 -47539
rect -5897 -47607 -5777 -47573
rect -5897 -47641 -5854 -47607
rect -5820 -47641 -5777 -47607
rect -5897 -47675 -5777 -47641
rect -5897 -47709 -5854 -47675
rect -5820 -47709 -5777 -47675
rect -5897 -47743 -5777 -47709
rect -5897 -47777 -5854 -47743
rect -5820 -47777 -5777 -47743
rect -5897 -47811 -5777 -47777
rect -5897 -47845 -5854 -47811
rect -5820 -47845 -5777 -47811
rect -5897 -47879 -5777 -47845
rect -5897 -47913 -5854 -47879
rect -5820 -47913 -5777 -47879
rect -5897 -47947 -5777 -47913
rect -5897 -47981 -5854 -47947
rect -5820 -47981 -5777 -47947
rect -5897 -48015 -5777 -47981
rect -5897 -48049 -5854 -48015
rect -5820 -48049 -5777 -48015
rect -5897 -48083 -5777 -48049
rect -5897 -48117 -5854 -48083
rect -5820 -48117 -5777 -48083
rect -5897 -48176 -5777 -48117
rect -5747 -47234 -5627 -47176
rect -5747 -47268 -5704 -47234
rect -5670 -47268 -5627 -47234
rect -5747 -47345 -5627 -47268
rect -5747 -47379 -5704 -47345
rect -5670 -47379 -5627 -47345
rect -5747 -47413 -5627 -47379
rect -5747 -47447 -5704 -47413
rect -5670 -47447 -5627 -47413
rect -5747 -47481 -5627 -47447
rect -5747 -47515 -5704 -47481
rect -5670 -47515 -5627 -47481
rect -5747 -47549 -5627 -47515
rect -5747 -47583 -5704 -47549
rect -5670 -47583 -5627 -47549
rect -5747 -47617 -5627 -47583
rect -5747 -47651 -5704 -47617
rect -5670 -47651 -5627 -47617
rect -5747 -47685 -5627 -47651
rect -5747 -47719 -5704 -47685
rect -5670 -47719 -5627 -47685
rect -5747 -47753 -5627 -47719
rect -5747 -47787 -5704 -47753
rect -5670 -47787 -5627 -47753
rect -5747 -47821 -5627 -47787
rect -5747 -47855 -5704 -47821
rect -5670 -47855 -5627 -47821
rect -5747 -47889 -5627 -47855
rect -5747 -47923 -5704 -47889
rect -5670 -47923 -5627 -47889
rect -5747 -47957 -5627 -47923
rect -5747 -47991 -5704 -47957
rect -5670 -47991 -5627 -47957
rect -5747 -48025 -5627 -47991
rect -5747 -48059 -5704 -48025
rect -5670 -48059 -5627 -48025
rect -5747 -48093 -5627 -48059
rect -5747 -48127 -5704 -48093
rect -5670 -48127 -5627 -48093
rect -5747 -48176 -5627 -48127
rect -5597 -47234 -5477 -47176
rect -5597 -47268 -5554 -47234
rect -5520 -47268 -5477 -47234
rect -5597 -47335 -5477 -47268
rect -5597 -47369 -5554 -47335
rect -5520 -47369 -5477 -47335
rect -5597 -47403 -5477 -47369
rect -5597 -47437 -5554 -47403
rect -5520 -47437 -5477 -47403
rect -5597 -47471 -5477 -47437
rect -5597 -47505 -5554 -47471
rect -5520 -47505 -5477 -47471
rect -5597 -47539 -5477 -47505
rect -5597 -47573 -5554 -47539
rect -5520 -47573 -5477 -47539
rect -5597 -47607 -5477 -47573
rect -5597 -47641 -5554 -47607
rect -5520 -47641 -5477 -47607
rect -5597 -47675 -5477 -47641
rect -5597 -47709 -5554 -47675
rect -5520 -47709 -5477 -47675
rect -5597 -47743 -5477 -47709
rect -5597 -47777 -5554 -47743
rect -5520 -47777 -5477 -47743
rect -5597 -47811 -5477 -47777
rect -5597 -47845 -5554 -47811
rect -5520 -47845 -5477 -47811
rect -5597 -47879 -5477 -47845
rect -5597 -47913 -5554 -47879
rect -5520 -47913 -5477 -47879
rect -5597 -47947 -5477 -47913
rect -5597 -47981 -5554 -47947
rect -5520 -47981 -5477 -47947
rect -5597 -48015 -5477 -47981
rect -5597 -48049 -5554 -48015
rect -5520 -48049 -5477 -48015
rect -5597 -48083 -5477 -48049
rect -5597 -48117 -5554 -48083
rect -5520 -48117 -5477 -48083
rect -5597 -48176 -5477 -48117
rect -5447 -47234 -5327 -47176
rect -5447 -47268 -5404 -47234
rect -5370 -47268 -5327 -47234
rect -5447 -47335 -5327 -47268
rect -5447 -47369 -5404 -47335
rect -5370 -47369 -5327 -47335
rect -5447 -47403 -5327 -47369
rect -5447 -47437 -5404 -47403
rect -5370 -47437 -5327 -47403
rect -5447 -47471 -5327 -47437
rect -5447 -47505 -5404 -47471
rect -5370 -47505 -5327 -47471
rect -5447 -47539 -5327 -47505
rect -5447 -47573 -5404 -47539
rect -5370 -47573 -5327 -47539
rect -5447 -47607 -5327 -47573
rect -5447 -47641 -5404 -47607
rect -5370 -47641 -5327 -47607
rect -5447 -47675 -5327 -47641
rect -5447 -47709 -5404 -47675
rect -5370 -47709 -5327 -47675
rect -5447 -47743 -5327 -47709
rect -5447 -47777 -5404 -47743
rect -5370 -47777 -5327 -47743
rect -5447 -47811 -5327 -47777
rect -5447 -47845 -5404 -47811
rect -5370 -47845 -5327 -47811
rect -5447 -47879 -5327 -47845
rect -5447 -47913 -5404 -47879
rect -5370 -47913 -5327 -47879
rect -5447 -47947 -5327 -47913
rect -5447 -47981 -5404 -47947
rect -5370 -47981 -5327 -47947
rect -5447 -48015 -5327 -47981
rect -5447 -48049 -5404 -48015
rect -5370 -48049 -5327 -48015
rect -5447 -48083 -5327 -48049
rect -5447 -48117 -5404 -48083
rect -5370 -48117 -5327 -48083
rect -5447 -48176 -5327 -48117
rect -5297 -47234 -5177 -47176
rect -5297 -47268 -5254 -47234
rect -5220 -47268 -5177 -47234
rect -5297 -47335 -5177 -47268
rect -5297 -47369 -5254 -47335
rect -5220 -47369 -5177 -47335
rect -5297 -47403 -5177 -47369
rect -5297 -47437 -5254 -47403
rect -5220 -47437 -5177 -47403
rect -5297 -47471 -5177 -47437
rect -5297 -47505 -5254 -47471
rect -5220 -47505 -5177 -47471
rect -5297 -47539 -5177 -47505
rect -5297 -47573 -5254 -47539
rect -5220 -47573 -5177 -47539
rect -5297 -47607 -5177 -47573
rect -5297 -47641 -5254 -47607
rect -5220 -47641 -5177 -47607
rect -5297 -47675 -5177 -47641
rect -5297 -47709 -5254 -47675
rect -5220 -47709 -5177 -47675
rect -5297 -47743 -5177 -47709
rect -5297 -47777 -5254 -47743
rect -5220 -47777 -5177 -47743
rect -5297 -47811 -5177 -47777
rect -5297 -47845 -5254 -47811
rect -5220 -47845 -5177 -47811
rect -5297 -47879 -5177 -47845
rect -5297 -47913 -5254 -47879
rect -5220 -47913 -5177 -47879
rect -5297 -47947 -5177 -47913
rect -5297 -47981 -5254 -47947
rect -5220 -47981 -5177 -47947
rect -5297 -48015 -5177 -47981
rect -5297 -48049 -5254 -48015
rect -5220 -48049 -5177 -48015
rect -5297 -48083 -5177 -48049
rect -5297 -48117 -5254 -48083
rect -5220 -48117 -5177 -48083
rect -5297 -48176 -5177 -48117
<< ndiffc >>
rect -9485 -44084 -9451 -44050
rect -9485 -44152 -9451 -44118
rect -9485 -44220 -9451 -44186
rect -9485 -44288 -9451 -44254
rect -9485 -44356 -9451 -44322
rect -9485 -44424 -9451 -44390
rect -9485 -44492 -9451 -44458
rect -9485 -44560 -9451 -44526
rect -9485 -44628 -9451 -44594
rect -9485 -44696 -9451 -44662
rect -9485 -44764 -9451 -44730
rect -9485 -44832 -9451 -44798
rect -9335 -44084 -9301 -44050
rect -9335 -44152 -9301 -44118
rect -9335 -44220 -9301 -44186
rect -9335 -44288 -9301 -44254
rect -9335 -44356 -9301 -44322
rect -9335 -44424 -9301 -44390
rect -9335 -44492 -9301 -44458
rect -9335 -44560 -9301 -44526
rect -9335 -44628 -9301 -44594
rect -9335 -44696 -9301 -44662
rect -9335 -44764 -9301 -44730
rect -9335 -44832 -9301 -44798
rect -9185 -44084 -9151 -44050
rect -9185 -44152 -9151 -44118
rect -9185 -44220 -9151 -44186
rect -9185 -44288 -9151 -44254
rect -9185 -44356 -9151 -44322
rect -9185 -44424 -9151 -44390
rect -9185 -44492 -9151 -44458
rect -9185 -44560 -9151 -44526
rect -9185 -44628 -9151 -44594
rect -9185 -44696 -9151 -44662
rect -9185 -44764 -9151 -44730
rect -9185 -44832 -9151 -44798
rect -9035 -44084 -9001 -44050
rect -9035 -44152 -9001 -44118
rect -9035 -44220 -9001 -44186
rect -9035 -44288 -9001 -44254
rect -9035 -44356 -9001 -44322
rect -9035 -44424 -9001 -44390
rect -9035 -44492 -9001 -44458
rect -9035 -44560 -9001 -44526
rect -9035 -44628 -9001 -44594
rect -9035 -44696 -9001 -44662
rect -9035 -44764 -9001 -44730
rect -9035 -44832 -9001 -44798
rect -8885 -44084 -8851 -44050
rect -8885 -44152 -8851 -44118
rect -8885 -44220 -8851 -44186
rect -8885 -44288 -8851 -44254
rect -8885 -44356 -8851 -44322
rect -8885 -44424 -8851 -44390
rect -8885 -44492 -8851 -44458
rect -8885 -44560 -8851 -44526
rect -8885 -44628 -8851 -44594
rect -8885 -44696 -8851 -44662
rect -8885 -44764 -8851 -44730
rect -8885 -44832 -8851 -44798
rect -8735 -44084 -8701 -44050
rect -8735 -44152 -8701 -44118
rect -8735 -44220 -8701 -44186
rect -8735 -44288 -8701 -44254
rect -8735 -44356 -8701 -44322
rect -8735 -44424 -8701 -44390
rect -8735 -44492 -8701 -44458
rect -8735 -44560 -8701 -44526
rect -8735 -44628 -8701 -44594
rect -8735 -44696 -8701 -44662
rect -8735 -44764 -8701 -44730
rect -8735 -44832 -8701 -44798
rect -8585 -44084 -8551 -44050
rect -8585 -44152 -8551 -44118
rect -8585 -44220 -8551 -44186
rect -8585 -44288 -8551 -44254
rect -8585 -44356 -8551 -44322
rect -8585 -44424 -8551 -44390
rect -8585 -44492 -8551 -44458
rect -8585 -44560 -8551 -44526
rect -8585 -44628 -8551 -44594
rect -8585 -44696 -8551 -44662
rect -8585 -44764 -8551 -44730
rect -8585 -44832 -8551 -44798
rect -8435 -44084 -8401 -44050
rect -8435 -44152 -8401 -44118
rect -8435 -44220 -8401 -44186
rect -8435 -44288 -8401 -44254
rect -8435 -44356 -8401 -44322
rect -8435 -44424 -8401 -44390
rect -8435 -44492 -8401 -44458
rect -8435 -44560 -8401 -44526
rect -8435 -44628 -8401 -44594
rect -8435 -44696 -8401 -44662
rect -8435 -44764 -8401 -44730
rect -8435 -44832 -8401 -44798
rect -8285 -44084 -8251 -44050
rect -8285 -44152 -8251 -44118
rect -8285 -44220 -8251 -44186
rect -8285 -44288 -8251 -44254
rect -8285 -44356 -8251 -44322
rect -8285 -44424 -8251 -44390
rect -8285 -44492 -8251 -44458
rect -8285 -44560 -8251 -44526
rect -8285 -44628 -8251 -44594
rect -8285 -44696 -8251 -44662
rect -8285 -44764 -8251 -44730
rect -8285 -44832 -8251 -44798
rect -8135 -44094 -8101 -44060
rect -8135 -44162 -8101 -44128
rect -8135 -44230 -8101 -44196
rect -8135 -44298 -8101 -44264
rect -8135 -44366 -8101 -44332
rect -8135 -44434 -8101 -44400
rect -8135 -44502 -8101 -44468
rect -8135 -44570 -8101 -44536
rect -8135 -44638 -8101 -44604
rect -8135 -44706 -8101 -44672
rect -8135 -44774 -8101 -44740
rect -8135 -44842 -8101 -44808
rect -7985 -44084 -7951 -44050
rect -7985 -44152 -7951 -44118
rect -7985 -44220 -7951 -44186
rect -7985 -44288 -7951 -44254
rect -7985 -44356 -7951 -44322
rect -7985 -44424 -7951 -44390
rect -7985 -44492 -7951 -44458
rect -7985 -44560 -7951 -44526
rect -7985 -44628 -7951 -44594
rect -7985 -44696 -7951 -44662
rect -7985 -44764 -7951 -44730
rect -7985 -44832 -7951 -44798
rect -7835 -44084 -7801 -44050
rect -7835 -44152 -7801 -44118
rect -7835 -44220 -7801 -44186
rect -7835 -44288 -7801 -44254
rect -7835 -44356 -7801 -44322
rect -7835 -44424 -7801 -44390
rect -7835 -44492 -7801 -44458
rect -7835 -44560 -7801 -44526
rect -7835 -44628 -7801 -44594
rect -7835 -44696 -7801 -44662
rect -7835 -44764 -7801 -44730
rect -7835 -44832 -7801 -44798
rect -7685 -44084 -7651 -44050
rect -7685 -44152 -7651 -44118
rect -7685 -44220 -7651 -44186
rect -7685 -44288 -7651 -44254
rect -7685 -44356 -7651 -44322
rect -7685 -44424 -7651 -44390
rect -7685 -44492 -7651 -44458
rect -7685 -44560 -7651 -44526
rect -7685 -44628 -7651 -44594
rect -7685 -44696 -7651 -44662
rect -7685 -44764 -7651 -44730
rect -7685 -44832 -7651 -44798
rect -7535 -44084 -7501 -44050
rect -7535 -44152 -7501 -44118
rect -7535 -44220 -7501 -44186
rect -7535 -44288 -7501 -44254
rect -7535 -44356 -7501 -44322
rect -7535 -44424 -7501 -44390
rect -7535 -44492 -7501 -44458
rect -7535 -44560 -7501 -44526
rect -7535 -44628 -7501 -44594
rect -7535 -44696 -7501 -44662
rect -7535 -44764 -7501 -44730
rect -7535 -44832 -7501 -44798
rect -7385 -44084 -7351 -44050
rect -7385 -44152 -7351 -44118
rect -7385 -44220 -7351 -44186
rect -7385 -44288 -7351 -44254
rect -7385 -44356 -7351 -44322
rect -7385 -44424 -7351 -44390
rect -7385 -44492 -7351 -44458
rect -7385 -44560 -7351 -44526
rect -7385 -44628 -7351 -44594
rect -7385 -44696 -7351 -44662
rect -7385 -44764 -7351 -44730
rect -7385 -44832 -7351 -44798
rect -7235 -44084 -7201 -44050
rect -7235 -44152 -7201 -44118
rect -7235 -44220 -7201 -44186
rect -7235 -44288 -7201 -44254
rect -7235 -44356 -7201 -44322
rect -7235 -44424 -7201 -44390
rect -7235 -44492 -7201 -44458
rect -7235 -44560 -7201 -44526
rect -7235 -44628 -7201 -44594
rect -7235 -44696 -7201 -44662
rect -7235 -44764 -7201 -44730
rect -7235 -44832 -7201 -44798
rect -7085 -44084 -7051 -44050
rect -7085 -44152 -7051 -44118
rect -7085 -44220 -7051 -44186
rect -7085 -44288 -7051 -44254
rect -7085 -44356 -7051 -44322
rect -7085 -44424 -7051 -44390
rect -7085 -44492 -7051 -44458
rect -7085 -44560 -7051 -44526
rect -7085 -44628 -7051 -44594
rect -7085 -44696 -7051 -44662
rect -7085 -44764 -7051 -44730
rect -7085 -44832 -7051 -44798
rect -6935 -44084 -6901 -44050
rect -6935 -44152 -6901 -44118
rect -6935 -44220 -6901 -44186
rect -6935 -44288 -6901 -44254
rect -6935 -44356 -6901 -44322
rect -6935 -44424 -6901 -44390
rect -6935 -44492 -6901 -44458
rect -6935 -44560 -6901 -44526
rect -6935 -44628 -6901 -44594
rect -6935 -44696 -6901 -44662
rect -6935 -44764 -6901 -44730
rect -6935 -44832 -6901 -44798
rect -6785 -44084 -6751 -44050
rect -6785 -44152 -6751 -44118
rect -6785 -44220 -6751 -44186
rect -6785 -44288 -6751 -44254
rect -6785 -44356 -6751 -44322
rect -6785 -44424 -6751 -44390
rect -6785 -44492 -6751 -44458
rect -6785 -44560 -6751 -44526
rect -6785 -44628 -6751 -44594
rect -6785 -44696 -6751 -44662
rect -6785 -44764 -6751 -44730
rect -6785 -44832 -6751 -44798
rect -6635 -44094 -6601 -44060
rect -6635 -44162 -6601 -44128
rect -6635 -44230 -6601 -44196
rect -6635 -44298 -6601 -44264
rect -6635 -44366 -6601 -44332
rect -6635 -44434 -6601 -44400
rect -6635 -44502 -6601 -44468
rect -6635 -44570 -6601 -44536
rect -6635 -44638 -6601 -44604
rect -6635 -44706 -6601 -44672
rect -6635 -44774 -6601 -44740
rect -6635 -44842 -6601 -44808
rect -6485 -44084 -6451 -44050
rect -6485 -44152 -6451 -44118
rect -6485 -44220 -6451 -44186
rect -6485 -44288 -6451 -44254
rect -6485 -44356 -6451 -44322
rect -6485 -44424 -6451 -44390
rect -6485 -44492 -6451 -44458
rect -6485 -44560 -6451 -44526
rect -6485 -44628 -6451 -44594
rect -6485 -44696 -6451 -44662
rect -6485 -44764 -6451 -44730
rect -6485 -44832 -6451 -44798
rect -5379 -44084 -5345 -44050
rect -5379 -44152 -5345 -44118
rect -5379 -44220 -5345 -44186
rect -5379 -44288 -5345 -44254
rect -5379 -44356 -5345 -44322
rect -5379 -44424 -5345 -44390
rect -5379 -44492 -5345 -44458
rect -5379 -44560 -5345 -44526
rect -5379 -44628 -5345 -44594
rect -5379 -44696 -5345 -44662
rect -5379 -44764 -5345 -44730
rect -5379 -44832 -5345 -44798
rect -5229 -44094 -5195 -44060
rect -5229 -44162 -5195 -44128
rect -5229 -44230 -5195 -44196
rect -5229 -44298 -5195 -44264
rect -5229 -44366 -5195 -44332
rect -5229 -44434 -5195 -44400
rect -5229 -44502 -5195 -44468
rect -5229 -44570 -5195 -44536
rect -5229 -44638 -5195 -44604
rect -5229 -44706 -5195 -44672
rect -5229 -44774 -5195 -44740
rect -5229 -44842 -5195 -44808
rect -5079 -44084 -5045 -44050
rect -5079 -44152 -5045 -44118
rect -5079 -44220 -5045 -44186
rect -5079 -44288 -5045 -44254
rect -5079 -44356 -5045 -44322
rect -5079 -44424 -5045 -44390
rect -5079 -44492 -5045 -44458
rect -5079 -44560 -5045 -44526
rect -5079 -44628 -5045 -44594
rect -5079 -44696 -5045 -44662
rect -5079 -44764 -5045 -44730
rect -5079 -44832 -5045 -44798
rect -4929 -44084 -4895 -44050
rect -4929 -44152 -4895 -44118
rect -4929 -44220 -4895 -44186
rect -4929 -44288 -4895 -44254
rect -4929 -44356 -4895 -44322
rect -4929 -44424 -4895 -44390
rect -4929 -44492 -4895 -44458
rect -4929 -44560 -4895 -44526
rect -4929 -44628 -4895 -44594
rect -4929 -44696 -4895 -44662
rect -4929 -44764 -4895 -44730
rect -4929 -44832 -4895 -44798
rect -4779 -44084 -4745 -44050
rect -4779 -44152 -4745 -44118
rect -4779 -44220 -4745 -44186
rect -4779 -44288 -4745 -44254
rect -4779 -44356 -4745 -44322
rect -4779 -44424 -4745 -44390
rect -4779 -44492 -4745 -44458
rect -4779 -44560 -4745 -44526
rect -4779 -44628 -4745 -44594
rect -4779 -44696 -4745 -44662
rect -4779 -44764 -4745 -44730
rect -4779 -44832 -4745 -44798
rect -4629 -44084 -4595 -44050
rect -4629 -44152 -4595 -44118
rect -4629 -44220 -4595 -44186
rect -4629 -44288 -4595 -44254
rect -4629 -44356 -4595 -44322
rect -4629 -44424 -4595 -44390
rect -4629 -44492 -4595 -44458
rect -4629 -44560 -4595 -44526
rect -4629 -44628 -4595 -44594
rect -4629 -44696 -4595 -44662
rect -4629 -44764 -4595 -44730
rect -4629 -44832 -4595 -44798
rect -4479 -44084 -4445 -44050
rect -4479 -44152 -4445 -44118
rect -4479 -44220 -4445 -44186
rect -4479 -44288 -4445 -44254
rect -4479 -44356 -4445 -44322
rect -4479 -44424 -4445 -44390
rect -4479 -44492 -4445 -44458
rect -4479 -44560 -4445 -44526
rect -4479 -44628 -4445 -44594
rect -4479 -44696 -4445 -44662
rect -4479 -44764 -4445 -44730
rect -4479 -44832 -4445 -44798
rect -4329 -44084 -4295 -44050
rect -4329 -44152 -4295 -44118
rect -4329 -44220 -4295 -44186
rect -4329 -44288 -4295 -44254
rect -4329 -44356 -4295 -44322
rect -4329 -44424 -4295 -44390
rect -4329 -44492 -4295 -44458
rect -4329 -44560 -4295 -44526
rect -4329 -44628 -4295 -44594
rect -4329 -44696 -4295 -44662
rect -4329 -44764 -4295 -44730
rect -4329 -44832 -4295 -44798
rect -4179 -44084 -4145 -44050
rect -4179 -44152 -4145 -44118
rect -4179 -44220 -4145 -44186
rect -4179 -44288 -4145 -44254
rect -4179 -44356 -4145 -44322
rect -4179 -44424 -4145 -44390
rect -4179 -44492 -4145 -44458
rect -4179 -44560 -4145 -44526
rect -4179 -44628 -4145 -44594
rect -4179 -44696 -4145 -44662
rect -4179 -44764 -4145 -44730
rect -4179 -44832 -4145 -44798
rect -4029 -44084 -3995 -44050
rect -4029 -44152 -3995 -44118
rect -4029 -44220 -3995 -44186
rect -4029 -44288 -3995 -44254
rect -4029 -44356 -3995 -44322
rect -4029 -44424 -3995 -44390
rect -4029 -44492 -3995 -44458
rect -4029 -44560 -3995 -44526
rect -4029 -44628 -3995 -44594
rect -4029 -44696 -3995 -44662
rect -4029 -44764 -3995 -44730
rect -4029 -44832 -3995 -44798
rect -3879 -44084 -3845 -44050
rect -3879 -44152 -3845 -44118
rect -3879 -44220 -3845 -44186
rect -3879 -44288 -3845 -44254
rect -3879 -44356 -3845 -44322
rect -3879 -44424 -3845 -44390
rect -3879 -44492 -3845 -44458
rect -3879 -44560 -3845 -44526
rect -3879 -44628 -3845 -44594
rect -3879 -44696 -3845 -44662
rect -3879 -44764 -3845 -44730
rect -3879 -44832 -3845 -44798
rect -3729 -44094 -3695 -44060
rect -3729 -44162 -3695 -44128
rect -3729 -44230 -3695 -44196
rect -3729 -44298 -3695 -44264
rect -3729 -44366 -3695 -44332
rect -3729 -44434 -3695 -44400
rect -3729 -44502 -3695 -44468
rect -3729 -44570 -3695 -44536
rect -3729 -44638 -3695 -44604
rect -3729 -44706 -3695 -44672
rect -3729 -44774 -3695 -44740
rect -3729 -44842 -3695 -44808
rect -3579 -44084 -3545 -44050
rect -3579 -44152 -3545 -44118
rect -3579 -44220 -3545 -44186
rect -3579 -44288 -3545 -44254
rect -3579 -44356 -3545 -44322
rect -3579 -44424 -3545 -44390
rect -3579 -44492 -3545 -44458
rect -3579 -44560 -3545 -44526
rect -3579 -44628 -3545 -44594
rect -3579 -44696 -3545 -44662
rect -3579 -44764 -3545 -44730
rect -3579 -44832 -3545 -44798
rect -3429 -44084 -3395 -44050
rect -3429 -44152 -3395 -44118
rect -3429 -44220 -3395 -44186
rect -3429 -44288 -3395 -44254
rect -3429 -44356 -3395 -44322
rect -3429 -44424 -3395 -44390
rect -3429 -44492 -3395 -44458
rect -3429 -44560 -3395 -44526
rect -3429 -44628 -3395 -44594
rect -3429 -44696 -3395 -44662
rect -3429 -44764 -3395 -44730
rect -3429 -44832 -3395 -44798
rect -3279 -44084 -3245 -44050
rect -3279 -44152 -3245 -44118
rect -3279 -44220 -3245 -44186
rect -3279 -44288 -3245 -44254
rect -3279 -44356 -3245 -44322
rect -3279 -44424 -3245 -44390
rect -3279 -44492 -3245 -44458
rect -3279 -44560 -3245 -44526
rect -3279 -44628 -3245 -44594
rect -3279 -44696 -3245 -44662
rect -3279 -44764 -3245 -44730
rect -3279 -44832 -3245 -44798
rect -3129 -44084 -3095 -44050
rect -3129 -44152 -3095 -44118
rect -3129 -44220 -3095 -44186
rect -3129 -44288 -3095 -44254
rect -3129 -44356 -3095 -44322
rect -3129 -44424 -3095 -44390
rect -3129 -44492 -3095 -44458
rect -3129 -44560 -3095 -44526
rect -3129 -44628 -3095 -44594
rect -3129 -44696 -3095 -44662
rect -3129 -44764 -3095 -44730
rect -3129 -44832 -3095 -44798
rect -2979 -44084 -2945 -44050
rect -2979 -44152 -2945 -44118
rect -2979 -44220 -2945 -44186
rect -2979 -44288 -2945 -44254
rect -2979 -44356 -2945 -44322
rect -2979 -44424 -2945 -44390
rect -2979 -44492 -2945 -44458
rect -2979 -44560 -2945 -44526
rect -2979 -44628 -2945 -44594
rect -2979 -44696 -2945 -44662
rect -2979 -44764 -2945 -44730
rect -2979 -44832 -2945 -44798
rect -2829 -44084 -2795 -44050
rect -2829 -44152 -2795 -44118
rect -2829 -44220 -2795 -44186
rect -2829 -44288 -2795 -44254
rect -2829 -44356 -2795 -44322
rect -2829 -44424 -2795 -44390
rect -2829 -44492 -2795 -44458
rect -2829 -44560 -2795 -44526
rect -2829 -44628 -2795 -44594
rect -2829 -44696 -2795 -44662
rect -2829 -44764 -2795 -44730
rect -2829 -44832 -2795 -44798
rect -2679 -44084 -2645 -44050
rect -2679 -44152 -2645 -44118
rect -2679 -44220 -2645 -44186
rect -2679 -44288 -2645 -44254
rect -2679 -44356 -2645 -44322
rect -2679 -44424 -2645 -44390
rect -2679 -44492 -2645 -44458
rect -2679 -44560 -2645 -44526
rect -2679 -44628 -2645 -44594
rect -2679 -44696 -2645 -44662
rect -2679 -44764 -2645 -44730
rect -2679 -44832 -2645 -44798
rect -2529 -44084 -2495 -44050
rect -2529 -44152 -2495 -44118
rect -2529 -44220 -2495 -44186
rect -2529 -44288 -2495 -44254
rect -2529 -44356 -2495 -44322
rect -2529 -44424 -2495 -44390
rect -2529 -44492 -2495 -44458
rect -2529 -44560 -2495 -44526
rect -2529 -44628 -2495 -44594
rect -2529 -44696 -2495 -44662
rect -2529 -44764 -2495 -44730
rect -2529 -44832 -2495 -44798
rect -2379 -44084 -2345 -44050
rect -2379 -44152 -2345 -44118
rect -2379 -44220 -2345 -44186
rect -2379 -44288 -2345 -44254
rect -2379 -44356 -2345 -44322
rect -2379 -44424 -2345 -44390
rect -2379 -44492 -2345 -44458
rect -2379 -44560 -2345 -44526
rect -2379 -44628 -2345 -44594
rect -2379 -44696 -2345 -44662
rect -2379 -44764 -2345 -44730
rect -2379 -44832 -2345 -44798
rect -6454 -47268 -6420 -47234
rect -6454 -47369 -6420 -47335
rect -6454 -47437 -6420 -47403
rect -6454 -47505 -6420 -47471
rect -6454 -47573 -6420 -47539
rect -6454 -47641 -6420 -47607
rect -6454 -47709 -6420 -47675
rect -6454 -47777 -6420 -47743
rect -6454 -47845 -6420 -47811
rect -6454 -47913 -6420 -47879
rect -6454 -47981 -6420 -47947
rect -6454 -48049 -6420 -48015
rect -6454 -48117 -6420 -48083
rect -6304 -47268 -6270 -47234
rect -6304 -47379 -6270 -47345
rect -6304 -47447 -6270 -47413
rect -6304 -47515 -6270 -47481
rect -6304 -47583 -6270 -47549
rect -6304 -47651 -6270 -47617
rect -6304 -47719 -6270 -47685
rect -6304 -47787 -6270 -47753
rect -6304 -47855 -6270 -47821
rect -6304 -47923 -6270 -47889
rect -6304 -47991 -6270 -47957
rect -6304 -48059 -6270 -48025
rect -6304 -48127 -6270 -48093
rect -6154 -47268 -6120 -47234
rect -6154 -47369 -6120 -47335
rect -6154 -47437 -6120 -47403
rect -6154 -47505 -6120 -47471
rect -6154 -47573 -6120 -47539
rect -6154 -47641 -6120 -47607
rect -6154 -47709 -6120 -47675
rect -6154 -47777 -6120 -47743
rect -6154 -47845 -6120 -47811
rect -6154 -47913 -6120 -47879
rect -6154 -47981 -6120 -47947
rect -6154 -48049 -6120 -48015
rect -6154 -48117 -6120 -48083
rect -6004 -47268 -5970 -47234
rect -6004 -47369 -5970 -47335
rect -6004 -47437 -5970 -47403
rect -6004 -47505 -5970 -47471
rect -6004 -47573 -5970 -47539
rect -6004 -47641 -5970 -47607
rect -6004 -47709 -5970 -47675
rect -6004 -47777 -5970 -47743
rect -6004 -47845 -5970 -47811
rect -6004 -47913 -5970 -47879
rect -6004 -47981 -5970 -47947
rect -6004 -48049 -5970 -48015
rect -6004 -48117 -5970 -48083
rect -5854 -47268 -5820 -47234
rect -5854 -47369 -5820 -47335
rect -5854 -47437 -5820 -47403
rect -5854 -47505 -5820 -47471
rect -5854 -47573 -5820 -47539
rect -5854 -47641 -5820 -47607
rect -5854 -47709 -5820 -47675
rect -5854 -47777 -5820 -47743
rect -5854 -47845 -5820 -47811
rect -5854 -47913 -5820 -47879
rect -5854 -47981 -5820 -47947
rect -5854 -48049 -5820 -48015
rect -5854 -48117 -5820 -48083
rect -5704 -47268 -5670 -47234
rect -5704 -47379 -5670 -47345
rect -5704 -47447 -5670 -47413
rect -5704 -47515 -5670 -47481
rect -5704 -47583 -5670 -47549
rect -5704 -47651 -5670 -47617
rect -5704 -47719 -5670 -47685
rect -5704 -47787 -5670 -47753
rect -5704 -47855 -5670 -47821
rect -5704 -47923 -5670 -47889
rect -5704 -47991 -5670 -47957
rect -5704 -48059 -5670 -48025
rect -5704 -48127 -5670 -48093
rect -5554 -47268 -5520 -47234
rect -5554 -47369 -5520 -47335
rect -5554 -47437 -5520 -47403
rect -5554 -47505 -5520 -47471
rect -5554 -47573 -5520 -47539
rect -5554 -47641 -5520 -47607
rect -5554 -47709 -5520 -47675
rect -5554 -47777 -5520 -47743
rect -5554 -47845 -5520 -47811
rect -5554 -47913 -5520 -47879
rect -5554 -47981 -5520 -47947
rect -5554 -48049 -5520 -48015
rect -5554 -48117 -5520 -48083
rect -5404 -47268 -5370 -47234
rect -5404 -47369 -5370 -47335
rect -5404 -47437 -5370 -47403
rect -5404 -47505 -5370 -47471
rect -5404 -47573 -5370 -47539
rect -5404 -47641 -5370 -47607
rect -5404 -47709 -5370 -47675
rect -5404 -47777 -5370 -47743
rect -5404 -47845 -5370 -47811
rect -5404 -47913 -5370 -47879
rect -5404 -47981 -5370 -47947
rect -5404 -48049 -5370 -48015
rect -5404 -48117 -5370 -48083
rect -5254 -47268 -5220 -47234
rect -5254 -47369 -5220 -47335
rect -5254 -47437 -5220 -47403
rect -5254 -47505 -5220 -47471
rect -5254 -47573 -5220 -47539
rect -5254 -47641 -5220 -47607
rect -5254 -47709 -5220 -47675
rect -5254 -47777 -5220 -47743
rect -5254 -47845 -5220 -47811
rect -5254 -47913 -5220 -47879
rect -5254 -47981 -5220 -47947
rect -5254 -48049 -5220 -48015
rect -5254 -48117 -5220 -48083
<< psubdiff >>
rect -9648 -44050 -9528 -43991
rect -9648 -44084 -9605 -44050
rect -9571 -44084 -9528 -44050
rect -9648 -44118 -9528 -44084
rect -9648 -44152 -9605 -44118
rect -9571 -44152 -9528 -44118
rect -9648 -44186 -9528 -44152
rect -9648 -44220 -9605 -44186
rect -9571 -44220 -9528 -44186
rect -9648 -44254 -9528 -44220
rect -9648 -44288 -9605 -44254
rect -9571 -44288 -9528 -44254
rect -9648 -44322 -9528 -44288
rect -9648 -44356 -9605 -44322
rect -9571 -44356 -9528 -44322
rect -9648 -44390 -9528 -44356
rect -9648 -44424 -9605 -44390
rect -9571 -44424 -9528 -44390
rect -9648 -44458 -9528 -44424
rect -9648 -44492 -9605 -44458
rect -9571 -44492 -9528 -44458
rect -9648 -44526 -9528 -44492
rect -9648 -44560 -9605 -44526
rect -9571 -44560 -9528 -44526
rect -9648 -44594 -9528 -44560
rect -9648 -44628 -9605 -44594
rect -9571 -44628 -9528 -44594
rect -9648 -44662 -9528 -44628
rect -9648 -44696 -9605 -44662
rect -9571 -44696 -9528 -44662
rect -9648 -44730 -9528 -44696
rect -9648 -44764 -9605 -44730
rect -9571 -44764 -9528 -44730
rect -9648 -44798 -9528 -44764
rect -9648 -44832 -9605 -44798
rect -9571 -44832 -9528 -44798
rect -9648 -44891 -9528 -44832
rect -6408 -44050 -6288 -43991
rect -6408 -44084 -6365 -44050
rect -6331 -44084 -6288 -44050
rect -6408 -44118 -6288 -44084
rect -6408 -44152 -6365 -44118
rect -6331 -44152 -6288 -44118
rect -6408 -44186 -6288 -44152
rect -6408 -44220 -6365 -44186
rect -6331 -44220 -6288 -44186
rect -6408 -44254 -6288 -44220
rect -6408 -44288 -6365 -44254
rect -6331 -44288 -6288 -44254
rect -6408 -44322 -6288 -44288
rect -6408 -44356 -6365 -44322
rect -6331 -44356 -6288 -44322
rect -6408 -44390 -6288 -44356
rect -6408 -44424 -6365 -44390
rect -6331 -44424 -6288 -44390
rect -6408 -44458 -6288 -44424
rect -6408 -44492 -6365 -44458
rect -6331 -44492 -6288 -44458
rect -6408 -44526 -6288 -44492
rect -6408 -44560 -6365 -44526
rect -6331 -44560 -6288 -44526
rect -6408 -44594 -6288 -44560
rect -6408 -44628 -6365 -44594
rect -6331 -44628 -6288 -44594
rect -6408 -44662 -6288 -44628
rect -6408 -44696 -6365 -44662
rect -6331 -44696 -6288 -44662
rect -6408 -44730 -6288 -44696
rect -6408 -44764 -6365 -44730
rect -6331 -44764 -6288 -44730
rect -6408 -44798 -6288 -44764
rect -6408 -44832 -6365 -44798
rect -6331 -44832 -6288 -44798
rect -6408 -44891 -6288 -44832
rect -5542 -44050 -5422 -43991
rect -5542 -44084 -5499 -44050
rect -5465 -44084 -5422 -44050
rect -5542 -44118 -5422 -44084
rect -5542 -44152 -5499 -44118
rect -5465 -44152 -5422 -44118
rect -5542 -44186 -5422 -44152
rect -5542 -44220 -5499 -44186
rect -5465 -44220 -5422 -44186
rect -5542 -44254 -5422 -44220
rect -5542 -44288 -5499 -44254
rect -5465 -44288 -5422 -44254
rect -5542 -44322 -5422 -44288
rect -5542 -44356 -5499 -44322
rect -5465 -44356 -5422 -44322
rect -5542 -44390 -5422 -44356
rect -5542 -44424 -5499 -44390
rect -5465 -44424 -5422 -44390
rect -5542 -44458 -5422 -44424
rect -5542 -44492 -5499 -44458
rect -5465 -44492 -5422 -44458
rect -5542 -44526 -5422 -44492
rect -5542 -44560 -5499 -44526
rect -5465 -44560 -5422 -44526
rect -5542 -44594 -5422 -44560
rect -5542 -44628 -5499 -44594
rect -5465 -44628 -5422 -44594
rect -5542 -44662 -5422 -44628
rect -5542 -44696 -5499 -44662
rect -5465 -44696 -5422 -44662
rect -5542 -44730 -5422 -44696
rect -5542 -44764 -5499 -44730
rect -5465 -44764 -5422 -44730
rect -5542 -44798 -5422 -44764
rect -5542 -44832 -5499 -44798
rect -5465 -44832 -5422 -44798
rect -5542 -44891 -5422 -44832
rect -2302 -44050 -2182 -43991
rect -2302 -44084 -2259 -44050
rect -2225 -44084 -2182 -44050
rect -2302 -44118 -2182 -44084
rect -2302 -44152 -2259 -44118
rect -2225 -44152 -2182 -44118
rect -2302 -44186 -2182 -44152
rect -2302 -44220 -2259 -44186
rect -2225 -44220 -2182 -44186
rect -2302 -44254 -2182 -44220
rect -2302 -44288 -2259 -44254
rect -2225 -44288 -2182 -44254
rect -2302 -44322 -2182 -44288
rect -2302 -44356 -2259 -44322
rect -2225 -44356 -2182 -44322
rect -2302 -44390 -2182 -44356
rect -2302 -44424 -2259 -44390
rect -2225 -44424 -2182 -44390
rect -2302 -44458 -2182 -44424
rect -2302 -44492 -2259 -44458
rect -2225 -44492 -2182 -44458
rect -2302 -44526 -2182 -44492
rect -2302 -44560 -2259 -44526
rect -2225 -44560 -2182 -44526
rect -2302 -44594 -2182 -44560
rect -2302 -44628 -2259 -44594
rect -2225 -44628 -2182 -44594
rect -2302 -44662 -2182 -44628
rect -2302 -44696 -2259 -44662
rect -2225 -44696 -2182 -44662
rect -2302 -44730 -2182 -44696
rect -2302 -44764 -2259 -44730
rect -2225 -44764 -2182 -44730
rect -2302 -44798 -2182 -44764
rect -2302 -44832 -2259 -44798
rect -2225 -44832 -2182 -44798
rect -2302 -44891 -2182 -44832
rect -6617 -47234 -6497 -47176
rect -6617 -47268 -6574 -47234
rect -6540 -47268 -6497 -47234
rect -6617 -47335 -6497 -47268
rect -6617 -47369 -6574 -47335
rect -6540 -47369 -6497 -47335
rect -6617 -47403 -6497 -47369
rect -6617 -47437 -6574 -47403
rect -6540 -47437 -6497 -47403
rect -6617 -47471 -6497 -47437
rect -6617 -47505 -6574 -47471
rect -6540 -47505 -6497 -47471
rect -6617 -47539 -6497 -47505
rect -6617 -47573 -6574 -47539
rect -6540 -47573 -6497 -47539
rect -6617 -47607 -6497 -47573
rect -6617 -47641 -6574 -47607
rect -6540 -47641 -6497 -47607
rect -6617 -47675 -6497 -47641
rect -6617 -47709 -6574 -47675
rect -6540 -47709 -6497 -47675
rect -6617 -47743 -6497 -47709
rect -6617 -47777 -6574 -47743
rect -6540 -47777 -6497 -47743
rect -6617 -47811 -6497 -47777
rect -6617 -47845 -6574 -47811
rect -6540 -47845 -6497 -47811
rect -6617 -47879 -6497 -47845
rect -6617 -47913 -6574 -47879
rect -6540 -47913 -6497 -47879
rect -6617 -47947 -6497 -47913
rect -6617 -47981 -6574 -47947
rect -6540 -47981 -6497 -47947
rect -6617 -48015 -6497 -47981
rect -6617 -48049 -6574 -48015
rect -6540 -48049 -6497 -48015
rect -6617 -48083 -6497 -48049
rect -6617 -48117 -6574 -48083
rect -6540 -48117 -6497 -48083
rect -6617 -48176 -6497 -48117
<< psubdiffcont >>
rect -9605 -44084 -9571 -44050
rect -9605 -44152 -9571 -44118
rect -9605 -44220 -9571 -44186
rect -9605 -44288 -9571 -44254
rect -9605 -44356 -9571 -44322
rect -9605 -44424 -9571 -44390
rect -9605 -44492 -9571 -44458
rect -9605 -44560 -9571 -44526
rect -9605 -44628 -9571 -44594
rect -9605 -44696 -9571 -44662
rect -9605 -44764 -9571 -44730
rect -9605 -44832 -9571 -44798
rect -6365 -44084 -6331 -44050
rect -6365 -44152 -6331 -44118
rect -6365 -44220 -6331 -44186
rect -6365 -44288 -6331 -44254
rect -6365 -44356 -6331 -44322
rect -6365 -44424 -6331 -44390
rect -6365 -44492 -6331 -44458
rect -6365 -44560 -6331 -44526
rect -6365 -44628 -6331 -44594
rect -6365 -44696 -6331 -44662
rect -6365 -44764 -6331 -44730
rect -6365 -44832 -6331 -44798
rect -5499 -44084 -5465 -44050
rect -5499 -44152 -5465 -44118
rect -5499 -44220 -5465 -44186
rect -5499 -44288 -5465 -44254
rect -5499 -44356 -5465 -44322
rect -5499 -44424 -5465 -44390
rect -5499 -44492 -5465 -44458
rect -5499 -44560 -5465 -44526
rect -5499 -44628 -5465 -44594
rect -5499 -44696 -5465 -44662
rect -5499 -44764 -5465 -44730
rect -5499 -44832 -5465 -44798
rect -2259 -44084 -2225 -44050
rect -2259 -44152 -2225 -44118
rect -2259 -44220 -2225 -44186
rect -2259 -44288 -2225 -44254
rect -2259 -44356 -2225 -44322
rect -2259 -44424 -2225 -44390
rect -2259 -44492 -2225 -44458
rect -2259 -44560 -2225 -44526
rect -2259 -44628 -2225 -44594
rect -2259 -44696 -2225 -44662
rect -2259 -44764 -2225 -44730
rect -2259 -44832 -2225 -44798
rect -6574 -47268 -6540 -47234
rect -6574 -47369 -6540 -47335
rect -6574 -47437 -6540 -47403
rect -6574 -47505 -6540 -47471
rect -6574 -47573 -6540 -47539
rect -6574 -47641 -6540 -47607
rect -6574 -47709 -6540 -47675
rect -6574 -47777 -6540 -47743
rect -6574 -47845 -6540 -47811
rect -6574 -47913 -6540 -47879
rect -6574 -47981 -6540 -47947
rect -6574 -48049 -6540 -48015
rect -6574 -48117 -6540 -48083
<< poly >>
rect -9420 -43842 -9354 -43826
rect -9420 -43876 -9404 -43842
rect -9370 -43876 -9354 -43842
rect -9420 -43892 -9354 -43876
rect -5320 -43829 -5254 -43813
rect -5320 -43863 -5304 -43829
rect -5270 -43863 -5254 -43829
rect -5320 -43879 -5254 -43863
rect -3814 -43842 -3748 -43826
rect -3814 -43876 -3798 -43842
rect -3764 -43876 -3748 -43842
rect -9408 -43911 -9354 -43892
rect -9408 -43941 -8028 -43911
rect -9408 -43991 -9378 -43941
rect -9258 -43991 -9228 -43941
rect -9108 -43991 -9078 -43941
rect -8958 -43991 -8928 -43941
rect -8808 -43991 -8778 -43941
rect -8658 -43991 -8628 -43941
rect -8508 -43991 -8478 -43941
rect -8358 -43991 -8328 -43941
rect -8208 -43991 -8178 -43941
rect -8058 -43991 -8028 -43941
rect -7908 -43991 -7878 -43941
rect -7758 -43991 -7728 -43941
rect -7608 -43991 -7578 -43941
rect -7458 -43991 -7428 -43941
rect -7308 -43991 -7278 -43941
rect -7158 -43991 -7128 -43941
rect -7008 -43991 -6978 -43941
rect -6858 -43991 -6828 -43941
rect -6708 -43991 -6678 -43941
rect -6558 -43991 -6528 -43941
rect -5302 -43991 -5272 -43879
rect -3814 -43892 -3748 -43876
rect -3802 -43911 -3748 -43892
rect -3802 -43941 -2422 -43911
rect -5152 -43991 -5122 -43941
rect -5002 -43991 -4972 -43941
rect -4852 -43991 -4822 -43941
rect -4702 -43991 -4672 -43941
rect -4552 -43991 -4522 -43941
rect -4402 -43991 -4372 -43941
rect -4252 -43991 -4222 -43941
rect -4102 -43991 -4072 -43941
rect -3952 -43991 -3922 -43941
rect -3802 -43991 -3772 -43941
rect -3652 -43991 -3622 -43941
rect -3502 -43991 -3472 -43941
rect -3352 -43991 -3322 -43941
rect -3202 -43991 -3172 -43941
rect -3052 -43991 -3022 -43941
rect -2902 -43991 -2872 -43941
rect -2752 -43991 -2722 -43941
rect -2602 -43991 -2572 -43941
rect -2452 -43991 -2422 -43941
rect -9408 -44921 -9378 -44891
rect -9258 -44921 -9228 -44891
rect -9108 -44921 -9078 -44891
rect -8958 -44921 -8928 -44891
rect -8808 -44921 -8778 -44891
rect -8658 -44921 -8628 -44891
rect -8508 -44921 -8478 -44891
rect -8358 -44921 -8328 -44891
rect -8208 -44921 -8178 -44891
rect -8058 -44921 -8028 -44891
rect -7908 -44942 -7878 -44891
rect -7758 -44942 -7728 -44891
rect -7608 -44942 -7578 -44891
rect -7458 -44942 -7428 -44891
rect -7308 -44942 -7278 -44891
rect -7158 -44942 -7128 -44891
rect -7008 -44942 -6978 -44891
rect -6858 -44942 -6828 -44891
rect -6708 -44942 -6678 -44891
rect -6558 -44942 -6528 -44891
rect -7908 -44972 -6528 -44942
rect -5302 -44942 -5272 -44891
rect -5152 -44942 -5122 -44891
rect -5002 -44942 -4972 -44891
rect -4852 -44942 -4822 -44891
rect -4702 -44942 -4672 -44891
rect -4552 -44942 -4522 -44891
rect -4402 -44942 -4372 -44891
rect -4252 -44942 -4222 -44891
rect -4102 -44942 -4072 -44891
rect -3952 -44942 -3922 -44891
rect -3802 -44921 -3772 -44891
rect -3652 -44921 -3622 -44891
rect -3502 -44921 -3472 -44891
rect -3352 -44921 -3322 -44891
rect -3202 -44921 -3172 -44891
rect -3052 -44921 -3022 -44891
rect -2902 -44921 -2872 -44891
rect -2752 -44921 -2722 -44891
rect -2602 -44921 -2572 -44891
rect -2452 -44921 -2422 -44891
rect -5302 -44972 -3922 -44942
rect -7908 -45043 -7878 -44972
rect -7926 -45059 -7860 -45043
rect -7926 -45093 -7910 -45059
rect -7876 -45093 -7860 -45059
rect -7926 -45109 -7860 -45093
rect -6360 -47096 -6290 -47080
rect -6377 -47130 -6342 -47096
rect -6307 -47126 -5297 -47096
rect -6307 -47130 -6290 -47126
rect -6377 -47150 -6290 -47130
rect -6377 -47176 -6347 -47150
rect -6227 -47176 -6197 -47126
rect -6077 -47176 -6047 -47126
rect -5927 -47176 -5897 -47126
rect -5777 -47176 -5747 -47126
rect -5627 -47176 -5597 -47126
rect -5477 -47176 -5447 -47126
rect -5327 -47176 -5297 -47126
rect -6805 -47798 -6717 -47782
rect -6805 -47832 -6778 -47798
rect -6744 -47832 -6717 -47798
rect -6805 -47855 -6717 -47832
rect -6805 -48216 -6717 -48193
rect -6805 -48250 -6778 -48216
rect -6744 -48236 -6717 -48216
rect -6377 -48236 -6347 -48176
rect -6227 -48206 -6197 -48176
rect -6077 -48206 -6047 -48176
rect -5927 -48206 -5897 -48176
rect -5777 -48206 -5747 -48176
rect -5627 -48206 -5597 -48176
rect -5477 -48206 -5447 -48176
rect -5327 -48206 -5297 -48176
rect -6744 -48250 -6347 -48236
rect -6805 -48266 -6347 -48250
<< polycont >>
rect -9404 -43876 -9370 -43842
rect -5304 -43863 -5270 -43829
rect -3798 -43876 -3764 -43842
rect -7910 -45093 -7876 -45059
rect -6342 -47130 -6307 -47096
rect -6778 -47832 -6744 -47798
rect -6778 -48250 -6744 -48216
<< xpolycontact >>
rect -7859 -43122 -7789 -42690
rect -7859 -43692 -7789 -43260
rect -7541 -43122 -7471 -42690
rect -7541 -43692 -7471 -43260
rect -7223 -43122 -7153 -42690
rect -7223 -43692 -7153 -43260
rect -6905 -43122 -6835 -42690
rect -6905 -43692 -6835 -43260
rect -2314 -43123 -2244 -42691
rect -2314 -43693 -2244 -43261
rect -1996 -43123 -1926 -42691
rect -1996 -43693 -1926 -43261
rect -1678 -43123 -1608 -42691
rect -1678 -43693 -1608 -43261
rect -1360 -43123 -1290 -42691
rect -1360 -43693 -1290 -43261
<< npolyres >>
rect -6805 -48193 -6717 -47855
<< xpolyres >>
rect -7859 -43260 -7789 -43122
rect -7541 -43260 -7471 -43122
rect -7223 -43260 -7153 -43122
rect -6905 -43260 -6835 -43122
rect -2314 -43261 -2244 -43123
rect -1996 -43261 -1926 -43123
rect -1678 -43261 -1608 -43123
rect -1360 -43261 -1290 -43123
<< locali >>
rect -44468 -34599 31781 -34576
rect -44468 -34633 -44422 -34599
rect -44388 -34633 -44342 -34599
rect -44308 -34633 -44262 -34599
rect -44228 -34633 -44182 -34599
rect -44148 -34633 -44102 -34599
rect -44068 -34633 -44022 -34599
rect -43988 -34633 -43942 -34599
rect -43908 -34633 -43862 -34599
rect -43828 -34633 -43782 -34599
rect -43748 -34633 -43702 -34599
rect -43668 -34633 -43622 -34599
rect -43588 -34633 -43542 -34599
rect -43508 -34633 -43462 -34599
rect -43428 -34633 -43382 -34599
rect -43348 -34633 -43302 -34599
rect -43268 -34633 -43222 -34599
rect -43188 -34633 -43142 -34599
rect -43108 -34633 -43062 -34599
rect -43028 -34633 -42982 -34599
rect -42948 -34633 -42902 -34599
rect -42868 -34633 -42822 -34599
rect -42788 -34633 -42742 -34599
rect -42708 -34633 -42662 -34599
rect -42628 -34633 -42582 -34599
rect -42548 -34633 -42502 -34599
rect -42468 -34633 -42422 -34599
rect -42388 -34633 -42342 -34599
rect -42308 -34633 -42262 -34599
rect -42228 -34633 -42182 -34599
rect -42148 -34633 -42102 -34599
rect -42068 -34633 -42022 -34599
rect -41988 -34633 -41942 -34599
rect -41908 -34633 -41862 -34599
rect -41828 -34633 -41782 -34599
rect -41748 -34633 -41702 -34599
rect -41668 -34633 -41622 -34599
rect -41588 -34633 -41542 -34599
rect -41508 -34633 -41462 -34599
rect -41428 -34633 -41382 -34599
rect -41348 -34633 -41302 -34599
rect -41268 -34633 -41222 -34599
rect -41188 -34633 -41142 -34599
rect -41108 -34633 -41062 -34599
rect -41028 -34633 -40982 -34599
rect -40948 -34633 -40902 -34599
rect -40868 -34633 -40822 -34599
rect -40788 -34633 -40742 -34599
rect -40708 -34633 -40662 -34599
rect -40628 -34633 -40582 -34599
rect -40548 -34633 -40502 -34599
rect -40468 -34633 -40422 -34599
rect -40388 -34633 -40342 -34599
rect -40308 -34633 -40262 -34599
rect -40228 -34633 -40182 -34599
rect -40148 -34633 -40102 -34599
rect -40068 -34633 -40022 -34599
rect -39988 -34633 -39942 -34599
rect -39908 -34633 -39862 -34599
rect -39828 -34633 -39782 -34599
rect -39748 -34633 -39702 -34599
rect -39668 -34633 -39622 -34599
rect -39588 -34633 -39542 -34599
rect -39508 -34633 -39462 -34599
rect -39428 -34633 -39382 -34599
rect -39348 -34633 -39302 -34599
rect -39268 -34633 -39222 -34599
rect -39188 -34633 -39142 -34599
rect -39108 -34633 -39062 -34599
rect -39028 -34633 -38982 -34599
rect -38948 -34633 -38902 -34599
rect -38868 -34633 -38822 -34599
rect -38788 -34633 -38742 -34599
rect -38708 -34633 -38662 -34599
rect -38628 -34633 -38582 -34599
rect -38548 -34633 -38502 -34599
rect -38468 -34633 -38422 -34599
rect -38388 -34633 -38342 -34599
rect -38308 -34633 -38262 -34599
rect -38228 -34633 -38182 -34599
rect -38148 -34633 -38102 -34599
rect -38068 -34633 -38022 -34599
rect -37988 -34633 -37942 -34599
rect -37908 -34633 -37862 -34599
rect -37828 -34633 -37782 -34599
rect -37748 -34633 -37702 -34599
rect -37668 -34633 -37622 -34599
rect -37588 -34633 -37542 -34599
rect -37508 -34633 -37462 -34599
rect -37428 -34633 -37382 -34599
rect -37348 -34633 -37302 -34599
rect -37268 -34633 -37222 -34599
rect -37188 -34633 -37142 -34599
rect -37108 -34633 -37062 -34599
rect -37028 -34633 -36982 -34599
rect -36948 -34633 -36902 -34599
rect -36868 -34633 -36822 -34599
rect -36788 -34633 -36742 -34599
rect -36708 -34633 -36662 -34599
rect -36628 -34633 -36582 -34599
rect -36548 -34633 -36502 -34599
rect -36468 -34633 -36422 -34599
rect -36388 -34633 -36342 -34599
rect -36308 -34633 -36262 -34599
rect -36228 -34633 -36182 -34599
rect -36148 -34633 -36102 -34599
rect -36068 -34633 -36022 -34599
rect -35988 -34633 -35942 -34599
rect -35908 -34633 -35862 -34599
rect -35828 -34633 -35782 -34599
rect -35748 -34633 -35702 -34599
rect -35668 -34633 -35622 -34599
rect -35588 -34633 -35542 -34599
rect -35508 -34633 -35462 -34599
rect -35428 -34633 -35382 -34599
rect -35348 -34633 -35302 -34599
rect -35268 -34633 -35222 -34599
rect -35188 -34633 -35142 -34599
rect -35108 -34633 -35062 -34599
rect -35028 -34633 -34982 -34599
rect -34948 -34633 -34902 -34599
rect -34868 -34633 -34822 -34599
rect -34788 -34633 -34742 -34599
rect -34708 -34633 -34662 -34599
rect -34628 -34633 -34582 -34599
rect -34548 -34633 -34502 -34599
rect -34468 -34633 -34422 -34599
rect -34388 -34633 -34342 -34599
rect -34308 -34633 -34262 -34599
rect -34228 -34633 -34182 -34599
rect -34148 -34633 -34102 -34599
rect -34068 -34633 -34022 -34599
rect -33988 -34633 -33942 -34599
rect -33908 -34633 -33862 -34599
rect -33828 -34633 -33782 -34599
rect -33748 -34633 -33702 -34599
rect -33668 -34633 -33622 -34599
rect -33588 -34633 -33542 -34599
rect -33508 -34633 -33462 -34599
rect -33428 -34633 -33382 -34599
rect -33348 -34633 -33302 -34599
rect -33268 -34633 -33222 -34599
rect -33188 -34633 -33142 -34599
rect -33108 -34633 -33062 -34599
rect -33028 -34633 -32982 -34599
rect -32948 -34633 -32902 -34599
rect -32868 -34633 -32822 -34599
rect -32788 -34633 -32742 -34599
rect -32708 -34633 -32662 -34599
rect -32628 -34633 -32582 -34599
rect -32548 -34633 -32502 -34599
rect -32468 -34633 -32422 -34599
rect -32388 -34633 -32342 -34599
rect -32308 -34633 -32262 -34599
rect -32228 -34633 -32182 -34599
rect -32148 -34633 -32102 -34599
rect -32068 -34633 -32022 -34599
rect -31988 -34633 -31942 -34599
rect -31908 -34633 -31862 -34599
rect -31828 -34633 -31782 -34599
rect -31748 -34633 -31702 -34599
rect -31668 -34633 -31622 -34599
rect -31588 -34633 -31542 -34599
rect -31508 -34633 -31461 -34599
rect -31427 -34633 -31381 -34599
rect -31347 -34633 -31301 -34599
rect -31267 -34633 -31221 -34599
rect -31187 -34633 -31141 -34599
rect -31107 -34633 -31061 -34599
rect -31027 -34633 -30981 -34599
rect -30947 -34633 -30901 -34599
rect -30867 -34633 -30821 -34599
rect -30787 -34633 -30741 -34599
rect -30707 -34633 -30661 -34599
rect -30627 -34633 -30581 -34599
rect -30547 -34633 -30501 -34599
rect -30467 -34633 -30421 -34599
rect -30387 -34633 -30341 -34599
rect -30307 -34633 -30261 -34599
rect -30227 -34633 -30181 -34599
rect -30147 -34633 -30101 -34599
rect -30067 -34633 -30021 -34599
rect -29987 -34633 -29941 -34599
rect -29907 -34633 -29861 -34599
rect -29827 -34633 -29781 -34599
rect -29747 -34633 -29701 -34599
rect -29667 -34633 -29621 -34599
rect -29587 -34633 -29541 -34599
rect -29507 -34633 -29461 -34599
rect -29427 -34633 -29381 -34599
rect -29347 -34633 -29301 -34599
rect -29267 -34633 -29221 -34599
rect -29187 -34633 -29141 -34599
rect -29107 -34633 -29061 -34599
rect -29027 -34633 -28981 -34599
rect -28947 -34633 -28901 -34599
rect -28867 -34633 -28821 -34599
rect -28787 -34633 -28741 -34599
rect -28707 -34633 -28661 -34599
rect -28627 -34633 -28581 -34599
rect -28547 -34633 -28501 -34599
rect -28467 -34633 -28421 -34599
rect -28387 -34633 -28341 -34599
rect -28307 -34633 -28261 -34599
rect -28227 -34633 -28181 -34599
rect -28147 -34633 -28101 -34599
rect -28067 -34633 -28021 -34599
rect -27987 -34633 -27941 -34599
rect -27907 -34633 -27861 -34599
rect -27827 -34633 -27781 -34599
rect -27747 -34633 -27701 -34599
rect -27667 -34633 -27621 -34599
rect -27587 -34633 -27541 -34599
rect -27507 -34633 -27461 -34599
rect -27427 -34633 -27381 -34599
rect -27347 -34633 -27301 -34599
rect -27267 -34633 -27221 -34599
rect -27187 -34633 -27141 -34599
rect -27107 -34633 -27061 -34599
rect -27027 -34633 -26981 -34599
rect -26947 -34633 -26901 -34599
rect -26867 -34633 -26821 -34599
rect -26787 -34633 -26741 -34599
rect -26707 -34633 -26661 -34599
rect -26627 -34633 -26581 -34599
rect -26547 -34633 -26501 -34599
rect -26467 -34633 -26421 -34599
rect -26387 -34633 -26341 -34599
rect -26307 -34633 -26261 -34599
rect -26227 -34633 -26181 -34599
rect -26147 -34633 -26101 -34599
rect -26067 -34633 -26021 -34599
rect -25987 -34633 -25941 -34599
rect -25907 -34633 -25861 -34599
rect -25827 -34633 -25781 -34599
rect -25747 -34633 -25701 -34599
rect -25667 -34633 -25621 -34599
rect -25587 -34633 -25541 -34599
rect -25507 -34633 -25461 -34599
rect -25427 -34633 -25381 -34599
rect -25347 -34633 -25301 -34599
rect -25267 -34633 -25221 -34599
rect -25187 -34633 -25141 -34599
rect -25107 -34633 -25061 -34599
rect -25027 -34633 -24981 -34599
rect -24947 -34633 -24901 -34599
rect -24867 -34633 -24821 -34599
rect -24787 -34633 -24741 -34599
rect -24707 -34633 -24661 -34599
rect -24627 -34633 -24581 -34599
rect -24547 -34633 -24501 -34599
rect -24467 -34633 -24421 -34599
rect -24387 -34633 -24341 -34599
rect -24307 -34633 -24261 -34599
rect -24227 -34633 -24181 -34599
rect -24147 -34633 -24101 -34599
rect -24067 -34633 -24021 -34599
rect -23987 -34633 -23941 -34599
rect -23907 -34633 -23861 -34599
rect -23827 -34633 -23781 -34599
rect -23747 -34633 -23701 -34599
rect -23667 -34633 -23621 -34599
rect -23587 -34633 -23541 -34599
rect -23507 -34633 -23461 -34599
rect -23427 -34633 -23381 -34599
rect -23347 -34633 -23301 -34599
rect -23267 -34633 -23221 -34599
rect -23187 -34633 -23141 -34599
rect -23107 -34633 -23061 -34599
rect -23027 -34633 -22981 -34599
rect -22947 -34633 -22901 -34599
rect -22867 -34633 -22821 -34599
rect -22787 -34633 -22741 -34599
rect -22707 -34633 -22661 -34599
rect -22627 -34633 -22581 -34599
rect -22547 -34633 -22501 -34599
rect -22467 -34633 -22421 -34599
rect -22387 -34633 -22341 -34599
rect -22307 -34633 -22261 -34599
rect -22227 -34633 -22181 -34599
rect -22147 -34633 -22101 -34599
rect -22067 -34633 -22021 -34599
rect -21987 -34633 -21941 -34599
rect -21907 -34633 -21861 -34599
rect -21827 -34633 -21781 -34599
rect -21747 -34633 -21701 -34599
rect -21667 -34633 -21621 -34599
rect -21587 -34633 -21541 -34599
rect -21507 -34633 -21461 -34599
rect -21427 -34633 -21381 -34599
rect -21347 -34633 -21301 -34599
rect -21267 -34633 -21221 -34599
rect -21187 -34633 -21141 -34599
rect -21107 -34633 -21061 -34599
rect -21027 -34633 -20981 -34599
rect -20947 -34633 -20901 -34599
rect -20867 -34633 -20821 -34599
rect -20787 -34633 -20741 -34599
rect -20707 -34633 -20661 -34599
rect -20627 -34633 -20581 -34599
rect -20547 -34633 -20501 -34599
rect -20467 -34633 -20421 -34599
rect -20387 -34633 -20341 -34599
rect -20307 -34633 -20261 -34599
rect -20227 -34633 -20181 -34599
rect -20147 -34633 -20101 -34599
rect -20067 -34633 -20021 -34599
rect -19987 -34633 -19941 -34599
rect -19907 -34633 -19861 -34599
rect -19827 -34633 -19781 -34599
rect -19747 -34633 -19701 -34599
rect -19667 -34633 -19621 -34599
rect -19587 -34633 -19541 -34599
rect -19507 -34633 -19461 -34599
rect -19427 -34633 -19381 -34599
rect -19347 -34633 -19301 -34599
rect -19267 -34633 -19221 -34599
rect -19187 -34633 -19141 -34599
rect -19107 -34633 -19061 -34599
rect -19027 -34633 -18981 -34599
rect -18947 -34633 -18901 -34599
rect -18867 -34633 -18821 -34599
rect -18787 -34633 -18741 -34599
rect -18707 -34633 -18661 -34599
rect -18627 -34633 -18581 -34599
rect -18547 -34633 -18500 -34599
rect -18466 -34633 -18420 -34599
rect -18386 -34633 -18340 -34599
rect -18306 -34633 -18260 -34599
rect -18226 -34633 -18180 -34599
rect -18146 -34633 -18100 -34599
rect -18066 -34633 -18020 -34599
rect -17986 -34633 -17940 -34599
rect -17906 -34633 -17860 -34599
rect -17826 -34633 -17780 -34599
rect -17746 -34633 -17700 -34599
rect -17666 -34633 -17620 -34599
rect -17586 -34633 -17540 -34599
rect -17506 -34633 -17460 -34599
rect -17426 -34633 -17380 -34599
rect -17346 -34633 -17300 -34599
rect -17266 -34633 -17220 -34599
rect -17186 -34633 -17140 -34599
rect -17106 -34633 -17060 -34599
rect -17026 -34633 -16980 -34599
rect -16946 -34633 -16900 -34599
rect -16866 -34633 -16820 -34599
rect -16786 -34633 -16740 -34599
rect -16706 -34633 -16660 -34599
rect -16626 -34633 -16580 -34599
rect -16546 -34633 -16500 -34599
rect -16466 -34633 -16420 -34599
rect -16386 -34633 -16340 -34599
rect -16306 -34633 -16260 -34599
rect -16226 -34633 -16180 -34599
rect -16146 -34633 -16100 -34599
rect -16066 -34633 -16020 -34599
rect -15986 -34633 -15940 -34599
rect -15906 -34633 -15860 -34599
rect -15826 -34633 -15780 -34599
rect -15746 -34633 -15700 -34599
rect -15666 -34633 -15620 -34599
rect -15586 -34633 -15540 -34599
rect -15506 -34633 -15460 -34599
rect -15426 -34633 -15380 -34599
rect -15346 -34633 -15300 -34599
rect -15266 -34633 -15220 -34599
rect -15186 -34633 -15140 -34599
rect -15106 -34633 -15060 -34599
rect -15026 -34633 -14980 -34599
rect -14946 -34633 -14900 -34599
rect -14866 -34633 -14820 -34599
rect -14786 -34633 -14740 -34599
rect -14706 -34633 -14660 -34599
rect -14626 -34633 -14580 -34599
rect -14546 -34633 -14500 -34599
rect -14466 -34633 -14420 -34599
rect -14386 -34633 -14340 -34599
rect -14306 -34633 -14260 -34599
rect -14226 -34633 -14180 -34599
rect -14146 -34633 -14100 -34599
rect -14066 -34633 -14020 -34599
rect -13986 -34633 -13940 -34599
rect -13906 -34633 -13860 -34599
rect -13826 -34633 -13780 -34599
rect -13746 -34633 -13700 -34599
rect -13666 -34633 -13620 -34599
rect -13586 -34633 -13540 -34599
rect -13506 -34633 -13460 -34599
rect -13426 -34633 -13380 -34599
rect -13346 -34633 -13300 -34599
rect -13266 -34633 -13220 -34599
rect -13186 -34633 -13140 -34599
rect -13106 -34633 -13060 -34599
rect -13026 -34633 -12980 -34599
rect -12946 -34633 -12900 -34599
rect -12866 -34633 -12820 -34599
rect -12786 -34633 -12740 -34599
rect -12706 -34633 -12660 -34599
rect -12626 -34633 -12580 -34599
rect -12546 -34633 -12500 -34599
rect -12466 -34633 -12420 -34599
rect -12386 -34633 -12340 -34599
rect -12306 -34633 -12260 -34599
rect -12226 -34633 -12180 -34599
rect -12146 -34633 -12100 -34599
rect -12066 -34633 -12020 -34599
rect -11986 -34633 -11940 -34599
rect -11906 -34633 -11860 -34599
rect -11826 -34633 -11780 -34599
rect -11746 -34633 -11700 -34599
rect -11666 -34633 -11620 -34599
rect -11586 -34633 -11540 -34599
rect -11506 -34633 -11460 -34599
rect -11426 -34633 -11380 -34599
rect -11346 -34633 -11300 -34599
rect -11266 -34633 -11220 -34599
rect -11186 -34633 -11140 -34599
rect -11106 -34633 -11060 -34599
rect -11026 -34633 -10980 -34599
rect -10946 -34633 -10900 -34599
rect -10866 -34633 -10820 -34599
rect -10786 -34633 -10740 -34599
rect -10706 -34633 -10660 -34599
rect -10626 -34633 -10580 -34599
rect -10546 -34633 -10500 -34599
rect -10466 -34633 -10420 -34599
rect -10386 -34633 -10340 -34599
rect -10306 -34633 -10260 -34599
rect -10226 -34633 -10180 -34599
rect -10146 -34633 -10100 -34599
rect -10066 -34633 -10020 -34599
rect -9986 -34633 -9940 -34599
rect -9906 -34633 -9859 -34599
rect -9825 -34633 -9779 -34599
rect -9745 -34633 -9699 -34599
rect -9665 -34633 -9619 -34599
rect -9585 -34633 -9539 -34599
rect -9505 -34633 -9459 -34599
rect -9425 -34633 -9379 -34599
rect -9345 -34633 -9299 -34599
rect -9265 -34633 -9219 -34599
rect -9185 -34633 -9139 -34599
rect -9105 -34633 -9059 -34599
rect -9025 -34633 -8979 -34599
rect -8945 -34633 -8899 -34599
rect -8865 -34633 -8819 -34599
rect -8785 -34633 -8739 -34599
rect -8705 -34633 -8659 -34599
rect -8625 -34633 -8579 -34599
rect -8545 -34633 -8499 -34599
rect -8465 -34633 -8419 -34599
rect -8385 -34633 -8339 -34599
rect -8305 -34633 -8259 -34599
rect -8225 -34633 -8179 -34599
rect -8145 -34633 -8099 -34599
rect -8065 -34633 -8019 -34599
rect -7985 -34633 -7939 -34599
rect -7905 -34633 -7859 -34599
rect -7825 -34633 -7779 -34599
rect -7745 -34633 -7699 -34599
rect -7665 -34633 -7619 -34599
rect -7585 -34633 -7539 -34599
rect -7505 -34633 -7459 -34599
rect -7425 -34633 -7379 -34599
rect -7345 -34633 -7299 -34599
rect -7265 -34633 -7219 -34599
rect -7185 -34633 -7139 -34599
rect -7105 -34633 -7059 -34599
rect -7025 -34633 -6979 -34599
rect -6945 -34633 -6899 -34599
rect -6865 -34633 -6819 -34599
rect -6785 -34633 -6739 -34599
rect -6705 -34633 -6659 -34599
rect -6625 -34633 -6579 -34599
rect -6545 -34633 -6499 -34599
rect -6465 -34633 -6419 -34599
rect -6385 -34633 -6339 -34599
rect -6305 -34633 -6259 -34599
rect -6225 -34633 -6179 -34599
rect -6145 -34633 -6099 -34599
rect -6065 -34633 -6019 -34599
rect -5985 -34633 -5939 -34599
rect -5905 -34633 -5859 -34599
rect -5825 -34633 -5779 -34599
rect -5745 -34633 -5699 -34599
rect -5665 -34633 -5619 -34599
rect -5585 -34633 -5539 -34599
rect -5505 -34633 -5459 -34599
rect -5425 -34633 -5379 -34599
rect -5345 -34633 -5299 -34599
rect -5265 -34633 -5219 -34599
rect -5185 -34633 -5139 -34599
rect -5105 -34633 -5059 -34599
rect -5025 -34633 -4979 -34599
rect -4945 -34633 -4899 -34599
rect -4865 -34633 -4819 -34599
rect -4785 -34633 -4739 -34599
rect -4705 -34633 -4659 -34599
rect -4625 -34633 -4579 -34599
rect -4545 -34633 -4499 -34599
rect -4465 -34633 -4419 -34599
rect -4385 -34633 -4339 -34599
rect -4305 -34633 -4259 -34599
rect -4225 -34633 -4140 -34599
rect -4106 -34633 -4060 -34599
rect -4026 -34633 -3980 -34599
rect -3946 -34633 -3900 -34599
rect -3866 -34633 -3820 -34599
rect -3786 -34633 -3740 -34599
rect -3706 -34633 -3660 -34599
rect -3626 -34633 -3580 -34599
rect -3546 -34633 -3500 -34599
rect -3466 -34633 -3420 -34599
rect -3386 -34633 -3340 -34599
rect -3306 -34633 -3260 -34599
rect -3226 -34633 -3180 -34599
rect -3146 -34633 -3100 -34599
rect -3066 -34633 -3020 -34599
rect -2986 -34633 -2940 -34599
rect -2906 -34633 -2860 -34599
rect -2826 -34633 -2780 -34599
rect -2746 -34633 -2700 -34599
rect -2666 -34633 -2620 -34599
rect -2586 -34633 -2540 -34599
rect -2506 -34633 -2460 -34599
rect -2426 -34633 -2380 -34599
rect -2346 -34633 -2300 -34599
rect -2266 -34633 -2220 -34599
rect -2186 -34633 -2140 -34599
rect -2106 -34633 -2060 -34599
rect -2026 -34633 -1980 -34599
rect -1946 -34633 -1900 -34599
rect -1866 -34633 -1820 -34599
rect -1786 -34633 -1740 -34599
rect -1706 -34633 -1660 -34599
rect -1626 -34633 -1580 -34599
rect -1546 -34633 -1500 -34599
rect -1466 -34633 -1420 -34599
rect -1386 -34633 -1340 -34599
rect -1306 -34633 -1260 -34599
rect -1226 -34633 -1180 -34599
rect -1146 -34633 -1100 -34599
rect -1066 -34633 -1020 -34599
rect -986 -34633 -940 -34599
rect -906 -34633 -860 -34599
rect -826 -34633 -780 -34599
rect -746 -34633 -700 -34599
rect -666 -34633 -620 -34599
rect -586 -34633 -540 -34599
rect -506 -34633 -460 -34599
rect -426 -34633 -380 -34599
rect -346 -34633 -300 -34599
rect -266 -34633 -220 -34599
rect -186 -34633 -140 -34599
rect -106 -34633 -60 -34599
rect -26 -34633 20 -34599
rect 54 -34633 100 -34599
rect 134 -34633 180 -34599
rect 214 -34633 260 -34599
rect 294 -34633 340 -34599
rect 374 -34633 420 -34599
rect 454 -34633 500 -34599
rect 534 -34633 580 -34599
rect 614 -34633 660 -34599
rect 694 -34633 740 -34599
rect 774 -34633 820 -34599
rect 854 -34633 900 -34599
rect 934 -34633 980 -34599
rect 1014 -34633 1060 -34599
rect 1094 -34633 1140 -34599
rect 1174 -34633 1220 -34599
rect 1254 -34633 1300 -34599
rect 1334 -34633 1380 -34599
rect 1414 -34633 1460 -34599
rect 1494 -34633 1540 -34599
rect 1574 -34633 1620 -34599
rect 1654 -34633 1700 -34599
rect 1734 -34633 1780 -34599
rect 1814 -34633 1860 -34599
rect 1894 -34633 1940 -34599
rect 1974 -34633 2020 -34599
rect 2054 -34633 2100 -34599
rect 2134 -34633 2180 -34599
rect 2214 -34633 2260 -34599
rect 2294 -34633 2340 -34599
rect 2374 -34633 2420 -34599
rect 2454 -34633 2500 -34599
rect 2534 -34633 2580 -34599
rect 2614 -34633 2660 -34599
rect 2694 -34633 2740 -34599
rect 2774 -34633 2820 -34599
rect 2854 -34633 2900 -34599
rect 2934 -34633 2980 -34599
rect 3014 -34633 3060 -34599
rect 3094 -34633 3140 -34599
rect 3174 -34633 3220 -34599
rect 3254 -34633 3300 -34599
rect 3334 -34633 3380 -34599
rect 3414 -34633 3460 -34599
rect 3494 -34633 3540 -34599
rect 3574 -34633 3620 -34599
rect 3654 -34633 3700 -34599
rect 3734 -34633 3780 -34599
rect 3814 -34633 3860 -34599
rect 3894 -34633 3940 -34599
rect 3974 -34633 4020 -34599
rect 4054 -34633 4100 -34599
rect 4134 -34633 4180 -34599
rect 4214 -34633 4260 -34599
rect 4294 -34633 4340 -34599
rect 4374 -34633 4420 -34599
rect 4454 -34633 4500 -34599
rect 4534 -34633 4580 -34599
rect 4614 -34633 4660 -34599
rect 4694 -34633 4740 -34599
rect 4774 -34633 4820 -34599
rect 4854 -34633 4900 -34599
rect 4934 -34633 4980 -34599
rect 5014 -34633 5060 -34599
rect 5094 -34633 5140 -34599
rect 5174 -34633 5220 -34599
rect 5254 -34633 5300 -34599
rect 5334 -34633 5380 -34599
rect 5414 -34633 5460 -34599
rect 5494 -34633 5540 -34599
rect 5574 -34633 5620 -34599
rect 5654 -34633 5700 -34599
rect 5734 -34633 5780 -34599
rect 5814 -34633 5860 -34599
rect 5894 -34633 5940 -34599
rect 5974 -34633 6020 -34599
rect 6054 -34633 6100 -34599
rect 6134 -34633 6180 -34599
rect 6214 -34633 6260 -34599
rect 6294 -34633 6340 -34599
rect 6374 -34633 6420 -34599
rect 6454 -34633 6500 -34599
rect 6534 -34633 6580 -34599
rect 6614 -34633 6660 -34599
rect 6694 -34633 6740 -34599
rect 6774 -34633 6820 -34599
rect 6854 -34633 6900 -34599
rect 6934 -34633 6980 -34599
rect 7014 -34633 7060 -34599
rect 7094 -34633 7140 -34599
rect 7174 -34633 7220 -34599
rect 7254 -34633 7300 -34599
rect 7334 -34633 7380 -34599
rect 7414 -34633 7460 -34599
rect 7494 -34633 7540 -34599
rect 7574 -34633 7620 -34599
rect 7654 -34633 7700 -34599
rect 7734 -34633 7780 -34599
rect 7814 -34633 7860 -34599
rect 7894 -34633 7940 -34599
rect 7974 -34633 8020 -34599
rect 8054 -34633 8100 -34599
rect 8134 -34633 8180 -34599
rect 8214 -34633 8260 -34599
rect 8294 -34633 8340 -34599
rect 8374 -34633 8420 -34599
rect 8454 -34633 8500 -34599
rect 8534 -34633 8580 -34599
rect 8614 -34633 8660 -34599
rect 8694 -34633 8740 -34599
rect 8774 -34633 8820 -34599
rect 8854 -34633 8900 -34599
rect 8934 -34633 8980 -34599
rect 9014 -34633 9060 -34599
rect 9094 -34633 9140 -34599
rect 9174 -34633 9220 -34599
rect 9254 -34633 9300 -34599
rect 9334 -34633 9380 -34599
rect 9414 -34633 9460 -34599
rect 9494 -34633 9540 -34599
rect 9574 -34633 9620 -34599
rect 9654 -34633 9700 -34599
rect 9734 -34633 9780 -34599
rect 9814 -34633 9860 -34599
rect 9894 -34633 9940 -34599
rect 9974 -34633 10020 -34599
rect 10054 -34633 10100 -34599
rect 10134 -34633 10181 -34599
rect 10215 -34633 10261 -34599
rect 10295 -34633 10341 -34599
rect 10375 -34633 10421 -34599
rect 10455 -34633 10501 -34599
rect 10535 -34633 10581 -34599
rect 10615 -34633 10661 -34599
rect 10695 -34633 10741 -34599
rect 10775 -34633 10821 -34599
rect 10855 -34633 10901 -34599
rect 10935 -34633 10981 -34599
rect 11015 -34633 11061 -34599
rect 11095 -34633 11141 -34599
rect 11175 -34633 11221 -34599
rect 11255 -34633 11301 -34599
rect 11335 -34633 11381 -34599
rect 11415 -34633 11461 -34599
rect 11495 -34633 11541 -34599
rect 11575 -34633 11621 -34599
rect 11655 -34633 11701 -34599
rect 11735 -34633 11781 -34599
rect 11815 -34633 11861 -34599
rect 11895 -34633 11941 -34599
rect 11975 -34633 12021 -34599
rect 12055 -34633 12101 -34599
rect 12135 -34633 12181 -34599
rect 12215 -34633 12261 -34599
rect 12295 -34633 12341 -34599
rect 12375 -34633 12421 -34599
rect 12455 -34633 12501 -34599
rect 12535 -34633 12581 -34599
rect 12615 -34633 12661 -34599
rect 12695 -34633 12741 -34599
rect 12775 -34633 12821 -34599
rect 12855 -34633 12901 -34599
rect 12935 -34633 12981 -34599
rect 13015 -34633 13061 -34599
rect 13095 -34633 13141 -34599
rect 13175 -34633 13221 -34599
rect 13255 -34633 13301 -34599
rect 13335 -34633 13381 -34599
rect 13415 -34633 13461 -34599
rect 13495 -34633 13541 -34599
rect 13575 -34633 13621 -34599
rect 13655 -34633 13701 -34599
rect 13735 -34633 13781 -34599
rect 13815 -34633 13861 -34599
rect 13895 -34633 13941 -34599
rect 13975 -34633 14021 -34599
rect 14055 -34633 14101 -34599
rect 14135 -34633 14181 -34599
rect 14215 -34633 14261 -34599
rect 14295 -34633 14341 -34599
rect 14375 -34633 14421 -34599
rect 14455 -34633 14501 -34599
rect 14535 -34633 14581 -34599
rect 14615 -34633 14661 -34599
rect 14695 -34633 14741 -34599
rect 14775 -34633 14821 -34599
rect 14855 -34633 14901 -34599
rect 14935 -34633 14981 -34599
rect 15015 -34633 15061 -34599
rect 15095 -34633 15141 -34599
rect 15175 -34633 15221 -34599
rect 15255 -34633 15301 -34599
rect 15335 -34633 15381 -34599
rect 15415 -34633 15461 -34599
rect 15495 -34633 15541 -34599
rect 15575 -34633 15621 -34599
rect 15655 -34633 15701 -34599
rect 15735 -34633 15781 -34599
rect 15815 -34633 15861 -34599
rect 15895 -34633 15941 -34599
rect 15975 -34633 16021 -34599
rect 16055 -34633 16101 -34599
rect 16135 -34633 16181 -34599
rect 16215 -34633 16261 -34599
rect 16295 -34633 16341 -34599
rect 16375 -34633 16421 -34599
rect 16455 -34633 16501 -34599
rect 16535 -34633 16581 -34599
rect 16615 -34633 16661 -34599
rect 16695 -34633 16741 -34599
rect 16775 -34633 16821 -34599
rect 16855 -34633 16901 -34599
rect 16935 -34633 16981 -34599
rect 17015 -34633 17061 -34599
rect 17095 -34633 17141 -34599
rect 17175 -34633 17221 -34599
rect 17255 -34633 17301 -34599
rect 17335 -34633 17381 -34599
rect 17415 -34633 17461 -34599
rect 17495 -34633 17541 -34599
rect 17575 -34633 17621 -34599
rect 17655 -34633 17701 -34599
rect 17735 -34633 17781 -34599
rect 17815 -34633 17861 -34599
rect 17895 -34633 17941 -34599
rect 17975 -34633 18021 -34599
rect 18055 -34633 18101 -34599
rect 18135 -34633 18181 -34599
rect 18215 -34633 18261 -34599
rect 18295 -34633 18341 -34599
rect 18375 -34633 18421 -34599
rect 18455 -34633 18501 -34599
rect 18535 -34633 18581 -34599
rect 18615 -34633 18661 -34599
rect 18695 -34633 18741 -34599
rect 18775 -34633 18821 -34599
rect 18855 -34633 18901 -34599
rect 18935 -34633 18981 -34599
rect 19015 -34633 19061 -34599
rect 19095 -34633 19141 -34599
rect 19175 -34633 19221 -34599
rect 19255 -34633 19301 -34599
rect 19335 -34633 19381 -34599
rect 19415 -34633 19461 -34599
rect 19495 -34633 19541 -34599
rect 19575 -34633 19621 -34599
rect 19655 -34633 19701 -34599
rect 19735 -34633 19781 -34599
rect 19815 -34633 19861 -34599
rect 19895 -34633 19941 -34599
rect 19975 -34633 20021 -34599
rect 20055 -34633 20101 -34599
rect 20135 -34633 20181 -34599
rect 20215 -34633 20261 -34599
rect 20295 -34633 20341 -34599
rect 20375 -34633 20421 -34599
rect 20455 -34633 20501 -34599
rect 20535 -34633 20581 -34599
rect 20615 -34633 20661 -34599
rect 20695 -34633 20741 -34599
rect 20775 -34633 20821 -34599
rect 20855 -34633 20901 -34599
rect 20935 -34633 20981 -34599
rect 21015 -34633 21061 -34599
rect 21095 -34633 21141 -34599
rect 21175 -34633 21221 -34599
rect 21255 -34633 21301 -34599
rect 21335 -34633 21381 -34599
rect 21415 -34633 21461 -34599
rect 21495 -34633 21541 -34599
rect 21575 -34633 21621 -34599
rect 21655 -34633 21701 -34599
rect 21735 -34633 21781 -34599
rect 21815 -34633 21861 -34599
rect 21895 -34633 21941 -34599
rect 21975 -34633 22021 -34599
rect 22055 -34633 22101 -34599
rect 22135 -34633 22181 -34599
rect 22215 -34633 22261 -34599
rect 22295 -34633 22341 -34599
rect 22375 -34633 22421 -34599
rect 22455 -34633 22501 -34599
rect 22535 -34633 22581 -34599
rect 22615 -34633 22661 -34599
rect 22695 -34633 22741 -34599
rect 22775 -34633 22821 -34599
rect 22855 -34633 22901 -34599
rect 22935 -34633 22981 -34599
rect 23015 -34633 23061 -34599
rect 23095 -34633 23141 -34599
rect 23175 -34633 23221 -34599
rect 23255 -34633 23301 -34599
rect 23335 -34633 23381 -34599
rect 23415 -34633 23461 -34599
rect 23495 -34633 23541 -34599
rect 23575 -34633 23621 -34599
rect 23655 -34633 23701 -34599
rect 23735 -34633 23781 -34599
rect 23815 -34633 23861 -34599
rect 23895 -34633 23941 -34599
rect 23975 -34633 24021 -34599
rect 24055 -34633 24101 -34599
rect 24135 -34633 24181 -34599
rect 24215 -34633 24261 -34599
rect 24295 -34633 24341 -34599
rect 24375 -34633 24421 -34599
rect 24455 -34633 24501 -34599
rect 24535 -34633 24581 -34599
rect 24615 -34633 24661 -34599
rect 24695 -34633 24741 -34599
rect 24775 -34633 24821 -34599
rect 24855 -34633 24901 -34599
rect 24935 -34633 24981 -34599
rect 25015 -34633 25061 -34599
rect 25095 -34633 25141 -34599
rect 25175 -34633 25221 -34599
rect 25255 -34633 25301 -34599
rect 25335 -34633 25381 -34599
rect 25415 -34633 25461 -34599
rect 25495 -34633 25541 -34599
rect 25575 -34633 25621 -34599
rect 25655 -34633 25701 -34599
rect 25735 -34633 25781 -34599
rect 25815 -34633 25861 -34599
rect 25895 -34633 25941 -34599
rect 25975 -34633 26021 -34599
rect 26055 -34633 26101 -34599
rect 26135 -34633 26181 -34599
rect 26215 -34633 26261 -34599
rect 26295 -34633 26341 -34599
rect 26375 -34633 26421 -34599
rect 26455 -34633 26501 -34599
rect 26535 -34633 26581 -34599
rect 26615 -34633 26661 -34599
rect 26695 -34633 26741 -34599
rect 26775 -34633 26821 -34599
rect 26855 -34633 26901 -34599
rect 26935 -34633 26981 -34599
rect 27015 -34633 27061 -34599
rect 27095 -34633 27141 -34599
rect 27175 -34633 27221 -34599
rect 27255 -34633 27301 -34599
rect 27335 -34633 27381 -34599
rect 27415 -34633 27461 -34599
rect 27495 -34633 27541 -34599
rect 27575 -34633 27621 -34599
rect 27655 -34633 27701 -34599
rect 27735 -34633 27781 -34599
rect 27815 -34633 27861 -34599
rect 27895 -34633 27941 -34599
rect 27975 -34633 28021 -34599
rect 28055 -34633 28101 -34599
rect 28135 -34633 28181 -34599
rect 28215 -34633 28261 -34599
rect 28295 -34633 28341 -34599
rect 28375 -34633 28421 -34599
rect 28455 -34633 28501 -34599
rect 28535 -34633 28581 -34599
rect 28615 -34633 28661 -34599
rect 28695 -34633 28741 -34599
rect 28775 -34633 28821 -34599
rect 28855 -34633 28901 -34599
rect 28935 -34633 28981 -34599
rect 29015 -34633 29061 -34599
rect 29095 -34633 29141 -34599
rect 29175 -34633 29221 -34599
rect 29255 -34633 29301 -34599
rect 29335 -34633 29381 -34599
rect 29415 -34633 29461 -34599
rect 29495 -34633 29541 -34599
rect 29575 -34633 29621 -34599
rect 29655 -34633 29701 -34599
rect 29735 -34633 29781 -34599
rect 29815 -34633 29861 -34599
rect 29895 -34633 29941 -34599
rect 29975 -34633 30021 -34599
rect 30055 -34633 30101 -34599
rect 30135 -34633 30181 -34599
rect 30215 -34633 30261 -34599
rect 30295 -34633 30341 -34599
rect 30375 -34633 30421 -34599
rect 30455 -34633 30501 -34599
rect 30535 -34633 30581 -34599
rect 30615 -34633 30661 -34599
rect 30695 -34633 30741 -34599
rect 30775 -34633 30821 -34599
rect 30855 -34633 30901 -34599
rect 30935 -34633 30981 -34599
rect 31015 -34633 31061 -34599
rect 31095 -34633 31141 -34599
rect 31175 -34633 31221 -34599
rect 31255 -34633 31301 -34599
rect 31335 -34633 31381 -34599
rect 31415 -34633 31461 -34599
rect 31495 -34633 31541 -34599
rect 31575 -34633 31621 -34599
rect 31655 -34633 31701 -34599
rect 31735 -34633 31781 -34599
rect -44468 -34656 31781 -34633
rect -27254 -34719 -27174 -34696
rect -27254 -34753 -27231 -34719
rect -27197 -34753 -27174 -34719
rect -27254 -34776 -27174 -34753
rect -27134 -34719 -27054 -34696
rect -27134 -34753 -27111 -34719
rect -27077 -34753 -27054 -34719
rect -27134 -34776 -27054 -34753
rect 12081 -34720 12161 -34697
rect 12081 -34754 12104 -34720
rect 12138 -34754 12161 -34720
rect 12081 -34777 12161 -34754
rect 12201 -34720 12281 -34697
rect 12201 -34754 12224 -34720
rect 12258 -34754 12281 -34720
rect 12201 -34777 12281 -34754
rect -27254 -34839 -27174 -34816
rect -27254 -34873 -27231 -34839
rect -27197 -34873 -27174 -34839
rect -27254 -34896 -27174 -34873
rect -27134 -34839 -27054 -34816
rect -27134 -34873 -27111 -34839
rect -27077 -34873 -27054 -34839
rect -27134 -34896 -27054 -34873
rect 12081 -34840 12161 -34817
rect 12081 -34874 12104 -34840
rect 12138 -34874 12161 -34840
rect 12081 -34897 12161 -34874
rect 12201 -34840 12281 -34817
rect 12201 -34874 12224 -34840
rect 12258 -34874 12281 -34840
rect 12201 -34897 12281 -34874
rect -44468 -42458 -624 -42435
rect -44468 -42492 -44422 -42458
rect -44388 -42492 -44342 -42458
rect -44308 -42492 -44262 -42458
rect -44228 -42492 -44182 -42458
rect -44148 -42492 -44102 -42458
rect -44068 -42492 -44022 -42458
rect -43988 -42492 -43942 -42458
rect -43908 -42492 -43862 -42458
rect -43828 -42492 -43782 -42458
rect -43748 -42492 -43702 -42458
rect -43668 -42492 -43622 -42458
rect -43588 -42492 -43542 -42458
rect -43508 -42492 -43462 -42458
rect -43428 -42492 -43382 -42458
rect -43348 -42492 -43302 -42458
rect -43268 -42492 -43222 -42458
rect -43188 -42492 -43142 -42458
rect -43108 -42492 -43062 -42458
rect -43028 -42492 -42982 -42458
rect -42948 -42492 -42902 -42458
rect -42868 -42492 -42822 -42458
rect -42788 -42492 -42742 -42458
rect -42708 -42492 -42662 -42458
rect -42628 -42492 -42582 -42458
rect -42548 -42492 -42502 -42458
rect -42468 -42492 -42422 -42458
rect -42388 -42492 -42342 -42458
rect -42308 -42492 -42262 -42458
rect -42228 -42492 -42182 -42458
rect -42148 -42492 -42102 -42458
rect -42068 -42492 -42022 -42458
rect -41988 -42492 -41942 -42458
rect -41908 -42492 -41862 -42458
rect -41828 -42492 -41782 -42458
rect -41748 -42492 -41702 -42458
rect -41668 -42492 -41622 -42458
rect -41588 -42492 -41542 -42458
rect -41508 -42492 -41462 -42458
rect -41428 -42492 -41382 -42458
rect -41348 -42492 -41302 -42458
rect -41268 -42492 -41222 -42458
rect -41188 -42492 -41142 -42458
rect -41108 -42492 -41062 -42458
rect -41028 -42492 -40982 -42458
rect -40948 -42492 -40902 -42458
rect -40868 -42492 -40822 -42458
rect -40788 -42492 -40742 -42458
rect -40708 -42492 -40662 -42458
rect -40628 -42492 -40582 -42458
rect -40548 -42492 -40502 -42458
rect -40468 -42492 -40422 -42458
rect -40388 -42492 -40342 -42458
rect -40308 -42492 -40262 -42458
rect -40228 -42492 -40182 -42458
rect -40148 -42492 -40102 -42458
rect -40068 -42492 -40022 -42458
rect -39988 -42492 -39942 -42458
rect -39908 -42492 -39862 -42458
rect -39828 -42492 -39782 -42458
rect -39748 -42492 -39702 -42458
rect -39668 -42492 -39622 -42458
rect -39588 -42492 -39542 -42458
rect -39508 -42492 -39462 -42458
rect -39428 -42492 -39382 -42458
rect -39348 -42492 -39302 -42458
rect -39268 -42492 -39222 -42458
rect -39188 -42492 -39142 -42458
rect -39108 -42492 -39062 -42458
rect -39028 -42492 -38982 -42458
rect -38948 -42492 -38902 -42458
rect -38868 -42492 -38822 -42458
rect -38788 -42492 -38742 -42458
rect -38708 -42492 -38662 -42458
rect -38628 -42492 -38582 -42458
rect -38548 -42492 -38502 -42458
rect -38468 -42492 -38422 -42458
rect -38388 -42492 -38342 -42458
rect -38308 -42492 -38262 -42458
rect -38228 -42492 -38182 -42458
rect -38148 -42492 -38102 -42458
rect -38068 -42492 -38022 -42458
rect -37988 -42492 -37942 -42458
rect -37908 -42492 -37862 -42458
rect -37828 -42492 -37782 -42458
rect -37748 -42492 -37702 -42458
rect -37668 -42492 -37622 -42458
rect -37588 -42492 -37542 -42458
rect -37508 -42492 -37462 -42458
rect -37428 -42492 -37382 -42458
rect -37348 -42492 -37302 -42458
rect -37268 -42492 -37222 -42458
rect -37188 -42492 -37142 -42458
rect -37108 -42492 -37062 -42458
rect -37028 -42492 -36982 -42458
rect -36948 -42492 -36902 -42458
rect -36868 -42492 -36822 -42458
rect -36788 -42492 -36742 -42458
rect -36708 -42492 -36662 -42458
rect -36628 -42492 -36582 -42458
rect -36548 -42492 -36502 -42458
rect -36468 -42492 -36422 -42458
rect -36388 -42492 -36342 -42458
rect -36308 -42492 -36262 -42458
rect -36228 -42492 -36182 -42458
rect -36148 -42492 -36102 -42458
rect -36068 -42492 -36022 -42458
rect -35988 -42492 -35942 -42458
rect -35908 -42492 -35862 -42458
rect -35828 -42492 -35782 -42458
rect -35748 -42492 -35702 -42458
rect -35668 -42492 -35622 -42458
rect -35588 -42492 -35542 -42458
rect -35508 -42492 -35462 -42458
rect -35428 -42492 -35382 -42458
rect -35348 -42492 -35302 -42458
rect -35268 -42492 -35222 -42458
rect -35188 -42492 -35142 -42458
rect -35108 -42492 -35062 -42458
rect -35028 -42492 -34982 -42458
rect -34948 -42492 -34902 -42458
rect -34868 -42492 -34822 -42458
rect -34788 -42492 -34742 -42458
rect -34708 -42492 -34662 -42458
rect -34628 -42492 -34582 -42458
rect -34548 -42492 -34502 -42458
rect -34468 -42492 -34422 -42458
rect -34388 -42492 -34342 -42458
rect -34308 -42492 -34262 -42458
rect -34228 -42492 -34182 -42458
rect -34148 -42492 -34102 -42458
rect -34068 -42492 -34022 -42458
rect -33988 -42492 -33942 -42458
rect -33908 -42492 -33862 -42458
rect -33828 -42492 -33782 -42458
rect -33748 -42492 -33702 -42458
rect -33668 -42492 -33622 -42458
rect -33588 -42492 -33542 -42458
rect -33508 -42492 -33462 -42458
rect -33428 -42492 -33382 -42458
rect -33348 -42492 -33302 -42458
rect -33268 -42492 -33222 -42458
rect -33188 -42492 -33142 -42458
rect -33108 -42492 -33062 -42458
rect -33028 -42492 -32982 -42458
rect -32948 -42492 -32902 -42458
rect -32868 -42492 -32822 -42458
rect -32788 -42492 -32742 -42458
rect -32708 -42492 -32662 -42458
rect -32628 -42492 -32582 -42458
rect -32548 -42492 -32502 -42458
rect -32468 -42492 -32422 -42458
rect -32388 -42492 -32342 -42458
rect -32308 -42492 -32262 -42458
rect -32228 -42492 -32182 -42458
rect -32148 -42492 -32102 -42458
rect -32068 -42492 -32022 -42458
rect -31988 -42492 -31942 -42458
rect -31908 -42492 -31862 -42458
rect -31828 -42492 -31782 -42458
rect -31748 -42492 -31702 -42458
rect -31668 -42492 -31622 -42458
rect -31588 -42492 -31542 -42458
rect -31508 -42492 -31461 -42458
rect -31427 -42492 -31381 -42458
rect -31347 -42492 -31301 -42458
rect -31267 -42492 -31221 -42458
rect -31187 -42492 -31141 -42458
rect -31107 -42492 -31061 -42458
rect -31027 -42492 -30981 -42458
rect -30947 -42492 -30901 -42458
rect -30867 -42492 -30821 -42458
rect -30787 -42492 -30741 -42458
rect -30707 -42492 -30661 -42458
rect -30627 -42492 -30581 -42458
rect -30547 -42492 -30501 -42458
rect -30467 -42492 -30421 -42458
rect -30387 -42492 -30341 -42458
rect -30307 -42492 -30261 -42458
rect -30227 -42492 -30181 -42458
rect -30147 -42492 -30101 -42458
rect -30067 -42492 -30021 -42458
rect -29987 -42492 -29941 -42458
rect -29907 -42492 -29861 -42458
rect -29827 -42492 -29781 -42458
rect -29747 -42492 -29701 -42458
rect -29667 -42492 -29621 -42458
rect -29587 -42492 -29541 -42458
rect -29507 -42492 -29461 -42458
rect -29427 -42492 -29381 -42458
rect -29347 -42492 -29301 -42458
rect -29267 -42492 -29221 -42458
rect -29187 -42492 -29141 -42458
rect -29107 -42492 -29061 -42458
rect -29027 -42492 -28981 -42458
rect -28947 -42492 -28901 -42458
rect -28867 -42492 -28821 -42458
rect -28787 -42492 -28741 -42458
rect -28707 -42492 -28661 -42458
rect -28627 -42492 -28581 -42458
rect -28547 -42492 -28501 -42458
rect -28467 -42492 -28421 -42458
rect -28387 -42492 -28341 -42458
rect -28307 -42492 -28261 -42458
rect -28227 -42492 -28181 -42458
rect -28147 -42492 -28101 -42458
rect -28067 -42492 -28021 -42458
rect -27987 -42492 -27941 -42458
rect -27907 -42492 -27861 -42458
rect -27827 -42492 -27781 -42458
rect -27747 -42492 -27701 -42458
rect -27667 -42492 -27621 -42458
rect -27587 -42492 -27541 -42458
rect -27507 -42492 -27461 -42458
rect -27427 -42492 -27381 -42458
rect -27347 -42492 -27301 -42458
rect -27267 -42492 -27221 -42458
rect -27187 -42492 -27141 -42458
rect -27107 -42492 -27061 -42458
rect -27027 -42492 -26981 -42458
rect -26947 -42492 -26901 -42458
rect -26867 -42492 -26821 -42458
rect -26787 -42492 -26741 -42458
rect -26707 -42492 -26661 -42458
rect -26627 -42492 -26581 -42458
rect -26547 -42492 -26501 -42458
rect -26467 -42492 -26421 -42458
rect -26387 -42492 -26341 -42458
rect -26307 -42492 -26261 -42458
rect -26227 -42492 -26181 -42458
rect -26147 -42492 -26101 -42458
rect -26067 -42492 -26021 -42458
rect -25987 -42492 -25941 -42458
rect -25907 -42492 -25861 -42458
rect -25827 -42492 -25781 -42458
rect -25747 -42492 -25701 -42458
rect -25667 -42492 -25621 -42458
rect -25587 -42492 -25541 -42458
rect -25507 -42492 -25461 -42458
rect -25427 -42492 -25381 -42458
rect -25347 -42492 -25301 -42458
rect -25267 -42492 -25221 -42458
rect -25187 -42492 -25141 -42458
rect -25107 -42492 -25061 -42458
rect -25027 -42492 -24981 -42458
rect -24947 -42492 -24901 -42458
rect -24867 -42492 -24821 -42458
rect -24787 -42492 -24741 -42458
rect -24707 -42492 -24661 -42458
rect -24627 -42492 -24581 -42458
rect -24547 -42492 -24501 -42458
rect -24467 -42492 -24421 -42458
rect -24387 -42492 -24341 -42458
rect -24307 -42492 -24261 -42458
rect -24227 -42492 -24181 -42458
rect -24147 -42492 -24101 -42458
rect -24067 -42492 -24021 -42458
rect -23987 -42492 -23941 -42458
rect -23907 -42492 -23861 -42458
rect -23827 -42492 -23781 -42458
rect -23747 -42492 -23701 -42458
rect -23667 -42492 -23621 -42458
rect -23587 -42492 -23541 -42458
rect -23507 -42492 -23461 -42458
rect -23427 -42492 -23381 -42458
rect -23347 -42492 -23301 -42458
rect -23267 -42492 -23221 -42458
rect -23187 -42492 -23141 -42458
rect -23107 -42492 -23061 -42458
rect -23027 -42492 -22981 -42458
rect -22947 -42492 -22901 -42458
rect -22867 -42492 -22821 -42458
rect -22787 -42492 -22741 -42458
rect -22707 -42492 -22661 -42458
rect -22627 -42492 -22581 -42458
rect -22547 -42492 -22501 -42458
rect -22467 -42492 -22421 -42458
rect -22387 -42492 -22341 -42458
rect -22307 -42492 -22261 -42458
rect -22227 -42492 -22181 -42458
rect -22147 -42492 -22101 -42458
rect -22067 -42492 -22021 -42458
rect -21987 -42492 -21941 -42458
rect -21907 -42492 -21861 -42458
rect -21827 -42492 -21781 -42458
rect -21747 -42492 -21701 -42458
rect -21667 -42492 -21621 -42458
rect -21587 -42492 -21541 -42458
rect -21507 -42492 -21461 -42458
rect -21427 -42492 -21381 -42458
rect -21347 -42492 -21301 -42458
rect -21267 -42492 -21221 -42458
rect -21187 -42492 -21141 -42458
rect -21107 -42492 -21061 -42458
rect -21027 -42492 -20981 -42458
rect -20947 -42492 -20901 -42458
rect -20867 -42492 -20821 -42458
rect -20787 -42492 -20741 -42458
rect -20707 -42492 -20661 -42458
rect -20627 -42492 -20581 -42458
rect -20547 -42492 -20501 -42458
rect -20467 -42492 -20421 -42458
rect -20387 -42492 -20341 -42458
rect -20307 -42492 -20261 -42458
rect -20227 -42492 -20181 -42458
rect -20147 -42492 -20101 -42458
rect -20067 -42492 -20021 -42458
rect -19987 -42492 -19941 -42458
rect -19907 -42492 -19861 -42458
rect -19827 -42492 -19781 -42458
rect -19747 -42492 -19701 -42458
rect -19667 -42492 -19621 -42458
rect -19587 -42492 -19541 -42458
rect -19507 -42492 -19461 -42458
rect -19427 -42492 -19381 -42458
rect -19347 -42492 -19301 -42458
rect -19267 -42492 -19221 -42458
rect -19187 -42492 -19141 -42458
rect -19107 -42492 -19061 -42458
rect -19027 -42492 -18981 -42458
rect -18947 -42492 -18901 -42458
rect -18867 -42492 -18821 -42458
rect -18787 -42492 -18741 -42458
rect -18707 -42492 -18661 -42458
rect -18627 -42492 -18581 -42458
rect -18547 -42492 -18500 -42458
rect -18466 -42492 -18420 -42458
rect -18386 -42492 -18340 -42458
rect -18306 -42492 -18260 -42458
rect -18226 -42492 -18180 -42458
rect -18146 -42492 -18100 -42458
rect -18066 -42492 -18020 -42458
rect -17986 -42492 -17940 -42458
rect -17906 -42492 -17860 -42458
rect -17826 -42492 -17780 -42458
rect -17746 -42492 -17700 -42458
rect -17666 -42492 -17620 -42458
rect -17586 -42492 -17540 -42458
rect -17506 -42492 -17460 -42458
rect -17426 -42492 -17380 -42458
rect -17346 -42492 -17300 -42458
rect -17266 -42492 -17220 -42458
rect -17186 -42492 -17140 -42458
rect -17106 -42492 -17060 -42458
rect -17026 -42492 -16980 -42458
rect -16946 -42492 -16900 -42458
rect -16866 -42492 -16820 -42458
rect -16786 -42492 -16740 -42458
rect -16706 -42492 -16660 -42458
rect -16626 -42492 -16580 -42458
rect -16546 -42492 -16500 -42458
rect -16466 -42492 -16420 -42458
rect -16386 -42492 -16340 -42458
rect -16306 -42492 -16260 -42458
rect -16226 -42492 -16180 -42458
rect -16146 -42492 -16100 -42458
rect -16066 -42492 -16020 -42458
rect -15986 -42492 -15940 -42458
rect -15906 -42492 -15860 -42458
rect -15826 -42492 -15780 -42458
rect -15746 -42492 -15700 -42458
rect -15666 -42492 -15620 -42458
rect -15586 -42492 -15540 -42458
rect -15506 -42492 -15460 -42458
rect -15426 -42492 -15380 -42458
rect -15346 -42492 -15300 -42458
rect -15266 -42492 -15220 -42458
rect -15186 -42492 -15140 -42458
rect -15106 -42492 -15060 -42458
rect -15026 -42492 -14980 -42458
rect -14946 -42492 -14900 -42458
rect -14866 -42492 -14820 -42458
rect -14786 -42492 -14740 -42458
rect -14706 -42492 -14660 -42458
rect -14626 -42492 -14580 -42458
rect -14546 -42492 -14500 -42458
rect -14466 -42492 -14420 -42458
rect -14386 -42492 -14340 -42458
rect -14306 -42492 -14260 -42458
rect -14226 -42492 -14180 -42458
rect -14146 -42492 -14100 -42458
rect -14066 -42492 -14020 -42458
rect -13986 -42492 -13940 -42458
rect -13906 -42492 -13860 -42458
rect -13826 -42492 -13780 -42458
rect -13746 -42492 -13700 -42458
rect -13666 -42492 -13620 -42458
rect -13586 -42492 -13540 -42458
rect -13506 -42492 -13460 -42458
rect -13426 -42492 -13380 -42458
rect -13346 -42492 -13300 -42458
rect -13266 -42492 -13220 -42458
rect -13186 -42492 -13140 -42458
rect -13106 -42492 -13060 -42458
rect -13026 -42492 -12980 -42458
rect -12946 -42492 -12900 -42458
rect -12866 -42492 -12820 -42458
rect -12786 -42492 -12740 -42458
rect -12706 -42492 -12660 -42458
rect -12626 -42492 -12580 -42458
rect -12546 -42492 -12500 -42458
rect -12466 -42492 -12420 -42458
rect -12386 -42492 -12340 -42458
rect -12306 -42492 -12260 -42458
rect -12226 -42492 -12180 -42458
rect -12146 -42492 -12100 -42458
rect -12066 -42492 -12020 -42458
rect -11986 -42492 -11940 -42458
rect -11906 -42492 -11860 -42458
rect -11826 -42492 -11780 -42458
rect -11746 -42492 -11700 -42458
rect -11666 -42492 -11620 -42458
rect -11586 -42492 -11540 -42458
rect -11506 -42492 -11460 -42458
rect -11426 -42492 -11380 -42458
rect -11346 -42492 -11300 -42458
rect -11266 -42492 -11220 -42458
rect -11186 -42492 -11140 -42458
rect -11106 -42492 -11060 -42458
rect -11026 -42492 -10980 -42458
rect -10946 -42492 -10900 -42458
rect -10866 -42492 -10820 -42458
rect -10786 -42492 -10740 -42458
rect -10706 -42492 -10660 -42458
rect -10626 -42492 -10580 -42458
rect -10546 -42492 -10500 -42458
rect -10466 -42492 -10420 -42458
rect -10386 -42492 -10340 -42458
rect -10306 -42492 -10260 -42458
rect -10226 -42492 -10180 -42458
rect -10146 -42492 -10100 -42458
rect -10066 -42492 -10020 -42458
rect -9986 -42492 -9940 -42458
rect -9906 -42492 -9859 -42458
rect -9825 -42492 -9779 -42458
rect -9745 -42492 -9699 -42458
rect -9665 -42492 -9619 -42458
rect -9585 -42492 -9539 -42458
rect -9505 -42492 -9459 -42458
rect -9425 -42492 -9379 -42458
rect -9345 -42492 -9299 -42458
rect -9265 -42492 -9219 -42458
rect -9185 -42492 -9139 -42458
rect -9105 -42492 -9059 -42458
rect -9025 -42492 -8979 -42458
rect -8945 -42492 -8899 -42458
rect -8865 -42492 -8819 -42458
rect -8785 -42492 -8739 -42458
rect -8705 -42492 -8659 -42458
rect -8625 -42492 -8579 -42458
rect -8545 -42492 -8499 -42458
rect -8465 -42492 -8419 -42458
rect -8385 -42492 -8339 -42458
rect -8305 -42492 -8259 -42458
rect -8225 -42492 -8179 -42458
rect -8145 -42492 -8099 -42458
rect -8065 -42492 -8019 -42458
rect -7985 -42492 -7939 -42458
rect -7905 -42492 -7859 -42458
rect -7825 -42492 -7779 -42458
rect -7745 -42492 -7699 -42458
rect -7665 -42492 -7619 -42458
rect -7585 -42492 -7539 -42458
rect -7505 -42492 -7459 -42458
rect -7425 -42492 -7379 -42458
rect -7345 -42492 -7299 -42458
rect -7265 -42492 -7219 -42458
rect -7185 -42492 -7139 -42458
rect -7105 -42492 -7059 -42458
rect -7025 -42492 -6979 -42458
rect -6945 -42492 -6899 -42458
rect -6865 -42492 -6819 -42458
rect -6785 -42492 -6739 -42458
rect -6705 -42492 -6659 -42458
rect -6625 -42492 -6579 -42458
rect -6545 -42492 -6499 -42458
rect -6465 -42492 -6419 -42458
rect -6385 -42492 -6339 -42458
rect -6305 -42492 -6259 -42458
rect -6225 -42492 -6179 -42458
rect -6145 -42492 -6099 -42458
rect -6065 -42492 -6019 -42458
rect -5985 -42492 -5939 -42458
rect -5905 -42492 -5859 -42458
rect -5825 -42492 -5779 -42458
rect -5745 -42492 -5699 -42458
rect -5665 -42492 -5619 -42458
rect -5585 -42492 -5539 -42458
rect -5505 -42492 -5459 -42458
rect -5425 -42492 -5379 -42458
rect -5345 -42492 -5299 -42458
rect -5265 -42492 -5219 -42458
rect -5185 -42492 -5139 -42458
rect -5105 -42492 -5059 -42458
rect -5025 -42492 -4979 -42458
rect -4945 -42492 -4899 -42458
rect -4865 -42492 -4819 -42458
rect -4785 -42492 -4739 -42458
rect -4705 -42492 -4659 -42458
rect -4625 -42492 -4579 -42458
rect -4545 -42492 -4499 -42458
rect -4465 -42492 -4419 -42458
rect -4385 -42492 -4339 -42458
rect -4305 -42492 -4259 -42458
rect -4225 -42492 -4140 -42458
rect -4106 -42492 -4060 -42458
rect -4026 -42492 -3980 -42458
rect -3946 -42492 -3900 -42458
rect -3866 -42492 -3820 -42458
rect -3786 -42492 -3740 -42458
rect -3706 -42492 -3660 -42458
rect -3626 -42492 -3580 -42458
rect -3546 -42492 -3500 -42458
rect -3466 -42492 -3420 -42458
rect -3386 -42492 -3340 -42458
rect -3306 -42492 -3260 -42458
rect -3226 -42492 -3180 -42458
rect -3146 -42492 -3100 -42458
rect -3066 -42492 -3020 -42458
rect -2986 -42492 -2940 -42458
rect -2906 -42492 -2860 -42458
rect -2826 -42492 -2780 -42458
rect -2746 -42492 -2700 -42458
rect -2666 -42492 -2620 -42458
rect -2586 -42492 -2540 -42458
rect -2506 -42492 -2460 -42458
rect -2426 -42492 -2380 -42458
rect -2346 -42492 -2300 -42458
rect -2266 -42492 -2220 -42458
rect -2186 -42492 -2140 -42458
rect -2106 -42492 -2060 -42458
rect -2026 -42492 -1980 -42458
rect -1946 -42492 -1900 -42458
rect -1866 -42492 -1820 -42458
rect -1786 -42492 -1740 -42458
rect -1706 -42492 -1660 -42458
rect -1626 -42492 -1580 -42458
rect -1546 -42492 -1500 -42458
rect -1466 -42492 -1420 -42458
rect -1386 -42492 -1340 -42458
rect -1306 -42492 -1260 -42458
rect -1226 -42492 -1180 -42458
rect -1146 -42492 -1100 -42458
rect -1066 -42492 -1020 -42458
rect -986 -42492 -940 -42458
rect -906 -42492 -860 -42458
rect -826 -42492 -780 -42458
rect -746 -42492 -700 -42458
rect -666 -42492 -624 -42458
rect -44468 -42515 -624 -42492
rect -10430 -43763 -10170 -43710
rect -10430 -43766 -10377 -43763
rect -10343 -43766 -10257 -43763
rect -10430 -43800 -10379 -43766
rect -10343 -43797 -10259 -43766
rect -10223 -43797 -10170 -43763
rect -10345 -43800 -10259 -43797
rect -10225 -43800 -10170 -43797
rect -10430 -43883 -10170 -43800
rect -10430 -43886 -10377 -43883
rect -10343 -43886 -10257 -43883
rect -10430 -43920 -10379 -43886
rect -10343 -43917 -10259 -43886
rect -10223 -43917 -10170 -43883
rect -9420 -43842 -9354 -42515
rect -6887 -42690 -6853 -42515
rect -8155 -43053 -8075 -43030
rect -8155 -43087 -8132 -43053
rect -8098 -43087 -7859 -43053
rect -8155 -43110 -8075 -43087
rect -8758 -43234 -8558 -43211
rect -8758 -43268 -8735 -43234
rect -8701 -43268 -8615 -43234
rect -8581 -43268 -8558 -43234
rect -8757 -43354 -8557 -43268
rect -8758 -43388 -8735 -43354
rect -8701 -43388 -8615 -43354
rect -8581 -43388 -8558 -43354
rect -8758 -43411 -8558 -43388
rect -8742 -43441 -8582 -43411
rect -8701 -43650 -8621 -43630
rect -8701 -43690 -8681 -43650
rect -8641 -43690 -8621 -43650
rect -8701 -43701 -8621 -43690
rect -9420 -43876 -9404 -43842
rect -9370 -43876 -9354 -43842
rect -9420 -43892 -9354 -43876
rect -10345 -43920 -10259 -43917
rect -10225 -43920 -10170 -43917
rect -10430 -43970 -10170 -43920
rect -8742 -43931 -8582 -43701
rect -8132 -43931 -8098 -43110
rect -5320 -43829 -5254 -43813
rect -5320 -43863 -5304 -43829
rect -5270 -43863 -5254 -43829
rect -5320 -43879 -5254 -43863
rect -3814 -43842 -3748 -42515
rect -1340 -42691 -1306 -42515
rect -2526 -43069 -2314 -43035
rect -2526 -43138 -2492 -43069
rect -2549 -43161 -2469 -43138
rect -2549 -43195 -2526 -43161
rect -2492 -43195 -2469 -43161
rect -3173 -43233 -2973 -43210
rect -2549 -43218 -2469 -43195
rect -3173 -43267 -3150 -43233
rect -3116 -43267 -3030 -43233
rect -2996 -43267 -2973 -43233
rect -3173 -43353 -2973 -43267
rect -3173 -43387 -3150 -43353
rect -3116 -43387 -3030 -43353
rect -2996 -43387 -2973 -43353
rect -3173 -43410 -2973 -43387
rect -3157 -43440 -2997 -43410
rect -3116 -43649 -3036 -43629
rect -3116 -43689 -3096 -43649
rect -3056 -43689 -3036 -43649
rect -3116 -43700 -3036 -43689
rect -3814 -43876 -3798 -43842
rect -3764 -43876 -3748 -43842
rect -3814 -43892 -3748 -43876
rect -3157 -43931 -2997 -43700
rect -2526 -43931 -2492 -43218
rect -9338 -43971 -8098 -43931
rect -9338 -44011 -9298 -43971
rect -9038 -44011 -8998 -43971
rect -8738 -44011 -8698 -43971
rect -8438 -44011 -8398 -43971
rect -8138 -44011 -8098 -43971
rect -7984 -43977 -6450 -43943
rect -7984 -44011 -7950 -43977
rect -7683 -44011 -7649 -43977
rect -7384 -44011 -7350 -43977
rect -7083 -44011 -7049 -43977
rect -6784 -44011 -6750 -43977
rect -6484 -44011 -6450 -43977
rect -5380 -43977 -3846 -43943
rect -5380 -44011 -5346 -43977
rect -5080 -44011 -5046 -43977
rect -4781 -44011 -4747 -43977
rect -4480 -44011 -4446 -43977
rect -4181 -44011 -4147 -43977
rect -3880 -44011 -3846 -43977
rect -3732 -43971 -2492 -43931
rect -3732 -44011 -3692 -43971
rect -3432 -44011 -3392 -43971
rect -3132 -44011 -3092 -43971
rect -2832 -44011 -2792 -43971
rect -2532 -44011 -2492 -43971
rect -9628 -44050 -9548 -44011
rect -9628 -44084 -9605 -44050
rect -9571 -44084 -9548 -44050
rect -9628 -44118 -9548 -44084
rect -9628 -44152 -9605 -44118
rect -9571 -44152 -9548 -44118
rect -9628 -44186 -9548 -44152
rect -9628 -44220 -9605 -44186
rect -9571 -44220 -9548 -44186
rect -9628 -44254 -9548 -44220
rect -9628 -44288 -9605 -44254
rect -9571 -44288 -9548 -44254
rect -9628 -44322 -9548 -44288
rect -9628 -44356 -9605 -44322
rect -9571 -44356 -9548 -44322
rect -9628 -44390 -9548 -44356
rect -9628 -44424 -9605 -44390
rect -9571 -44424 -9548 -44390
rect -9628 -44458 -9548 -44424
rect -9628 -44492 -9605 -44458
rect -9571 -44492 -9548 -44458
rect -9628 -44526 -9548 -44492
rect -9628 -44560 -9605 -44526
rect -9571 -44560 -9548 -44526
rect -9628 -44594 -9548 -44560
rect -9628 -44628 -9605 -44594
rect -9571 -44628 -9548 -44594
rect -9628 -44662 -9548 -44628
rect -9628 -44696 -9605 -44662
rect -9571 -44696 -9548 -44662
rect -9628 -44730 -9548 -44696
rect -9628 -44764 -9605 -44730
rect -9571 -44764 -9548 -44730
rect -9628 -44798 -9548 -44764
rect -9628 -44832 -9605 -44798
rect -9571 -44832 -9548 -44798
rect -10430 -44998 -10170 -44948
rect -10430 -45004 -10378 -44998
rect -10344 -45001 -10258 -44998
rect -10224 -45001 -10170 -44998
rect -10343 -45004 -10258 -45001
rect -10430 -45038 -10379 -45004
rect -10343 -45035 -10259 -45004
rect -10223 -45035 -10170 -45001
rect -10345 -45038 -10259 -45035
rect -10225 -45038 -10170 -45035
rect -10430 -45118 -10170 -45038
rect -10430 -45124 -10378 -45118
rect -10344 -45121 -10258 -45118
rect -10224 -45121 -10170 -45118
rect -10343 -45124 -10258 -45121
rect -10430 -45158 -10379 -45124
rect -10343 -45155 -10259 -45124
rect -10223 -45155 -10170 -45121
rect -10345 -45158 -10259 -45155
rect -10225 -45158 -10170 -45155
rect -10430 -45208 -10170 -45158
rect -9628 -45413 -9548 -44832
rect -9508 -44050 -9428 -44011
rect -9508 -44084 -9485 -44050
rect -9451 -44084 -9428 -44050
rect -9508 -44118 -9428 -44084
rect -9508 -44152 -9485 -44118
rect -9451 -44152 -9428 -44118
rect -9508 -44186 -9428 -44152
rect -9508 -44220 -9485 -44186
rect -9451 -44220 -9428 -44186
rect -9508 -44254 -9428 -44220
rect -9508 -44288 -9485 -44254
rect -9451 -44288 -9428 -44254
rect -9508 -44322 -9428 -44288
rect -9508 -44356 -9485 -44322
rect -9451 -44356 -9428 -44322
rect -9508 -44390 -9428 -44356
rect -9508 -44424 -9485 -44390
rect -9451 -44424 -9428 -44390
rect -9508 -44458 -9428 -44424
rect -9508 -44492 -9485 -44458
rect -9451 -44492 -9428 -44458
rect -9508 -44526 -9428 -44492
rect -9508 -44560 -9485 -44526
rect -9451 -44560 -9428 -44526
rect -9508 -44594 -9428 -44560
rect -9508 -44628 -9485 -44594
rect -9451 -44628 -9428 -44594
rect -9508 -44662 -9428 -44628
rect -9508 -44696 -9485 -44662
rect -9451 -44696 -9428 -44662
rect -9508 -44730 -9428 -44696
rect -9508 -44764 -9485 -44730
rect -9451 -44764 -9428 -44730
rect -9508 -44798 -9428 -44764
rect -9508 -44832 -9485 -44798
rect -9451 -44832 -9428 -44798
rect -9508 -44871 -9428 -44832
rect -9358 -44050 -9278 -44011
rect -9358 -44084 -9335 -44050
rect -9301 -44084 -9278 -44050
rect -9358 -44118 -9278 -44084
rect -9358 -44152 -9335 -44118
rect -9301 -44152 -9278 -44118
rect -9358 -44186 -9278 -44152
rect -9358 -44220 -9335 -44186
rect -9301 -44220 -9278 -44186
rect -9358 -44254 -9278 -44220
rect -9358 -44288 -9335 -44254
rect -9301 -44288 -9278 -44254
rect -9358 -44322 -9278 -44288
rect -9358 -44356 -9335 -44322
rect -9301 -44356 -9278 -44322
rect -9358 -44390 -9278 -44356
rect -9358 -44424 -9335 -44390
rect -9301 -44424 -9278 -44390
rect -9358 -44458 -9278 -44424
rect -9358 -44492 -9335 -44458
rect -9301 -44492 -9278 -44458
rect -9358 -44526 -9278 -44492
rect -9358 -44560 -9335 -44526
rect -9301 -44560 -9278 -44526
rect -9358 -44594 -9278 -44560
rect -9358 -44628 -9335 -44594
rect -9301 -44628 -9278 -44594
rect -9358 -44662 -9278 -44628
rect -9358 -44696 -9335 -44662
rect -9301 -44696 -9278 -44662
rect -9358 -44730 -9278 -44696
rect -9358 -44764 -9335 -44730
rect -9301 -44764 -9278 -44730
rect -9358 -44798 -9278 -44764
rect -9358 -44832 -9335 -44798
rect -9301 -44832 -9278 -44798
rect -9358 -44871 -9278 -44832
rect -9208 -44050 -9128 -44011
rect -9208 -44084 -9185 -44050
rect -9151 -44084 -9128 -44050
rect -9208 -44118 -9128 -44084
rect -9208 -44152 -9185 -44118
rect -9151 -44152 -9128 -44118
rect -9208 -44186 -9128 -44152
rect -9208 -44220 -9185 -44186
rect -9151 -44220 -9128 -44186
rect -9208 -44254 -9128 -44220
rect -9208 -44288 -9185 -44254
rect -9151 -44288 -9128 -44254
rect -9208 -44322 -9128 -44288
rect -9208 -44356 -9185 -44322
rect -9151 -44356 -9128 -44322
rect -9208 -44390 -9128 -44356
rect -9208 -44424 -9185 -44390
rect -9151 -44424 -9128 -44390
rect -9208 -44458 -9128 -44424
rect -9208 -44492 -9185 -44458
rect -9151 -44492 -9128 -44458
rect -9208 -44526 -9128 -44492
rect -9208 -44560 -9185 -44526
rect -9151 -44560 -9128 -44526
rect -9208 -44594 -9128 -44560
rect -9208 -44628 -9185 -44594
rect -9151 -44628 -9128 -44594
rect -9208 -44662 -9128 -44628
rect -9208 -44696 -9185 -44662
rect -9151 -44696 -9128 -44662
rect -9208 -44730 -9128 -44696
rect -9208 -44764 -9185 -44730
rect -9151 -44764 -9128 -44730
rect -9208 -44798 -9128 -44764
rect -9208 -44832 -9185 -44798
rect -9151 -44832 -9128 -44798
rect -9208 -44871 -9128 -44832
rect -9058 -44050 -8978 -44011
rect -9058 -44084 -9035 -44050
rect -9001 -44084 -8978 -44050
rect -9058 -44118 -8978 -44084
rect -9058 -44152 -9035 -44118
rect -9001 -44152 -8978 -44118
rect -9058 -44186 -8978 -44152
rect -9058 -44220 -9035 -44186
rect -9001 -44220 -8978 -44186
rect -9058 -44254 -8978 -44220
rect -9058 -44288 -9035 -44254
rect -9001 -44288 -8978 -44254
rect -9058 -44322 -8978 -44288
rect -9058 -44356 -9035 -44322
rect -9001 -44356 -8978 -44322
rect -9058 -44390 -8978 -44356
rect -9058 -44424 -9035 -44390
rect -9001 -44424 -8978 -44390
rect -9058 -44458 -8978 -44424
rect -9058 -44492 -9035 -44458
rect -9001 -44492 -8978 -44458
rect -9058 -44526 -8978 -44492
rect -9058 -44560 -9035 -44526
rect -9001 -44560 -8978 -44526
rect -9058 -44594 -8978 -44560
rect -9058 -44628 -9035 -44594
rect -9001 -44628 -8978 -44594
rect -9058 -44662 -8978 -44628
rect -9058 -44696 -9035 -44662
rect -9001 -44696 -8978 -44662
rect -9058 -44730 -8978 -44696
rect -9058 -44764 -9035 -44730
rect -9001 -44764 -8978 -44730
rect -9058 -44798 -8978 -44764
rect -9058 -44832 -9035 -44798
rect -9001 -44832 -8978 -44798
rect -9058 -44871 -8978 -44832
rect -8908 -44050 -8828 -44011
rect -8908 -44084 -8885 -44050
rect -8851 -44084 -8828 -44050
rect -8908 -44118 -8828 -44084
rect -8908 -44152 -8885 -44118
rect -8851 -44152 -8828 -44118
rect -8908 -44186 -8828 -44152
rect -8908 -44220 -8885 -44186
rect -8851 -44220 -8828 -44186
rect -8908 -44254 -8828 -44220
rect -8908 -44288 -8885 -44254
rect -8851 -44288 -8828 -44254
rect -8908 -44322 -8828 -44288
rect -8908 -44356 -8885 -44322
rect -8851 -44356 -8828 -44322
rect -8908 -44390 -8828 -44356
rect -8908 -44424 -8885 -44390
rect -8851 -44424 -8828 -44390
rect -8908 -44458 -8828 -44424
rect -8908 -44492 -8885 -44458
rect -8851 -44492 -8828 -44458
rect -8908 -44526 -8828 -44492
rect -8908 -44560 -8885 -44526
rect -8851 -44560 -8828 -44526
rect -8908 -44594 -8828 -44560
rect -8908 -44628 -8885 -44594
rect -8851 -44628 -8828 -44594
rect -8908 -44662 -8828 -44628
rect -8908 -44696 -8885 -44662
rect -8851 -44696 -8828 -44662
rect -8908 -44730 -8828 -44696
rect -8908 -44764 -8885 -44730
rect -8851 -44764 -8828 -44730
rect -8908 -44798 -8828 -44764
rect -8908 -44832 -8885 -44798
rect -8851 -44832 -8828 -44798
rect -8908 -44871 -8828 -44832
rect -8758 -44050 -8678 -44011
rect -8758 -44084 -8735 -44050
rect -8701 -44084 -8678 -44050
rect -8758 -44118 -8678 -44084
rect -8758 -44152 -8735 -44118
rect -8701 -44152 -8678 -44118
rect -8758 -44186 -8678 -44152
rect -8758 -44220 -8735 -44186
rect -8701 -44220 -8678 -44186
rect -8758 -44254 -8678 -44220
rect -8758 -44288 -8735 -44254
rect -8701 -44288 -8678 -44254
rect -8758 -44322 -8678 -44288
rect -8758 -44356 -8735 -44322
rect -8701 -44356 -8678 -44322
rect -8758 -44390 -8678 -44356
rect -8758 -44424 -8735 -44390
rect -8701 -44424 -8678 -44390
rect -8758 -44458 -8678 -44424
rect -8758 -44492 -8735 -44458
rect -8701 -44492 -8678 -44458
rect -8758 -44526 -8678 -44492
rect -8758 -44560 -8735 -44526
rect -8701 -44560 -8678 -44526
rect -8758 -44594 -8678 -44560
rect -8758 -44628 -8735 -44594
rect -8701 -44628 -8678 -44594
rect -8758 -44662 -8678 -44628
rect -8758 -44696 -8735 -44662
rect -8701 -44696 -8678 -44662
rect -8758 -44730 -8678 -44696
rect -8758 -44764 -8735 -44730
rect -8701 -44764 -8678 -44730
rect -8758 -44798 -8678 -44764
rect -8758 -44832 -8735 -44798
rect -8701 -44832 -8678 -44798
rect -8758 -44871 -8678 -44832
rect -8608 -44050 -8528 -44011
rect -8608 -44084 -8585 -44050
rect -8551 -44084 -8528 -44050
rect -8608 -44118 -8528 -44084
rect -8608 -44152 -8585 -44118
rect -8551 -44152 -8528 -44118
rect -8608 -44186 -8528 -44152
rect -8608 -44220 -8585 -44186
rect -8551 -44220 -8528 -44186
rect -8608 -44254 -8528 -44220
rect -8608 -44288 -8585 -44254
rect -8551 -44288 -8528 -44254
rect -8608 -44322 -8528 -44288
rect -8608 -44356 -8585 -44322
rect -8551 -44356 -8528 -44322
rect -8608 -44390 -8528 -44356
rect -8608 -44424 -8585 -44390
rect -8551 -44424 -8528 -44390
rect -8608 -44458 -8528 -44424
rect -8608 -44492 -8585 -44458
rect -8551 -44492 -8528 -44458
rect -8608 -44526 -8528 -44492
rect -8608 -44560 -8585 -44526
rect -8551 -44560 -8528 -44526
rect -8608 -44594 -8528 -44560
rect -8608 -44628 -8585 -44594
rect -8551 -44628 -8528 -44594
rect -8608 -44662 -8528 -44628
rect -8608 -44696 -8585 -44662
rect -8551 -44696 -8528 -44662
rect -8608 -44730 -8528 -44696
rect -8608 -44764 -8585 -44730
rect -8551 -44764 -8528 -44730
rect -8608 -44798 -8528 -44764
rect -8608 -44832 -8585 -44798
rect -8551 -44832 -8528 -44798
rect -8608 -44871 -8528 -44832
rect -8458 -44050 -8378 -44011
rect -8458 -44084 -8435 -44050
rect -8401 -44084 -8378 -44050
rect -8458 -44118 -8378 -44084
rect -8458 -44152 -8435 -44118
rect -8401 -44152 -8378 -44118
rect -8458 -44186 -8378 -44152
rect -8458 -44220 -8435 -44186
rect -8401 -44220 -8378 -44186
rect -8458 -44254 -8378 -44220
rect -8458 -44288 -8435 -44254
rect -8401 -44288 -8378 -44254
rect -8458 -44322 -8378 -44288
rect -8458 -44356 -8435 -44322
rect -8401 -44356 -8378 -44322
rect -8458 -44390 -8378 -44356
rect -8458 -44424 -8435 -44390
rect -8401 -44424 -8378 -44390
rect -8458 -44458 -8378 -44424
rect -8458 -44492 -8435 -44458
rect -8401 -44492 -8378 -44458
rect -8458 -44526 -8378 -44492
rect -8458 -44560 -8435 -44526
rect -8401 -44560 -8378 -44526
rect -8458 -44594 -8378 -44560
rect -8458 -44628 -8435 -44594
rect -8401 -44628 -8378 -44594
rect -8458 -44662 -8378 -44628
rect -8458 -44696 -8435 -44662
rect -8401 -44696 -8378 -44662
rect -8458 -44730 -8378 -44696
rect -8458 -44764 -8435 -44730
rect -8401 -44764 -8378 -44730
rect -8458 -44798 -8378 -44764
rect -8458 -44832 -8435 -44798
rect -8401 -44832 -8378 -44798
rect -8458 -44871 -8378 -44832
rect -8308 -44050 -8228 -44011
rect -8308 -44084 -8285 -44050
rect -8251 -44084 -8228 -44050
rect -8308 -44118 -8228 -44084
rect -8308 -44152 -8285 -44118
rect -8251 -44152 -8228 -44118
rect -8308 -44186 -8228 -44152
rect -8308 -44220 -8285 -44186
rect -8251 -44220 -8228 -44186
rect -8308 -44254 -8228 -44220
rect -8308 -44288 -8285 -44254
rect -8251 -44288 -8228 -44254
rect -8308 -44322 -8228 -44288
rect -8308 -44356 -8285 -44322
rect -8251 -44356 -8228 -44322
rect -8308 -44390 -8228 -44356
rect -8308 -44424 -8285 -44390
rect -8251 -44424 -8228 -44390
rect -8308 -44458 -8228 -44424
rect -8308 -44492 -8285 -44458
rect -8251 -44492 -8228 -44458
rect -8308 -44526 -8228 -44492
rect -8308 -44560 -8285 -44526
rect -8251 -44560 -8228 -44526
rect -8308 -44594 -8228 -44560
rect -8308 -44628 -8285 -44594
rect -8251 -44628 -8228 -44594
rect -8308 -44662 -8228 -44628
rect -8308 -44696 -8285 -44662
rect -8251 -44696 -8228 -44662
rect -8308 -44730 -8228 -44696
rect -8308 -44764 -8285 -44730
rect -8251 -44764 -8228 -44730
rect -8308 -44798 -8228 -44764
rect -8308 -44832 -8285 -44798
rect -8251 -44832 -8228 -44798
rect -8308 -44871 -8228 -44832
rect -8158 -44060 -8078 -44011
rect -8158 -44094 -8135 -44060
rect -8101 -44094 -8078 -44060
rect -8158 -44128 -8078 -44094
rect -8158 -44162 -8135 -44128
rect -8101 -44162 -8078 -44128
rect -8158 -44196 -8078 -44162
rect -8158 -44230 -8135 -44196
rect -8101 -44230 -8078 -44196
rect -8158 -44264 -8078 -44230
rect -8158 -44298 -8135 -44264
rect -8101 -44298 -8078 -44264
rect -8158 -44332 -8078 -44298
rect -8158 -44366 -8135 -44332
rect -8101 -44366 -8078 -44332
rect -8158 -44400 -8078 -44366
rect -8158 -44434 -8135 -44400
rect -8101 -44434 -8078 -44400
rect -8158 -44468 -8078 -44434
rect -8158 -44502 -8135 -44468
rect -8101 -44502 -8078 -44468
rect -8158 -44536 -8078 -44502
rect -8158 -44570 -8135 -44536
rect -8101 -44570 -8078 -44536
rect -8158 -44604 -8078 -44570
rect -8158 -44638 -8135 -44604
rect -8101 -44638 -8078 -44604
rect -8158 -44672 -8078 -44638
rect -8158 -44706 -8135 -44672
rect -8101 -44706 -8078 -44672
rect -8158 -44740 -8078 -44706
rect -8158 -44774 -8135 -44740
rect -8101 -44774 -8078 -44740
rect -8158 -44808 -8078 -44774
rect -8158 -44842 -8135 -44808
rect -8101 -44842 -8078 -44808
rect -8158 -44871 -8078 -44842
rect -8008 -44050 -7928 -44011
rect -8008 -44084 -7985 -44050
rect -7951 -44084 -7928 -44050
rect -8008 -44118 -7928 -44084
rect -8008 -44152 -7985 -44118
rect -7951 -44152 -7928 -44118
rect -8008 -44186 -7928 -44152
rect -8008 -44220 -7985 -44186
rect -7951 -44220 -7928 -44186
rect -8008 -44254 -7928 -44220
rect -8008 -44288 -7985 -44254
rect -7951 -44288 -7928 -44254
rect -8008 -44322 -7928 -44288
rect -8008 -44356 -7985 -44322
rect -7951 -44356 -7928 -44322
rect -8008 -44390 -7928 -44356
rect -8008 -44424 -7985 -44390
rect -7951 -44424 -7928 -44390
rect -8008 -44458 -7928 -44424
rect -8008 -44492 -7985 -44458
rect -7951 -44492 -7928 -44458
rect -8008 -44526 -7928 -44492
rect -8008 -44560 -7985 -44526
rect -7951 -44560 -7928 -44526
rect -8008 -44594 -7928 -44560
rect -8008 -44628 -7985 -44594
rect -7951 -44628 -7928 -44594
rect -8008 -44662 -7928 -44628
rect -8008 -44696 -7985 -44662
rect -7951 -44696 -7928 -44662
rect -8008 -44730 -7928 -44696
rect -8008 -44764 -7985 -44730
rect -7951 -44764 -7928 -44730
rect -8008 -44798 -7928 -44764
rect -8008 -44832 -7985 -44798
rect -7951 -44832 -7928 -44798
rect -8008 -44871 -7928 -44832
rect -7858 -44050 -7778 -44011
rect -7858 -44084 -7835 -44050
rect -7801 -44084 -7778 -44050
rect -7858 -44118 -7778 -44084
rect -7858 -44152 -7835 -44118
rect -7801 -44152 -7778 -44118
rect -7858 -44186 -7778 -44152
rect -7858 -44220 -7835 -44186
rect -7801 -44220 -7778 -44186
rect -7858 -44254 -7778 -44220
rect -7858 -44288 -7835 -44254
rect -7801 -44288 -7778 -44254
rect -7858 -44322 -7778 -44288
rect -7858 -44356 -7835 -44322
rect -7801 -44356 -7778 -44322
rect -7858 -44390 -7778 -44356
rect -7858 -44424 -7835 -44390
rect -7801 -44424 -7778 -44390
rect -7858 -44458 -7778 -44424
rect -7858 -44492 -7835 -44458
rect -7801 -44492 -7778 -44458
rect -7858 -44526 -7778 -44492
rect -7858 -44560 -7835 -44526
rect -7801 -44560 -7778 -44526
rect -7858 -44594 -7778 -44560
rect -7858 -44628 -7835 -44594
rect -7801 -44628 -7778 -44594
rect -7858 -44662 -7778 -44628
rect -7858 -44696 -7835 -44662
rect -7801 -44696 -7778 -44662
rect -7858 -44730 -7778 -44696
rect -7858 -44764 -7835 -44730
rect -7801 -44764 -7778 -44730
rect -7858 -44798 -7778 -44764
rect -7858 -44832 -7835 -44798
rect -7801 -44832 -7778 -44798
rect -7858 -44871 -7778 -44832
rect -7708 -44050 -7628 -44011
rect -7708 -44084 -7685 -44050
rect -7651 -44084 -7628 -44050
rect -7708 -44118 -7628 -44084
rect -7708 -44152 -7685 -44118
rect -7651 -44152 -7628 -44118
rect -7708 -44186 -7628 -44152
rect -7708 -44220 -7685 -44186
rect -7651 -44220 -7628 -44186
rect -7708 -44254 -7628 -44220
rect -7708 -44288 -7685 -44254
rect -7651 -44288 -7628 -44254
rect -7708 -44322 -7628 -44288
rect -7708 -44356 -7685 -44322
rect -7651 -44356 -7628 -44322
rect -7708 -44390 -7628 -44356
rect -7708 -44424 -7685 -44390
rect -7651 -44424 -7628 -44390
rect -7708 -44458 -7628 -44424
rect -7708 -44492 -7685 -44458
rect -7651 -44492 -7628 -44458
rect -7708 -44526 -7628 -44492
rect -7708 -44560 -7685 -44526
rect -7651 -44560 -7628 -44526
rect -7708 -44594 -7628 -44560
rect -7708 -44628 -7685 -44594
rect -7651 -44628 -7628 -44594
rect -7708 -44662 -7628 -44628
rect -7708 -44696 -7685 -44662
rect -7651 -44696 -7628 -44662
rect -7708 -44730 -7628 -44696
rect -7708 -44764 -7685 -44730
rect -7651 -44764 -7628 -44730
rect -7708 -44798 -7628 -44764
rect -7708 -44832 -7685 -44798
rect -7651 -44832 -7628 -44798
rect -7708 -44871 -7628 -44832
rect -7558 -44050 -7478 -44011
rect -7558 -44084 -7535 -44050
rect -7501 -44084 -7478 -44050
rect -7558 -44118 -7478 -44084
rect -7558 -44152 -7535 -44118
rect -7501 -44152 -7478 -44118
rect -7558 -44186 -7478 -44152
rect -7558 -44220 -7535 -44186
rect -7501 -44220 -7478 -44186
rect -7558 -44254 -7478 -44220
rect -7558 -44288 -7535 -44254
rect -7501 -44288 -7478 -44254
rect -7558 -44322 -7478 -44288
rect -7558 -44356 -7535 -44322
rect -7501 -44356 -7478 -44322
rect -7558 -44390 -7478 -44356
rect -7558 -44424 -7535 -44390
rect -7501 -44424 -7478 -44390
rect -7558 -44458 -7478 -44424
rect -7558 -44492 -7535 -44458
rect -7501 -44492 -7478 -44458
rect -7558 -44526 -7478 -44492
rect -7558 -44560 -7535 -44526
rect -7501 -44560 -7478 -44526
rect -7558 -44594 -7478 -44560
rect -7558 -44628 -7535 -44594
rect -7501 -44628 -7478 -44594
rect -7558 -44662 -7478 -44628
rect -7558 -44696 -7535 -44662
rect -7501 -44696 -7478 -44662
rect -7558 -44730 -7478 -44696
rect -7558 -44764 -7535 -44730
rect -7501 -44764 -7478 -44730
rect -7558 -44798 -7478 -44764
rect -7558 -44832 -7535 -44798
rect -7501 -44832 -7478 -44798
rect -7558 -44871 -7478 -44832
rect -7408 -44050 -7328 -44011
rect -7408 -44084 -7385 -44050
rect -7351 -44084 -7328 -44050
rect -7408 -44118 -7328 -44084
rect -7408 -44152 -7385 -44118
rect -7351 -44152 -7328 -44118
rect -7408 -44186 -7328 -44152
rect -7408 -44220 -7385 -44186
rect -7351 -44220 -7328 -44186
rect -7408 -44254 -7328 -44220
rect -7408 -44288 -7385 -44254
rect -7351 -44288 -7328 -44254
rect -7408 -44322 -7328 -44288
rect -7408 -44356 -7385 -44322
rect -7351 -44356 -7328 -44322
rect -7408 -44390 -7328 -44356
rect -7408 -44424 -7385 -44390
rect -7351 -44424 -7328 -44390
rect -7408 -44458 -7328 -44424
rect -7408 -44492 -7385 -44458
rect -7351 -44492 -7328 -44458
rect -7408 -44526 -7328 -44492
rect -7408 -44560 -7385 -44526
rect -7351 -44560 -7328 -44526
rect -7408 -44594 -7328 -44560
rect -7408 -44628 -7385 -44594
rect -7351 -44628 -7328 -44594
rect -7408 -44662 -7328 -44628
rect -7408 -44696 -7385 -44662
rect -7351 -44696 -7328 -44662
rect -7408 -44730 -7328 -44696
rect -7408 -44764 -7385 -44730
rect -7351 -44764 -7328 -44730
rect -7408 -44798 -7328 -44764
rect -7408 -44832 -7385 -44798
rect -7351 -44832 -7328 -44798
rect -7408 -44871 -7328 -44832
rect -7258 -44050 -7178 -44011
rect -7258 -44084 -7235 -44050
rect -7201 -44084 -7178 -44050
rect -7258 -44118 -7178 -44084
rect -7258 -44152 -7235 -44118
rect -7201 -44152 -7178 -44118
rect -7258 -44186 -7178 -44152
rect -7258 -44220 -7235 -44186
rect -7201 -44220 -7178 -44186
rect -7258 -44254 -7178 -44220
rect -7258 -44288 -7235 -44254
rect -7201 -44288 -7178 -44254
rect -7258 -44322 -7178 -44288
rect -7258 -44356 -7235 -44322
rect -7201 -44356 -7178 -44322
rect -7258 -44390 -7178 -44356
rect -7258 -44424 -7235 -44390
rect -7201 -44424 -7178 -44390
rect -7258 -44458 -7178 -44424
rect -7258 -44492 -7235 -44458
rect -7201 -44492 -7178 -44458
rect -7258 -44526 -7178 -44492
rect -7258 -44560 -7235 -44526
rect -7201 -44560 -7178 -44526
rect -7258 -44594 -7178 -44560
rect -7258 -44628 -7235 -44594
rect -7201 -44628 -7178 -44594
rect -7258 -44662 -7178 -44628
rect -7258 -44696 -7235 -44662
rect -7201 -44696 -7178 -44662
rect -7258 -44730 -7178 -44696
rect -7258 -44764 -7235 -44730
rect -7201 -44764 -7178 -44730
rect -7258 -44798 -7178 -44764
rect -7258 -44832 -7235 -44798
rect -7201 -44832 -7178 -44798
rect -7258 -44871 -7178 -44832
rect -7108 -44050 -7028 -44011
rect -7108 -44084 -7085 -44050
rect -7051 -44084 -7028 -44050
rect -7108 -44118 -7028 -44084
rect -7108 -44152 -7085 -44118
rect -7051 -44152 -7028 -44118
rect -7108 -44186 -7028 -44152
rect -7108 -44220 -7085 -44186
rect -7051 -44220 -7028 -44186
rect -7108 -44254 -7028 -44220
rect -7108 -44288 -7085 -44254
rect -7051 -44288 -7028 -44254
rect -7108 -44322 -7028 -44288
rect -7108 -44356 -7085 -44322
rect -7051 -44356 -7028 -44322
rect -7108 -44390 -7028 -44356
rect -7108 -44424 -7085 -44390
rect -7051 -44424 -7028 -44390
rect -7108 -44458 -7028 -44424
rect -7108 -44492 -7085 -44458
rect -7051 -44492 -7028 -44458
rect -7108 -44526 -7028 -44492
rect -7108 -44560 -7085 -44526
rect -7051 -44560 -7028 -44526
rect -7108 -44594 -7028 -44560
rect -7108 -44628 -7085 -44594
rect -7051 -44628 -7028 -44594
rect -7108 -44662 -7028 -44628
rect -7108 -44696 -7085 -44662
rect -7051 -44696 -7028 -44662
rect -7108 -44730 -7028 -44696
rect -7108 -44764 -7085 -44730
rect -7051 -44764 -7028 -44730
rect -7108 -44798 -7028 -44764
rect -7108 -44832 -7085 -44798
rect -7051 -44832 -7028 -44798
rect -7108 -44871 -7028 -44832
rect -6958 -44050 -6878 -44011
rect -6958 -44084 -6935 -44050
rect -6901 -44084 -6878 -44050
rect -6958 -44118 -6878 -44084
rect -6958 -44152 -6935 -44118
rect -6901 -44152 -6878 -44118
rect -6958 -44186 -6878 -44152
rect -6958 -44220 -6935 -44186
rect -6901 -44220 -6878 -44186
rect -6958 -44254 -6878 -44220
rect -6958 -44288 -6935 -44254
rect -6901 -44288 -6878 -44254
rect -6958 -44322 -6878 -44288
rect -6958 -44356 -6935 -44322
rect -6901 -44356 -6878 -44322
rect -6958 -44390 -6878 -44356
rect -6958 -44424 -6935 -44390
rect -6901 -44424 -6878 -44390
rect -6958 -44458 -6878 -44424
rect -6958 -44492 -6935 -44458
rect -6901 -44492 -6878 -44458
rect -6958 -44526 -6878 -44492
rect -6958 -44560 -6935 -44526
rect -6901 -44560 -6878 -44526
rect -6958 -44594 -6878 -44560
rect -6958 -44628 -6935 -44594
rect -6901 -44628 -6878 -44594
rect -6958 -44662 -6878 -44628
rect -6958 -44696 -6935 -44662
rect -6901 -44696 -6878 -44662
rect -6958 -44730 -6878 -44696
rect -6958 -44764 -6935 -44730
rect -6901 -44764 -6878 -44730
rect -6958 -44798 -6878 -44764
rect -6958 -44832 -6935 -44798
rect -6901 -44832 -6878 -44798
rect -6958 -44871 -6878 -44832
rect -6808 -44050 -6728 -44011
rect -6808 -44084 -6785 -44050
rect -6751 -44084 -6728 -44050
rect -6808 -44118 -6728 -44084
rect -6808 -44152 -6785 -44118
rect -6751 -44152 -6728 -44118
rect -6808 -44186 -6728 -44152
rect -6808 -44220 -6785 -44186
rect -6751 -44220 -6728 -44186
rect -6808 -44254 -6728 -44220
rect -6808 -44288 -6785 -44254
rect -6751 -44288 -6728 -44254
rect -6808 -44322 -6728 -44288
rect -6808 -44356 -6785 -44322
rect -6751 -44356 -6728 -44322
rect -6808 -44390 -6728 -44356
rect -6808 -44424 -6785 -44390
rect -6751 -44424 -6728 -44390
rect -6808 -44458 -6728 -44424
rect -6808 -44492 -6785 -44458
rect -6751 -44492 -6728 -44458
rect -6808 -44526 -6728 -44492
rect -6808 -44560 -6785 -44526
rect -6751 -44560 -6728 -44526
rect -6808 -44594 -6728 -44560
rect -6808 -44628 -6785 -44594
rect -6751 -44628 -6728 -44594
rect -6808 -44662 -6728 -44628
rect -6808 -44696 -6785 -44662
rect -6751 -44696 -6728 -44662
rect -6808 -44730 -6728 -44696
rect -6808 -44764 -6785 -44730
rect -6751 -44764 -6728 -44730
rect -6808 -44798 -6728 -44764
rect -6808 -44832 -6785 -44798
rect -6751 -44832 -6728 -44798
rect -6808 -44871 -6728 -44832
rect -6658 -44060 -6578 -44011
rect -6658 -44094 -6635 -44060
rect -6601 -44094 -6578 -44060
rect -6658 -44128 -6578 -44094
rect -6658 -44162 -6635 -44128
rect -6601 -44162 -6578 -44128
rect -6658 -44196 -6578 -44162
rect -6658 -44230 -6635 -44196
rect -6601 -44230 -6578 -44196
rect -6658 -44264 -6578 -44230
rect -6658 -44298 -6635 -44264
rect -6601 -44298 -6578 -44264
rect -6658 -44332 -6578 -44298
rect -6658 -44366 -6635 -44332
rect -6601 -44366 -6578 -44332
rect -6658 -44400 -6578 -44366
rect -6658 -44434 -6635 -44400
rect -6601 -44434 -6578 -44400
rect -6658 -44468 -6578 -44434
rect -6658 -44502 -6635 -44468
rect -6601 -44502 -6578 -44468
rect -6658 -44536 -6578 -44502
rect -6658 -44570 -6635 -44536
rect -6601 -44570 -6578 -44536
rect -6658 -44604 -6578 -44570
rect -6658 -44638 -6635 -44604
rect -6601 -44638 -6578 -44604
rect -6658 -44672 -6578 -44638
rect -6658 -44706 -6635 -44672
rect -6601 -44706 -6578 -44672
rect -6658 -44740 -6578 -44706
rect -6658 -44774 -6635 -44740
rect -6601 -44774 -6578 -44740
rect -6658 -44808 -6578 -44774
rect -6658 -44842 -6635 -44808
rect -6601 -44842 -6578 -44808
rect -6658 -44871 -6578 -44842
rect -6508 -44050 -6428 -44011
rect -6508 -44084 -6485 -44050
rect -6451 -44084 -6428 -44050
rect -6508 -44118 -6428 -44084
rect -6508 -44152 -6485 -44118
rect -6451 -44152 -6428 -44118
rect -6508 -44186 -6428 -44152
rect -6508 -44220 -6485 -44186
rect -6451 -44220 -6428 -44186
rect -6508 -44254 -6428 -44220
rect -6508 -44288 -6485 -44254
rect -6451 -44288 -6428 -44254
rect -6508 -44322 -6428 -44288
rect -6508 -44356 -6485 -44322
rect -6451 -44356 -6428 -44322
rect -6508 -44390 -6428 -44356
rect -6508 -44424 -6485 -44390
rect -6451 -44424 -6428 -44390
rect -6508 -44458 -6428 -44424
rect -6508 -44492 -6485 -44458
rect -6451 -44492 -6428 -44458
rect -6508 -44526 -6428 -44492
rect -6508 -44560 -6485 -44526
rect -6451 -44560 -6428 -44526
rect -6508 -44594 -6428 -44560
rect -6508 -44628 -6485 -44594
rect -6451 -44628 -6428 -44594
rect -6508 -44662 -6428 -44628
rect -6508 -44696 -6485 -44662
rect -6451 -44696 -6428 -44662
rect -6508 -44730 -6428 -44696
rect -6508 -44764 -6485 -44730
rect -6451 -44764 -6428 -44730
rect -6508 -44798 -6428 -44764
rect -6508 -44832 -6485 -44798
rect -6451 -44832 -6428 -44798
rect -6508 -44871 -6428 -44832
rect -6388 -44050 -6308 -44011
rect -6388 -44084 -6365 -44050
rect -6331 -44084 -6308 -44050
rect -6388 -44118 -6308 -44084
rect -6388 -44152 -6365 -44118
rect -6331 -44152 -6308 -44118
rect -6388 -44186 -6308 -44152
rect -6388 -44220 -6365 -44186
rect -6331 -44220 -6308 -44186
rect -6388 -44254 -6308 -44220
rect -6388 -44288 -6365 -44254
rect -6331 -44288 -6308 -44254
rect -6388 -44322 -6308 -44288
rect -6388 -44356 -6365 -44322
rect -6331 -44356 -6308 -44322
rect -6388 -44390 -6308 -44356
rect -6388 -44424 -6365 -44390
rect -6331 -44424 -6308 -44390
rect -6388 -44458 -6308 -44424
rect -6388 -44492 -6365 -44458
rect -6331 -44492 -6308 -44458
rect -6388 -44526 -6308 -44492
rect -6388 -44560 -6365 -44526
rect -6331 -44560 -6308 -44526
rect -6388 -44594 -6308 -44560
rect -6388 -44628 -6365 -44594
rect -6331 -44628 -6308 -44594
rect -6388 -44662 -6308 -44628
rect -6388 -44696 -6365 -44662
rect -6331 -44696 -6308 -44662
rect -6388 -44730 -6308 -44696
rect -6388 -44764 -6365 -44730
rect -6331 -44764 -6308 -44730
rect -6388 -44798 -6308 -44764
rect -6388 -44832 -6365 -44798
rect -6331 -44832 -6308 -44798
rect -9488 -44911 -9448 -44871
rect -9188 -44911 -9148 -44871
rect -8888 -44911 -8848 -44871
rect -8588 -44911 -8548 -44871
rect -8288 -44911 -8248 -44871
rect -7988 -44911 -7948 -44871
rect -9488 -44951 -7948 -44911
rect -7838 -44911 -7798 -44871
rect -7539 -44911 -7499 -44871
rect -7239 -44911 -7199 -44871
rect -6939 -44911 -6899 -44871
rect -6638 -44911 -6598 -44871
rect -7838 -44951 -6598 -44911
rect -7926 -45059 -7860 -45043
rect -7926 -45093 -7910 -45059
rect -7876 -45093 -7860 -45059
rect -7926 -45109 -7860 -45093
rect -6858 -45090 -6598 -44951
rect -6858 -45096 -6807 -45090
rect -6773 -45093 -6687 -45090
rect -6653 -45093 -6598 -45090
rect -6772 -45096 -6687 -45093
rect -6858 -45130 -6808 -45096
rect -6772 -45127 -6688 -45096
rect -6652 -45127 -6598 -45093
rect -6773 -45130 -6688 -45127
rect -6858 -45131 -6807 -45130
rect -6773 -45131 -6687 -45130
rect -6653 -45131 -6598 -45127
rect -6858 -45210 -6598 -45131
rect -6858 -45216 -6807 -45210
rect -6773 -45213 -6687 -45210
rect -6653 -45213 -6598 -45210
rect -6772 -45216 -6687 -45213
rect -6858 -45250 -6808 -45216
rect -6772 -45247 -6688 -45216
rect -6652 -45247 -6598 -45213
rect -6773 -45250 -6688 -45247
rect -6858 -45251 -6807 -45250
rect -6773 -45251 -6687 -45250
rect -6653 -45251 -6598 -45247
rect -6858 -45303 -6598 -45251
rect -6388 -45413 -6308 -44832
rect -5522 -44050 -5442 -44011
rect -5522 -44084 -5499 -44050
rect -5465 -44084 -5442 -44050
rect -5522 -44118 -5442 -44084
rect -5522 -44152 -5499 -44118
rect -5465 -44152 -5442 -44118
rect -5522 -44186 -5442 -44152
rect -5522 -44220 -5499 -44186
rect -5465 -44220 -5442 -44186
rect -5522 -44254 -5442 -44220
rect -5522 -44288 -5499 -44254
rect -5465 -44288 -5442 -44254
rect -5522 -44322 -5442 -44288
rect -5522 -44356 -5499 -44322
rect -5465 -44356 -5442 -44322
rect -5522 -44390 -5442 -44356
rect -5522 -44424 -5499 -44390
rect -5465 -44424 -5442 -44390
rect -5522 -44458 -5442 -44424
rect -5522 -44492 -5499 -44458
rect -5465 -44492 -5442 -44458
rect -5522 -44526 -5442 -44492
rect -5522 -44560 -5499 -44526
rect -5465 -44560 -5442 -44526
rect -5522 -44594 -5442 -44560
rect -5522 -44628 -5499 -44594
rect -5465 -44628 -5442 -44594
rect -5522 -44662 -5442 -44628
rect -5522 -44696 -5499 -44662
rect -5465 -44696 -5442 -44662
rect -5522 -44730 -5442 -44696
rect -5522 -44764 -5499 -44730
rect -5465 -44764 -5442 -44730
rect -5522 -44798 -5442 -44764
rect -5522 -44832 -5499 -44798
rect -5465 -44832 -5442 -44798
rect -5522 -45413 -5442 -44832
rect -5402 -44050 -5322 -44011
rect -5402 -44084 -5379 -44050
rect -5345 -44084 -5322 -44050
rect -5402 -44118 -5322 -44084
rect -5402 -44152 -5379 -44118
rect -5345 -44152 -5322 -44118
rect -5402 -44186 -5322 -44152
rect -5402 -44220 -5379 -44186
rect -5345 -44220 -5322 -44186
rect -5402 -44254 -5322 -44220
rect -5402 -44288 -5379 -44254
rect -5345 -44288 -5322 -44254
rect -5402 -44322 -5322 -44288
rect -5402 -44356 -5379 -44322
rect -5345 -44356 -5322 -44322
rect -5402 -44390 -5322 -44356
rect -5402 -44424 -5379 -44390
rect -5345 -44424 -5322 -44390
rect -5402 -44458 -5322 -44424
rect -5402 -44492 -5379 -44458
rect -5345 -44492 -5322 -44458
rect -5402 -44526 -5322 -44492
rect -5402 -44560 -5379 -44526
rect -5345 -44560 -5322 -44526
rect -5402 -44594 -5322 -44560
rect -5402 -44628 -5379 -44594
rect -5345 -44628 -5322 -44594
rect -5402 -44662 -5322 -44628
rect -5402 -44696 -5379 -44662
rect -5345 -44696 -5322 -44662
rect -5402 -44730 -5322 -44696
rect -5402 -44764 -5379 -44730
rect -5345 -44764 -5322 -44730
rect -5402 -44798 -5322 -44764
rect -5402 -44832 -5379 -44798
rect -5345 -44832 -5322 -44798
rect -5402 -44871 -5322 -44832
rect -5252 -44060 -5172 -44011
rect -5252 -44094 -5229 -44060
rect -5195 -44094 -5172 -44060
rect -5252 -44128 -5172 -44094
rect -5252 -44162 -5229 -44128
rect -5195 -44162 -5172 -44128
rect -5252 -44196 -5172 -44162
rect -5252 -44230 -5229 -44196
rect -5195 -44230 -5172 -44196
rect -5252 -44264 -5172 -44230
rect -5252 -44298 -5229 -44264
rect -5195 -44298 -5172 -44264
rect -5252 -44332 -5172 -44298
rect -5252 -44366 -5229 -44332
rect -5195 -44366 -5172 -44332
rect -5252 -44400 -5172 -44366
rect -5252 -44434 -5229 -44400
rect -5195 -44434 -5172 -44400
rect -5252 -44468 -5172 -44434
rect -5252 -44502 -5229 -44468
rect -5195 -44502 -5172 -44468
rect -5252 -44536 -5172 -44502
rect -5252 -44570 -5229 -44536
rect -5195 -44570 -5172 -44536
rect -5252 -44604 -5172 -44570
rect -5252 -44638 -5229 -44604
rect -5195 -44638 -5172 -44604
rect -5252 -44672 -5172 -44638
rect -5252 -44706 -5229 -44672
rect -5195 -44706 -5172 -44672
rect -5252 -44740 -5172 -44706
rect -5252 -44774 -5229 -44740
rect -5195 -44774 -5172 -44740
rect -5252 -44808 -5172 -44774
rect -5252 -44842 -5229 -44808
rect -5195 -44842 -5172 -44808
rect -5252 -44871 -5172 -44842
rect -5102 -44050 -5022 -44011
rect -5102 -44084 -5079 -44050
rect -5045 -44084 -5022 -44050
rect -5102 -44118 -5022 -44084
rect -5102 -44152 -5079 -44118
rect -5045 -44152 -5022 -44118
rect -5102 -44186 -5022 -44152
rect -5102 -44220 -5079 -44186
rect -5045 -44220 -5022 -44186
rect -5102 -44254 -5022 -44220
rect -5102 -44288 -5079 -44254
rect -5045 -44288 -5022 -44254
rect -5102 -44322 -5022 -44288
rect -5102 -44356 -5079 -44322
rect -5045 -44356 -5022 -44322
rect -5102 -44390 -5022 -44356
rect -5102 -44424 -5079 -44390
rect -5045 -44424 -5022 -44390
rect -5102 -44458 -5022 -44424
rect -5102 -44492 -5079 -44458
rect -5045 -44492 -5022 -44458
rect -5102 -44526 -5022 -44492
rect -5102 -44560 -5079 -44526
rect -5045 -44560 -5022 -44526
rect -5102 -44594 -5022 -44560
rect -5102 -44628 -5079 -44594
rect -5045 -44628 -5022 -44594
rect -5102 -44662 -5022 -44628
rect -5102 -44696 -5079 -44662
rect -5045 -44696 -5022 -44662
rect -5102 -44730 -5022 -44696
rect -5102 -44764 -5079 -44730
rect -5045 -44764 -5022 -44730
rect -5102 -44798 -5022 -44764
rect -5102 -44832 -5079 -44798
rect -5045 -44832 -5022 -44798
rect -5102 -44871 -5022 -44832
rect -4952 -44050 -4872 -44011
rect -4952 -44084 -4929 -44050
rect -4895 -44084 -4872 -44050
rect -4952 -44118 -4872 -44084
rect -4952 -44152 -4929 -44118
rect -4895 -44152 -4872 -44118
rect -4952 -44186 -4872 -44152
rect -4952 -44220 -4929 -44186
rect -4895 -44220 -4872 -44186
rect -4952 -44254 -4872 -44220
rect -4952 -44288 -4929 -44254
rect -4895 -44288 -4872 -44254
rect -4952 -44322 -4872 -44288
rect -4952 -44356 -4929 -44322
rect -4895 -44356 -4872 -44322
rect -4952 -44390 -4872 -44356
rect -4952 -44424 -4929 -44390
rect -4895 -44424 -4872 -44390
rect -4952 -44458 -4872 -44424
rect -4952 -44492 -4929 -44458
rect -4895 -44492 -4872 -44458
rect -4952 -44526 -4872 -44492
rect -4952 -44560 -4929 -44526
rect -4895 -44560 -4872 -44526
rect -4952 -44594 -4872 -44560
rect -4952 -44628 -4929 -44594
rect -4895 -44628 -4872 -44594
rect -4952 -44662 -4872 -44628
rect -4952 -44696 -4929 -44662
rect -4895 -44696 -4872 -44662
rect -4952 -44730 -4872 -44696
rect -4952 -44764 -4929 -44730
rect -4895 -44764 -4872 -44730
rect -4952 -44798 -4872 -44764
rect -4952 -44832 -4929 -44798
rect -4895 -44832 -4872 -44798
rect -4952 -44871 -4872 -44832
rect -4802 -44050 -4722 -44011
rect -4802 -44084 -4779 -44050
rect -4745 -44084 -4722 -44050
rect -4802 -44118 -4722 -44084
rect -4802 -44152 -4779 -44118
rect -4745 -44152 -4722 -44118
rect -4802 -44186 -4722 -44152
rect -4802 -44220 -4779 -44186
rect -4745 -44220 -4722 -44186
rect -4802 -44254 -4722 -44220
rect -4802 -44288 -4779 -44254
rect -4745 -44288 -4722 -44254
rect -4802 -44322 -4722 -44288
rect -4802 -44356 -4779 -44322
rect -4745 -44356 -4722 -44322
rect -4802 -44390 -4722 -44356
rect -4802 -44424 -4779 -44390
rect -4745 -44424 -4722 -44390
rect -4802 -44458 -4722 -44424
rect -4802 -44492 -4779 -44458
rect -4745 -44492 -4722 -44458
rect -4802 -44526 -4722 -44492
rect -4802 -44560 -4779 -44526
rect -4745 -44560 -4722 -44526
rect -4802 -44594 -4722 -44560
rect -4802 -44628 -4779 -44594
rect -4745 -44628 -4722 -44594
rect -4802 -44662 -4722 -44628
rect -4802 -44696 -4779 -44662
rect -4745 -44696 -4722 -44662
rect -4802 -44730 -4722 -44696
rect -4802 -44764 -4779 -44730
rect -4745 -44764 -4722 -44730
rect -4802 -44798 -4722 -44764
rect -4802 -44832 -4779 -44798
rect -4745 -44832 -4722 -44798
rect -4802 -44871 -4722 -44832
rect -4652 -44050 -4572 -44011
rect -4652 -44084 -4629 -44050
rect -4595 -44084 -4572 -44050
rect -4652 -44118 -4572 -44084
rect -4652 -44152 -4629 -44118
rect -4595 -44152 -4572 -44118
rect -4652 -44186 -4572 -44152
rect -4652 -44220 -4629 -44186
rect -4595 -44220 -4572 -44186
rect -4652 -44254 -4572 -44220
rect -4652 -44288 -4629 -44254
rect -4595 -44288 -4572 -44254
rect -4652 -44322 -4572 -44288
rect -4652 -44356 -4629 -44322
rect -4595 -44356 -4572 -44322
rect -4652 -44390 -4572 -44356
rect -4652 -44424 -4629 -44390
rect -4595 -44424 -4572 -44390
rect -4652 -44458 -4572 -44424
rect -4652 -44492 -4629 -44458
rect -4595 -44492 -4572 -44458
rect -4652 -44526 -4572 -44492
rect -4652 -44560 -4629 -44526
rect -4595 -44560 -4572 -44526
rect -4652 -44594 -4572 -44560
rect -4652 -44628 -4629 -44594
rect -4595 -44628 -4572 -44594
rect -4652 -44662 -4572 -44628
rect -4652 -44696 -4629 -44662
rect -4595 -44696 -4572 -44662
rect -4652 -44730 -4572 -44696
rect -4652 -44764 -4629 -44730
rect -4595 -44764 -4572 -44730
rect -4652 -44798 -4572 -44764
rect -4652 -44832 -4629 -44798
rect -4595 -44832 -4572 -44798
rect -4652 -44871 -4572 -44832
rect -4502 -44050 -4422 -44011
rect -4502 -44084 -4479 -44050
rect -4445 -44084 -4422 -44050
rect -4502 -44118 -4422 -44084
rect -4502 -44152 -4479 -44118
rect -4445 -44152 -4422 -44118
rect -4502 -44186 -4422 -44152
rect -4502 -44220 -4479 -44186
rect -4445 -44220 -4422 -44186
rect -4502 -44254 -4422 -44220
rect -4502 -44288 -4479 -44254
rect -4445 -44288 -4422 -44254
rect -4502 -44322 -4422 -44288
rect -4502 -44356 -4479 -44322
rect -4445 -44356 -4422 -44322
rect -4502 -44390 -4422 -44356
rect -4502 -44424 -4479 -44390
rect -4445 -44424 -4422 -44390
rect -4502 -44458 -4422 -44424
rect -4502 -44492 -4479 -44458
rect -4445 -44492 -4422 -44458
rect -4502 -44526 -4422 -44492
rect -4502 -44560 -4479 -44526
rect -4445 -44560 -4422 -44526
rect -4502 -44594 -4422 -44560
rect -4502 -44628 -4479 -44594
rect -4445 -44628 -4422 -44594
rect -4502 -44662 -4422 -44628
rect -4502 -44696 -4479 -44662
rect -4445 -44696 -4422 -44662
rect -4502 -44730 -4422 -44696
rect -4502 -44764 -4479 -44730
rect -4445 -44764 -4422 -44730
rect -4502 -44798 -4422 -44764
rect -4502 -44832 -4479 -44798
rect -4445 -44832 -4422 -44798
rect -4502 -44871 -4422 -44832
rect -4352 -44050 -4272 -44011
rect -4352 -44084 -4329 -44050
rect -4295 -44084 -4272 -44050
rect -4352 -44118 -4272 -44084
rect -4352 -44152 -4329 -44118
rect -4295 -44152 -4272 -44118
rect -4352 -44186 -4272 -44152
rect -4352 -44220 -4329 -44186
rect -4295 -44220 -4272 -44186
rect -4352 -44254 -4272 -44220
rect -4352 -44288 -4329 -44254
rect -4295 -44288 -4272 -44254
rect -4352 -44322 -4272 -44288
rect -4352 -44356 -4329 -44322
rect -4295 -44356 -4272 -44322
rect -4352 -44390 -4272 -44356
rect -4352 -44424 -4329 -44390
rect -4295 -44424 -4272 -44390
rect -4352 -44458 -4272 -44424
rect -4352 -44492 -4329 -44458
rect -4295 -44492 -4272 -44458
rect -4352 -44526 -4272 -44492
rect -4352 -44560 -4329 -44526
rect -4295 -44560 -4272 -44526
rect -4352 -44594 -4272 -44560
rect -4352 -44628 -4329 -44594
rect -4295 -44628 -4272 -44594
rect -4352 -44662 -4272 -44628
rect -4352 -44696 -4329 -44662
rect -4295 -44696 -4272 -44662
rect -4352 -44730 -4272 -44696
rect -4352 -44764 -4329 -44730
rect -4295 -44764 -4272 -44730
rect -4352 -44798 -4272 -44764
rect -4352 -44832 -4329 -44798
rect -4295 -44832 -4272 -44798
rect -4352 -44871 -4272 -44832
rect -4202 -44050 -4122 -44011
rect -4202 -44084 -4179 -44050
rect -4145 -44084 -4122 -44050
rect -4202 -44118 -4122 -44084
rect -4202 -44152 -4179 -44118
rect -4145 -44152 -4122 -44118
rect -4202 -44186 -4122 -44152
rect -4202 -44220 -4179 -44186
rect -4145 -44220 -4122 -44186
rect -4202 -44254 -4122 -44220
rect -4202 -44288 -4179 -44254
rect -4145 -44288 -4122 -44254
rect -4202 -44322 -4122 -44288
rect -4202 -44356 -4179 -44322
rect -4145 -44356 -4122 -44322
rect -4202 -44390 -4122 -44356
rect -4202 -44424 -4179 -44390
rect -4145 -44424 -4122 -44390
rect -4202 -44458 -4122 -44424
rect -4202 -44492 -4179 -44458
rect -4145 -44492 -4122 -44458
rect -4202 -44526 -4122 -44492
rect -4202 -44560 -4179 -44526
rect -4145 -44560 -4122 -44526
rect -4202 -44594 -4122 -44560
rect -4202 -44628 -4179 -44594
rect -4145 -44628 -4122 -44594
rect -4202 -44662 -4122 -44628
rect -4202 -44696 -4179 -44662
rect -4145 -44696 -4122 -44662
rect -4202 -44730 -4122 -44696
rect -4202 -44764 -4179 -44730
rect -4145 -44764 -4122 -44730
rect -4202 -44798 -4122 -44764
rect -4202 -44832 -4179 -44798
rect -4145 -44832 -4122 -44798
rect -4202 -44871 -4122 -44832
rect -4052 -44050 -3972 -44011
rect -4052 -44084 -4029 -44050
rect -3995 -44084 -3972 -44050
rect -4052 -44118 -3972 -44084
rect -4052 -44152 -4029 -44118
rect -3995 -44152 -3972 -44118
rect -4052 -44186 -3972 -44152
rect -4052 -44220 -4029 -44186
rect -3995 -44220 -3972 -44186
rect -4052 -44254 -3972 -44220
rect -4052 -44288 -4029 -44254
rect -3995 -44288 -3972 -44254
rect -4052 -44322 -3972 -44288
rect -4052 -44356 -4029 -44322
rect -3995 -44356 -3972 -44322
rect -4052 -44390 -3972 -44356
rect -4052 -44424 -4029 -44390
rect -3995 -44424 -3972 -44390
rect -4052 -44458 -3972 -44424
rect -4052 -44492 -4029 -44458
rect -3995 -44492 -3972 -44458
rect -4052 -44526 -3972 -44492
rect -4052 -44560 -4029 -44526
rect -3995 -44560 -3972 -44526
rect -4052 -44594 -3972 -44560
rect -4052 -44628 -4029 -44594
rect -3995 -44628 -3972 -44594
rect -4052 -44662 -3972 -44628
rect -4052 -44696 -4029 -44662
rect -3995 -44696 -3972 -44662
rect -4052 -44730 -3972 -44696
rect -4052 -44764 -4029 -44730
rect -3995 -44764 -3972 -44730
rect -4052 -44798 -3972 -44764
rect -4052 -44832 -4029 -44798
rect -3995 -44832 -3972 -44798
rect -4052 -44871 -3972 -44832
rect -3902 -44050 -3822 -44011
rect -3902 -44084 -3879 -44050
rect -3845 -44084 -3822 -44050
rect -3902 -44118 -3822 -44084
rect -3902 -44152 -3879 -44118
rect -3845 -44152 -3822 -44118
rect -3902 -44186 -3822 -44152
rect -3902 -44220 -3879 -44186
rect -3845 -44220 -3822 -44186
rect -3902 -44254 -3822 -44220
rect -3902 -44288 -3879 -44254
rect -3845 -44288 -3822 -44254
rect -3902 -44322 -3822 -44288
rect -3902 -44356 -3879 -44322
rect -3845 -44356 -3822 -44322
rect -3902 -44390 -3822 -44356
rect -3902 -44424 -3879 -44390
rect -3845 -44424 -3822 -44390
rect -3902 -44458 -3822 -44424
rect -3902 -44492 -3879 -44458
rect -3845 -44492 -3822 -44458
rect -3902 -44526 -3822 -44492
rect -3902 -44560 -3879 -44526
rect -3845 -44560 -3822 -44526
rect -3902 -44594 -3822 -44560
rect -3902 -44628 -3879 -44594
rect -3845 -44628 -3822 -44594
rect -3902 -44662 -3822 -44628
rect -3902 -44696 -3879 -44662
rect -3845 -44696 -3822 -44662
rect -3902 -44730 -3822 -44696
rect -3902 -44764 -3879 -44730
rect -3845 -44764 -3822 -44730
rect -3902 -44798 -3822 -44764
rect -3902 -44832 -3879 -44798
rect -3845 -44832 -3822 -44798
rect -3902 -44871 -3822 -44832
rect -3752 -44060 -3672 -44011
rect -3752 -44094 -3729 -44060
rect -3695 -44094 -3672 -44060
rect -3752 -44128 -3672 -44094
rect -3752 -44162 -3729 -44128
rect -3695 -44162 -3672 -44128
rect -3752 -44196 -3672 -44162
rect -3752 -44230 -3729 -44196
rect -3695 -44230 -3672 -44196
rect -3752 -44264 -3672 -44230
rect -3752 -44298 -3729 -44264
rect -3695 -44298 -3672 -44264
rect -3752 -44332 -3672 -44298
rect -3752 -44366 -3729 -44332
rect -3695 -44366 -3672 -44332
rect -3752 -44400 -3672 -44366
rect -3752 -44434 -3729 -44400
rect -3695 -44434 -3672 -44400
rect -3752 -44468 -3672 -44434
rect -3752 -44502 -3729 -44468
rect -3695 -44502 -3672 -44468
rect -3752 -44536 -3672 -44502
rect -3752 -44570 -3729 -44536
rect -3695 -44570 -3672 -44536
rect -3752 -44604 -3672 -44570
rect -3752 -44638 -3729 -44604
rect -3695 -44638 -3672 -44604
rect -3752 -44672 -3672 -44638
rect -3752 -44706 -3729 -44672
rect -3695 -44706 -3672 -44672
rect -3752 -44740 -3672 -44706
rect -3752 -44774 -3729 -44740
rect -3695 -44774 -3672 -44740
rect -3752 -44808 -3672 -44774
rect -3752 -44842 -3729 -44808
rect -3695 -44842 -3672 -44808
rect -3752 -44871 -3672 -44842
rect -3602 -44050 -3522 -44011
rect -3602 -44084 -3579 -44050
rect -3545 -44084 -3522 -44050
rect -3602 -44118 -3522 -44084
rect -3602 -44152 -3579 -44118
rect -3545 -44152 -3522 -44118
rect -3602 -44186 -3522 -44152
rect -3602 -44220 -3579 -44186
rect -3545 -44220 -3522 -44186
rect -3602 -44254 -3522 -44220
rect -3602 -44288 -3579 -44254
rect -3545 -44288 -3522 -44254
rect -3602 -44322 -3522 -44288
rect -3602 -44356 -3579 -44322
rect -3545 -44356 -3522 -44322
rect -3602 -44390 -3522 -44356
rect -3602 -44424 -3579 -44390
rect -3545 -44424 -3522 -44390
rect -3602 -44458 -3522 -44424
rect -3602 -44492 -3579 -44458
rect -3545 -44492 -3522 -44458
rect -3602 -44526 -3522 -44492
rect -3602 -44560 -3579 -44526
rect -3545 -44560 -3522 -44526
rect -3602 -44594 -3522 -44560
rect -3602 -44628 -3579 -44594
rect -3545 -44628 -3522 -44594
rect -3602 -44662 -3522 -44628
rect -3602 -44696 -3579 -44662
rect -3545 -44696 -3522 -44662
rect -3602 -44730 -3522 -44696
rect -3602 -44764 -3579 -44730
rect -3545 -44764 -3522 -44730
rect -3602 -44798 -3522 -44764
rect -3602 -44832 -3579 -44798
rect -3545 -44832 -3522 -44798
rect -3602 -44871 -3522 -44832
rect -3452 -44050 -3372 -44011
rect -3452 -44084 -3429 -44050
rect -3395 -44084 -3372 -44050
rect -3452 -44118 -3372 -44084
rect -3452 -44152 -3429 -44118
rect -3395 -44152 -3372 -44118
rect -3452 -44186 -3372 -44152
rect -3452 -44220 -3429 -44186
rect -3395 -44220 -3372 -44186
rect -3452 -44254 -3372 -44220
rect -3452 -44288 -3429 -44254
rect -3395 -44288 -3372 -44254
rect -3452 -44322 -3372 -44288
rect -3452 -44356 -3429 -44322
rect -3395 -44356 -3372 -44322
rect -3452 -44390 -3372 -44356
rect -3452 -44424 -3429 -44390
rect -3395 -44424 -3372 -44390
rect -3452 -44458 -3372 -44424
rect -3452 -44492 -3429 -44458
rect -3395 -44492 -3372 -44458
rect -3452 -44526 -3372 -44492
rect -3452 -44560 -3429 -44526
rect -3395 -44560 -3372 -44526
rect -3452 -44594 -3372 -44560
rect -3452 -44628 -3429 -44594
rect -3395 -44628 -3372 -44594
rect -3452 -44662 -3372 -44628
rect -3452 -44696 -3429 -44662
rect -3395 -44696 -3372 -44662
rect -3452 -44730 -3372 -44696
rect -3452 -44764 -3429 -44730
rect -3395 -44764 -3372 -44730
rect -3452 -44798 -3372 -44764
rect -3452 -44832 -3429 -44798
rect -3395 -44832 -3372 -44798
rect -3452 -44871 -3372 -44832
rect -3302 -44050 -3222 -44011
rect -3302 -44084 -3279 -44050
rect -3245 -44084 -3222 -44050
rect -3302 -44118 -3222 -44084
rect -3302 -44152 -3279 -44118
rect -3245 -44152 -3222 -44118
rect -3302 -44186 -3222 -44152
rect -3302 -44220 -3279 -44186
rect -3245 -44220 -3222 -44186
rect -3302 -44254 -3222 -44220
rect -3302 -44288 -3279 -44254
rect -3245 -44288 -3222 -44254
rect -3302 -44322 -3222 -44288
rect -3302 -44356 -3279 -44322
rect -3245 -44356 -3222 -44322
rect -3302 -44390 -3222 -44356
rect -3302 -44424 -3279 -44390
rect -3245 -44424 -3222 -44390
rect -3302 -44458 -3222 -44424
rect -3302 -44492 -3279 -44458
rect -3245 -44492 -3222 -44458
rect -3302 -44526 -3222 -44492
rect -3302 -44560 -3279 -44526
rect -3245 -44560 -3222 -44526
rect -3302 -44594 -3222 -44560
rect -3302 -44628 -3279 -44594
rect -3245 -44628 -3222 -44594
rect -3302 -44662 -3222 -44628
rect -3302 -44696 -3279 -44662
rect -3245 -44696 -3222 -44662
rect -3302 -44730 -3222 -44696
rect -3302 -44764 -3279 -44730
rect -3245 -44764 -3222 -44730
rect -3302 -44798 -3222 -44764
rect -3302 -44832 -3279 -44798
rect -3245 -44832 -3222 -44798
rect -3302 -44871 -3222 -44832
rect -3152 -44050 -3072 -44011
rect -3152 -44084 -3129 -44050
rect -3095 -44084 -3072 -44050
rect -3152 -44118 -3072 -44084
rect -3152 -44152 -3129 -44118
rect -3095 -44152 -3072 -44118
rect -3152 -44186 -3072 -44152
rect -3152 -44220 -3129 -44186
rect -3095 -44220 -3072 -44186
rect -3152 -44254 -3072 -44220
rect -3152 -44288 -3129 -44254
rect -3095 -44288 -3072 -44254
rect -3152 -44322 -3072 -44288
rect -3152 -44356 -3129 -44322
rect -3095 -44356 -3072 -44322
rect -3152 -44390 -3072 -44356
rect -3152 -44424 -3129 -44390
rect -3095 -44424 -3072 -44390
rect -3152 -44458 -3072 -44424
rect -3152 -44492 -3129 -44458
rect -3095 -44492 -3072 -44458
rect -3152 -44526 -3072 -44492
rect -3152 -44560 -3129 -44526
rect -3095 -44560 -3072 -44526
rect -3152 -44594 -3072 -44560
rect -3152 -44628 -3129 -44594
rect -3095 -44628 -3072 -44594
rect -3152 -44662 -3072 -44628
rect -3152 -44696 -3129 -44662
rect -3095 -44696 -3072 -44662
rect -3152 -44730 -3072 -44696
rect -3152 -44764 -3129 -44730
rect -3095 -44764 -3072 -44730
rect -3152 -44798 -3072 -44764
rect -3152 -44832 -3129 -44798
rect -3095 -44832 -3072 -44798
rect -3152 -44871 -3072 -44832
rect -3002 -44050 -2922 -44011
rect -3002 -44084 -2979 -44050
rect -2945 -44084 -2922 -44050
rect -3002 -44118 -2922 -44084
rect -3002 -44152 -2979 -44118
rect -2945 -44152 -2922 -44118
rect -3002 -44186 -2922 -44152
rect -3002 -44220 -2979 -44186
rect -2945 -44220 -2922 -44186
rect -3002 -44254 -2922 -44220
rect -3002 -44288 -2979 -44254
rect -2945 -44288 -2922 -44254
rect -3002 -44322 -2922 -44288
rect -3002 -44356 -2979 -44322
rect -2945 -44356 -2922 -44322
rect -3002 -44390 -2922 -44356
rect -3002 -44424 -2979 -44390
rect -2945 -44424 -2922 -44390
rect -3002 -44458 -2922 -44424
rect -3002 -44492 -2979 -44458
rect -2945 -44492 -2922 -44458
rect -3002 -44526 -2922 -44492
rect -3002 -44560 -2979 -44526
rect -2945 -44560 -2922 -44526
rect -3002 -44594 -2922 -44560
rect -3002 -44628 -2979 -44594
rect -2945 -44628 -2922 -44594
rect -3002 -44662 -2922 -44628
rect -3002 -44696 -2979 -44662
rect -2945 -44696 -2922 -44662
rect -3002 -44730 -2922 -44696
rect -3002 -44764 -2979 -44730
rect -2945 -44764 -2922 -44730
rect -3002 -44798 -2922 -44764
rect -3002 -44832 -2979 -44798
rect -2945 -44832 -2922 -44798
rect -3002 -44871 -2922 -44832
rect -2852 -44050 -2772 -44011
rect -2852 -44084 -2829 -44050
rect -2795 -44084 -2772 -44050
rect -2852 -44118 -2772 -44084
rect -2852 -44152 -2829 -44118
rect -2795 -44152 -2772 -44118
rect -2852 -44186 -2772 -44152
rect -2852 -44220 -2829 -44186
rect -2795 -44220 -2772 -44186
rect -2852 -44254 -2772 -44220
rect -2852 -44288 -2829 -44254
rect -2795 -44288 -2772 -44254
rect -2852 -44322 -2772 -44288
rect -2852 -44356 -2829 -44322
rect -2795 -44356 -2772 -44322
rect -2852 -44390 -2772 -44356
rect -2852 -44424 -2829 -44390
rect -2795 -44424 -2772 -44390
rect -2852 -44458 -2772 -44424
rect -2852 -44492 -2829 -44458
rect -2795 -44492 -2772 -44458
rect -2852 -44526 -2772 -44492
rect -2852 -44560 -2829 -44526
rect -2795 -44560 -2772 -44526
rect -2852 -44594 -2772 -44560
rect -2852 -44628 -2829 -44594
rect -2795 -44628 -2772 -44594
rect -2852 -44662 -2772 -44628
rect -2852 -44696 -2829 -44662
rect -2795 -44696 -2772 -44662
rect -2852 -44730 -2772 -44696
rect -2852 -44764 -2829 -44730
rect -2795 -44764 -2772 -44730
rect -2852 -44798 -2772 -44764
rect -2852 -44832 -2829 -44798
rect -2795 -44832 -2772 -44798
rect -2852 -44871 -2772 -44832
rect -2702 -44050 -2622 -44011
rect -2702 -44084 -2679 -44050
rect -2645 -44084 -2622 -44050
rect -2702 -44118 -2622 -44084
rect -2702 -44152 -2679 -44118
rect -2645 -44152 -2622 -44118
rect -2702 -44186 -2622 -44152
rect -2702 -44220 -2679 -44186
rect -2645 -44220 -2622 -44186
rect -2702 -44254 -2622 -44220
rect -2702 -44288 -2679 -44254
rect -2645 -44288 -2622 -44254
rect -2702 -44322 -2622 -44288
rect -2702 -44356 -2679 -44322
rect -2645 -44356 -2622 -44322
rect -2702 -44390 -2622 -44356
rect -2702 -44424 -2679 -44390
rect -2645 -44424 -2622 -44390
rect -2702 -44458 -2622 -44424
rect -2702 -44492 -2679 -44458
rect -2645 -44492 -2622 -44458
rect -2702 -44526 -2622 -44492
rect -2702 -44560 -2679 -44526
rect -2645 -44560 -2622 -44526
rect -2702 -44594 -2622 -44560
rect -2702 -44628 -2679 -44594
rect -2645 -44628 -2622 -44594
rect -2702 -44662 -2622 -44628
rect -2702 -44696 -2679 -44662
rect -2645 -44696 -2622 -44662
rect -2702 -44730 -2622 -44696
rect -2702 -44764 -2679 -44730
rect -2645 -44764 -2622 -44730
rect -2702 -44798 -2622 -44764
rect -2702 -44832 -2679 -44798
rect -2645 -44832 -2622 -44798
rect -2702 -44871 -2622 -44832
rect -2552 -44050 -2472 -44011
rect -2552 -44084 -2529 -44050
rect -2495 -44084 -2472 -44050
rect -2552 -44118 -2472 -44084
rect -2552 -44152 -2529 -44118
rect -2495 -44152 -2472 -44118
rect -2552 -44186 -2472 -44152
rect -2552 -44220 -2529 -44186
rect -2495 -44220 -2472 -44186
rect -2552 -44254 -2472 -44220
rect -2552 -44288 -2529 -44254
rect -2495 -44288 -2472 -44254
rect -2552 -44322 -2472 -44288
rect -2552 -44356 -2529 -44322
rect -2495 -44356 -2472 -44322
rect -2552 -44390 -2472 -44356
rect -2552 -44424 -2529 -44390
rect -2495 -44424 -2472 -44390
rect -2552 -44458 -2472 -44424
rect -2552 -44492 -2529 -44458
rect -2495 -44492 -2472 -44458
rect -2552 -44526 -2472 -44492
rect -2552 -44560 -2529 -44526
rect -2495 -44560 -2472 -44526
rect -2552 -44594 -2472 -44560
rect -2552 -44628 -2529 -44594
rect -2495 -44628 -2472 -44594
rect -2552 -44662 -2472 -44628
rect -2552 -44696 -2529 -44662
rect -2495 -44696 -2472 -44662
rect -2552 -44730 -2472 -44696
rect -2552 -44764 -2529 -44730
rect -2495 -44764 -2472 -44730
rect -2552 -44798 -2472 -44764
rect -2552 -44832 -2529 -44798
rect -2495 -44832 -2472 -44798
rect -2552 -44871 -2472 -44832
rect -2402 -44050 -2322 -44011
rect -2402 -44084 -2379 -44050
rect -2345 -44084 -2322 -44050
rect -2402 -44118 -2322 -44084
rect -2402 -44152 -2379 -44118
rect -2345 -44152 -2322 -44118
rect -2402 -44186 -2322 -44152
rect -2402 -44220 -2379 -44186
rect -2345 -44220 -2322 -44186
rect -2402 -44254 -2322 -44220
rect -2402 -44288 -2379 -44254
rect -2345 -44288 -2322 -44254
rect -2402 -44322 -2322 -44288
rect -2402 -44356 -2379 -44322
rect -2345 -44356 -2322 -44322
rect -2402 -44390 -2322 -44356
rect -2402 -44424 -2379 -44390
rect -2345 -44424 -2322 -44390
rect -2402 -44458 -2322 -44424
rect -2402 -44492 -2379 -44458
rect -2345 -44492 -2322 -44458
rect -2402 -44526 -2322 -44492
rect -2402 -44560 -2379 -44526
rect -2345 -44560 -2322 -44526
rect -2402 -44594 -2322 -44560
rect -2402 -44628 -2379 -44594
rect -2345 -44628 -2322 -44594
rect -2402 -44662 -2322 -44628
rect -2402 -44696 -2379 -44662
rect -2345 -44696 -2322 -44662
rect -2402 -44730 -2322 -44696
rect -2402 -44764 -2379 -44730
rect -2345 -44764 -2322 -44730
rect -2402 -44798 -2322 -44764
rect -2402 -44832 -2379 -44798
rect -2345 -44832 -2322 -44798
rect -2402 -44871 -2322 -44832
rect -2282 -44050 -2202 -44011
rect -2282 -44084 -2259 -44050
rect -2225 -44084 -2202 -44050
rect -2282 -44118 -2202 -44084
rect -2282 -44152 -2259 -44118
rect -2225 -44152 -2202 -44118
rect -2282 -44186 -2202 -44152
rect -2282 -44220 -2259 -44186
rect -2225 -44220 -2202 -44186
rect -2282 -44254 -2202 -44220
rect -2282 -44288 -2259 -44254
rect -2225 -44288 -2202 -44254
rect -2282 -44322 -2202 -44288
rect -2282 -44356 -2259 -44322
rect -2225 -44356 -2202 -44322
rect -2282 -44390 -2202 -44356
rect -2282 -44424 -2259 -44390
rect -2225 -44424 -2202 -44390
rect -2282 -44458 -2202 -44424
rect -2282 -44492 -2259 -44458
rect -2225 -44492 -2202 -44458
rect -2282 -44526 -2202 -44492
rect -2282 -44560 -2259 -44526
rect -2225 -44560 -2202 -44526
rect -2282 -44594 -2202 -44560
rect -2282 -44628 -2259 -44594
rect -2225 -44628 -2202 -44594
rect -2282 -44662 -2202 -44628
rect -2282 -44696 -2259 -44662
rect -2225 -44696 -2202 -44662
rect -2282 -44730 -2202 -44696
rect -2282 -44764 -2259 -44730
rect -2225 -44764 -2202 -44730
rect -2282 -44798 -2202 -44764
rect -2282 -44832 -2259 -44798
rect -2225 -44832 -2202 -44798
rect -5232 -44911 -5192 -44871
rect -4931 -44911 -4891 -44871
rect -4631 -44911 -4591 -44871
rect -4331 -44911 -4291 -44871
rect -4032 -44911 -3992 -44871
rect -5232 -44951 -3992 -44911
rect -3882 -44911 -3842 -44871
rect -3582 -44911 -3542 -44871
rect -3282 -44911 -3242 -44871
rect -2982 -44911 -2942 -44871
rect -2682 -44911 -2642 -44871
rect -2382 -44911 -2342 -44871
rect -3882 -44951 -2342 -44911
rect -5232 -45096 -4972 -44951
rect -5232 -45130 -5179 -45096
rect -5145 -45130 -5059 -45096
rect -5025 -45130 -4972 -45096
rect -5232 -45216 -4972 -45130
rect -5232 -45250 -5179 -45216
rect -5145 -45250 -5059 -45216
rect -5025 -45250 -4972 -45216
rect -5232 -45303 -4972 -45250
rect -2282 -45413 -2202 -44832
rect -11742 -45436 -2100 -45413
rect -11742 -45470 -11699 -45436
rect -11665 -45470 -11619 -45436
rect -11585 -45470 -11539 -45436
rect -11505 -45470 -11459 -45436
rect -11425 -45470 -11379 -45436
rect -11345 -45470 -11299 -45436
rect -11265 -45470 -11219 -45436
rect -11185 -45470 -11139 -45436
rect -11105 -45470 -11059 -45436
rect -11025 -45470 -10979 -45436
rect -10945 -45470 -10899 -45436
rect -10865 -45470 -10819 -45436
rect -10785 -45470 -10739 -45436
rect -10705 -45470 -10659 -45436
rect -10625 -45470 -10579 -45436
rect -10545 -45470 -10499 -45436
rect -10465 -45470 -10419 -45436
rect -10385 -45470 -10339 -45436
rect -10305 -45470 -10259 -45436
rect -10225 -45470 -10179 -45436
rect -10145 -45470 -10099 -45436
rect -10065 -45470 -10019 -45436
rect -9985 -45470 -9939 -45436
rect -9905 -45470 -9859 -45436
rect -9825 -45470 -9779 -45436
rect -9745 -45470 -9699 -45436
rect -9665 -45470 -9619 -45436
rect -9585 -45470 -9539 -45436
rect -9505 -45470 -9459 -45436
rect -9425 -45470 -9379 -45436
rect -9345 -45470 -9299 -45436
rect -9265 -45470 -9219 -45436
rect -9185 -45470 -9139 -45436
rect -9105 -45470 -9059 -45436
rect -9025 -45470 -8979 -45436
rect -8945 -45470 -8899 -45436
rect -8865 -45470 -8819 -45436
rect -8785 -45470 -8739 -45436
rect -8705 -45470 -8659 -45436
rect -8625 -45470 -8579 -45436
rect -8545 -45470 -8499 -45436
rect -8465 -45470 -8419 -45436
rect -8385 -45470 -8339 -45436
rect -8305 -45470 -8259 -45436
rect -8225 -45470 -8179 -45436
rect -8145 -45470 -8099 -45436
rect -8065 -45470 -8019 -45436
rect -7985 -45470 -7939 -45436
rect -7905 -45470 -7859 -45436
rect -7825 -45470 -7779 -45436
rect -7745 -45470 -7699 -45436
rect -7665 -45470 -7619 -45436
rect -7585 -45470 -7539 -45436
rect -7505 -45470 -7459 -45436
rect -7425 -45470 -7379 -45436
rect -7345 -45470 -7299 -45436
rect -7265 -45470 -7219 -45436
rect -7185 -45470 -7139 -45436
rect -7105 -45470 -7059 -45436
rect -7025 -45470 -6979 -45436
rect -6945 -45470 -6899 -45436
rect -6865 -45470 -6819 -45436
rect -6785 -45470 -6739 -45436
rect -6705 -45470 -6659 -45436
rect -6625 -45470 -6579 -45436
rect -6545 -45470 -6499 -45436
rect -6465 -45470 -6419 -45436
rect -6385 -45470 -6339 -45436
rect -6305 -45470 -6259 -45436
rect -6225 -45470 -6179 -45436
rect -6145 -45470 -6099 -45436
rect -6065 -45470 -6019 -45436
rect -5985 -45470 -5939 -45436
rect -5905 -45470 -5859 -45436
rect -5825 -45470 -5779 -45436
rect -5745 -45470 -5699 -45436
rect -5665 -45470 -5619 -45436
rect -5585 -45470 -5539 -45436
rect -5505 -45470 -5459 -45436
rect -5425 -45470 -5379 -45436
rect -5345 -45470 -5299 -45436
rect -5265 -45470 -5219 -45436
rect -5185 -45470 -5139 -45436
rect -5105 -45470 -5059 -45436
rect -5025 -45470 -4979 -45436
rect -4945 -45470 -4899 -45436
rect -4865 -45470 -4819 -45436
rect -4785 -45470 -4739 -45436
rect -4705 -45470 -4659 -45436
rect -4625 -45470 -4579 -45436
rect -4545 -45470 -4499 -45436
rect -4465 -45470 -4419 -45436
rect -4385 -45470 -4339 -45436
rect -4305 -45470 -4259 -45436
rect -4225 -45470 -4179 -45436
rect -4145 -45470 -4099 -45436
rect -4065 -45470 -4019 -45436
rect -3985 -45470 -3939 -45436
rect -3905 -45470 -3859 -45436
rect -3825 -45470 -3779 -45436
rect -3745 -45470 -3699 -45436
rect -3665 -45470 -3619 -45436
rect -3585 -45470 -3539 -45436
rect -3505 -45470 -3459 -45436
rect -3425 -45470 -3379 -45436
rect -3345 -45470 -3299 -45436
rect -3265 -45470 -3219 -45436
rect -3185 -45470 -3139 -45436
rect -3105 -45470 -3059 -45436
rect -3025 -45470 -2979 -45436
rect -2945 -45470 -2899 -45436
rect -2865 -45470 -2819 -45436
rect -2785 -45470 -2739 -45436
rect -2705 -45470 -2659 -45436
rect -2625 -45470 -2579 -45436
rect -2545 -45470 -2499 -45436
rect -2465 -45470 -2419 -45436
rect -2385 -45470 -2339 -45436
rect -2305 -45470 -2259 -45436
rect -2225 -45470 -2179 -45436
rect -2145 -45470 -2100 -45436
rect -11742 -45493 -2100 -45470
rect -6855 -45958 -6595 -45905
rect -6855 -45992 -6802 -45958
rect -6768 -45992 -6682 -45958
rect -6648 -45992 -6595 -45958
rect -6855 -46078 -6595 -45992
rect -6855 -46112 -6802 -46078
rect -6768 -46112 -6682 -46078
rect -6648 -46112 -6595 -46078
rect -6855 -46165 -6595 -46112
rect -5229 -45958 -4969 -45905
rect -5229 -45992 -5176 -45958
rect -5142 -45992 -5056 -45958
rect -5022 -45992 -4969 -45958
rect -5229 -46078 -4969 -45992
rect -5229 -46112 -5176 -46078
rect -5142 -46112 -5056 -46078
rect -5022 -46112 -4969 -46078
rect -5229 -46165 -4969 -46112
rect -44481 -46975 -4170 -46952
rect -44481 -47009 -44435 -46975
rect -44401 -47009 -44355 -46975
rect -44321 -47009 -44275 -46975
rect -44241 -47009 -44195 -46975
rect -44161 -47009 -44115 -46975
rect -44081 -47009 -44035 -46975
rect -44001 -47009 -43955 -46975
rect -43921 -47009 -43875 -46975
rect -43841 -47009 -43795 -46975
rect -43761 -47009 -43715 -46975
rect -43681 -47009 -43635 -46975
rect -43601 -47009 -43555 -46975
rect -43521 -47009 -43475 -46975
rect -43441 -47009 -43395 -46975
rect -43361 -47009 -43315 -46975
rect -43281 -47009 -43235 -46975
rect -43201 -47009 -43155 -46975
rect -43121 -47009 -43075 -46975
rect -43041 -47009 -42995 -46975
rect -42961 -47009 -42915 -46975
rect -42881 -47009 -42835 -46975
rect -42801 -47009 -42755 -46975
rect -42721 -47009 -42675 -46975
rect -42641 -47009 -42595 -46975
rect -42561 -47009 -42515 -46975
rect -42481 -47009 -42435 -46975
rect -42401 -47009 -42355 -46975
rect -42321 -47009 -42275 -46975
rect -42241 -47009 -42195 -46975
rect -42161 -47009 -42115 -46975
rect -42081 -47009 -42035 -46975
rect -42001 -47009 -41955 -46975
rect -41921 -47009 -41875 -46975
rect -41841 -47009 -41795 -46975
rect -41761 -47009 -41715 -46975
rect -41681 -47009 -41635 -46975
rect -41601 -47009 -41555 -46975
rect -41521 -47009 -41475 -46975
rect -41441 -47009 -41395 -46975
rect -41361 -47009 -41315 -46975
rect -41281 -47009 -41235 -46975
rect -41201 -47009 -41155 -46975
rect -41121 -47009 -41075 -46975
rect -41041 -47009 -40995 -46975
rect -40961 -47009 -40915 -46975
rect -40881 -47009 -40835 -46975
rect -40801 -47009 -40755 -46975
rect -40721 -47009 -40675 -46975
rect -40641 -47009 -40595 -46975
rect -40561 -47009 -40515 -46975
rect -40481 -47009 -40435 -46975
rect -40401 -47009 -40355 -46975
rect -40321 -47009 -40275 -46975
rect -40241 -47009 -40195 -46975
rect -40161 -47009 -40115 -46975
rect -40081 -47009 -40035 -46975
rect -40001 -47009 -39955 -46975
rect -39921 -47009 -39875 -46975
rect -39841 -47009 -39795 -46975
rect -39761 -47009 -39715 -46975
rect -39681 -47009 -39635 -46975
rect -39601 -47009 -39555 -46975
rect -39521 -47009 -39475 -46975
rect -39441 -47009 -39395 -46975
rect -39361 -47009 -39315 -46975
rect -39281 -47009 -39235 -46975
rect -39201 -47009 -39155 -46975
rect -39121 -47009 -39075 -46975
rect -39041 -47009 -38995 -46975
rect -38961 -47009 -38915 -46975
rect -38881 -47009 -38835 -46975
rect -38801 -47009 -38755 -46975
rect -38721 -47009 -38675 -46975
rect -38641 -47009 -38595 -46975
rect -38561 -47009 -38515 -46975
rect -38481 -47009 -38435 -46975
rect -38401 -47009 -38355 -46975
rect -38321 -47009 -38275 -46975
rect -38241 -47009 -38195 -46975
rect -38161 -47009 -38115 -46975
rect -38081 -47009 -38035 -46975
rect -38001 -47009 -37955 -46975
rect -37921 -47009 -37875 -46975
rect -37841 -47009 -37795 -46975
rect -37761 -47009 -37715 -46975
rect -37681 -47009 -37635 -46975
rect -37601 -47009 -37555 -46975
rect -37521 -47009 -37475 -46975
rect -37441 -47009 -37395 -46975
rect -37361 -47009 -37315 -46975
rect -37281 -47009 -37235 -46975
rect -37201 -47009 -37155 -46975
rect -37121 -47009 -37075 -46975
rect -37041 -47009 -36995 -46975
rect -36961 -47009 -36915 -46975
rect -36881 -47009 -36835 -46975
rect -36801 -47009 -36755 -46975
rect -36721 -47009 -36675 -46975
rect -36641 -47009 -36595 -46975
rect -36561 -47009 -36515 -46975
rect -36481 -47009 -36435 -46975
rect -36401 -47009 -36355 -46975
rect -36321 -47009 -36275 -46975
rect -36241 -47009 -36195 -46975
rect -36161 -47009 -36115 -46975
rect -36081 -47009 -36035 -46975
rect -36001 -47009 -35955 -46975
rect -35921 -47009 -35875 -46975
rect -35841 -47009 -35795 -46975
rect -35761 -47009 -35715 -46975
rect -35681 -47009 -35635 -46975
rect -35601 -47009 -35555 -46975
rect -35521 -47009 -35475 -46975
rect -35441 -47009 -35395 -46975
rect -35361 -47009 -35315 -46975
rect -35281 -47009 -35235 -46975
rect -35201 -47009 -35155 -46975
rect -35121 -47009 -35075 -46975
rect -35041 -47009 -34995 -46975
rect -34961 -47009 -34915 -46975
rect -34881 -47009 -34835 -46975
rect -34801 -47009 -34755 -46975
rect -34721 -47009 -34675 -46975
rect -34641 -47009 -34595 -46975
rect -34561 -47009 -34515 -46975
rect -34481 -47009 -34435 -46975
rect -34401 -47009 -34355 -46975
rect -34321 -47009 -34275 -46975
rect -34241 -47009 -34195 -46975
rect -34161 -47009 -34115 -46975
rect -34081 -47009 -34035 -46975
rect -34001 -47009 -33955 -46975
rect -33921 -47009 -33875 -46975
rect -33841 -47009 -33795 -46975
rect -33761 -47009 -33715 -46975
rect -33681 -47009 -33635 -46975
rect -33601 -47009 -33555 -46975
rect -33521 -47009 -33475 -46975
rect -33441 -47009 -33395 -46975
rect -33361 -47009 -33315 -46975
rect -33281 -47009 -33235 -46975
rect -33201 -47009 -33155 -46975
rect -33121 -47009 -33075 -46975
rect -33041 -47009 -32995 -46975
rect -32961 -47009 -32915 -46975
rect -32881 -47009 -32835 -46975
rect -32801 -47009 -32755 -46975
rect -32721 -47009 -32675 -46975
rect -32641 -47009 -32595 -46975
rect -32561 -47009 -32515 -46975
rect -32481 -47009 -32435 -46975
rect -32401 -47009 -32355 -46975
rect -32321 -47009 -32275 -46975
rect -32241 -47009 -32195 -46975
rect -32161 -47009 -32115 -46975
rect -32081 -47009 -32035 -46975
rect -32001 -47009 -31955 -46975
rect -31921 -47009 -31875 -46975
rect -31841 -47009 -31795 -46975
rect -31761 -47009 -31715 -46975
rect -31681 -47009 -31635 -46975
rect -31601 -47009 -31555 -46975
rect -31521 -47009 -31475 -46975
rect -31441 -47009 -31395 -46975
rect -31361 -47009 -31315 -46975
rect -31281 -47009 -31235 -46975
rect -31201 -47009 -31155 -46975
rect -31121 -47009 -31075 -46975
rect -31041 -47009 -30995 -46975
rect -30961 -47009 -30915 -46975
rect -30881 -47009 -30835 -46975
rect -30801 -47009 -30755 -46975
rect -30721 -47009 -30675 -46975
rect -30641 -47009 -30595 -46975
rect -30561 -47009 -30515 -46975
rect -30481 -47009 -30435 -46975
rect -30401 -47009 -30355 -46975
rect -30321 -47009 -30275 -46975
rect -30241 -47009 -30195 -46975
rect -30161 -47009 -30115 -46975
rect -30081 -47009 -30035 -46975
rect -30001 -47009 -29955 -46975
rect -29921 -47009 -29875 -46975
rect -29841 -47009 -29795 -46975
rect -29761 -47009 -29715 -46975
rect -29681 -47009 -29635 -46975
rect -29601 -47009 -29555 -46975
rect -29521 -47009 -29475 -46975
rect -29441 -47009 -29395 -46975
rect -29361 -47009 -29315 -46975
rect -29281 -47009 -29235 -46975
rect -29201 -47009 -29155 -46975
rect -29121 -47009 -29075 -46975
rect -29041 -47009 -28995 -46975
rect -28961 -47009 -28915 -46975
rect -28881 -47009 -28835 -46975
rect -28801 -47009 -28755 -46975
rect -28721 -47009 -28675 -46975
rect -28641 -47009 -28595 -46975
rect -28561 -47009 -28514 -46975
rect -28480 -47009 -28434 -46975
rect -28400 -47009 -28354 -46975
rect -28320 -47009 -28274 -46975
rect -28240 -47009 -28194 -46975
rect -28160 -47009 -28114 -46975
rect -28080 -47009 -28034 -46975
rect -28000 -47009 -27954 -46975
rect -27920 -47009 -27874 -46975
rect -27840 -47009 -27794 -46975
rect -27760 -47009 -27714 -46975
rect -27680 -47009 -27634 -46975
rect -27600 -47009 -27554 -46975
rect -27520 -47009 -27474 -46975
rect -27440 -47009 -27394 -46975
rect -27360 -47009 -27314 -46975
rect -27280 -47009 -27234 -46975
rect -27200 -47009 -27154 -46975
rect -27120 -47009 -27074 -46975
rect -27040 -47009 -26994 -46975
rect -26960 -47009 -26914 -46975
rect -26880 -47009 -26834 -46975
rect -26800 -47009 -26754 -46975
rect -26720 -47009 -26674 -46975
rect -26640 -47009 -26594 -46975
rect -26560 -47009 -26514 -46975
rect -26480 -47009 -26434 -46975
rect -26400 -47009 -26354 -46975
rect -26320 -47009 -26274 -46975
rect -26240 -47009 -26194 -46975
rect -26160 -47009 -26114 -46975
rect -26080 -47009 -26034 -46975
rect -26000 -47009 -25954 -46975
rect -25920 -47009 -25874 -46975
rect -25840 -47009 -25794 -46975
rect -25760 -47009 -25714 -46975
rect -25680 -47009 -25634 -46975
rect -25600 -47009 -25554 -46975
rect -25520 -47009 -25474 -46975
rect -25440 -47009 -25394 -46975
rect -25360 -47009 -25314 -46975
rect -25280 -47009 -25234 -46975
rect -25200 -47009 -25154 -46975
rect -25120 -47009 -25074 -46975
rect -25040 -47009 -24994 -46975
rect -24960 -47009 -24914 -46975
rect -24880 -47009 -24834 -46975
rect -24800 -47009 -24754 -46975
rect -24720 -47009 -24674 -46975
rect -24640 -47009 -24594 -46975
rect -24560 -47009 -24514 -46975
rect -24480 -47009 -24434 -46975
rect -24400 -47009 -24354 -46975
rect -24320 -47009 -24274 -46975
rect -24240 -47009 -24194 -46975
rect -24160 -47009 -24114 -46975
rect -24080 -47009 -24034 -46975
rect -24000 -47009 -23954 -46975
rect -23920 -47009 -23874 -46975
rect -23840 -47009 -23794 -46975
rect -23760 -47009 -23714 -46975
rect -23680 -47009 -23634 -46975
rect -23600 -47009 -23554 -46975
rect -23520 -47009 -23474 -46975
rect -23440 -47009 -23394 -46975
rect -23360 -47009 -23314 -46975
rect -23280 -47009 -23234 -46975
rect -23200 -47009 -23154 -46975
rect -23120 -47009 -23074 -46975
rect -23040 -47009 -22994 -46975
rect -22960 -47009 -22914 -46975
rect -22880 -47009 -22834 -46975
rect -22800 -47009 -22754 -46975
rect -22720 -47009 -22674 -46975
rect -22640 -47009 -22594 -46975
rect -22560 -47009 -22514 -46975
rect -22480 -47009 -22434 -46975
rect -22400 -47009 -22354 -46975
rect -22320 -47009 -22274 -46975
rect -22240 -47009 -22194 -46975
rect -22160 -47009 -22114 -46975
rect -22080 -47009 -22034 -46975
rect -22000 -47009 -21954 -46975
rect -21920 -47009 -21874 -46975
rect -21840 -47009 -21794 -46975
rect -21760 -47009 -21714 -46975
rect -21680 -47009 -21634 -46975
rect -21600 -47009 -21554 -46975
rect -21520 -47009 -21474 -46975
rect -21440 -47009 -21394 -46975
rect -21360 -47009 -21314 -46975
rect -21280 -47009 -21234 -46975
rect -21200 -47009 -21154 -46975
rect -21120 -47009 -21074 -46975
rect -21040 -47009 -20994 -46975
rect -20960 -47009 -20914 -46975
rect -20880 -47009 -20834 -46975
rect -20800 -47009 -20754 -46975
rect -20720 -47009 -20674 -46975
rect -20640 -47009 -20594 -46975
rect -20560 -47009 -20514 -46975
rect -20480 -47009 -20434 -46975
rect -20400 -47009 -20354 -46975
rect -20320 -47009 -20274 -46975
rect -20240 -47009 -20194 -46975
rect -20160 -47009 -20114 -46975
rect -20080 -47009 -20034 -46975
rect -20000 -47009 -19954 -46975
rect -19920 -47009 -19874 -46975
rect -19840 -47009 -19794 -46975
rect -19760 -47009 -19714 -46975
rect -19680 -47009 -19634 -46975
rect -19600 -47009 -19554 -46975
rect -19520 -47009 -19474 -46975
rect -19440 -47009 -19394 -46975
rect -19360 -47009 -19314 -46975
rect -19280 -47009 -19234 -46975
rect -19200 -47009 -19154 -46975
rect -19120 -47009 -19074 -46975
rect -19040 -47009 -18994 -46975
rect -18960 -47009 -18914 -46975
rect -18880 -47009 -18834 -46975
rect -18800 -47009 -18754 -46975
rect -18720 -47009 -18674 -46975
rect -18640 -47009 -18594 -46975
rect -18560 -47009 -18514 -46975
rect -18480 -47009 -18434 -46975
rect -18400 -47009 -18354 -46975
rect -18320 -47009 -18274 -46975
rect -18240 -47009 -18194 -46975
rect -18160 -47009 -18114 -46975
rect -18080 -47009 -18034 -46975
rect -18000 -47009 -17954 -46975
rect -17920 -47009 -17874 -46975
rect -17840 -47009 -17794 -46975
rect -17760 -47009 -17714 -46975
rect -17680 -47009 -17634 -46975
rect -17600 -47009 -17554 -46975
rect -17520 -47009 -17474 -46975
rect -17440 -47009 -17394 -46975
rect -17360 -47009 -17314 -46975
rect -17280 -47009 -17234 -46975
rect -17200 -47009 -17154 -46975
rect -17120 -47009 -17074 -46975
rect -17040 -47009 -16994 -46975
rect -16960 -47009 -16914 -46975
rect -16880 -47009 -16834 -46975
rect -16800 -47009 -16754 -46975
rect -16720 -47009 -16674 -46975
rect -16640 -47009 -16594 -46975
rect -16560 -47009 -16514 -46975
rect -16480 -47009 -16434 -46975
rect -16400 -47009 -16354 -46975
rect -16320 -47009 -16274 -46975
rect -16240 -47009 -16194 -46975
rect -16160 -47009 -16114 -46975
rect -16080 -47009 -16034 -46975
rect -16000 -47009 -15954 -46975
rect -15920 -47009 -15874 -46975
rect -15840 -47009 -15794 -46975
rect -15760 -47009 -15714 -46975
rect -15680 -47009 -15634 -46975
rect -15600 -47009 -15553 -46975
rect -15519 -47009 -15473 -46975
rect -15439 -47009 -15393 -46975
rect -15359 -47009 -15313 -46975
rect -15279 -47009 -15233 -46975
rect -15199 -47009 -15153 -46975
rect -15119 -47009 -15073 -46975
rect -15039 -47009 -14993 -46975
rect -14959 -47009 -14913 -46975
rect -14879 -47009 -14833 -46975
rect -14799 -47009 -14753 -46975
rect -14719 -47009 -14673 -46975
rect -14639 -47009 -14593 -46975
rect -14559 -47009 -14513 -46975
rect -14479 -47009 -14433 -46975
rect -14399 -47009 -14353 -46975
rect -14319 -47009 -14273 -46975
rect -14239 -47009 -14193 -46975
rect -14159 -47009 -14113 -46975
rect -14079 -47009 -14033 -46975
rect -13999 -47009 -13953 -46975
rect -13919 -47009 -13873 -46975
rect -13839 -47009 -13793 -46975
rect -13759 -47009 -13713 -46975
rect -13679 -47009 -13633 -46975
rect -13599 -47009 -13553 -46975
rect -13519 -47009 -13473 -46975
rect -13439 -47009 -13393 -46975
rect -13359 -47009 -13313 -46975
rect -13279 -47009 -13233 -46975
rect -13199 -47009 -13153 -46975
rect -13119 -47009 -13073 -46975
rect -13039 -47009 -12993 -46975
rect -12959 -47009 -12913 -46975
rect -12879 -47009 -12833 -46975
rect -12799 -47009 -12753 -46975
rect -12719 -47009 -12673 -46975
rect -12639 -47009 -12593 -46975
rect -12559 -47009 -12513 -46975
rect -12479 -47009 -12433 -46975
rect -12399 -47009 -12353 -46975
rect -12319 -47009 -12273 -46975
rect -12239 -47009 -12193 -46975
rect -12159 -47009 -12113 -46975
rect -12079 -47009 -12033 -46975
rect -11999 -47009 -11953 -46975
rect -11919 -47009 -11873 -46975
rect -11839 -47009 -11793 -46975
rect -11759 -47009 -11713 -46975
rect -11679 -47009 -11633 -46975
rect -11599 -47009 -11553 -46975
rect -11519 -47009 -11473 -46975
rect -11439 -47009 -11393 -46975
rect -11359 -47009 -11313 -46975
rect -11279 -47009 -11233 -46975
rect -11199 -47009 -11153 -46975
rect -11119 -47009 -11073 -46975
rect -11039 -47009 -10993 -46975
rect -10959 -47009 -10913 -46975
rect -10879 -47009 -10833 -46975
rect -10799 -47009 -10753 -46975
rect -10719 -47009 -10673 -46975
rect -10639 -47009 -10593 -46975
rect -10559 -47009 -10513 -46975
rect -10479 -47009 -10433 -46975
rect -10399 -47009 -10353 -46975
rect -10319 -47009 -10273 -46975
rect -10239 -47009 -10193 -46975
rect -10159 -47009 -10113 -46975
rect -10079 -47009 -10033 -46975
rect -9999 -47009 -9953 -46975
rect -9919 -47009 -9873 -46975
rect -9839 -47009 -9793 -46975
rect -9759 -47009 -9713 -46975
rect -9679 -47009 -9633 -46975
rect -9599 -47009 -9553 -46975
rect -9519 -47009 -9473 -46975
rect -9439 -47009 -9393 -46975
rect -9359 -47009 -9313 -46975
rect -9279 -47009 -9233 -46975
rect -9199 -47009 -9153 -46975
rect -9119 -47009 -9073 -46975
rect -9039 -47009 -8993 -46975
rect -8959 -47009 -8913 -46975
rect -8879 -47009 -8833 -46975
rect -8799 -47009 -8753 -46975
rect -8719 -47009 -8673 -46975
rect -8639 -47009 -8593 -46975
rect -8559 -47009 -8513 -46975
rect -8479 -47009 -8433 -46975
rect -8399 -47009 -8353 -46975
rect -8319 -47009 -8273 -46975
rect -8239 -47009 -8193 -46975
rect -8159 -47009 -8113 -46975
rect -8079 -47009 -8033 -46975
rect -7999 -47009 -7953 -46975
rect -7919 -47009 -7873 -46975
rect -7839 -47009 -7793 -46975
rect -7759 -47009 -7713 -46975
rect -7679 -47009 -7633 -46975
rect -7599 -47009 -7553 -46975
rect -7519 -47009 -7473 -46975
rect -7439 -47009 -7393 -46975
rect -7359 -47009 -7313 -46975
rect -7279 -47009 -7233 -46975
rect -7199 -47009 -7153 -46975
rect -7119 -47009 -7073 -46975
rect -7039 -47009 -6993 -46975
rect -6959 -47009 -6913 -46975
rect -6879 -47009 -6841 -46975
rect -6807 -47009 -6769 -46975
rect -6735 -47009 -6697 -46975
rect -6663 -47009 -6625 -46975
rect -6591 -47009 -6553 -46975
rect -6519 -47009 -6481 -46975
rect -6447 -47009 -6409 -46975
rect -6375 -47009 -6337 -46975
rect -6303 -47009 -6265 -46975
rect -6231 -47009 -6193 -46975
rect -6159 -47009 -6121 -46975
rect -6087 -47009 -6049 -46975
rect -6015 -47009 -5977 -46975
rect -5943 -47009 -5905 -46975
rect -5871 -47009 -5833 -46975
rect -5799 -47009 -5761 -46975
rect -5727 -47009 -5689 -46975
rect -5655 -47009 -5617 -46975
rect -5583 -47009 -5545 -46975
rect -5511 -47009 -5473 -46975
rect -5439 -47009 -5401 -46975
rect -5367 -47009 -5329 -46975
rect -5295 -47009 -5257 -46975
rect -5223 -47009 -5185 -46975
rect -5151 -47009 -5113 -46975
rect -5079 -47009 -5041 -46975
rect -5007 -47009 -4969 -46975
rect -4935 -47009 -4889 -46975
rect -4855 -47009 -4809 -46975
rect -4775 -47009 -4729 -46975
rect -4695 -47009 -4649 -46975
rect -4615 -47009 -4569 -46975
rect -4535 -47009 -4489 -46975
rect -4455 -47009 -4409 -46975
rect -4375 -47009 -4329 -46975
rect -4295 -47009 -4249 -46975
rect -4215 -47009 -4170 -46975
rect -44481 -47032 -4170 -47009
rect -6805 -47798 -6715 -47032
rect -6360 -47096 -6290 -47080
rect -6360 -47130 -6342 -47096
rect -6307 -47116 -6290 -47096
rect -4956 -47116 -4876 -47096
rect -6307 -47130 -5967 -47116
rect -6360 -47150 -5967 -47130
rect -6307 -47156 -5967 -47150
rect -6307 -47196 -6267 -47156
rect -6007 -47196 -5967 -47156
rect -5707 -47119 -4876 -47116
rect -5707 -47153 -4933 -47119
rect -4899 -47153 -4876 -47119
rect -5707 -47156 -4876 -47153
rect -5707 -47196 -5667 -47156
rect -5407 -47196 -5367 -47156
rect -4956 -47176 -4876 -47156
rect -6805 -47835 -6778 -47798
rect -6744 -47835 -6715 -47798
rect -6805 -47856 -6715 -47835
rect -6597 -47234 -6397 -47196
rect -6597 -47268 -6574 -47234
rect -6540 -47268 -6454 -47234
rect -6420 -47268 -6397 -47234
rect -6597 -47335 -6397 -47268
rect -6597 -47369 -6574 -47335
rect -6540 -47369 -6454 -47335
rect -6420 -47369 -6397 -47335
rect -6597 -47403 -6397 -47369
rect -6597 -47437 -6574 -47403
rect -6540 -47437 -6454 -47403
rect -6420 -47437 -6397 -47403
rect -6597 -47471 -6397 -47437
rect -6597 -47505 -6574 -47471
rect -6540 -47505 -6454 -47471
rect -6420 -47505 -6397 -47471
rect -6597 -47539 -6397 -47505
rect -6597 -47573 -6574 -47539
rect -6540 -47573 -6454 -47539
rect -6420 -47573 -6397 -47539
rect -6597 -47607 -6397 -47573
rect -6597 -47641 -6574 -47607
rect -6540 -47641 -6454 -47607
rect -6420 -47641 -6397 -47607
rect -6597 -47675 -6397 -47641
rect -6597 -47709 -6574 -47675
rect -6540 -47709 -6454 -47675
rect -6420 -47709 -6397 -47675
rect -6597 -47743 -6397 -47709
rect -6597 -47777 -6574 -47743
rect -6540 -47777 -6454 -47743
rect -6420 -47777 -6397 -47743
rect -6597 -47811 -6397 -47777
rect -6597 -47845 -6574 -47811
rect -6540 -47845 -6454 -47811
rect -6420 -47845 -6397 -47811
rect -6597 -47879 -6397 -47845
rect -6597 -47913 -6574 -47879
rect -6540 -47913 -6454 -47879
rect -6420 -47913 -6397 -47879
rect -6597 -47947 -6397 -47913
rect -6597 -47981 -6574 -47947
rect -6540 -47981 -6454 -47947
rect -6420 -47981 -6397 -47947
rect -6597 -48015 -6397 -47981
rect -6597 -48049 -6574 -48015
rect -6540 -48049 -6454 -48015
rect -6420 -48049 -6397 -48015
rect -6597 -48083 -6397 -48049
rect -6597 -48117 -6574 -48083
rect -6540 -48117 -6454 -48083
rect -6420 -48117 -6397 -48083
rect -6597 -48156 -6397 -48117
rect -6327 -47234 -6247 -47196
rect -6327 -47268 -6304 -47234
rect -6270 -47268 -6247 -47234
rect -6327 -47345 -6247 -47268
rect -6327 -47379 -6304 -47345
rect -6270 -47379 -6247 -47345
rect -6327 -47413 -6247 -47379
rect -6327 -47447 -6304 -47413
rect -6270 -47447 -6247 -47413
rect -6327 -47481 -6247 -47447
rect -6327 -47515 -6304 -47481
rect -6270 -47515 -6247 -47481
rect -6327 -47549 -6247 -47515
rect -6327 -47583 -6304 -47549
rect -6270 -47583 -6247 -47549
rect -6327 -47617 -6247 -47583
rect -6327 -47651 -6304 -47617
rect -6270 -47651 -6247 -47617
rect -6327 -47685 -6247 -47651
rect -6327 -47719 -6304 -47685
rect -6270 -47719 -6247 -47685
rect -6327 -47753 -6247 -47719
rect -6327 -47787 -6304 -47753
rect -6270 -47787 -6247 -47753
rect -6327 -47821 -6247 -47787
rect -6327 -47855 -6304 -47821
rect -6270 -47855 -6247 -47821
rect -6327 -47889 -6247 -47855
rect -6327 -47923 -6304 -47889
rect -6270 -47923 -6247 -47889
rect -6327 -47957 -6247 -47923
rect -6327 -47991 -6304 -47957
rect -6270 -47991 -6247 -47957
rect -6327 -48025 -6247 -47991
rect -6327 -48059 -6304 -48025
rect -6270 -48059 -6247 -48025
rect -6327 -48093 -6247 -48059
rect -6327 -48127 -6304 -48093
rect -6270 -48127 -6247 -48093
rect -6327 -48156 -6247 -48127
rect -6177 -47234 -6097 -47196
rect -6177 -47268 -6154 -47234
rect -6120 -47268 -6097 -47234
rect -6177 -47335 -6097 -47268
rect -6177 -47369 -6154 -47335
rect -6120 -47369 -6097 -47335
rect -6177 -47403 -6097 -47369
rect -6177 -47437 -6154 -47403
rect -6120 -47437 -6097 -47403
rect -6177 -47471 -6097 -47437
rect -6177 -47505 -6154 -47471
rect -6120 -47505 -6097 -47471
rect -6177 -47539 -6097 -47505
rect -6177 -47573 -6154 -47539
rect -6120 -47573 -6097 -47539
rect -6177 -47607 -6097 -47573
rect -6177 -47641 -6154 -47607
rect -6120 -47641 -6097 -47607
rect -6177 -47675 -6097 -47641
rect -6177 -47709 -6154 -47675
rect -6120 -47709 -6097 -47675
rect -6177 -47743 -6097 -47709
rect -6177 -47777 -6154 -47743
rect -6120 -47777 -6097 -47743
rect -6177 -47811 -6097 -47777
rect -6177 -47845 -6154 -47811
rect -6120 -47845 -6097 -47811
rect -6177 -47879 -6097 -47845
rect -6177 -47913 -6154 -47879
rect -6120 -47913 -6097 -47879
rect -6177 -47947 -6097 -47913
rect -6177 -47981 -6154 -47947
rect -6120 -47981 -6097 -47947
rect -6177 -48015 -6097 -47981
rect -6177 -48049 -6154 -48015
rect -6120 -48049 -6097 -48015
rect -6177 -48083 -6097 -48049
rect -6177 -48117 -6154 -48083
rect -6120 -48117 -6097 -48083
rect -6177 -48156 -6097 -48117
rect -6027 -47234 -5947 -47196
rect -6027 -47268 -6004 -47234
rect -5970 -47268 -5947 -47234
rect -6027 -47335 -5947 -47268
rect -6027 -47369 -6004 -47335
rect -5970 -47369 -5947 -47335
rect -6027 -47403 -5947 -47369
rect -6027 -47437 -6004 -47403
rect -5970 -47437 -5947 -47403
rect -6027 -47471 -5947 -47437
rect -6027 -47505 -6004 -47471
rect -5970 -47505 -5947 -47471
rect -6027 -47539 -5947 -47505
rect -6027 -47573 -6004 -47539
rect -5970 -47573 -5947 -47539
rect -6027 -47607 -5947 -47573
rect -6027 -47641 -6004 -47607
rect -5970 -47641 -5947 -47607
rect -6027 -47675 -5947 -47641
rect -6027 -47709 -6004 -47675
rect -5970 -47709 -5947 -47675
rect -6027 -47743 -5947 -47709
rect -6027 -47777 -6004 -47743
rect -5970 -47777 -5947 -47743
rect -6027 -47811 -5947 -47777
rect -6027 -47845 -6004 -47811
rect -5970 -47845 -5947 -47811
rect -6027 -47879 -5947 -47845
rect -6027 -47913 -6004 -47879
rect -5970 -47913 -5947 -47879
rect -6027 -47947 -5947 -47913
rect -6027 -47981 -6004 -47947
rect -5970 -47981 -5947 -47947
rect -6027 -48015 -5947 -47981
rect -6027 -48049 -6004 -48015
rect -5970 -48049 -5947 -48015
rect -6027 -48083 -5947 -48049
rect -6027 -48117 -6004 -48083
rect -5970 -48117 -5947 -48083
rect -6027 -48156 -5947 -48117
rect -5877 -47234 -5797 -47196
rect -5877 -47268 -5854 -47234
rect -5820 -47268 -5797 -47234
rect -5877 -47335 -5797 -47268
rect -5877 -47369 -5854 -47335
rect -5820 -47369 -5797 -47335
rect -5877 -47403 -5797 -47369
rect -5877 -47437 -5854 -47403
rect -5820 -47437 -5797 -47403
rect -5877 -47471 -5797 -47437
rect -5877 -47505 -5854 -47471
rect -5820 -47505 -5797 -47471
rect -5877 -47539 -5797 -47505
rect -5877 -47573 -5854 -47539
rect -5820 -47573 -5797 -47539
rect -5877 -47607 -5797 -47573
rect -5877 -47641 -5854 -47607
rect -5820 -47641 -5797 -47607
rect -5877 -47675 -5797 -47641
rect -5877 -47709 -5854 -47675
rect -5820 -47709 -5797 -47675
rect -5877 -47743 -5797 -47709
rect -5877 -47777 -5854 -47743
rect -5820 -47777 -5797 -47743
rect -5877 -47811 -5797 -47777
rect -5877 -47845 -5854 -47811
rect -5820 -47845 -5797 -47811
rect -5877 -47879 -5797 -47845
rect -5877 -47913 -5854 -47879
rect -5820 -47913 -5797 -47879
rect -5877 -47947 -5797 -47913
rect -5877 -47981 -5854 -47947
rect -5820 -47981 -5797 -47947
rect -5877 -48015 -5797 -47981
rect -5877 -48049 -5854 -48015
rect -5820 -48049 -5797 -48015
rect -5877 -48083 -5797 -48049
rect -5877 -48117 -5854 -48083
rect -5820 -48117 -5797 -48083
rect -5877 -48156 -5797 -48117
rect -5727 -47234 -5647 -47196
rect -5727 -47268 -5704 -47234
rect -5670 -47268 -5647 -47234
rect -5727 -47345 -5647 -47268
rect -5727 -47379 -5704 -47345
rect -5670 -47379 -5647 -47345
rect -5727 -47413 -5647 -47379
rect -5727 -47447 -5704 -47413
rect -5670 -47447 -5647 -47413
rect -5727 -47481 -5647 -47447
rect -5727 -47515 -5704 -47481
rect -5670 -47515 -5647 -47481
rect -5727 -47549 -5647 -47515
rect -5727 -47583 -5704 -47549
rect -5670 -47583 -5647 -47549
rect -5727 -47617 -5647 -47583
rect -5727 -47651 -5704 -47617
rect -5670 -47651 -5647 -47617
rect -5727 -47685 -5647 -47651
rect -5727 -47719 -5704 -47685
rect -5670 -47719 -5647 -47685
rect -5727 -47753 -5647 -47719
rect -5727 -47787 -5704 -47753
rect -5670 -47787 -5647 -47753
rect -5727 -47821 -5647 -47787
rect -5727 -47855 -5704 -47821
rect -5670 -47855 -5647 -47821
rect -5727 -47889 -5647 -47855
rect -5727 -47923 -5704 -47889
rect -5670 -47923 -5647 -47889
rect -5727 -47957 -5647 -47923
rect -5727 -47991 -5704 -47957
rect -5670 -47991 -5647 -47957
rect -5727 -48025 -5647 -47991
rect -5727 -48059 -5704 -48025
rect -5670 -48059 -5647 -48025
rect -5727 -48093 -5647 -48059
rect -5727 -48127 -5704 -48093
rect -5670 -48127 -5647 -48093
rect -5727 -48156 -5647 -48127
rect -5577 -47234 -5497 -47196
rect -5577 -47268 -5554 -47234
rect -5520 -47268 -5497 -47234
rect -5577 -47335 -5497 -47268
rect -5577 -47369 -5554 -47335
rect -5520 -47369 -5497 -47335
rect -5577 -47403 -5497 -47369
rect -5577 -47437 -5554 -47403
rect -5520 -47437 -5497 -47403
rect -5577 -47471 -5497 -47437
rect -5577 -47505 -5554 -47471
rect -5520 -47505 -5497 -47471
rect -5577 -47539 -5497 -47505
rect -5577 -47573 -5554 -47539
rect -5520 -47573 -5497 -47539
rect -5577 -47607 -5497 -47573
rect -5577 -47641 -5554 -47607
rect -5520 -47641 -5497 -47607
rect -5577 -47675 -5497 -47641
rect -5577 -47709 -5554 -47675
rect -5520 -47709 -5497 -47675
rect -5577 -47743 -5497 -47709
rect -5577 -47777 -5554 -47743
rect -5520 -47777 -5497 -47743
rect -5577 -47811 -5497 -47777
rect -5577 -47845 -5554 -47811
rect -5520 -47845 -5497 -47811
rect -5577 -47879 -5497 -47845
rect -5577 -47913 -5554 -47879
rect -5520 -47913 -5497 -47879
rect -5577 -47947 -5497 -47913
rect -5577 -47981 -5554 -47947
rect -5520 -47981 -5497 -47947
rect -5577 -48015 -5497 -47981
rect -5577 -48049 -5554 -48015
rect -5520 -48049 -5497 -48015
rect -5577 -48083 -5497 -48049
rect -5577 -48117 -5554 -48083
rect -5520 -48117 -5497 -48083
rect -5577 -48156 -5497 -48117
rect -5427 -47234 -5347 -47196
rect -5427 -47268 -5404 -47234
rect -5370 -47268 -5347 -47234
rect -5427 -47335 -5347 -47268
rect -5427 -47369 -5404 -47335
rect -5370 -47369 -5347 -47335
rect -5427 -47403 -5347 -47369
rect -5427 -47437 -5404 -47403
rect -5370 -47437 -5347 -47403
rect -5427 -47471 -5347 -47437
rect -5427 -47505 -5404 -47471
rect -5370 -47505 -5347 -47471
rect -5427 -47539 -5347 -47505
rect -5427 -47573 -5404 -47539
rect -5370 -47573 -5347 -47539
rect -5427 -47607 -5347 -47573
rect -5427 -47641 -5404 -47607
rect -5370 -47641 -5347 -47607
rect -5427 -47675 -5347 -47641
rect -5427 -47709 -5404 -47675
rect -5370 -47709 -5347 -47675
rect -5427 -47743 -5347 -47709
rect -5427 -47777 -5404 -47743
rect -5370 -47777 -5347 -47743
rect -5427 -47811 -5347 -47777
rect -5427 -47845 -5404 -47811
rect -5370 -47845 -5347 -47811
rect -5427 -47879 -5347 -47845
rect -5427 -47913 -5404 -47879
rect -5370 -47913 -5347 -47879
rect -5427 -47947 -5347 -47913
rect -5427 -47981 -5404 -47947
rect -5370 -47981 -5347 -47947
rect -5427 -48015 -5347 -47981
rect -5427 -48049 -5404 -48015
rect -5370 -48049 -5347 -48015
rect -5427 -48083 -5347 -48049
rect -5427 -48117 -5404 -48083
rect -5370 -48117 -5347 -48083
rect -5427 -48156 -5347 -48117
rect -5277 -47234 -5197 -47196
rect -5277 -47268 -5254 -47234
rect -5220 -47268 -5197 -47234
rect -5277 -47335 -5197 -47268
rect -5277 -47369 -5254 -47335
rect -5220 -47369 -5197 -47335
rect -5277 -47403 -5197 -47369
rect -5277 -47437 -5254 -47403
rect -5220 -47437 -5197 -47403
rect -5277 -47471 -5197 -47437
rect -5277 -47505 -5254 -47471
rect -5220 -47505 -5197 -47471
rect -5277 -47539 -5197 -47505
rect -5277 -47573 -5254 -47539
rect -5220 -47573 -5197 -47539
rect -5277 -47607 -5197 -47573
rect -5277 -47641 -5254 -47607
rect -5220 -47641 -5197 -47607
rect -5277 -47675 -5197 -47641
rect -5277 -47709 -5254 -47675
rect -5220 -47709 -5197 -47675
rect -5277 -47743 -5197 -47709
rect -5277 -47777 -5254 -47743
rect -5220 -47777 -5197 -47743
rect -5277 -47811 -5197 -47777
rect -5277 -47845 -5254 -47811
rect -5220 -47845 -5197 -47811
rect -5277 -47879 -5197 -47845
rect -5277 -47913 -5254 -47879
rect -5220 -47913 -5197 -47879
rect -5277 -47947 -5197 -47913
rect -5277 -47981 -5254 -47947
rect -5220 -47981 -5197 -47947
rect -5277 -48015 -5197 -47981
rect -5277 -48049 -5254 -48015
rect -5220 -48049 -5197 -48015
rect -5277 -48083 -5197 -48049
rect -5277 -48117 -5254 -48083
rect -5220 -48117 -5197 -48083
rect -5277 -48156 -5197 -48117
rect -6457 -48196 -6417 -48156
rect -6157 -48196 -6117 -48156
rect -5857 -48196 -5817 -48156
rect -5557 -48196 -5517 -48156
rect -5257 -48196 -5217 -48156
rect -6789 -48213 -6733 -48210
rect -6789 -48216 -6778 -48213
rect -6744 -48216 -6733 -48213
rect -6805 -48250 -6778 -48216
rect -6744 -48250 -6717 -48216
rect -6457 -48236 -5217 -48196
rect -6457 -48322 -6423 -48236
rect -10124 -48345 -2087 -48322
rect -10124 -48379 -10087 -48345
rect -10053 -48379 -10007 -48345
rect -9973 -48379 -9927 -48345
rect -9893 -48379 -9847 -48345
rect -9813 -48379 -9767 -48345
rect -9733 -48379 -9687 -48345
rect -9653 -48379 -9607 -48345
rect -9573 -48379 -9527 -48345
rect -9493 -48379 -9447 -48345
rect -9413 -48379 -9367 -48345
rect -9333 -48379 -9287 -48345
rect -9253 -48379 -9207 -48345
rect -9173 -48379 -9127 -48345
rect -9093 -48379 -9047 -48345
rect -9013 -48379 -8967 -48345
rect -8933 -48379 -8887 -48345
rect -8853 -48379 -8807 -48345
rect -8773 -48379 -8727 -48345
rect -8693 -48379 -8647 -48345
rect -8613 -48379 -8567 -48345
rect -8533 -48379 -8487 -48345
rect -8453 -48379 -8407 -48345
rect -8373 -48379 -8327 -48345
rect -8293 -48379 -8247 -48345
rect -8213 -48379 -8167 -48345
rect -8133 -48379 -8087 -48345
rect -8053 -48379 -8007 -48345
rect -7973 -48379 -7927 -48345
rect -7893 -48379 -7847 -48345
rect -7813 -48379 -7767 -48345
rect -7733 -48379 -7687 -48345
rect -7653 -48379 -7607 -48345
rect -7573 -48379 -7527 -48345
rect -7493 -48379 -7447 -48345
rect -7413 -48379 -7367 -48345
rect -7333 -48379 -7287 -48345
rect -7253 -48379 -7207 -48345
rect -7173 -48379 -7127 -48345
rect -7093 -48379 -7047 -48345
rect -7013 -48379 -6967 -48345
rect -6933 -48379 -6887 -48345
rect -6853 -48379 -6807 -48345
rect -6773 -48379 -6727 -48345
rect -6693 -48379 -6647 -48345
rect -6613 -48379 -6567 -48345
rect -6533 -48379 -6487 -48345
rect -6453 -48379 -6407 -48345
rect -6373 -48379 -6327 -48345
rect -6293 -48379 -6247 -48345
rect -6213 -48379 -6167 -48345
rect -6133 -48379 -6087 -48345
rect -6053 -48379 -6007 -48345
rect -5973 -48379 -5927 -48345
rect -5893 -48379 -5847 -48345
rect -5813 -48379 -5767 -48345
rect -5733 -48379 -5687 -48345
rect -5653 -48379 -5607 -48345
rect -5573 -48379 -5527 -48345
rect -5493 -48379 -5447 -48345
rect -5413 -48379 -5367 -48345
rect -5333 -48379 -5287 -48345
rect -5253 -48379 -5207 -48345
rect -5173 -48379 -5127 -48345
rect -5093 -48379 -5047 -48345
rect -5013 -48379 -4967 -48345
rect -4933 -48379 -4887 -48345
rect -4853 -48379 -4807 -48345
rect -4773 -48379 -4727 -48345
rect -4693 -48379 -4647 -48345
rect -4613 -48379 -4567 -48345
rect -4533 -48379 -4487 -48345
rect -4453 -48379 -4407 -48345
rect -4373 -48379 -4327 -48345
rect -4293 -48379 -4247 -48345
rect -4213 -48379 -4167 -48345
rect -4133 -48379 -4087 -48345
rect -4053 -48379 -4007 -48345
rect -3973 -48379 -3927 -48345
rect -3893 -48379 -3847 -48345
rect -3813 -48379 -3767 -48345
rect -3733 -48379 -3687 -48345
rect -3653 -48379 -3607 -48345
rect -3573 -48379 -3527 -48345
rect -3493 -48379 -3447 -48345
rect -3413 -48379 -3367 -48345
rect -3333 -48379 -3287 -48345
rect -3253 -48379 -3207 -48345
rect -3173 -48379 -3127 -48345
rect -3093 -48379 -3047 -48345
rect -3013 -48379 -2967 -48345
rect -2933 -48379 -2887 -48345
rect -2853 -48379 -2807 -48345
rect -2773 -48379 -2727 -48345
rect -2693 -48379 -2647 -48345
rect -2613 -48379 -2567 -48345
rect -2533 -48379 -2487 -48345
rect -2453 -48379 -2407 -48345
rect -2373 -48379 -2327 -48345
rect -2293 -48379 -2247 -48345
rect -2213 -48379 -2167 -48345
rect -2133 -48379 -2087 -48345
rect -10124 -48402 -2087 -48379
<< viali >>
rect -44422 -34633 -44388 -34599
rect -44342 -34633 -44308 -34599
rect -44262 -34633 -44228 -34599
rect -44182 -34633 -44148 -34599
rect -44102 -34633 -44068 -34599
rect -44022 -34633 -43988 -34599
rect -43942 -34633 -43908 -34599
rect -43862 -34633 -43828 -34599
rect -43782 -34633 -43748 -34599
rect -43702 -34633 -43668 -34599
rect -43622 -34633 -43588 -34599
rect -43542 -34633 -43508 -34599
rect -43462 -34633 -43428 -34599
rect -43382 -34633 -43348 -34599
rect -43302 -34633 -43268 -34599
rect -43222 -34633 -43188 -34599
rect -43142 -34633 -43108 -34599
rect -43062 -34633 -43028 -34599
rect -42982 -34633 -42948 -34599
rect -42902 -34633 -42868 -34599
rect -42822 -34633 -42788 -34599
rect -42742 -34633 -42708 -34599
rect -42662 -34633 -42628 -34599
rect -42582 -34633 -42548 -34599
rect -42502 -34633 -42468 -34599
rect -42422 -34633 -42388 -34599
rect -42342 -34633 -42308 -34599
rect -42262 -34633 -42228 -34599
rect -42182 -34633 -42148 -34599
rect -42102 -34633 -42068 -34599
rect -42022 -34633 -41988 -34599
rect -41942 -34633 -41908 -34599
rect -41862 -34633 -41828 -34599
rect -41782 -34633 -41748 -34599
rect -41702 -34633 -41668 -34599
rect -41622 -34633 -41588 -34599
rect -41542 -34633 -41508 -34599
rect -41462 -34633 -41428 -34599
rect -41382 -34633 -41348 -34599
rect -41302 -34633 -41268 -34599
rect -41222 -34633 -41188 -34599
rect -41142 -34633 -41108 -34599
rect -41062 -34633 -41028 -34599
rect -40982 -34633 -40948 -34599
rect -40902 -34633 -40868 -34599
rect -40822 -34633 -40788 -34599
rect -40742 -34633 -40708 -34599
rect -40662 -34633 -40628 -34599
rect -40582 -34633 -40548 -34599
rect -40502 -34633 -40468 -34599
rect -40422 -34633 -40388 -34599
rect -40342 -34633 -40308 -34599
rect -40262 -34633 -40228 -34599
rect -40182 -34633 -40148 -34599
rect -40102 -34633 -40068 -34599
rect -40022 -34633 -39988 -34599
rect -39942 -34633 -39908 -34599
rect -39862 -34633 -39828 -34599
rect -39782 -34633 -39748 -34599
rect -39702 -34633 -39668 -34599
rect -39622 -34633 -39588 -34599
rect -39542 -34633 -39508 -34599
rect -39462 -34633 -39428 -34599
rect -39382 -34633 -39348 -34599
rect -39302 -34633 -39268 -34599
rect -39222 -34633 -39188 -34599
rect -39142 -34633 -39108 -34599
rect -39062 -34633 -39028 -34599
rect -38982 -34633 -38948 -34599
rect -38902 -34633 -38868 -34599
rect -38822 -34633 -38788 -34599
rect -38742 -34633 -38708 -34599
rect -38662 -34633 -38628 -34599
rect -38582 -34633 -38548 -34599
rect -38502 -34633 -38468 -34599
rect -38422 -34633 -38388 -34599
rect -38342 -34633 -38308 -34599
rect -38262 -34633 -38228 -34599
rect -38182 -34633 -38148 -34599
rect -38102 -34633 -38068 -34599
rect -38022 -34633 -37988 -34599
rect -37942 -34633 -37908 -34599
rect -37862 -34633 -37828 -34599
rect -37782 -34633 -37748 -34599
rect -37702 -34633 -37668 -34599
rect -37622 -34633 -37588 -34599
rect -37542 -34633 -37508 -34599
rect -37462 -34633 -37428 -34599
rect -37382 -34633 -37348 -34599
rect -37302 -34633 -37268 -34599
rect -37222 -34633 -37188 -34599
rect -37142 -34633 -37108 -34599
rect -37062 -34633 -37028 -34599
rect -36982 -34633 -36948 -34599
rect -36902 -34633 -36868 -34599
rect -36822 -34633 -36788 -34599
rect -36742 -34633 -36708 -34599
rect -36662 -34633 -36628 -34599
rect -36582 -34633 -36548 -34599
rect -36502 -34633 -36468 -34599
rect -36422 -34633 -36388 -34599
rect -36342 -34633 -36308 -34599
rect -36262 -34633 -36228 -34599
rect -36182 -34633 -36148 -34599
rect -36102 -34633 -36068 -34599
rect -36022 -34633 -35988 -34599
rect -35942 -34633 -35908 -34599
rect -35862 -34633 -35828 -34599
rect -35782 -34633 -35748 -34599
rect -35702 -34633 -35668 -34599
rect -35622 -34633 -35588 -34599
rect -35542 -34633 -35508 -34599
rect -35462 -34633 -35428 -34599
rect -35382 -34633 -35348 -34599
rect -35302 -34633 -35268 -34599
rect -35222 -34633 -35188 -34599
rect -35142 -34633 -35108 -34599
rect -35062 -34633 -35028 -34599
rect -34982 -34633 -34948 -34599
rect -34902 -34633 -34868 -34599
rect -34822 -34633 -34788 -34599
rect -34742 -34633 -34708 -34599
rect -34662 -34633 -34628 -34599
rect -34582 -34633 -34548 -34599
rect -34502 -34633 -34468 -34599
rect -34422 -34633 -34388 -34599
rect -34342 -34633 -34308 -34599
rect -34262 -34633 -34228 -34599
rect -34182 -34633 -34148 -34599
rect -34102 -34633 -34068 -34599
rect -34022 -34633 -33988 -34599
rect -33942 -34633 -33908 -34599
rect -33862 -34633 -33828 -34599
rect -33782 -34633 -33748 -34599
rect -33702 -34633 -33668 -34599
rect -33622 -34633 -33588 -34599
rect -33542 -34633 -33508 -34599
rect -33462 -34633 -33428 -34599
rect -33382 -34633 -33348 -34599
rect -33302 -34633 -33268 -34599
rect -33222 -34633 -33188 -34599
rect -33142 -34633 -33108 -34599
rect -33062 -34633 -33028 -34599
rect -32982 -34633 -32948 -34599
rect -32902 -34633 -32868 -34599
rect -32822 -34633 -32788 -34599
rect -32742 -34633 -32708 -34599
rect -32662 -34633 -32628 -34599
rect -32582 -34633 -32548 -34599
rect -32502 -34633 -32468 -34599
rect -32422 -34633 -32388 -34599
rect -32342 -34633 -32308 -34599
rect -32262 -34633 -32228 -34599
rect -32182 -34633 -32148 -34599
rect -32102 -34633 -32068 -34599
rect -32022 -34633 -31988 -34599
rect -31942 -34633 -31908 -34599
rect -31862 -34633 -31828 -34599
rect -31782 -34633 -31748 -34599
rect -31702 -34633 -31668 -34599
rect -31622 -34633 -31588 -34599
rect -31542 -34633 -31508 -34599
rect -31461 -34633 -31427 -34599
rect -31381 -34633 -31347 -34599
rect -31301 -34633 -31267 -34599
rect -31221 -34633 -31187 -34599
rect -31141 -34633 -31107 -34599
rect -31061 -34633 -31027 -34599
rect -30981 -34633 -30947 -34599
rect -30901 -34633 -30867 -34599
rect -30821 -34633 -30787 -34599
rect -30741 -34633 -30707 -34599
rect -30661 -34633 -30627 -34599
rect -30581 -34633 -30547 -34599
rect -30501 -34633 -30467 -34599
rect -30421 -34633 -30387 -34599
rect -30341 -34633 -30307 -34599
rect -30261 -34633 -30227 -34599
rect -30181 -34633 -30147 -34599
rect -30101 -34633 -30067 -34599
rect -30021 -34633 -29987 -34599
rect -29941 -34633 -29907 -34599
rect -29861 -34633 -29827 -34599
rect -29781 -34633 -29747 -34599
rect -29701 -34633 -29667 -34599
rect -29621 -34633 -29587 -34599
rect -29541 -34633 -29507 -34599
rect -29461 -34633 -29427 -34599
rect -29381 -34633 -29347 -34599
rect -29301 -34633 -29267 -34599
rect -29221 -34633 -29187 -34599
rect -29141 -34633 -29107 -34599
rect -29061 -34633 -29027 -34599
rect -28981 -34633 -28947 -34599
rect -28901 -34633 -28867 -34599
rect -28821 -34633 -28787 -34599
rect -28741 -34633 -28707 -34599
rect -28661 -34633 -28627 -34599
rect -28581 -34633 -28547 -34599
rect -28501 -34633 -28467 -34599
rect -28421 -34633 -28387 -34599
rect -28341 -34633 -28307 -34599
rect -28261 -34633 -28227 -34599
rect -28181 -34633 -28147 -34599
rect -28101 -34633 -28067 -34599
rect -28021 -34633 -27987 -34599
rect -27941 -34633 -27907 -34599
rect -27861 -34633 -27827 -34599
rect -27781 -34633 -27747 -34599
rect -27701 -34633 -27667 -34599
rect -27621 -34633 -27587 -34599
rect -27541 -34633 -27507 -34599
rect -27461 -34633 -27427 -34599
rect -27381 -34633 -27347 -34599
rect -27301 -34633 -27267 -34599
rect -27221 -34633 -27187 -34599
rect -27141 -34633 -27107 -34599
rect -27061 -34633 -27027 -34599
rect -26981 -34633 -26947 -34599
rect -26901 -34633 -26867 -34599
rect -26821 -34633 -26787 -34599
rect -26741 -34633 -26707 -34599
rect -26661 -34633 -26627 -34599
rect -26581 -34633 -26547 -34599
rect -26501 -34633 -26467 -34599
rect -26421 -34633 -26387 -34599
rect -26341 -34633 -26307 -34599
rect -26261 -34633 -26227 -34599
rect -26181 -34633 -26147 -34599
rect -26101 -34633 -26067 -34599
rect -26021 -34633 -25987 -34599
rect -25941 -34633 -25907 -34599
rect -25861 -34633 -25827 -34599
rect -25781 -34633 -25747 -34599
rect -25701 -34633 -25667 -34599
rect -25621 -34633 -25587 -34599
rect -25541 -34633 -25507 -34599
rect -25461 -34633 -25427 -34599
rect -25381 -34633 -25347 -34599
rect -25301 -34633 -25267 -34599
rect -25221 -34633 -25187 -34599
rect -25141 -34633 -25107 -34599
rect -25061 -34633 -25027 -34599
rect -24981 -34633 -24947 -34599
rect -24901 -34633 -24867 -34599
rect -24821 -34633 -24787 -34599
rect -24741 -34633 -24707 -34599
rect -24661 -34633 -24627 -34599
rect -24581 -34633 -24547 -34599
rect -24501 -34633 -24467 -34599
rect -24421 -34633 -24387 -34599
rect -24341 -34633 -24307 -34599
rect -24261 -34633 -24227 -34599
rect -24181 -34633 -24147 -34599
rect -24101 -34633 -24067 -34599
rect -24021 -34633 -23987 -34599
rect -23941 -34633 -23907 -34599
rect -23861 -34633 -23827 -34599
rect -23781 -34633 -23747 -34599
rect -23701 -34633 -23667 -34599
rect -23621 -34633 -23587 -34599
rect -23541 -34633 -23507 -34599
rect -23461 -34633 -23427 -34599
rect -23381 -34633 -23347 -34599
rect -23301 -34633 -23267 -34599
rect -23221 -34633 -23187 -34599
rect -23141 -34633 -23107 -34599
rect -23061 -34633 -23027 -34599
rect -22981 -34633 -22947 -34599
rect -22901 -34633 -22867 -34599
rect -22821 -34633 -22787 -34599
rect -22741 -34633 -22707 -34599
rect -22661 -34633 -22627 -34599
rect -22581 -34633 -22547 -34599
rect -22501 -34633 -22467 -34599
rect -22421 -34633 -22387 -34599
rect -22341 -34633 -22307 -34599
rect -22261 -34633 -22227 -34599
rect -22181 -34633 -22147 -34599
rect -22101 -34633 -22067 -34599
rect -22021 -34633 -21987 -34599
rect -21941 -34633 -21907 -34599
rect -21861 -34633 -21827 -34599
rect -21781 -34633 -21747 -34599
rect -21701 -34633 -21667 -34599
rect -21621 -34633 -21587 -34599
rect -21541 -34633 -21507 -34599
rect -21461 -34633 -21427 -34599
rect -21381 -34633 -21347 -34599
rect -21301 -34633 -21267 -34599
rect -21221 -34633 -21187 -34599
rect -21141 -34633 -21107 -34599
rect -21061 -34633 -21027 -34599
rect -20981 -34633 -20947 -34599
rect -20901 -34633 -20867 -34599
rect -20821 -34633 -20787 -34599
rect -20741 -34633 -20707 -34599
rect -20661 -34633 -20627 -34599
rect -20581 -34633 -20547 -34599
rect -20501 -34633 -20467 -34599
rect -20421 -34633 -20387 -34599
rect -20341 -34633 -20307 -34599
rect -20261 -34633 -20227 -34599
rect -20181 -34633 -20147 -34599
rect -20101 -34633 -20067 -34599
rect -20021 -34633 -19987 -34599
rect -19941 -34633 -19907 -34599
rect -19861 -34633 -19827 -34599
rect -19781 -34633 -19747 -34599
rect -19701 -34633 -19667 -34599
rect -19621 -34633 -19587 -34599
rect -19541 -34633 -19507 -34599
rect -19461 -34633 -19427 -34599
rect -19381 -34633 -19347 -34599
rect -19301 -34633 -19267 -34599
rect -19221 -34633 -19187 -34599
rect -19141 -34633 -19107 -34599
rect -19061 -34633 -19027 -34599
rect -18981 -34633 -18947 -34599
rect -18901 -34633 -18867 -34599
rect -18821 -34633 -18787 -34599
rect -18741 -34633 -18707 -34599
rect -18661 -34633 -18627 -34599
rect -18581 -34633 -18547 -34599
rect -18500 -34633 -18466 -34599
rect -18420 -34633 -18386 -34599
rect -18340 -34633 -18306 -34599
rect -18260 -34633 -18226 -34599
rect -18180 -34633 -18146 -34599
rect -18100 -34633 -18066 -34599
rect -18020 -34633 -17986 -34599
rect -17940 -34633 -17906 -34599
rect -17860 -34633 -17826 -34599
rect -17780 -34633 -17746 -34599
rect -17700 -34633 -17666 -34599
rect -17620 -34633 -17586 -34599
rect -17540 -34633 -17506 -34599
rect -17460 -34633 -17426 -34599
rect -17380 -34633 -17346 -34599
rect -17300 -34633 -17266 -34599
rect -17220 -34633 -17186 -34599
rect -17140 -34633 -17106 -34599
rect -17060 -34633 -17026 -34599
rect -16980 -34633 -16946 -34599
rect -16900 -34633 -16866 -34599
rect -16820 -34633 -16786 -34599
rect -16740 -34633 -16706 -34599
rect -16660 -34633 -16626 -34599
rect -16580 -34633 -16546 -34599
rect -16500 -34633 -16466 -34599
rect -16420 -34633 -16386 -34599
rect -16340 -34633 -16306 -34599
rect -16260 -34633 -16226 -34599
rect -16180 -34633 -16146 -34599
rect -16100 -34633 -16066 -34599
rect -16020 -34633 -15986 -34599
rect -15940 -34633 -15906 -34599
rect -15860 -34633 -15826 -34599
rect -15780 -34633 -15746 -34599
rect -15700 -34633 -15666 -34599
rect -15620 -34633 -15586 -34599
rect -15540 -34633 -15506 -34599
rect -15460 -34633 -15426 -34599
rect -15380 -34633 -15346 -34599
rect -15300 -34633 -15266 -34599
rect -15220 -34633 -15186 -34599
rect -15140 -34633 -15106 -34599
rect -15060 -34633 -15026 -34599
rect -14980 -34633 -14946 -34599
rect -14900 -34633 -14866 -34599
rect -14820 -34633 -14786 -34599
rect -14740 -34633 -14706 -34599
rect -14660 -34633 -14626 -34599
rect -14580 -34633 -14546 -34599
rect -14500 -34633 -14466 -34599
rect -14420 -34633 -14386 -34599
rect -14340 -34633 -14306 -34599
rect -14260 -34633 -14226 -34599
rect -14180 -34633 -14146 -34599
rect -14100 -34633 -14066 -34599
rect -14020 -34633 -13986 -34599
rect -13940 -34633 -13906 -34599
rect -13860 -34633 -13826 -34599
rect -13780 -34633 -13746 -34599
rect -13700 -34633 -13666 -34599
rect -13620 -34633 -13586 -34599
rect -13540 -34633 -13506 -34599
rect -13460 -34633 -13426 -34599
rect -13380 -34633 -13346 -34599
rect -13300 -34633 -13266 -34599
rect -13220 -34633 -13186 -34599
rect -13140 -34633 -13106 -34599
rect -13060 -34633 -13026 -34599
rect -12980 -34633 -12946 -34599
rect -12900 -34633 -12866 -34599
rect -12820 -34633 -12786 -34599
rect -12740 -34633 -12706 -34599
rect -12660 -34633 -12626 -34599
rect -12580 -34633 -12546 -34599
rect -12500 -34633 -12466 -34599
rect -12420 -34633 -12386 -34599
rect -12340 -34633 -12306 -34599
rect -12260 -34633 -12226 -34599
rect -12180 -34633 -12146 -34599
rect -12100 -34633 -12066 -34599
rect -12020 -34633 -11986 -34599
rect -11940 -34633 -11906 -34599
rect -11860 -34633 -11826 -34599
rect -11780 -34633 -11746 -34599
rect -11700 -34633 -11666 -34599
rect -11620 -34633 -11586 -34599
rect -11540 -34633 -11506 -34599
rect -11460 -34633 -11426 -34599
rect -11380 -34633 -11346 -34599
rect -11300 -34633 -11266 -34599
rect -11220 -34633 -11186 -34599
rect -11140 -34633 -11106 -34599
rect -11060 -34633 -11026 -34599
rect -10980 -34633 -10946 -34599
rect -10900 -34633 -10866 -34599
rect -10820 -34633 -10786 -34599
rect -10740 -34633 -10706 -34599
rect -10660 -34633 -10626 -34599
rect -10580 -34633 -10546 -34599
rect -10500 -34633 -10466 -34599
rect -10420 -34633 -10386 -34599
rect -10340 -34633 -10306 -34599
rect -10260 -34633 -10226 -34599
rect -10180 -34633 -10146 -34599
rect -10100 -34633 -10066 -34599
rect -10020 -34633 -9986 -34599
rect -9940 -34633 -9906 -34599
rect -9859 -34633 -9825 -34599
rect -9779 -34633 -9745 -34599
rect -9699 -34633 -9665 -34599
rect -9619 -34633 -9585 -34599
rect -9539 -34633 -9505 -34599
rect -9459 -34633 -9425 -34599
rect -9379 -34633 -9345 -34599
rect -9299 -34633 -9265 -34599
rect -9219 -34633 -9185 -34599
rect -9139 -34633 -9105 -34599
rect -9059 -34633 -9025 -34599
rect -8979 -34633 -8945 -34599
rect -8899 -34633 -8865 -34599
rect -8819 -34633 -8785 -34599
rect -8739 -34633 -8705 -34599
rect -8659 -34633 -8625 -34599
rect -8579 -34633 -8545 -34599
rect -8499 -34633 -8465 -34599
rect -8419 -34633 -8385 -34599
rect -8339 -34633 -8305 -34599
rect -8259 -34633 -8225 -34599
rect -8179 -34633 -8145 -34599
rect -8099 -34633 -8065 -34599
rect -8019 -34633 -7985 -34599
rect -7939 -34633 -7905 -34599
rect -7859 -34633 -7825 -34599
rect -7779 -34633 -7745 -34599
rect -7699 -34633 -7665 -34599
rect -7619 -34633 -7585 -34599
rect -7539 -34633 -7505 -34599
rect -7459 -34633 -7425 -34599
rect -7379 -34633 -7345 -34599
rect -7299 -34633 -7265 -34599
rect -7219 -34633 -7185 -34599
rect -7139 -34633 -7105 -34599
rect -7059 -34633 -7025 -34599
rect -6979 -34633 -6945 -34599
rect -6899 -34633 -6865 -34599
rect -6819 -34633 -6785 -34599
rect -6739 -34633 -6705 -34599
rect -6659 -34633 -6625 -34599
rect -6579 -34633 -6545 -34599
rect -6499 -34633 -6465 -34599
rect -6419 -34633 -6385 -34599
rect -6339 -34633 -6305 -34599
rect -6259 -34633 -6225 -34599
rect -6179 -34633 -6145 -34599
rect -6099 -34633 -6065 -34599
rect -6019 -34633 -5985 -34599
rect -5939 -34633 -5905 -34599
rect -5859 -34633 -5825 -34599
rect -5779 -34633 -5745 -34599
rect -5699 -34633 -5665 -34599
rect -5619 -34633 -5585 -34599
rect -5539 -34633 -5505 -34599
rect -5459 -34633 -5425 -34599
rect -5379 -34633 -5345 -34599
rect -5299 -34633 -5265 -34599
rect -5219 -34633 -5185 -34599
rect -5139 -34633 -5105 -34599
rect -5059 -34633 -5025 -34599
rect -4979 -34633 -4945 -34599
rect -4899 -34633 -4865 -34599
rect -4819 -34633 -4785 -34599
rect -4739 -34633 -4705 -34599
rect -4659 -34633 -4625 -34599
rect -4579 -34633 -4545 -34599
rect -4499 -34633 -4465 -34599
rect -4419 -34633 -4385 -34599
rect -4339 -34633 -4305 -34599
rect -4259 -34633 -4225 -34599
rect -4140 -34633 -4106 -34599
rect -4060 -34633 -4026 -34599
rect -3980 -34633 -3946 -34599
rect -3900 -34633 -3866 -34599
rect -3820 -34633 -3786 -34599
rect -3740 -34633 -3706 -34599
rect -3660 -34633 -3626 -34599
rect -3580 -34633 -3546 -34599
rect -3500 -34633 -3466 -34599
rect -3420 -34633 -3386 -34599
rect -3340 -34633 -3306 -34599
rect -3260 -34633 -3226 -34599
rect -3180 -34633 -3146 -34599
rect -3100 -34633 -3066 -34599
rect -3020 -34633 -2986 -34599
rect -2940 -34633 -2906 -34599
rect -2860 -34633 -2826 -34599
rect -2780 -34633 -2746 -34599
rect -2700 -34633 -2666 -34599
rect -2620 -34633 -2586 -34599
rect -2540 -34633 -2506 -34599
rect -2460 -34633 -2426 -34599
rect -2380 -34633 -2346 -34599
rect -2300 -34633 -2266 -34599
rect -2220 -34633 -2186 -34599
rect -2140 -34633 -2106 -34599
rect -2060 -34633 -2026 -34599
rect -1980 -34633 -1946 -34599
rect -1900 -34633 -1866 -34599
rect -1820 -34633 -1786 -34599
rect -1740 -34633 -1706 -34599
rect -1660 -34633 -1626 -34599
rect -1580 -34633 -1546 -34599
rect -1500 -34633 -1466 -34599
rect -1420 -34633 -1386 -34599
rect -1340 -34633 -1306 -34599
rect -1260 -34633 -1226 -34599
rect -1180 -34633 -1146 -34599
rect -1100 -34633 -1066 -34599
rect -1020 -34633 -986 -34599
rect -940 -34633 -906 -34599
rect -860 -34633 -826 -34599
rect -780 -34633 -746 -34599
rect -700 -34633 -666 -34599
rect -620 -34633 -586 -34599
rect -540 -34633 -506 -34599
rect -460 -34633 -426 -34599
rect -380 -34633 -346 -34599
rect -300 -34633 -266 -34599
rect -220 -34633 -186 -34599
rect -140 -34633 -106 -34599
rect -60 -34633 -26 -34599
rect 20 -34633 54 -34599
rect 100 -34633 134 -34599
rect 180 -34633 214 -34599
rect 260 -34633 294 -34599
rect 340 -34633 374 -34599
rect 420 -34633 454 -34599
rect 500 -34633 534 -34599
rect 580 -34633 614 -34599
rect 660 -34633 694 -34599
rect 740 -34633 774 -34599
rect 820 -34633 854 -34599
rect 900 -34633 934 -34599
rect 980 -34633 1014 -34599
rect 1060 -34633 1094 -34599
rect 1140 -34633 1174 -34599
rect 1220 -34633 1254 -34599
rect 1300 -34633 1334 -34599
rect 1380 -34633 1414 -34599
rect 1460 -34633 1494 -34599
rect 1540 -34633 1574 -34599
rect 1620 -34633 1654 -34599
rect 1700 -34633 1734 -34599
rect 1780 -34633 1814 -34599
rect 1860 -34633 1894 -34599
rect 1940 -34633 1974 -34599
rect 2020 -34633 2054 -34599
rect 2100 -34633 2134 -34599
rect 2180 -34633 2214 -34599
rect 2260 -34633 2294 -34599
rect 2340 -34633 2374 -34599
rect 2420 -34633 2454 -34599
rect 2500 -34633 2534 -34599
rect 2580 -34633 2614 -34599
rect 2660 -34633 2694 -34599
rect 2740 -34633 2774 -34599
rect 2820 -34633 2854 -34599
rect 2900 -34633 2934 -34599
rect 2980 -34633 3014 -34599
rect 3060 -34633 3094 -34599
rect 3140 -34633 3174 -34599
rect 3220 -34633 3254 -34599
rect 3300 -34633 3334 -34599
rect 3380 -34633 3414 -34599
rect 3460 -34633 3494 -34599
rect 3540 -34633 3574 -34599
rect 3620 -34633 3654 -34599
rect 3700 -34633 3734 -34599
rect 3780 -34633 3814 -34599
rect 3860 -34633 3894 -34599
rect 3940 -34633 3974 -34599
rect 4020 -34633 4054 -34599
rect 4100 -34633 4134 -34599
rect 4180 -34633 4214 -34599
rect 4260 -34633 4294 -34599
rect 4340 -34633 4374 -34599
rect 4420 -34633 4454 -34599
rect 4500 -34633 4534 -34599
rect 4580 -34633 4614 -34599
rect 4660 -34633 4694 -34599
rect 4740 -34633 4774 -34599
rect 4820 -34633 4854 -34599
rect 4900 -34633 4934 -34599
rect 4980 -34633 5014 -34599
rect 5060 -34633 5094 -34599
rect 5140 -34633 5174 -34599
rect 5220 -34633 5254 -34599
rect 5300 -34633 5334 -34599
rect 5380 -34633 5414 -34599
rect 5460 -34633 5494 -34599
rect 5540 -34633 5574 -34599
rect 5620 -34633 5654 -34599
rect 5700 -34633 5734 -34599
rect 5780 -34633 5814 -34599
rect 5860 -34633 5894 -34599
rect 5940 -34633 5974 -34599
rect 6020 -34633 6054 -34599
rect 6100 -34633 6134 -34599
rect 6180 -34633 6214 -34599
rect 6260 -34633 6294 -34599
rect 6340 -34633 6374 -34599
rect 6420 -34633 6454 -34599
rect 6500 -34633 6534 -34599
rect 6580 -34633 6614 -34599
rect 6660 -34633 6694 -34599
rect 6740 -34633 6774 -34599
rect 6820 -34633 6854 -34599
rect 6900 -34633 6934 -34599
rect 6980 -34633 7014 -34599
rect 7060 -34633 7094 -34599
rect 7140 -34633 7174 -34599
rect 7220 -34633 7254 -34599
rect 7300 -34633 7334 -34599
rect 7380 -34633 7414 -34599
rect 7460 -34633 7494 -34599
rect 7540 -34633 7574 -34599
rect 7620 -34633 7654 -34599
rect 7700 -34633 7734 -34599
rect 7780 -34633 7814 -34599
rect 7860 -34633 7894 -34599
rect 7940 -34633 7974 -34599
rect 8020 -34633 8054 -34599
rect 8100 -34633 8134 -34599
rect 8180 -34633 8214 -34599
rect 8260 -34633 8294 -34599
rect 8340 -34633 8374 -34599
rect 8420 -34633 8454 -34599
rect 8500 -34633 8534 -34599
rect 8580 -34633 8614 -34599
rect 8660 -34633 8694 -34599
rect 8740 -34633 8774 -34599
rect 8820 -34633 8854 -34599
rect 8900 -34633 8934 -34599
rect 8980 -34633 9014 -34599
rect 9060 -34633 9094 -34599
rect 9140 -34633 9174 -34599
rect 9220 -34633 9254 -34599
rect 9300 -34633 9334 -34599
rect 9380 -34633 9414 -34599
rect 9460 -34633 9494 -34599
rect 9540 -34633 9574 -34599
rect 9620 -34633 9654 -34599
rect 9700 -34633 9734 -34599
rect 9780 -34633 9814 -34599
rect 9860 -34633 9894 -34599
rect 9940 -34633 9974 -34599
rect 10020 -34633 10054 -34599
rect 10100 -34633 10134 -34599
rect 10181 -34633 10215 -34599
rect 10261 -34633 10295 -34599
rect 10341 -34633 10375 -34599
rect 10421 -34633 10455 -34599
rect 10501 -34633 10535 -34599
rect 10581 -34633 10615 -34599
rect 10661 -34633 10695 -34599
rect 10741 -34633 10775 -34599
rect 10821 -34633 10855 -34599
rect 10901 -34633 10935 -34599
rect 10981 -34633 11015 -34599
rect 11061 -34633 11095 -34599
rect 11141 -34633 11175 -34599
rect 11221 -34633 11255 -34599
rect 11301 -34633 11335 -34599
rect 11381 -34633 11415 -34599
rect 11461 -34633 11495 -34599
rect 11541 -34633 11575 -34599
rect 11621 -34633 11655 -34599
rect 11701 -34633 11735 -34599
rect 11781 -34633 11815 -34599
rect 11861 -34633 11895 -34599
rect 11941 -34633 11975 -34599
rect 12021 -34633 12055 -34599
rect 12101 -34633 12135 -34599
rect 12181 -34633 12215 -34599
rect 12261 -34633 12295 -34599
rect 12341 -34633 12375 -34599
rect 12421 -34633 12455 -34599
rect 12501 -34633 12535 -34599
rect 12581 -34633 12615 -34599
rect 12661 -34633 12695 -34599
rect 12741 -34633 12775 -34599
rect 12821 -34633 12855 -34599
rect 12901 -34633 12935 -34599
rect 12981 -34633 13015 -34599
rect 13061 -34633 13095 -34599
rect 13141 -34633 13175 -34599
rect 13221 -34633 13255 -34599
rect 13301 -34633 13335 -34599
rect 13381 -34633 13415 -34599
rect 13461 -34633 13495 -34599
rect 13541 -34633 13575 -34599
rect 13621 -34633 13655 -34599
rect 13701 -34633 13735 -34599
rect 13781 -34633 13815 -34599
rect 13861 -34633 13895 -34599
rect 13941 -34633 13975 -34599
rect 14021 -34633 14055 -34599
rect 14101 -34633 14135 -34599
rect 14181 -34633 14215 -34599
rect 14261 -34633 14295 -34599
rect 14341 -34633 14375 -34599
rect 14421 -34633 14455 -34599
rect 14501 -34633 14535 -34599
rect 14581 -34633 14615 -34599
rect 14661 -34633 14695 -34599
rect 14741 -34633 14775 -34599
rect 14821 -34633 14855 -34599
rect 14901 -34633 14935 -34599
rect 14981 -34633 15015 -34599
rect 15061 -34633 15095 -34599
rect 15141 -34633 15175 -34599
rect 15221 -34633 15255 -34599
rect 15301 -34633 15335 -34599
rect 15381 -34633 15415 -34599
rect 15461 -34633 15495 -34599
rect 15541 -34633 15575 -34599
rect 15621 -34633 15655 -34599
rect 15701 -34633 15735 -34599
rect 15781 -34633 15815 -34599
rect 15861 -34633 15895 -34599
rect 15941 -34633 15975 -34599
rect 16021 -34633 16055 -34599
rect 16101 -34633 16135 -34599
rect 16181 -34633 16215 -34599
rect 16261 -34633 16295 -34599
rect 16341 -34633 16375 -34599
rect 16421 -34633 16455 -34599
rect 16501 -34633 16535 -34599
rect 16581 -34633 16615 -34599
rect 16661 -34633 16695 -34599
rect 16741 -34633 16775 -34599
rect 16821 -34633 16855 -34599
rect 16901 -34633 16935 -34599
rect 16981 -34633 17015 -34599
rect 17061 -34633 17095 -34599
rect 17141 -34633 17175 -34599
rect 17221 -34633 17255 -34599
rect 17301 -34633 17335 -34599
rect 17381 -34633 17415 -34599
rect 17461 -34633 17495 -34599
rect 17541 -34633 17575 -34599
rect 17621 -34633 17655 -34599
rect 17701 -34633 17735 -34599
rect 17781 -34633 17815 -34599
rect 17861 -34633 17895 -34599
rect 17941 -34633 17975 -34599
rect 18021 -34633 18055 -34599
rect 18101 -34633 18135 -34599
rect 18181 -34633 18215 -34599
rect 18261 -34633 18295 -34599
rect 18341 -34633 18375 -34599
rect 18421 -34633 18455 -34599
rect 18501 -34633 18535 -34599
rect 18581 -34633 18615 -34599
rect 18661 -34633 18695 -34599
rect 18741 -34633 18775 -34599
rect 18821 -34633 18855 -34599
rect 18901 -34633 18935 -34599
rect 18981 -34633 19015 -34599
rect 19061 -34633 19095 -34599
rect 19141 -34633 19175 -34599
rect 19221 -34633 19255 -34599
rect 19301 -34633 19335 -34599
rect 19381 -34633 19415 -34599
rect 19461 -34633 19495 -34599
rect 19541 -34633 19575 -34599
rect 19621 -34633 19655 -34599
rect 19701 -34633 19735 -34599
rect 19781 -34633 19815 -34599
rect 19861 -34633 19895 -34599
rect 19941 -34633 19975 -34599
rect 20021 -34633 20055 -34599
rect 20101 -34633 20135 -34599
rect 20181 -34633 20215 -34599
rect 20261 -34633 20295 -34599
rect 20341 -34633 20375 -34599
rect 20421 -34633 20455 -34599
rect 20501 -34633 20535 -34599
rect 20581 -34633 20615 -34599
rect 20661 -34633 20695 -34599
rect 20741 -34633 20775 -34599
rect 20821 -34633 20855 -34599
rect 20901 -34633 20935 -34599
rect 20981 -34633 21015 -34599
rect 21061 -34633 21095 -34599
rect 21141 -34633 21175 -34599
rect 21221 -34633 21255 -34599
rect 21301 -34633 21335 -34599
rect 21381 -34633 21415 -34599
rect 21461 -34633 21495 -34599
rect 21541 -34633 21575 -34599
rect 21621 -34633 21655 -34599
rect 21701 -34633 21735 -34599
rect 21781 -34633 21815 -34599
rect 21861 -34633 21895 -34599
rect 21941 -34633 21975 -34599
rect 22021 -34633 22055 -34599
rect 22101 -34633 22135 -34599
rect 22181 -34633 22215 -34599
rect 22261 -34633 22295 -34599
rect 22341 -34633 22375 -34599
rect 22421 -34633 22455 -34599
rect 22501 -34633 22535 -34599
rect 22581 -34633 22615 -34599
rect 22661 -34633 22695 -34599
rect 22741 -34633 22775 -34599
rect 22821 -34633 22855 -34599
rect 22901 -34633 22935 -34599
rect 22981 -34633 23015 -34599
rect 23061 -34633 23095 -34599
rect 23141 -34633 23175 -34599
rect 23221 -34633 23255 -34599
rect 23301 -34633 23335 -34599
rect 23381 -34633 23415 -34599
rect 23461 -34633 23495 -34599
rect 23541 -34633 23575 -34599
rect 23621 -34633 23655 -34599
rect 23701 -34633 23735 -34599
rect 23781 -34633 23815 -34599
rect 23861 -34633 23895 -34599
rect 23941 -34633 23975 -34599
rect 24021 -34633 24055 -34599
rect 24101 -34633 24135 -34599
rect 24181 -34633 24215 -34599
rect 24261 -34633 24295 -34599
rect 24341 -34633 24375 -34599
rect 24421 -34633 24455 -34599
rect 24501 -34633 24535 -34599
rect 24581 -34633 24615 -34599
rect 24661 -34633 24695 -34599
rect 24741 -34633 24775 -34599
rect 24821 -34633 24855 -34599
rect 24901 -34633 24935 -34599
rect 24981 -34633 25015 -34599
rect 25061 -34633 25095 -34599
rect 25141 -34633 25175 -34599
rect 25221 -34633 25255 -34599
rect 25301 -34633 25335 -34599
rect 25381 -34633 25415 -34599
rect 25461 -34633 25495 -34599
rect 25541 -34633 25575 -34599
rect 25621 -34633 25655 -34599
rect 25701 -34633 25735 -34599
rect 25781 -34633 25815 -34599
rect 25861 -34633 25895 -34599
rect 25941 -34633 25975 -34599
rect 26021 -34633 26055 -34599
rect 26101 -34633 26135 -34599
rect 26181 -34633 26215 -34599
rect 26261 -34633 26295 -34599
rect 26341 -34633 26375 -34599
rect 26421 -34633 26455 -34599
rect 26501 -34633 26535 -34599
rect 26581 -34633 26615 -34599
rect 26661 -34633 26695 -34599
rect 26741 -34633 26775 -34599
rect 26821 -34633 26855 -34599
rect 26901 -34633 26935 -34599
rect 26981 -34633 27015 -34599
rect 27061 -34633 27095 -34599
rect 27141 -34633 27175 -34599
rect 27221 -34633 27255 -34599
rect 27301 -34633 27335 -34599
rect 27381 -34633 27415 -34599
rect 27461 -34633 27495 -34599
rect 27541 -34633 27575 -34599
rect 27621 -34633 27655 -34599
rect 27701 -34633 27735 -34599
rect 27781 -34633 27815 -34599
rect 27861 -34633 27895 -34599
rect 27941 -34633 27975 -34599
rect 28021 -34633 28055 -34599
rect 28101 -34633 28135 -34599
rect 28181 -34633 28215 -34599
rect 28261 -34633 28295 -34599
rect 28341 -34633 28375 -34599
rect 28421 -34633 28455 -34599
rect 28501 -34633 28535 -34599
rect 28581 -34633 28615 -34599
rect 28661 -34633 28695 -34599
rect 28741 -34633 28775 -34599
rect 28821 -34633 28855 -34599
rect 28901 -34633 28935 -34599
rect 28981 -34633 29015 -34599
rect 29061 -34633 29095 -34599
rect 29141 -34633 29175 -34599
rect 29221 -34633 29255 -34599
rect 29301 -34633 29335 -34599
rect 29381 -34633 29415 -34599
rect 29461 -34633 29495 -34599
rect 29541 -34633 29575 -34599
rect 29621 -34633 29655 -34599
rect 29701 -34633 29735 -34599
rect 29781 -34633 29815 -34599
rect 29861 -34633 29895 -34599
rect 29941 -34633 29975 -34599
rect 30021 -34633 30055 -34599
rect 30101 -34633 30135 -34599
rect 30181 -34633 30215 -34599
rect 30261 -34633 30295 -34599
rect 30341 -34633 30375 -34599
rect 30421 -34633 30455 -34599
rect 30501 -34633 30535 -34599
rect 30581 -34633 30615 -34599
rect 30661 -34633 30695 -34599
rect 30741 -34633 30775 -34599
rect 30821 -34633 30855 -34599
rect 30901 -34633 30935 -34599
rect 30981 -34633 31015 -34599
rect 31061 -34633 31095 -34599
rect 31141 -34633 31175 -34599
rect 31221 -34633 31255 -34599
rect 31301 -34633 31335 -34599
rect 31381 -34633 31415 -34599
rect 31461 -34633 31495 -34599
rect 31541 -34633 31575 -34599
rect 31621 -34633 31655 -34599
rect 31701 -34633 31735 -34599
rect -27231 -34753 -27197 -34719
rect -27111 -34753 -27077 -34719
rect 12104 -34754 12138 -34720
rect 12224 -34754 12258 -34720
rect -27231 -34873 -27197 -34839
rect -27111 -34873 -27077 -34839
rect 12104 -34874 12138 -34840
rect 12224 -34874 12258 -34840
rect -44422 -42492 -44388 -42458
rect -44342 -42492 -44308 -42458
rect -44262 -42492 -44228 -42458
rect -44182 -42492 -44148 -42458
rect -44102 -42492 -44068 -42458
rect -44022 -42492 -43988 -42458
rect -43942 -42492 -43908 -42458
rect -43862 -42492 -43828 -42458
rect -43782 -42492 -43748 -42458
rect -43702 -42492 -43668 -42458
rect -43622 -42492 -43588 -42458
rect -43542 -42492 -43508 -42458
rect -43462 -42492 -43428 -42458
rect -43382 -42492 -43348 -42458
rect -43302 -42492 -43268 -42458
rect -43222 -42492 -43188 -42458
rect -43142 -42492 -43108 -42458
rect -43062 -42492 -43028 -42458
rect -42982 -42492 -42948 -42458
rect -42902 -42492 -42868 -42458
rect -42822 -42492 -42788 -42458
rect -42742 -42492 -42708 -42458
rect -42662 -42492 -42628 -42458
rect -42582 -42492 -42548 -42458
rect -42502 -42492 -42468 -42458
rect -42422 -42492 -42388 -42458
rect -42342 -42492 -42308 -42458
rect -42262 -42492 -42228 -42458
rect -42182 -42492 -42148 -42458
rect -42102 -42492 -42068 -42458
rect -42022 -42492 -41988 -42458
rect -41942 -42492 -41908 -42458
rect -41862 -42492 -41828 -42458
rect -41782 -42492 -41748 -42458
rect -41702 -42492 -41668 -42458
rect -41622 -42492 -41588 -42458
rect -41542 -42492 -41508 -42458
rect -41462 -42492 -41428 -42458
rect -41382 -42492 -41348 -42458
rect -41302 -42492 -41268 -42458
rect -41222 -42492 -41188 -42458
rect -41142 -42492 -41108 -42458
rect -41062 -42492 -41028 -42458
rect -40982 -42492 -40948 -42458
rect -40902 -42492 -40868 -42458
rect -40822 -42492 -40788 -42458
rect -40742 -42492 -40708 -42458
rect -40662 -42492 -40628 -42458
rect -40582 -42492 -40548 -42458
rect -40502 -42492 -40468 -42458
rect -40422 -42492 -40388 -42458
rect -40342 -42492 -40308 -42458
rect -40262 -42492 -40228 -42458
rect -40182 -42492 -40148 -42458
rect -40102 -42492 -40068 -42458
rect -40022 -42492 -39988 -42458
rect -39942 -42492 -39908 -42458
rect -39862 -42492 -39828 -42458
rect -39782 -42492 -39748 -42458
rect -39702 -42492 -39668 -42458
rect -39622 -42492 -39588 -42458
rect -39542 -42492 -39508 -42458
rect -39462 -42492 -39428 -42458
rect -39382 -42492 -39348 -42458
rect -39302 -42492 -39268 -42458
rect -39222 -42492 -39188 -42458
rect -39142 -42492 -39108 -42458
rect -39062 -42492 -39028 -42458
rect -38982 -42492 -38948 -42458
rect -38902 -42492 -38868 -42458
rect -38822 -42492 -38788 -42458
rect -38742 -42492 -38708 -42458
rect -38662 -42492 -38628 -42458
rect -38582 -42492 -38548 -42458
rect -38502 -42492 -38468 -42458
rect -38422 -42492 -38388 -42458
rect -38342 -42492 -38308 -42458
rect -38262 -42492 -38228 -42458
rect -38182 -42492 -38148 -42458
rect -38102 -42492 -38068 -42458
rect -38022 -42492 -37988 -42458
rect -37942 -42492 -37908 -42458
rect -37862 -42492 -37828 -42458
rect -37782 -42492 -37748 -42458
rect -37702 -42492 -37668 -42458
rect -37622 -42492 -37588 -42458
rect -37542 -42492 -37508 -42458
rect -37462 -42492 -37428 -42458
rect -37382 -42492 -37348 -42458
rect -37302 -42492 -37268 -42458
rect -37222 -42492 -37188 -42458
rect -37142 -42492 -37108 -42458
rect -37062 -42492 -37028 -42458
rect -36982 -42492 -36948 -42458
rect -36902 -42492 -36868 -42458
rect -36822 -42492 -36788 -42458
rect -36742 -42492 -36708 -42458
rect -36662 -42492 -36628 -42458
rect -36582 -42492 -36548 -42458
rect -36502 -42492 -36468 -42458
rect -36422 -42492 -36388 -42458
rect -36342 -42492 -36308 -42458
rect -36262 -42492 -36228 -42458
rect -36182 -42492 -36148 -42458
rect -36102 -42492 -36068 -42458
rect -36022 -42492 -35988 -42458
rect -35942 -42492 -35908 -42458
rect -35862 -42492 -35828 -42458
rect -35782 -42492 -35748 -42458
rect -35702 -42492 -35668 -42458
rect -35622 -42492 -35588 -42458
rect -35542 -42492 -35508 -42458
rect -35462 -42492 -35428 -42458
rect -35382 -42492 -35348 -42458
rect -35302 -42492 -35268 -42458
rect -35222 -42492 -35188 -42458
rect -35142 -42492 -35108 -42458
rect -35062 -42492 -35028 -42458
rect -34982 -42492 -34948 -42458
rect -34902 -42492 -34868 -42458
rect -34822 -42492 -34788 -42458
rect -34742 -42492 -34708 -42458
rect -34662 -42492 -34628 -42458
rect -34582 -42492 -34548 -42458
rect -34502 -42492 -34468 -42458
rect -34422 -42492 -34388 -42458
rect -34342 -42492 -34308 -42458
rect -34262 -42492 -34228 -42458
rect -34182 -42492 -34148 -42458
rect -34102 -42492 -34068 -42458
rect -34022 -42492 -33988 -42458
rect -33942 -42492 -33908 -42458
rect -33862 -42492 -33828 -42458
rect -33782 -42492 -33748 -42458
rect -33702 -42492 -33668 -42458
rect -33622 -42492 -33588 -42458
rect -33542 -42492 -33508 -42458
rect -33462 -42492 -33428 -42458
rect -33382 -42492 -33348 -42458
rect -33302 -42492 -33268 -42458
rect -33222 -42492 -33188 -42458
rect -33142 -42492 -33108 -42458
rect -33062 -42492 -33028 -42458
rect -32982 -42492 -32948 -42458
rect -32902 -42492 -32868 -42458
rect -32822 -42492 -32788 -42458
rect -32742 -42492 -32708 -42458
rect -32662 -42492 -32628 -42458
rect -32582 -42492 -32548 -42458
rect -32502 -42492 -32468 -42458
rect -32422 -42492 -32388 -42458
rect -32342 -42492 -32308 -42458
rect -32262 -42492 -32228 -42458
rect -32182 -42492 -32148 -42458
rect -32102 -42492 -32068 -42458
rect -32022 -42492 -31988 -42458
rect -31942 -42492 -31908 -42458
rect -31862 -42492 -31828 -42458
rect -31782 -42492 -31748 -42458
rect -31702 -42492 -31668 -42458
rect -31622 -42492 -31588 -42458
rect -31542 -42492 -31508 -42458
rect -31461 -42492 -31427 -42458
rect -31381 -42492 -31347 -42458
rect -31301 -42492 -31267 -42458
rect -31221 -42492 -31187 -42458
rect -31141 -42492 -31107 -42458
rect -31061 -42492 -31027 -42458
rect -30981 -42492 -30947 -42458
rect -30901 -42492 -30867 -42458
rect -30821 -42492 -30787 -42458
rect -30741 -42492 -30707 -42458
rect -30661 -42492 -30627 -42458
rect -30581 -42492 -30547 -42458
rect -30501 -42492 -30467 -42458
rect -30421 -42492 -30387 -42458
rect -30341 -42492 -30307 -42458
rect -30261 -42492 -30227 -42458
rect -30181 -42492 -30147 -42458
rect -30101 -42492 -30067 -42458
rect -30021 -42492 -29987 -42458
rect -29941 -42492 -29907 -42458
rect -29861 -42492 -29827 -42458
rect -29781 -42492 -29747 -42458
rect -29701 -42492 -29667 -42458
rect -29621 -42492 -29587 -42458
rect -29541 -42492 -29507 -42458
rect -29461 -42492 -29427 -42458
rect -29381 -42492 -29347 -42458
rect -29301 -42492 -29267 -42458
rect -29221 -42492 -29187 -42458
rect -29141 -42492 -29107 -42458
rect -29061 -42492 -29027 -42458
rect -28981 -42492 -28947 -42458
rect -28901 -42492 -28867 -42458
rect -28821 -42492 -28787 -42458
rect -28741 -42492 -28707 -42458
rect -28661 -42492 -28627 -42458
rect -28581 -42492 -28547 -42458
rect -28501 -42492 -28467 -42458
rect -28421 -42492 -28387 -42458
rect -28341 -42492 -28307 -42458
rect -28261 -42492 -28227 -42458
rect -28181 -42492 -28147 -42458
rect -28101 -42492 -28067 -42458
rect -28021 -42492 -27987 -42458
rect -27941 -42492 -27907 -42458
rect -27861 -42492 -27827 -42458
rect -27781 -42492 -27747 -42458
rect -27701 -42492 -27667 -42458
rect -27621 -42492 -27587 -42458
rect -27541 -42492 -27507 -42458
rect -27461 -42492 -27427 -42458
rect -27381 -42492 -27347 -42458
rect -27301 -42492 -27267 -42458
rect -27221 -42492 -27187 -42458
rect -27141 -42492 -27107 -42458
rect -27061 -42492 -27027 -42458
rect -26981 -42492 -26947 -42458
rect -26901 -42492 -26867 -42458
rect -26821 -42492 -26787 -42458
rect -26741 -42492 -26707 -42458
rect -26661 -42492 -26627 -42458
rect -26581 -42492 -26547 -42458
rect -26501 -42492 -26467 -42458
rect -26421 -42492 -26387 -42458
rect -26341 -42492 -26307 -42458
rect -26261 -42492 -26227 -42458
rect -26181 -42492 -26147 -42458
rect -26101 -42492 -26067 -42458
rect -26021 -42492 -25987 -42458
rect -25941 -42492 -25907 -42458
rect -25861 -42492 -25827 -42458
rect -25781 -42492 -25747 -42458
rect -25701 -42492 -25667 -42458
rect -25621 -42492 -25587 -42458
rect -25541 -42492 -25507 -42458
rect -25461 -42492 -25427 -42458
rect -25381 -42492 -25347 -42458
rect -25301 -42492 -25267 -42458
rect -25221 -42492 -25187 -42458
rect -25141 -42492 -25107 -42458
rect -25061 -42492 -25027 -42458
rect -24981 -42492 -24947 -42458
rect -24901 -42492 -24867 -42458
rect -24821 -42492 -24787 -42458
rect -24741 -42492 -24707 -42458
rect -24661 -42492 -24627 -42458
rect -24581 -42492 -24547 -42458
rect -24501 -42492 -24467 -42458
rect -24421 -42492 -24387 -42458
rect -24341 -42492 -24307 -42458
rect -24261 -42492 -24227 -42458
rect -24181 -42492 -24147 -42458
rect -24101 -42492 -24067 -42458
rect -24021 -42492 -23987 -42458
rect -23941 -42492 -23907 -42458
rect -23861 -42492 -23827 -42458
rect -23781 -42492 -23747 -42458
rect -23701 -42492 -23667 -42458
rect -23621 -42492 -23587 -42458
rect -23541 -42492 -23507 -42458
rect -23461 -42492 -23427 -42458
rect -23381 -42492 -23347 -42458
rect -23301 -42492 -23267 -42458
rect -23221 -42492 -23187 -42458
rect -23141 -42492 -23107 -42458
rect -23061 -42492 -23027 -42458
rect -22981 -42492 -22947 -42458
rect -22901 -42492 -22867 -42458
rect -22821 -42492 -22787 -42458
rect -22741 -42492 -22707 -42458
rect -22661 -42492 -22627 -42458
rect -22581 -42492 -22547 -42458
rect -22501 -42492 -22467 -42458
rect -22421 -42492 -22387 -42458
rect -22341 -42492 -22307 -42458
rect -22261 -42492 -22227 -42458
rect -22181 -42492 -22147 -42458
rect -22101 -42492 -22067 -42458
rect -22021 -42492 -21987 -42458
rect -21941 -42492 -21907 -42458
rect -21861 -42492 -21827 -42458
rect -21781 -42492 -21747 -42458
rect -21701 -42492 -21667 -42458
rect -21621 -42492 -21587 -42458
rect -21541 -42492 -21507 -42458
rect -21461 -42492 -21427 -42458
rect -21381 -42492 -21347 -42458
rect -21301 -42492 -21267 -42458
rect -21221 -42492 -21187 -42458
rect -21141 -42492 -21107 -42458
rect -21061 -42492 -21027 -42458
rect -20981 -42492 -20947 -42458
rect -20901 -42492 -20867 -42458
rect -20821 -42492 -20787 -42458
rect -20741 -42492 -20707 -42458
rect -20661 -42492 -20627 -42458
rect -20581 -42492 -20547 -42458
rect -20501 -42492 -20467 -42458
rect -20421 -42492 -20387 -42458
rect -20341 -42492 -20307 -42458
rect -20261 -42492 -20227 -42458
rect -20181 -42492 -20147 -42458
rect -20101 -42492 -20067 -42458
rect -20021 -42492 -19987 -42458
rect -19941 -42492 -19907 -42458
rect -19861 -42492 -19827 -42458
rect -19781 -42492 -19747 -42458
rect -19701 -42492 -19667 -42458
rect -19621 -42492 -19587 -42458
rect -19541 -42492 -19507 -42458
rect -19461 -42492 -19427 -42458
rect -19381 -42492 -19347 -42458
rect -19301 -42492 -19267 -42458
rect -19221 -42492 -19187 -42458
rect -19141 -42492 -19107 -42458
rect -19061 -42492 -19027 -42458
rect -18981 -42492 -18947 -42458
rect -18901 -42492 -18867 -42458
rect -18821 -42492 -18787 -42458
rect -18741 -42492 -18707 -42458
rect -18661 -42492 -18627 -42458
rect -18581 -42492 -18547 -42458
rect -18500 -42492 -18466 -42458
rect -18420 -42492 -18386 -42458
rect -18340 -42492 -18306 -42458
rect -18260 -42492 -18226 -42458
rect -18180 -42492 -18146 -42458
rect -18100 -42492 -18066 -42458
rect -18020 -42492 -17986 -42458
rect -17940 -42492 -17906 -42458
rect -17860 -42492 -17826 -42458
rect -17780 -42492 -17746 -42458
rect -17700 -42492 -17666 -42458
rect -17620 -42492 -17586 -42458
rect -17540 -42492 -17506 -42458
rect -17460 -42492 -17426 -42458
rect -17380 -42492 -17346 -42458
rect -17300 -42492 -17266 -42458
rect -17220 -42492 -17186 -42458
rect -17140 -42492 -17106 -42458
rect -17060 -42492 -17026 -42458
rect -16980 -42492 -16946 -42458
rect -16900 -42492 -16866 -42458
rect -16820 -42492 -16786 -42458
rect -16740 -42492 -16706 -42458
rect -16660 -42492 -16626 -42458
rect -16580 -42492 -16546 -42458
rect -16500 -42492 -16466 -42458
rect -16420 -42492 -16386 -42458
rect -16340 -42492 -16306 -42458
rect -16260 -42492 -16226 -42458
rect -16180 -42492 -16146 -42458
rect -16100 -42492 -16066 -42458
rect -16020 -42492 -15986 -42458
rect -15940 -42492 -15906 -42458
rect -15860 -42492 -15826 -42458
rect -15780 -42492 -15746 -42458
rect -15700 -42492 -15666 -42458
rect -15620 -42492 -15586 -42458
rect -15540 -42492 -15506 -42458
rect -15460 -42492 -15426 -42458
rect -15380 -42492 -15346 -42458
rect -15300 -42492 -15266 -42458
rect -15220 -42492 -15186 -42458
rect -15140 -42492 -15106 -42458
rect -15060 -42492 -15026 -42458
rect -14980 -42492 -14946 -42458
rect -14900 -42492 -14866 -42458
rect -14820 -42492 -14786 -42458
rect -14740 -42492 -14706 -42458
rect -14660 -42492 -14626 -42458
rect -14580 -42492 -14546 -42458
rect -14500 -42492 -14466 -42458
rect -14420 -42492 -14386 -42458
rect -14340 -42492 -14306 -42458
rect -14260 -42492 -14226 -42458
rect -14180 -42492 -14146 -42458
rect -14100 -42492 -14066 -42458
rect -14020 -42492 -13986 -42458
rect -13940 -42492 -13906 -42458
rect -13860 -42492 -13826 -42458
rect -13780 -42492 -13746 -42458
rect -13700 -42492 -13666 -42458
rect -13620 -42492 -13586 -42458
rect -13540 -42492 -13506 -42458
rect -13460 -42492 -13426 -42458
rect -13380 -42492 -13346 -42458
rect -13300 -42492 -13266 -42458
rect -13220 -42492 -13186 -42458
rect -13140 -42492 -13106 -42458
rect -13060 -42492 -13026 -42458
rect -12980 -42492 -12946 -42458
rect -12900 -42492 -12866 -42458
rect -12820 -42492 -12786 -42458
rect -12740 -42492 -12706 -42458
rect -12660 -42492 -12626 -42458
rect -12580 -42492 -12546 -42458
rect -12500 -42492 -12466 -42458
rect -12420 -42492 -12386 -42458
rect -12340 -42492 -12306 -42458
rect -12260 -42492 -12226 -42458
rect -12180 -42492 -12146 -42458
rect -12100 -42492 -12066 -42458
rect -12020 -42492 -11986 -42458
rect -11940 -42492 -11906 -42458
rect -11860 -42492 -11826 -42458
rect -11780 -42492 -11746 -42458
rect -11700 -42492 -11666 -42458
rect -11620 -42492 -11586 -42458
rect -11540 -42492 -11506 -42458
rect -11460 -42492 -11426 -42458
rect -11380 -42492 -11346 -42458
rect -11300 -42492 -11266 -42458
rect -11220 -42492 -11186 -42458
rect -11140 -42492 -11106 -42458
rect -11060 -42492 -11026 -42458
rect -10980 -42492 -10946 -42458
rect -10900 -42492 -10866 -42458
rect -10820 -42492 -10786 -42458
rect -10740 -42492 -10706 -42458
rect -10660 -42492 -10626 -42458
rect -10580 -42492 -10546 -42458
rect -10500 -42492 -10466 -42458
rect -10420 -42492 -10386 -42458
rect -10340 -42492 -10306 -42458
rect -10260 -42492 -10226 -42458
rect -10180 -42492 -10146 -42458
rect -10100 -42492 -10066 -42458
rect -10020 -42492 -9986 -42458
rect -9940 -42492 -9906 -42458
rect -9859 -42492 -9825 -42458
rect -9779 -42492 -9745 -42458
rect -9699 -42492 -9665 -42458
rect -9619 -42492 -9585 -42458
rect -9539 -42492 -9505 -42458
rect -9459 -42492 -9425 -42458
rect -9379 -42492 -9345 -42458
rect -9299 -42492 -9265 -42458
rect -9219 -42492 -9185 -42458
rect -9139 -42492 -9105 -42458
rect -9059 -42492 -9025 -42458
rect -8979 -42492 -8945 -42458
rect -8899 -42492 -8865 -42458
rect -8819 -42492 -8785 -42458
rect -8739 -42492 -8705 -42458
rect -8659 -42492 -8625 -42458
rect -8579 -42492 -8545 -42458
rect -8499 -42492 -8465 -42458
rect -8419 -42492 -8385 -42458
rect -8339 -42492 -8305 -42458
rect -8259 -42492 -8225 -42458
rect -8179 -42492 -8145 -42458
rect -8099 -42492 -8065 -42458
rect -8019 -42492 -7985 -42458
rect -7939 -42492 -7905 -42458
rect -7859 -42492 -7825 -42458
rect -7779 -42492 -7745 -42458
rect -7699 -42492 -7665 -42458
rect -7619 -42492 -7585 -42458
rect -7539 -42492 -7505 -42458
rect -7459 -42492 -7425 -42458
rect -7379 -42492 -7345 -42458
rect -7299 -42492 -7265 -42458
rect -7219 -42492 -7185 -42458
rect -7139 -42492 -7105 -42458
rect -7059 -42492 -7025 -42458
rect -6979 -42492 -6945 -42458
rect -6899 -42492 -6865 -42458
rect -6819 -42492 -6785 -42458
rect -6739 -42492 -6705 -42458
rect -6659 -42492 -6625 -42458
rect -6579 -42492 -6545 -42458
rect -6499 -42492 -6465 -42458
rect -6419 -42492 -6385 -42458
rect -6339 -42492 -6305 -42458
rect -6259 -42492 -6225 -42458
rect -6179 -42492 -6145 -42458
rect -6099 -42492 -6065 -42458
rect -6019 -42492 -5985 -42458
rect -5939 -42492 -5905 -42458
rect -5859 -42492 -5825 -42458
rect -5779 -42492 -5745 -42458
rect -5699 -42492 -5665 -42458
rect -5619 -42492 -5585 -42458
rect -5539 -42492 -5505 -42458
rect -5459 -42492 -5425 -42458
rect -5379 -42492 -5345 -42458
rect -5299 -42492 -5265 -42458
rect -5219 -42492 -5185 -42458
rect -5139 -42492 -5105 -42458
rect -5059 -42492 -5025 -42458
rect -4979 -42492 -4945 -42458
rect -4899 -42492 -4865 -42458
rect -4819 -42492 -4785 -42458
rect -4739 -42492 -4705 -42458
rect -4659 -42492 -4625 -42458
rect -4579 -42492 -4545 -42458
rect -4499 -42492 -4465 -42458
rect -4419 -42492 -4385 -42458
rect -4339 -42492 -4305 -42458
rect -4259 -42492 -4225 -42458
rect -4140 -42492 -4106 -42458
rect -4060 -42492 -4026 -42458
rect -3980 -42492 -3946 -42458
rect -3900 -42492 -3866 -42458
rect -3820 -42492 -3786 -42458
rect -3740 -42492 -3706 -42458
rect -3660 -42492 -3626 -42458
rect -3580 -42492 -3546 -42458
rect -3500 -42492 -3466 -42458
rect -3420 -42492 -3386 -42458
rect -3340 -42492 -3306 -42458
rect -3260 -42492 -3226 -42458
rect -3180 -42492 -3146 -42458
rect -3100 -42492 -3066 -42458
rect -3020 -42492 -2986 -42458
rect -2940 -42492 -2906 -42458
rect -2860 -42492 -2826 -42458
rect -2780 -42492 -2746 -42458
rect -2700 -42492 -2666 -42458
rect -2620 -42492 -2586 -42458
rect -2540 -42492 -2506 -42458
rect -2460 -42492 -2426 -42458
rect -2380 -42492 -2346 -42458
rect -2300 -42492 -2266 -42458
rect -2220 -42492 -2186 -42458
rect -2140 -42492 -2106 -42458
rect -2060 -42492 -2026 -42458
rect -1980 -42492 -1946 -42458
rect -1900 -42492 -1866 -42458
rect -1820 -42492 -1786 -42458
rect -1740 -42492 -1706 -42458
rect -1660 -42492 -1626 -42458
rect -1580 -42492 -1546 -42458
rect -1500 -42492 -1466 -42458
rect -1420 -42492 -1386 -42458
rect -1340 -42492 -1306 -42458
rect -1260 -42492 -1226 -42458
rect -1180 -42492 -1146 -42458
rect -1100 -42492 -1066 -42458
rect -1020 -42492 -986 -42458
rect -940 -42492 -906 -42458
rect -860 -42492 -826 -42458
rect -780 -42492 -746 -42458
rect -700 -42492 -666 -42458
rect -10377 -43766 -10343 -43763
rect -10257 -43766 -10223 -43763
rect -10379 -43797 -10343 -43766
rect -10259 -43797 -10223 -43766
rect -10379 -43800 -10345 -43797
rect -10259 -43800 -10225 -43797
rect -10377 -43886 -10343 -43883
rect -10257 -43886 -10223 -43883
rect -10379 -43917 -10343 -43886
rect -10259 -43917 -10223 -43886
rect -7841 -42744 -7807 -42710
rect -7841 -42816 -7807 -42782
rect -7841 -42888 -7807 -42854
rect -7841 -42960 -7807 -42926
rect -7841 -43032 -7807 -42998
rect -8132 -43087 -8098 -43053
rect -7841 -43104 -7807 -43070
rect -8735 -43268 -8701 -43234
rect -8615 -43268 -8581 -43234
rect -8735 -43388 -8701 -43354
rect -8615 -43388 -8581 -43354
rect -8681 -43690 -8641 -43650
rect -10379 -43920 -10345 -43917
rect -10259 -43920 -10225 -43917
rect -7523 -42744 -7489 -42710
rect -7523 -42816 -7489 -42782
rect -7523 -42888 -7489 -42854
rect -7523 -42960 -7489 -42926
rect -7523 -43032 -7489 -42998
rect -7523 -43104 -7489 -43070
rect -7205 -42744 -7171 -42710
rect -7205 -42816 -7171 -42782
rect -7205 -42888 -7171 -42854
rect -7205 -42960 -7171 -42926
rect -7205 -43032 -7171 -42998
rect -7205 -43104 -7171 -43070
rect -6887 -42744 -6853 -42710
rect -6887 -42816 -6853 -42782
rect -6887 -42888 -6853 -42854
rect -6887 -42960 -6853 -42926
rect -6887 -43032 -6853 -42998
rect -6887 -43104 -6853 -43070
rect -7841 -43313 -7807 -43279
rect -7841 -43385 -7807 -43351
rect -7841 -43457 -7807 -43423
rect -7841 -43529 -7807 -43495
rect -7841 -43601 -7807 -43567
rect -7841 -43673 -7807 -43639
rect -7523 -43313 -7489 -43279
rect -7523 -43385 -7489 -43351
rect -7523 -43457 -7489 -43423
rect -7523 -43529 -7489 -43495
rect -7523 -43601 -7489 -43567
rect -7523 -43673 -7489 -43639
rect -7205 -43313 -7171 -43279
rect -7205 -43385 -7171 -43351
rect -7205 -43457 -7171 -43423
rect -7205 -43529 -7171 -43495
rect -7205 -43601 -7171 -43567
rect -7205 -43673 -7171 -43639
rect -6887 -43313 -6853 -43279
rect -6887 -43385 -6853 -43351
rect -6887 -43457 -6853 -43423
rect -6887 -43529 -6853 -43495
rect -6887 -43601 -6853 -43567
rect -6887 -43673 -6853 -43639
rect -5304 -43863 -5270 -43829
rect -2296 -42745 -2262 -42711
rect -2296 -42817 -2262 -42783
rect -2296 -42889 -2262 -42855
rect -2296 -42961 -2262 -42927
rect -2296 -43033 -2262 -42999
rect -2296 -43105 -2262 -43071
rect -1978 -42745 -1944 -42711
rect -1978 -42817 -1944 -42783
rect -1978 -42889 -1944 -42855
rect -1978 -42961 -1944 -42927
rect -1978 -43033 -1944 -42999
rect -1978 -43105 -1944 -43071
rect -1660 -42745 -1626 -42711
rect -1660 -42817 -1626 -42783
rect -1660 -42889 -1626 -42855
rect -1660 -42961 -1626 -42927
rect -1660 -43033 -1626 -42999
rect -1660 -43105 -1626 -43071
rect -1342 -42745 -1308 -42711
rect -1342 -42817 -1308 -42783
rect -1342 -42889 -1308 -42855
rect -1342 -42961 -1308 -42927
rect -1342 -43033 -1308 -42999
rect -1342 -43105 -1308 -43071
rect -2526 -43195 -2492 -43161
rect -3150 -43267 -3116 -43233
rect -3030 -43267 -2996 -43233
rect -3150 -43387 -3116 -43353
rect -3030 -43387 -2996 -43353
rect -3096 -43689 -3056 -43649
rect -2296 -43314 -2262 -43280
rect -2296 -43386 -2262 -43352
rect -2296 -43458 -2262 -43424
rect -2296 -43530 -2262 -43496
rect -2296 -43602 -2262 -43568
rect -2296 -43674 -2262 -43640
rect -1978 -43314 -1944 -43280
rect -1978 -43386 -1944 -43352
rect -1978 -43458 -1944 -43424
rect -1978 -43530 -1944 -43496
rect -1978 -43602 -1944 -43568
rect -1978 -43674 -1944 -43640
rect -1660 -43314 -1626 -43280
rect -1660 -43386 -1626 -43352
rect -1660 -43458 -1626 -43424
rect -1660 -43530 -1626 -43496
rect -1660 -43602 -1626 -43568
rect -1660 -43674 -1626 -43640
rect -1342 -43314 -1308 -43280
rect -1342 -43386 -1308 -43352
rect -1342 -43458 -1308 -43424
rect -1342 -43530 -1308 -43496
rect -1342 -43602 -1308 -43568
rect -1342 -43674 -1308 -43640
rect -10378 -45001 -10344 -44998
rect -10258 -45001 -10224 -44998
rect -10378 -45004 -10343 -45001
rect -10258 -45004 -10223 -45001
rect -10379 -45035 -10343 -45004
rect -10259 -45035 -10223 -45004
rect -10379 -45038 -10345 -45035
rect -10259 -45038 -10225 -45035
rect -10378 -45121 -10344 -45118
rect -10258 -45121 -10224 -45118
rect -10378 -45124 -10343 -45121
rect -10258 -45124 -10223 -45121
rect -10379 -45155 -10343 -45124
rect -10259 -45155 -10223 -45124
rect -10379 -45158 -10345 -45155
rect -10259 -45158 -10225 -45155
rect -7910 -45093 -7876 -45059
rect -6807 -45093 -6773 -45090
rect -6687 -45093 -6653 -45090
rect -6807 -45096 -6772 -45093
rect -6687 -45096 -6652 -45093
rect -6808 -45127 -6772 -45096
rect -6688 -45127 -6652 -45096
rect -6808 -45130 -6773 -45127
rect -6688 -45130 -6653 -45127
rect -6807 -45131 -6773 -45130
rect -6687 -45131 -6653 -45130
rect -6807 -45213 -6773 -45210
rect -6687 -45213 -6653 -45210
rect -6807 -45216 -6772 -45213
rect -6687 -45216 -6652 -45213
rect -6808 -45247 -6772 -45216
rect -6688 -45247 -6652 -45216
rect -6808 -45250 -6773 -45247
rect -6688 -45250 -6653 -45247
rect -6807 -45251 -6773 -45250
rect -6687 -45251 -6653 -45250
rect -5179 -45130 -5145 -45096
rect -5059 -45130 -5025 -45096
rect -5179 -45250 -5145 -45216
rect -5059 -45250 -5025 -45216
rect -11699 -45470 -11665 -45436
rect -11619 -45470 -11585 -45436
rect -11539 -45470 -11505 -45436
rect -11459 -45470 -11425 -45436
rect -11379 -45470 -11345 -45436
rect -11299 -45470 -11265 -45436
rect -11219 -45470 -11185 -45436
rect -11139 -45470 -11105 -45436
rect -11059 -45470 -11025 -45436
rect -10979 -45470 -10945 -45436
rect -10899 -45470 -10865 -45436
rect -10819 -45470 -10785 -45436
rect -10739 -45470 -10705 -45436
rect -10659 -45470 -10625 -45436
rect -10579 -45470 -10545 -45436
rect -10499 -45470 -10465 -45436
rect -10419 -45470 -10385 -45436
rect -10339 -45470 -10305 -45436
rect -10259 -45470 -10225 -45436
rect -10179 -45470 -10145 -45436
rect -10099 -45470 -10065 -45436
rect -10019 -45470 -9985 -45436
rect -9939 -45470 -9905 -45436
rect -9859 -45470 -9825 -45436
rect -9779 -45470 -9745 -45436
rect -9699 -45470 -9665 -45436
rect -9619 -45470 -9585 -45436
rect -9539 -45470 -9505 -45436
rect -9459 -45470 -9425 -45436
rect -9379 -45470 -9345 -45436
rect -9299 -45470 -9265 -45436
rect -9219 -45470 -9185 -45436
rect -9139 -45470 -9105 -45436
rect -9059 -45470 -9025 -45436
rect -8979 -45470 -8945 -45436
rect -8899 -45470 -8865 -45436
rect -8819 -45470 -8785 -45436
rect -8739 -45470 -8705 -45436
rect -8659 -45470 -8625 -45436
rect -8579 -45470 -8545 -45436
rect -8499 -45470 -8465 -45436
rect -8419 -45470 -8385 -45436
rect -8339 -45470 -8305 -45436
rect -8259 -45470 -8225 -45436
rect -8179 -45470 -8145 -45436
rect -8099 -45470 -8065 -45436
rect -8019 -45470 -7985 -45436
rect -7939 -45470 -7905 -45436
rect -7859 -45470 -7825 -45436
rect -7779 -45470 -7745 -45436
rect -7699 -45470 -7665 -45436
rect -7619 -45470 -7585 -45436
rect -7539 -45470 -7505 -45436
rect -7459 -45470 -7425 -45436
rect -7379 -45470 -7345 -45436
rect -7299 -45470 -7265 -45436
rect -7219 -45470 -7185 -45436
rect -7139 -45470 -7105 -45436
rect -7059 -45470 -7025 -45436
rect -6979 -45470 -6945 -45436
rect -6899 -45470 -6865 -45436
rect -6819 -45470 -6785 -45436
rect -6739 -45470 -6705 -45436
rect -6659 -45470 -6625 -45436
rect -6579 -45470 -6545 -45436
rect -6499 -45470 -6465 -45436
rect -6419 -45470 -6385 -45436
rect -6339 -45470 -6305 -45436
rect -6259 -45470 -6225 -45436
rect -6179 -45470 -6145 -45436
rect -6099 -45470 -6065 -45436
rect -6019 -45470 -5985 -45436
rect -5939 -45470 -5905 -45436
rect -5859 -45470 -5825 -45436
rect -5779 -45470 -5745 -45436
rect -5699 -45470 -5665 -45436
rect -5619 -45470 -5585 -45436
rect -5539 -45470 -5505 -45436
rect -5459 -45470 -5425 -45436
rect -5379 -45470 -5345 -45436
rect -5299 -45470 -5265 -45436
rect -5219 -45470 -5185 -45436
rect -5139 -45470 -5105 -45436
rect -5059 -45470 -5025 -45436
rect -4979 -45470 -4945 -45436
rect -4899 -45470 -4865 -45436
rect -4819 -45470 -4785 -45436
rect -4739 -45470 -4705 -45436
rect -4659 -45470 -4625 -45436
rect -4579 -45470 -4545 -45436
rect -4499 -45470 -4465 -45436
rect -4419 -45470 -4385 -45436
rect -4339 -45470 -4305 -45436
rect -4259 -45470 -4225 -45436
rect -4179 -45470 -4145 -45436
rect -4099 -45470 -4065 -45436
rect -4019 -45470 -3985 -45436
rect -3939 -45470 -3905 -45436
rect -3859 -45470 -3825 -45436
rect -3779 -45470 -3745 -45436
rect -3699 -45470 -3665 -45436
rect -3619 -45470 -3585 -45436
rect -3539 -45470 -3505 -45436
rect -3459 -45470 -3425 -45436
rect -3379 -45470 -3345 -45436
rect -3299 -45470 -3265 -45436
rect -3219 -45470 -3185 -45436
rect -3139 -45470 -3105 -45436
rect -3059 -45470 -3025 -45436
rect -2979 -45470 -2945 -45436
rect -2899 -45470 -2865 -45436
rect -2819 -45470 -2785 -45436
rect -2739 -45470 -2705 -45436
rect -2659 -45470 -2625 -45436
rect -2579 -45470 -2545 -45436
rect -2499 -45470 -2465 -45436
rect -2419 -45470 -2385 -45436
rect -2339 -45470 -2305 -45436
rect -2259 -45470 -2225 -45436
rect -2179 -45470 -2145 -45436
rect -6802 -45992 -6768 -45958
rect -6682 -45992 -6648 -45958
rect -6802 -46112 -6768 -46078
rect -6682 -46112 -6648 -46078
rect -5176 -45992 -5142 -45958
rect -5056 -45992 -5022 -45958
rect -5176 -46112 -5142 -46078
rect -5056 -46112 -5022 -46078
rect -44435 -47009 -44401 -46975
rect -44355 -47009 -44321 -46975
rect -44275 -47009 -44241 -46975
rect -44195 -47009 -44161 -46975
rect -44115 -47009 -44081 -46975
rect -44035 -47009 -44001 -46975
rect -43955 -47009 -43921 -46975
rect -43875 -47009 -43841 -46975
rect -43795 -47009 -43761 -46975
rect -43715 -47009 -43681 -46975
rect -43635 -47009 -43601 -46975
rect -43555 -47009 -43521 -46975
rect -43475 -47009 -43441 -46975
rect -43395 -47009 -43361 -46975
rect -43315 -47009 -43281 -46975
rect -43235 -47009 -43201 -46975
rect -43155 -47009 -43121 -46975
rect -43075 -47009 -43041 -46975
rect -42995 -47009 -42961 -46975
rect -42915 -47009 -42881 -46975
rect -42835 -47009 -42801 -46975
rect -42755 -47009 -42721 -46975
rect -42675 -47009 -42641 -46975
rect -42595 -47009 -42561 -46975
rect -42515 -47009 -42481 -46975
rect -42435 -47009 -42401 -46975
rect -42355 -47009 -42321 -46975
rect -42275 -47009 -42241 -46975
rect -42195 -47009 -42161 -46975
rect -42115 -47009 -42081 -46975
rect -42035 -47009 -42001 -46975
rect -41955 -47009 -41921 -46975
rect -41875 -47009 -41841 -46975
rect -41795 -47009 -41761 -46975
rect -41715 -47009 -41681 -46975
rect -41635 -47009 -41601 -46975
rect -41555 -47009 -41521 -46975
rect -41475 -47009 -41441 -46975
rect -41395 -47009 -41361 -46975
rect -41315 -47009 -41281 -46975
rect -41235 -47009 -41201 -46975
rect -41155 -47009 -41121 -46975
rect -41075 -47009 -41041 -46975
rect -40995 -47009 -40961 -46975
rect -40915 -47009 -40881 -46975
rect -40835 -47009 -40801 -46975
rect -40755 -47009 -40721 -46975
rect -40675 -47009 -40641 -46975
rect -40595 -47009 -40561 -46975
rect -40515 -47009 -40481 -46975
rect -40435 -47009 -40401 -46975
rect -40355 -47009 -40321 -46975
rect -40275 -47009 -40241 -46975
rect -40195 -47009 -40161 -46975
rect -40115 -47009 -40081 -46975
rect -40035 -47009 -40001 -46975
rect -39955 -47009 -39921 -46975
rect -39875 -47009 -39841 -46975
rect -39795 -47009 -39761 -46975
rect -39715 -47009 -39681 -46975
rect -39635 -47009 -39601 -46975
rect -39555 -47009 -39521 -46975
rect -39475 -47009 -39441 -46975
rect -39395 -47009 -39361 -46975
rect -39315 -47009 -39281 -46975
rect -39235 -47009 -39201 -46975
rect -39155 -47009 -39121 -46975
rect -39075 -47009 -39041 -46975
rect -38995 -47009 -38961 -46975
rect -38915 -47009 -38881 -46975
rect -38835 -47009 -38801 -46975
rect -38755 -47009 -38721 -46975
rect -38675 -47009 -38641 -46975
rect -38595 -47009 -38561 -46975
rect -38515 -47009 -38481 -46975
rect -38435 -47009 -38401 -46975
rect -38355 -47009 -38321 -46975
rect -38275 -47009 -38241 -46975
rect -38195 -47009 -38161 -46975
rect -38115 -47009 -38081 -46975
rect -38035 -47009 -38001 -46975
rect -37955 -47009 -37921 -46975
rect -37875 -47009 -37841 -46975
rect -37795 -47009 -37761 -46975
rect -37715 -47009 -37681 -46975
rect -37635 -47009 -37601 -46975
rect -37555 -47009 -37521 -46975
rect -37475 -47009 -37441 -46975
rect -37395 -47009 -37361 -46975
rect -37315 -47009 -37281 -46975
rect -37235 -47009 -37201 -46975
rect -37155 -47009 -37121 -46975
rect -37075 -47009 -37041 -46975
rect -36995 -47009 -36961 -46975
rect -36915 -47009 -36881 -46975
rect -36835 -47009 -36801 -46975
rect -36755 -47009 -36721 -46975
rect -36675 -47009 -36641 -46975
rect -36595 -47009 -36561 -46975
rect -36515 -47009 -36481 -46975
rect -36435 -47009 -36401 -46975
rect -36355 -47009 -36321 -46975
rect -36275 -47009 -36241 -46975
rect -36195 -47009 -36161 -46975
rect -36115 -47009 -36081 -46975
rect -36035 -47009 -36001 -46975
rect -35955 -47009 -35921 -46975
rect -35875 -47009 -35841 -46975
rect -35795 -47009 -35761 -46975
rect -35715 -47009 -35681 -46975
rect -35635 -47009 -35601 -46975
rect -35555 -47009 -35521 -46975
rect -35475 -47009 -35441 -46975
rect -35395 -47009 -35361 -46975
rect -35315 -47009 -35281 -46975
rect -35235 -47009 -35201 -46975
rect -35155 -47009 -35121 -46975
rect -35075 -47009 -35041 -46975
rect -34995 -47009 -34961 -46975
rect -34915 -47009 -34881 -46975
rect -34835 -47009 -34801 -46975
rect -34755 -47009 -34721 -46975
rect -34675 -47009 -34641 -46975
rect -34595 -47009 -34561 -46975
rect -34515 -47009 -34481 -46975
rect -34435 -47009 -34401 -46975
rect -34355 -47009 -34321 -46975
rect -34275 -47009 -34241 -46975
rect -34195 -47009 -34161 -46975
rect -34115 -47009 -34081 -46975
rect -34035 -47009 -34001 -46975
rect -33955 -47009 -33921 -46975
rect -33875 -47009 -33841 -46975
rect -33795 -47009 -33761 -46975
rect -33715 -47009 -33681 -46975
rect -33635 -47009 -33601 -46975
rect -33555 -47009 -33521 -46975
rect -33475 -47009 -33441 -46975
rect -33395 -47009 -33361 -46975
rect -33315 -47009 -33281 -46975
rect -33235 -47009 -33201 -46975
rect -33155 -47009 -33121 -46975
rect -33075 -47009 -33041 -46975
rect -32995 -47009 -32961 -46975
rect -32915 -47009 -32881 -46975
rect -32835 -47009 -32801 -46975
rect -32755 -47009 -32721 -46975
rect -32675 -47009 -32641 -46975
rect -32595 -47009 -32561 -46975
rect -32515 -47009 -32481 -46975
rect -32435 -47009 -32401 -46975
rect -32355 -47009 -32321 -46975
rect -32275 -47009 -32241 -46975
rect -32195 -47009 -32161 -46975
rect -32115 -47009 -32081 -46975
rect -32035 -47009 -32001 -46975
rect -31955 -47009 -31921 -46975
rect -31875 -47009 -31841 -46975
rect -31795 -47009 -31761 -46975
rect -31715 -47009 -31681 -46975
rect -31635 -47009 -31601 -46975
rect -31555 -47009 -31521 -46975
rect -31475 -47009 -31441 -46975
rect -31395 -47009 -31361 -46975
rect -31315 -47009 -31281 -46975
rect -31235 -47009 -31201 -46975
rect -31155 -47009 -31121 -46975
rect -31075 -47009 -31041 -46975
rect -30995 -47009 -30961 -46975
rect -30915 -47009 -30881 -46975
rect -30835 -47009 -30801 -46975
rect -30755 -47009 -30721 -46975
rect -30675 -47009 -30641 -46975
rect -30595 -47009 -30561 -46975
rect -30515 -47009 -30481 -46975
rect -30435 -47009 -30401 -46975
rect -30355 -47009 -30321 -46975
rect -30275 -47009 -30241 -46975
rect -30195 -47009 -30161 -46975
rect -30115 -47009 -30081 -46975
rect -30035 -47009 -30001 -46975
rect -29955 -47009 -29921 -46975
rect -29875 -47009 -29841 -46975
rect -29795 -47009 -29761 -46975
rect -29715 -47009 -29681 -46975
rect -29635 -47009 -29601 -46975
rect -29555 -47009 -29521 -46975
rect -29475 -47009 -29441 -46975
rect -29395 -47009 -29361 -46975
rect -29315 -47009 -29281 -46975
rect -29235 -47009 -29201 -46975
rect -29155 -47009 -29121 -46975
rect -29075 -47009 -29041 -46975
rect -28995 -47009 -28961 -46975
rect -28915 -47009 -28881 -46975
rect -28835 -47009 -28801 -46975
rect -28755 -47009 -28721 -46975
rect -28675 -47009 -28641 -46975
rect -28595 -47009 -28561 -46975
rect -28514 -47009 -28480 -46975
rect -28434 -47009 -28400 -46975
rect -28354 -47009 -28320 -46975
rect -28274 -47009 -28240 -46975
rect -28194 -47009 -28160 -46975
rect -28114 -47009 -28080 -46975
rect -28034 -47009 -28000 -46975
rect -27954 -47009 -27920 -46975
rect -27874 -47009 -27840 -46975
rect -27794 -47009 -27760 -46975
rect -27714 -47009 -27680 -46975
rect -27634 -47009 -27600 -46975
rect -27554 -47009 -27520 -46975
rect -27474 -47009 -27440 -46975
rect -27394 -47009 -27360 -46975
rect -27314 -47009 -27280 -46975
rect -27234 -47009 -27200 -46975
rect -27154 -47009 -27120 -46975
rect -27074 -47009 -27040 -46975
rect -26994 -47009 -26960 -46975
rect -26914 -47009 -26880 -46975
rect -26834 -47009 -26800 -46975
rect -26754 -47009 -26720 -46975
rect -26674 -47009 -26640 -46975
rect -26594 -47009 -26560 -46975
rect -26514 -47009 -26480 -46975
rect -26434 -47009 -26400 -46975
rect -26354 -47009 -26320 -46975
rect -26274 -47009 -26240 -46975
rect -26194 -47009 -26160 -46975
rect -26114 -47009 -26080 -46975
rect -26034 -47009 -26000 -46975
rect -25954 -47009 -25920 -46975
rect -25874 -47009 -25840 -46975
rect -25794 -47009 -25760 -46975
rect -25714 -47009 -25680 -46975
rect -25634 -47009 -25600 -46975
rect -25554 -47009 -25520 -46975
rect -25474 -47009 -25440 -46975
rect -25394 -47009 -25360 -46975
rect -25314 -47009 -25280 -46975
rect -25234 -47009 -25200 -46975
rect -25154 -47009 -25120 -46975
rect -25074 -47009 -25040 -46975
rect -24994 -47009 -24960 -46975
rect -24914 -47009 -24880 -46975
rect -24834 -47009 -24800 -46975
rect -24754 -47009 -24720 -46975
rect -24674 -47009 -24640 -46975
rect -24594 -47009 -24560 -46975
rect -24514 -47009 -24480 -46975
rect -24434 -47009 -24400 -46975
rect -24354 -47009 -24320 -46975
rect -24274 -47009 -24240 -46975
rect -24194 -47009 -24160 -46975
rect -24114 -47009 -24080 -46975
rect -24034 -47009 -24000 -46975
rect -23954 -47009 -23920 -46975
rect -23874 -47009 -23840 -46975
rect -23794 -47009 -23760 -46975
rect -23714 -47009 -23680 -46975
rect -23634 -47009 -23600 -46975
rect -23554 -47009 -23520 -46975
rect -23474 -47009 -23440 -46975
rect -23394 -47009 -23360 -46975
rect -23314 -47009 -23280 -46975
rect -23234 -47009 -23200 -46975
rect -23154 -47009 -23120 -46975
rect -23074 -47009 -23040 -46975
rect -22994 -47009 -22960 -46975
rect -22914 -47009 -22880 -46975
rect -22834 -47009 -22800 -46975
rect -22754 -47009 -22720 -46975
rect -22674 -47009 -22640 -46975
rect -22594 -47009 -22560 -46975
rect -22514 -47009 -22480 -46975
rect -22434 -47009 -22400 -46975
rect -22354 -47009 -22320 -46975
rect -22274 -47009 -22240 -46975
rect -22194 -47009 -22160 -46975
rect -22114 -47009 -22080 -46975
rect -22034 -47009 -22000 -46975
rect -21954 -47009 -21920 -46975
rect -21874 -47009 -21840 -46975
rect -21794 -47009 -21760 -46975
rect -21714 -47009 -21680 -46975
rect -21634 -47009 -21600 -46975
rect -21554 -47009 -21520 -46975
rect -21474 -47009 -21440 -46975
rect -21394 -47009 -21360 -46975
rect -21314 -47009 -21280 -46975
rect -21234 -47009 -21200 -46975
rect -21154 -47009 -21120 -46975
rect -21074 -47009 -21040 -46975
rect -20994 -47009 -20960 -46975
rect -20914 -47009 -20880 -46975
rect -20834 -47009 -20800 -46975
rect -20754 -47009 -20720 -46975
rect -20674 -47009 -20640 -46975
rect -20594 -47009 -20560 -46975
rect -20514 -47009 -20480 -46975
rect -20434 -47009 -20400 -46975
rect -20354 -47009 -20320 -46975
rect -20274 -47009 -20240 -46975
rect -20194 -47009 -20160 -46975
rect -20114 -47009 -20080 -46975
rect -20034 -47009 -20000 -46975
rect -19954 -47009 -19920 -46975
rect -19874 -47009 -19840 -46975
rect -19794 -47009 -19760 -46975
rect -19714 -47009 -19680 -46975
rect -19634 -47009 -19600 -46975
rect -19554 -47009 -19520 -46975
rect -19474 -47009 -19440 -46975
rect -19394 -47009 -19360 -46975
rect -19314 -47009 -19280 -46975
rect -19234 -47009 -19200 -46975
rect -19154 -47009 -19120 -46975
rect -19074 -47009 -19040 -46975
rect -18994 -47009 -18960 -46975
rect -18914 -47009 -18880 -46975
rect -18834 -47009 -18800 -46975
rect -18754 -47009 -18720 -46975
rect -18674 -47009 -18640 -46975
rect -18594 -47009 -18560 -46975
rect -18514 -47009 -18480 -46975
rect -18434 -47009 -18400 -46975
rect -18354 -47009 -18320 -46975
rect -18274 -47009 -18240 -46975
rect -18194 -47009 -18160 -46975
rect -18114 -47009 -18080 -46975
rect -18034 -47009 -18000 -46975
rect -17954 -47009 -17920 -46975
rect -17874 -47009 -17840 -46975
rect -17794 -47009 -17760 -46975
rect -17714 -47009 -17680 -46975
rect -17634 -47009 -17600 -46975
rect -17554 -47009 -17520 -46975
rect -17474 -47009 -17440 -46975
rect -17394 -47009 -17360 -46975
rect -17314 -47009 -17280 -46975
rect -17234 -47009 -17200 -46975
rect -17154 -47009 -17120 -46975
rect -17074 -47009 -17040 -46975
rect -16994 -47009 -16960 -46975
rect -16914 -47009 -16880 -46975
rect -16834 -47009 -16800 -46975
rect -16754 -47009 -16720 -46975
rect -16674 -47009 -16640 -46975
rect -16594 -47009 -16560 -46975
rect -16514 -47009 -16480 -46975
rect -16434 -47009 -16400 -46975
rect -16354 -47009 -16320 -46975
rect -16274 -47009 -16240 -46975
rect -16194 -47009 -16160 -46975
rect -16114 -47009 -16080 -46975
rect -16034 -47009 -16000 -46975
rect -15954 -47009 -15920 -46975
rect -15874 -47009 -15840 -46975
rect -15794 -47009 -15760 -46975
rect -15714 -47009 -15680 -46975
rect -15634 -47009 -15600 -46975
rect -15553 -47009 -15519 -46975
rect -15473 -47009 -15439 -46975
rect -15393 -47009 -15359 -46975
rect -15313 -47009 -15279 -46975
rect -15233 -47009 -15199 -46975
rect -15153 -47009 -15119 -46975
rect -15073 -47009 -15039 -46975
rect -14993 -47009 -14959 -46975
rect -14913 -47009 -14879 -46975
rect -14833 -47009 -14799 -46975
rect -14753 -47009 -14719 -46975
rect -14673 -47009 -14639 -46975
rect -14593 -47009 -14559 -46975
rect -14513 -47009 -14479 -46975
rect -14433 -47009 -14399 -46975
rect -14353 -47009 -14319 -46975
rect -14273 -47009 -14239 -46975
rect -14193 -47009 -14159 -46975
rect -14113 -47009 -14079 -46975
rect -14033 -47009 -13999 -46975
rect -13953 -47009 -13919 -46975
rect -13873 -47009 -13839 -46975
rect -13793 -47009 -13759 -46975
rect -13713 -47009 -13679 -46975
rect -13633 -47009 -13599 -46975
rect -13553 -47009 -13519 -46975
rect -13473 -47009 -13439 -46975
rect -13393 -47009 -13359 -46975
rect -13313 -47009 -13279 -46975
rect -13233 -47009 -13199 -46975
rect -13153 -47009 -13119 -46975
rect -13073 -47009 -13039 -46975
rect -12993 -47009 -12959 -46975
rect -12913 -47009 -12879 -46975
rect -12833 -47009 -12799 -46975
rect -12753 -47009 -12719 -46975
rect -12673 -47009 -12639 -46975
rect -12593 -47009 -12559 -46975
rect -12513 -47009 -12479 -46975
rect -12433 -47009 -12399 -46975
rect -12353 -47009 -12319 -46975
rect -12273 -47009 -12239 -46975
rect -12193 -47009 -12159 -46975
rect -12113 -47009 -12079 -46975
rect -12033 -47009 -11999 -46975
rect -11953 -47009 -11919 -46975
rect -11873 -47009 -11839 -46975
rect -11793 -47009 -11759 -46975
rect -11713 -47009 -11679 -46975
rect -11633 -47009 -11599 -46975
rect -11553 -47009 -11519 -46975
rect -11473 -47009 -11439 -46975
rect -11393 -47009 -11359 -46975
rect -11313 -47009 -11279 -46975
rect -11233 -47009 -11199 -46975
rect -11153 -47009 -11119 -46975
rect -11073 -47009 -11039 -46975
rect -10993 -47009 -10959 -46975
rect -10913 -47009 -10879 -46975
rect -10833 -47009 -10799 -46975
rect -10753 -47009 -10719 -46975
rect -10673 -47009 -10639 -46975
rect -10593 -47009 -10559 -46975
rect -10513 -47009 -10479 -46975
rect -10433 -47009 -10399 -46975
rect -10353 -47009 -10319 -46975
rect -10273 -47009 -10239 -46975
rect -10193 -47009 -10159 -46975
rect -10113 -47009 -10079 -46975
rect -10033 -47009 -9999 -46975
rect -9953 -47009 -9919 -46975
rect -9873 -47009 -9839 -46975
rect -9793 -47009 -9759 -46975
rect -9713 -47009 -9679 -46975
rect -9633 -47009 -9599 -46975
rect -9553 -47009 -9519 -46975
rect -9473 -47009 -9439 -46975
rect -9393 -47009 -9359 -46975
rect -9313 -47009 -9279 -46975
rect -9233 -47009 -9199 -46975
rect -9153 -47009 -9119 -46975
rect -9073 -47009 -9039 -46975
rect -8993 -47009 -8959 -46975
rect -8913 -47009 -8879 -46975
rect -8833 -47009 -8799 -46975
rect -8753 -47009 -8719 -46975
rect -8673 -47009 -8639 -46975
rect -8593 -47009 -8559 -46975
rect -8513 -47009 -8479 -46975
rect -8433 -47009 -8399 -46975
rect -8353 -47009 -8319 -46975
rect -8273 -47009 -8239 -46975
rect -8193 -47009 -8159 -46975
rect -8113 -47009 -8079 -46975
rect -8033 -47009 -7999 -46975
rect -7953 -47009 -7919 -46975
rect -7873 -47009 -7839 -46975
rect -7793 -47009 -7759 -46975
rect -7713 -47009 -7679 -46975
rect -7633 -47009 -7599 -46975
rect -7553 -47009 -7519 -46975
rect -7473 -47009 -7439 -46975
rect -7393 -47009 -7359 -46975
rect -7313 -47009 -7279 -46975
rect -7233 -47009 -7199 -46975
rect -7153 -47009 -7119 -46975
rect -7073 -47009 -7039 -46975
rect -6993 -47009 -6959 -46975
rect -6913 -47009 -6879 -46975
rect -6841 -47009 -6807 -46975
rect -6769 -47009 -6735 -46975
rect -6697 -47009 -6663 -46975
rect -6625 -47009 -6591 -46975
rect -6553 -47009 -6519 -46975
rect -6481 -47009 -6447 -46975
rect -6409 -47009 -6375 -46975
rect -6337 -47009 -6303 -46975
rect -6265 -47009 -6231 -46975
rect -6193 -47009 -6159 -46975
rect -6121 -47009 -6087 -46975
rect -6049 -47009 -6015 -46975
rect -5977 -47009 -5943 -46975
rect -5905 -47009 -5871 -46975
rect -5833 -47009 -5799 -46975
rect -5761 -47009 -5727 -46975
rect -5689 -47009 -5655 -46975
rect -5617 -47009 -5583 -46975
rect -5545 -47009 -5511 -46975
rect -5473 -47009 -5439 -46975
rect -5401 -47009 -5367 -46975
rect -5329 -47009 -5295 -46975
rect -5257 -47009 -5223 -46975
rect -5185 -47009 -5151 -46975
rect -5113 -47009 -5079 -46975
rect -5041 -47009 -5007 -46975
rect -4969 -47009 -4935 -46975
rect -4889 -47009 -4855 -46975
rect -4809 -47009 -4775 -46975
rect -4729 -47009 -4695 -46975
rect -4649 -47009 -4615 -46975
rect -4569 -47009 -4535 -46975
rect -4489 -47009 -4455 -46975
rect -4409 -47009 -4375 -46975
rect -4329 -47009 -4295 -46975
rect -4249 -47009 -4215 -46975
rect -4933 -47153 -4899 -47119
rect -6778 -47832 -6744 -47801
rect -6778 -47835 -6744 -47832
rect -6778 -48216 -6744 -48213
rect -6778 -48247 -6744 -48216
rect -10087 -48379 -10053 -48345
rect -10007 -48379 -9973 -48345
rect -9927 -48379 -9893 -48345
rect -9847 -48379 -9813 -48345
rect -9767 -48379 -9733 -48345
rect -9687 -48379 -9653 -48345
rect -9607 -48379 -9573 -48345
rect -9527 -48379 -9493 -48345
rect -9447 -48379 -9413 -48345
rect -9367 -48379 -9333 -48345
rect -9287 -48379 -9253 -48345
rect -9207 -48379 -9173 -48345
rect -9127 -48379 -9093 -48345
rect -9047 -48379 -9013 -48345
rect -8967 -48379 -8933 -48345
rect -8887 -48379 -8853 -48345
rect -8807 -48379 -8773 -48345
rect -8727 -48379 -8693 -48345
rect -8647 -48379 -8613 -48345
rect -8567 -48379 -8533 -48345
rect -8487 -48379 -8453 -48345
rect -8407 -48379 -8373 -48345
rect -8327 -48379 -8293 -48345
rect -8247 -48379 -8213 -48345
rect -8167 -48379 -8133 -48345
rect -8087 -48379 -8053 -48345
rect -8007 -48379 -7973 -48345
rect -7927 -48379 -7893 -48345
rect -7847 -48379 -7813 -48345
rect -7767 -48379 -7733 -48345
rect -7687 -48379 -7653 -48345
rect -7607 -48379 -7573 -48345
rect -7527 -48379 -7493 -48345
rect -7447 -48379 -7413 -48345
rect -7367 -48379 -7333 -48345
rect -7287 -48379 -7253 -48345
rect -7207 -48379 -7173 -48345
rect -7127 -48379 -7093 -48345
rect -7047 -48379 -7013 -48345
rect -6967 -48379 -6933 -48345
rect -6887 -48379 -6853 -48345
rect -6807 -48379 -6773 -48345
rect -6727 -48379 -6693 -48345
rect -6647 -48379 -6613 -48345
rect -6567 -48379 -6533 -48345
rect -6487 -48379 -6453 -48345
rect -6407 -48379 -6373 -48345
rect -6327 -48379 -6293 -48345
rect -6247 -48379 -6213 -48345
rect -6167 -48379 -6133 -48345
rect -6087 -48379 -6053 -48345
rect -6007 -48379 -5973 -48345
rect -5927 -48379 -5893 -48345
rect -5847 -48379 -5813 -48345
rect -5767 -48379 -5733 -48345
rect -5687 -48379 -5653 -48345
rect -5607 -48379 -5573 -48345
rect -5527 -48379 -5493 -48345
rect -5447 -48379 -5413 -48345
rect -5367 -48379 -5333 -48345
rect -5287 -48379 -5253 -48345
rect -5207 -48379 -5173 -48345
rect -5127 -48379 -5093 -48345
rect -5047 -48379 -5013 -48345
rect -4967 -48379 -4933 -48345
rect -4887 -48379 -4853 -48345
rect -4807 -48379 -4773 -48345
rect -4727 -48379 -4693 -48345
rect -4647 -48379 -4613 -48345
rect -4567 -48379 -4533 -48345
rect -4487 -48379 -4453 -48345
rect -4407 -48379 -4373 -48345
rect -4327 -48379 -4293 -48345
rect -4247 -48379 -4213 -48345
rect -4167 -48379 -4133 -48345
rect -4087 -48379 -4053 -48345
rect -4007 -48379 -3973 -48345
rect -3927 -48379 -3893 -48345
rect -3847 -48379 -3813 -48345
rect -3767 -48379 -3733 -48345
rect -3687 -48379 -3653 -48345
rect -3607 -48379 -3573 -48345
rect -3527 -48379 -3493 -48345
rect -3447 -48379 -3413 -48345
rect -3367 -48379 -3333 -48345
rect -3287 -48379 -3253 -48345
rect -3207 -48379 -3173 -48345
rect -3127 -48379 -3093 -48345
rect -3047 -48379 -3013 -48345
rect -2967 -48379 -2933 -48345
rect -2887 -48379 -2853 -48345
rect -2807 -48379 -2773 -48345
rect -2727 -48379 -2693 -48345
rect -2647 -48379 -2613 -48345
rect -2567 -48379 -2533 -48345
rect -2487 -48379 -2453 -48345
rect -2407 -48379 -2373 -48345
rect -2327 -48379 -2293 -48345
rect -2247 -48379 -2213 -48345
rect -2167 -48379 -2133 -48345
<< metal1 >>
rect -44482 -34599 31781 -34566
rect -44482 -34633 -44422 -34599
rect -44388 -34633 -44342 -34599
rect -44308 -34633 -44262 -34599
rect -44228 -34633 -44182 -34599
rect -44148 -34633 -44102 -34599
rect -44068 -34633 -44022 -34599
rect -43988 -34633 -43942 -34599
rect -43908 -34633 -43862 -34599
rect -43828 -34633 -43782 -34599
rect -43748 -34633 -43702 -34599
rect -43668 -34633 -43622 -34599
rect -43588 -34633 -43542 -34599
rect -43508 -34633 -43462 -34599
rect -43428 -34633 -43382 -34599
rect -43348 -34633 -43302 -34599
rect -43268 -34633 -43222 -34599
rect -43188 -34633 -43142 -34599
rect -43108 -34633 -43062 -34599
rect -43028 -34633 -42982 -34599
rect -42948 -34633 -42902 -34599
rect -42868 -34633 -42822 -34599
rect -42788 -34633 -42742 -34599
rect -42708 -34633 -42662 -34599
rect -42628 -34633 -42582 -34599
rect -42548 -34633 -42502 -34599
rect -42468 -34633 -42422 -34599
rect -42388 -34633 -42342 -34599
rect -42308 -34633 -42262 -34599
rect -42228 -34633 -42182 -34599
rect -42148 -34633 -42102 -34599
rect -42068 -34633 -42022 -34599
rect -41988 -34633 -41942 -34599
rect -41908 -34633 -41862 -34599
rect -41828 -34633 -41782 -34599
rect -41748 -34633 -41702 -34599
rect -41668 -34633 -41622 -34599
rect -41588 -34633 -41542 -34599
rect -41508 -34633 -41462 -34599
rect -41428 -34633 -41382 -34599
rect -41348 -34633 -41302 -34599
rect -41268 -34633 -41222 -34599
rect -41188 -34633 -41142 -34599
rect -41108 -34633 -41062 -34599
rect -41028 -34633 -40982 -34599
rect -40948 -34633 -40902 -34599
rect -40868 -34633 -40822 -34599
rect -40788 -34633 -40742 -34599
rect -40708 -34633 -40662 -34599
rect -40628 -34633 -40582 -34599
rect -40548 -34633 -40502 -34599
rect -40468 -34633 -40422 -34599
rect -40388 -34633 -40342 -34599
rect -40308 -34633 -40262 -34599
rect -40228 -34633 -40182 -34599
rect -40148 -34633 -40102 -34599
rect -40068 -34633 -40022 -34599
rect -39988 -34633 -39942 -34599
rect -39908 -34633 -39862 -34599
rect -39828 -34633 -39782 -34599
rect -39748 -34633 -39702 -34599
rect -39668 -34633 -39622 -34599
rect -39588 -34633 -39542 -34599
rect -39508 -34633 -39462 -34599
rect -39428 -34633 -39382 -34599
rect -39348 -34633 -39302 -34599
rect -39268 -34633 -39222 -34599
rect -39188 -34633 -39142 -34599
rect -39108 -34633 -39062 -34599
rect -39028 -34633 -38982 -34599
rect -38948 -34633 -38902 -34599
rect -38868 -34633 -38822 -34599
rect -38788 -34633 -38742 -34599
rect -38708 -34633 -38662 -34599
rect -38628 -34633 -38582 -34599
rect -38548 -34633 -38502 -34599
rect -38468 -34633 -38422 -34599
rect -38388 -34633 -38342 -34599
rect -38308 -34633 -38262 -34599
rect -38228 -34633 -38182 -34599
rect -38148 -34633 -38102 -34599
rect -38068 -34633 -38022 -34599
rect -37988 -34633 -37942 -34599
rect -37908 -34633 -37862 -34599
rect -37828 -34633 -37782 -34599
rect -37748 -34633 -37702 -34599
rect -37668 -34633 -37622 -34599
rect -37588 -34633 -37542 -34599
rect -37508 -34633 -37462 -34599
rect -37428 -34633 -37382 -34599
rect -37348 -34633 -37302 -34599
rect -37268 -34633 -37222 -34599
rect -37188 -34633 -37142 -34599
rect -37108 -34633 -37062 -34599
rect -37028 -34633 -36982 -34599
rect -36948 -34633 -36902 -34599
rect -36868 -34633 -36822 -34599
rect -36788 -34633 -36742 -34599
rect -36708 -34633 -36662 -34599
rect -36628 -34633 -36582 -34599
rect -36548 -34633 -36502 -34599
rect -36468 -34633 -36422 -34599
rect -36388 -34633 -36342 -34599
rect -36308 -34633 -36262 -34599
rect -36228 -34633 -36182 -34599
rect -36148 -34633 -36102 -34599
rect -36068 -34633 -36022 -34599
rect -35988 -34633 -35942 -34599
rect -35908 -34633 -35862 -34599
rect -35828 -34633 -35782 -34599
rect -35748 -34633 -35702 -34599
rect -35668 -34633 -35622 -34599
rect -35588 -34633 -35542 -34599
rect -35508 -34633 -35462 -34599
rect -35428 -34633 -35382 -34599
rect -35348 -34633 -35302 -34599
rect -35268 -34633 -35222 -34599
rect -35188 -34633 -35142 -34599
rect -35108 -34633 -35062 -34599
rect -35028 -34633 -34982 -34599
rect -34948 -34633 -34902 -34599
rect -34868 -34633 -34822 -34599
rect -34788 -34633 -34742 -34599
rect -34708 -34633 -34662 -34599
rect -34628 -34633 -34582 -34599
rect -34548 -34633 -34502 -34599
rect -34468 -34633 -34422 -34599
rect -34388 -34633 -34342 -34599
rect -34308 -34633 -34262 -34599
rect -34228 -34633 -34182 -34599
rect -34148 -34633 -34102 -34599
rect -34068 -34633 -34022 -34599
rect -33988 -34633 -33942 -34599
rect -33908 -34633 -33862 -34599
rect -33828 -34633 -33782 -34599
rect -33748 -34633 -33702 -34599
rect -33668 -34633 -33622 -34599
rect -33588 -34633 -33542 -34599
rect -33508 -34633 -33462 -34599
rect -33428 -34633 -33382 -34599
rect -33348 -34633 -33302 -34599
rect -33268 -34633 -33222 -34599
rect -33188 -34633 -33142 -34599
rect -33108 -34633 -33062 -34599
rect -33028 -34633 -32982 -34599
rect -32948 -34633 -32902 -34599
rect -32868 -34633 -32822 -34599
rect -32788 -34633 -32742 -34599
rect -32708 -34633 -32662 -34599
rect -32628 -34633 -32582 -34599
rect -32548 -34633 -32502 -34599
rect -32468 -34633 -32422 -34599
rect -32388 -34633 -32342 -34599
rect -32308 -34633 -32262 -34599
rect -32228 -34633 -32182 -34599
rect -32148 -34633 -32102 -34599
rect -32068 -34633 -32022 -34599
rect -31988 -34633 -31942 -34599
rect -31908 -34633 -31862 -34599
rect -31828 -34633 -31782 -34599
rect -31748 -34633 -31702 -34599
rect -31668 -34633 -31622 -34599
rect -31588 -34633 -31542 -34599
rect -31508 -34633 -31461 -34599
rect -31427 -34633 -31381 -34599
rect -31347 -34633 -31301 -34599
rect -31267 -34633 -31221 -34599
rect -31187 -34633 -31141 -34599
rect -31107 -34633 -31061 -34599
rect -31027 -34633 -30981 -34599
rect -30947 -34633 -30901 -34599
rect -30867 -34633 -30821 -34599
rect -30787 -34633 -30741 -34599
rect -30707 -34633 -30661 -34599
rect -30627 -34633 -30581 -34599
rect -30547 -34633 -30501 -34599
rect -30467 -34633 -30421 -34599
rect -30387 -34633 -30341 -34599
rect -30307 -34633 -30261 -34599
rect -30227 -34633 -30181 -34599
rect -30147 -34633 -30101 -34599
rect -30067 -34633 -30021 -34599
rect -29987 -34633 -29941 -34599
rect -29907 -34633 -29861 -34599
rect -29827 -34633 -29781 -34599
rect -29747 -34633 -29701 -34599
rect -29667 -34633 -29621 -34599
rect -29587 -34633 -29541 -34599
rect -29507 -34633 -29461 -34599
rect -29427 -34633 -29381 -34599
rect -29347 -34633 -29301 -34599
rect -29267 -34633 -29221 -34599
rect -29187 -34633 -29141 -34599
rect -29107 -34633 -29061 -34599
rect -29027 -34633 -28981 -34599
rect -28947 -34633 -28901 -34599
rect -28867 -34633 -28821 -34599
rect -28787 -34633 -28741 -34599
rect -28707 -34633 -28661 -34599
rect -28627 -34633 -28581 -34599
rect -28547 -34633 -28501 -34599
rect -28467 -34633 -28421 -34599
rect -28387 -34633 -28341 -34599
rect -28307 -34633 -28261 -34599
rect -28227 -34633 -28181 -34599
rect -28147 -34633 -28101 -34599
rect -28067 -34633 -28021 -34599
rect -27987 -34633 -27941 -34599
rect -27907 -34633 -27861 -34599
rect -27827 -34633 -27781 -34599
rect -27747 -34633 -27701 -34599
rect -27667 -34633 -27621 -34599
rect -27587 -34633 -27541 -34599
rect -27507 -34633 -27461 -34599
rect -27427 -34633 -27381 -34599
rect -27347 -34633 -27301 -34599
rect -27267 -34633 -27221 -34599
rect -27187 -34633 -27141 -34599
rect -27107 -34633 -27061 -34599
rect -27027 -34633 -26981 -34599
rect -26947 -34633 -26901 -34599
rect -26867 -34633 -26821 -34599
rect -26787 -34633 -26741 -34599
rect -26707 -34633 -26661 -34599
rect -26627 -34633 -26581 -34599
rect -26547 -34633 -26501 -34599
rect -26467 -34633 -26421 -34599
rect -26387 -34633 -26341 -34599
rect -26307 -34633 -26261 -34599
rect -26227 -34633 -26181 -34599
rect -26147 -34633 -26101 -34599
rect -26067 -34633 -26021 -34599
rect -25987 -34633 -25941 -34599
rect -25907 -34633 -25861 -34599
rect -25827 -34633 -25781 -34599
rect -25747 -34633 -25701 -34599
rect -25667 -34633 -25621 -34599
rect -25587 -34633 -25541 -34599
rect -25507 -34633 -25461 -34599
rect -25427 -34633 -25381 -34599
rect -25347 -34633 -25301 -34599
rect -25267 -34633 -25221 -34599
rect -25187 -34633 -25141 -34599
rect -25107 -34633 -25061 -34599
rect -25027 -34633 -24981 -34599
rect -24947 -34633 -24901 -34599
rect -24867 -34633 -24821 -34599
rect -24787 -34633 -24741 -34599
rect -24707 -34633 -24661 -34599
rect -24627 -34633 -24581 -34599
rect -24547 -34633 -24501 -34599
rect -24467 -34633 -24421 -34599
rect -24387 -34633 -24341 -34599
rect -24307 -34633 -24261 -34599
rect -24227 -34633 -24181 -34599
rect -24147 -34633 -24101 -34599
rect -24067 -34633 -24021 -34599
rect -23987 -34633 -23941 -34599
rect -23907 -34633 -23861 -34599
rect -23827 -34633 -23781 -34599
rect -23747 -34633 -23701 -34599
rect -23667 -34633 -23621 -34599
rect -23587 -34633 -23541 -34599
rect -23507 -34633 -23461 -34599
rect -23427 -34633 -23381 -34599
rect -23347 -34633 -23301 -34599
rect -23267 -34633 -23221 -34599
rect -23187 -34633 -23141 -34599
rect -23107 -34633 -23061 -34599
rect -23027 -34633 -22981 -34599
rect -22947 -34633 -22901 -34599
rect -22867 -34633 -22821 -34599
rect -22787 -34633 -22741 -34599
rect -22707 -34633 -22661 -34599
rect -22627 -34633 -22581 -34599
rect -22547 -34633 -22501 -34599
rect -22467 -34633 -22421 -34599
rect -22387 -34633 -22341 -34599
rect -22307 -34633 -22261 -34599
rect -22227 -34633 -22181 -34599
rect -22147 -34633 -22101 -34599
rect -22067 -34633 -22021 -34599
rect -21987 -34633 -21941 -34599
rect -21907 -34633 -21861 -34599
rect -21827 -34633 -21781 -34599
rect -21747 -34633 -21701 -34599
rect -21667 -34633 -21621 -34599
rect -21587 -34633 -21541 -34599
rect -21507 -34633 -21461 -34599
rect -21427 -34633 -21381 -34599
rect -21347 -34633 -21301 -34599
rect -21267 -34633 -21221 -34599
rect -21187 -34633 -21141 -34599
rect -21107 -34633 -21061 -34599
rect -21027 -34633 -20981 -34599
rect -20947 -34633 -20901 -34599
rect -20867 -34633 -20821 -34599
rect -20787 -34633 -20741 -34599
rect -20707 -34633 -20661 -34599
rect -20627 -34633 -20581 -34599
rect -20547 -34633 -20501 -34599
rect -20467 -34633 -20421 -34599
rect -20387 -34633 -20341 -34599
rect -20307 -34633 -20261 -34599
rect -20227 -34633 -20181 -34599
rect -20147 -34633 -20101 -34599
rect -20067 -34633 -20021 -34599
rect -19987 -34633 -19941 -34599
rect -19907 -34633 -19861 -34599
rect -19827 -34633 -19781 -34599
rect -19747 -34633 -19701 -34599
rect -19667 -34633 -19621 -34599
rect -19587 -34633 -19541 -34599
rect -19507 -34633 -19461 -34599
rect -19427 -34633 -19381 -34599
rect -19347 -34633 -19301 -34599
rect -19267 -34633 -19221 -34599
rect -19187 -34633 -19141 -34599
rect -19107 -34633 -19061 -34599
rect -19027 -34633 -18981 -34599
rect -18947 -34633 -18901 -34599
rect -18867 -34633 -18821 -34599
rect -18787 -34633 -18741 -34599
rect -18707 -34633 -18661 -34599
rect -18627 -34633 -18581 -34599
rect -18547 -34633 -18500 -34599
rect -18466 -34633 -18420 -34599
rect -18386 -34633 -18340 -34599
rect -18306 -34633 -18260 -34599
rect -18226 -34633 -18180 -34599
rect -18146 -34633 -18100 -34599
rect -18066 -34633 -18020 -34599
rect -17986 -34633 -17940 -34599
rect -17906 -34633 -17860 -34599
rect -17826 -34633 -17780 -34599
rect -17746 -34633 -17700 -34599
rect -17666 -34633 -17620 -34599
rect -17586 -34633 -17540 -34599
rect -17506 -34633 -17460 -34599
rect -17426 -34633 -17380 -34599
rect -17346 -34633 -17300 -34599
rect -17266 -34633 -17220 -34599
rect -17186 -34633 -17140 -34599
rect -17106 -34633 -17060 -34599
rect -17026 -34633 -16980 -34599
rect -16946 -34633 -16900 -34599
rect -16866 -34633 -16820 -34599
rect -16786 -34633 -16740 -34599
rect -16706 -34633 -16660 -34599
rect -16626 -34633 -16580 -34599
rect -16546 -34633 -16500 -34599
rect -16466 -34633 -16420 -34599
rect -16386 -34633 -16340 -34599
rect -16306 -34633 -16260 -34599
rect -16226 -34633 -16180 -34599
rect -16146 -34633 -16100 -34599
rect -16066 -34633 -16020 -34599
rect -15986 -34633 -15940 -34599
rect -15906 -34633 -15860 -34599
rect -15826 -34633 -15780 -34599
rect -15746 -34633 -15700 -34599
rect -15666 -34633 -15620 -34599
rect -15586 -34633 -15540 -34599
rect -15506 -34633 -15460 -34599
rect -15426 -34633 -15380 -34599
rect -15346 -34633 -15300 -34599
rect -15266 -34633 -15220 -34599
rect -15186 -34633 -15140 -34599
rect -15106 -34633 -15060 -34599
rect -15026 -34633 -14980 -34599
rect -14946 -34633 -14900 -34599
rect -14866 -34633 -14820 -34599
rect -14786 -34633 -14740 -34599
rect -14706 -34633 -14660 -34599
rect -14626 -34633 -14580 -34599
rect -14546 -34633 -14500 -34599
rect -14466 -34633 -14420 -34599
rect -14386 -34633 -14340 -34599
rect -14306 -34633 -14260 -34599
rect -14226 -34633 -14180 -34599
rect -14146 -34633 -14100 -34599
rect -14066 -34633 -14020 -34599
rect -13986 -34633 -13940 -34599
rect -13906 -34633 -13860 -34599
rect -13826 -34633 -13780 -34599
rect -13746 -34633 -13700 -34599
rect -13666 -34633 -13620 -34599
rect -13586 -34633 -13540 -34599
rect -13506 -34633 -13460 -34599
rect -13426 -34633 -13380 -34599
rect -13346 -34633 -13300 -34599
rect -13266 -34633 -13220 -34599
rect -13186 -34633 -13140 -34599
rect -13106 -34633 -13060 -34599
rect -13026 -34633 -12980 -34599
rect -12946 -34633 -12900 -34599
rect -12866 -34633 -12820 -34599
rect -12786 -34633 -12740 -34599
rect -12706 -34633 -12660 -34599
rect -12626 -34633 -12580 -34599
rect -12546 -34633 -12500 -34599
rect -12466 -34633 -12420 -34599
rect -12386 -34633 -12340 -34599
rect -12306 -34633 -12260 -34599
rect -12226 -34633 -12180 -34599
rect -12146 -34633 -12100 -34599
rect -12066 -34633 -12020 -34599
rect -11986 -34633 -11940 -34599
rect -11906 -34633 -11860 -34599
rect -11826 -34633 -11780 -34599
rect -11746 -34633 -11700 -34599
rect -11666 -34633 -11620 -34599
rect -11586 -34633 -11540 -34599
rect -11506 -34633 -11460 -34599
rect -11426 -34633 -11380 -34599
rect -11346 -34633 -11300 -34599
rect -11266 -34633 -11220 -34599
rect -11186 -34633 -11140 -34599
rect -11106 -34633 -11060 -34599
rect -11026 -34633 -10980 -34599
rect -10946 -34633 -10900 -34599
rect -10866 -34633 -10820 -34599
rect -10786 -34633 -10740 -34599
rect -10706 -34633 -10660 -34599
rect -10626 -34633 -10580 -34599
rect -10546 -34633 -10500 -34599
rect -10466 -34633 -10420 -34599
rect -10386 -34633 -10340 -34599
rect -10306 -34633 -10260 -34599
rect -10226 -34633 -10180 -34599
rect -10146 -34633 -10100 -34599
rect -10066 -34633 -10020 -34599
rect -9986 -34633 -9940 -34599
rect -9906 -34633 -9859 -34599
rect -9825 -34633 -9779 -34599
rect -9745 -34633 -9699 -34599
rect -9665 -34633 -9619 -34599
rect -9585 -34633 -9539 -34599
rect -9505 -34633 -9459 -34599
rect -9425 -34633 -9379 -34599
rect -9345 -34633 -9299 -34599
rect -9265 -34633 -9219 -34599
rect -9185 -34633 -9139 -34599
rect -9105 -34633 -9059 -34599
rect -9025 -34633 -8979 -34599
rect -8945 -34633 -8899 -34599
rect -8865 -34633 -8819 -34599
rect -8785 -34633 -8739 -34599
rect -8705 -34633 -8659 -34599
rect -8625 -34633 -8579 -34599
rect -8545 -34633 -8499 -34599
rect -8465 -34633 -8419 -34599
rect -8385 -34633 -8339 -34599
rect -8305 -34633 -8259 -34599
rect -8225 -34633 -8179 -34599
rect -8145 -34633 -8099 -34599
rect -8065 -34633 -8019 -34599
rect -7985 -34633 -7939 -34599
rect -7905 -34633 -7859 -34599
rect -7825 -34633 -7779 -34599
rect -7745 -34633 -7699 -34599
rect -7665 -34633 -7619 -34599
rect -7585 -34633 -7539 -34599
rect -7505 -34633 -7459 -34599
rect -7425 -34633 -7379 -34599
rect -7345 -34633 -7299 -34599
rect -7265 -34633 -7219 -34599
rect -7185 -34633 -7139 -34599
rect -7105 -34633 -7059 -34599
rect -7025 -34633 -6979 -34599
rect -6945 -34633 -6899 -34599
rect -6865 -34633 -6819 -34599
rect -6785 -34633 -6739 -34599
rect -6705 -34633 -6659 -34599
rect -6625 -34633 -6579 -34599
rect -6545 -34633 -6499 -34599
rect -6465 -34633 -6419 -34599
rect -6385 -34633 -6339 -34599
rect -6305 -34633 -6259 -34599
rect -6225 -34633 -6179 -34599
rect -6145 -34633 -6099 -34599
rect -6065 -34633 -6019 -34599
rect -5985 -34633 -5939 -34599
rect -5905 -34633 -5859 -34599
rect -5825 -34633 -5779 -34599
rect -5745 -34633 -5699 -34599
rect -5665 -34633 -5619 -34599
rect -5585 -34633 -5539 -34599
rect -5505 -34633 -5459 -34599
rect -5425 -34633 -5379 -34599
rect -5345 -34633 -5299 -34599
rect -5265 -34633 -5219 -34599
rect -5185 -34633 -5139 -34599
rect -5105 -34633 -5059 -34599
rect -5025 -34633 -4979 -34599
rect -4945 -34633 -4899 -34599
rect -4865 -34633 -4819 -34599
rect -4785 -34633 -4739 -34599
rect -4705 -34633 -4659 -34599
rect -4625 -34633 -4579 -34599
rect -4545 -34633 -4499 -34599
rect -4465 -34633 -4419 -34599
rect -4385 -34633 -4339 -34599
rect -4305 -34633 -4259 -34599
rect -4225 -34633 -4140 -34599
rect -4106 -34633 -4060 -34599
rect -4026 -34633 -3980 -34599
rect -3946 -34633 -3900 -34599
rect -3866 -34633 -3820 -34599
rect -3786 -34633 -3740 -34599
rect -3706 -34633 -3660 -34599
rect -3626 -34633 -3580 -34599
rect -3546 -34633 -3500 -34599
rect -3466 -34633 -3420 -34599
rect -3386 -34633 -3340 -34599
rect -3306 -34633 -3260 -34599
rect -3226 -34633 -3180 -34599
rect -3146 -34633 -3100 -34599
rect -3066 -34633 -3020 -34599
rect -2986 -34633 -2940 -34599
rect -2906 -34633 -2860 -34599
rect -2826 -34633 -2780 -34599
rect -2746 -34633 -2700 -34599
rect -2666 -34633 -2620 -34599
rect -2586 -34633 -2540 -34599
rect -2506 -34633 -2460 -34599
rect -2426 -34633 -2380 -34599
rect -2346 -34633 -2300 -34599
rect -2266 -34633 -2220 -34599
rect -2186 -34633 -2140 -34599
rect -2106 -34633 -2060 -34599
rect -2026 -34633 -1980 -34599
rect -1946 -34633 -1900 -34599
rect -1866 -34633 -1820 -34599
rect -1786 -34633 -1740 -34599
rect -1706 -34633 -1660 -34599
rect -1626 -34633 -1580 -34599
rect -1546 -34633 -1500 -34599
rect -1466 -34633 -1420 -34599
rect -1386 -34633 -1340 -34599
rect -1306 -34633 -1260 -34599
rect -1226 -34633 -1180 -34599
rect -1146 -34633 -1100 -34599
rect -1066 -34633 -1020 -34599
rect -986 -34633 -940 -34599
rect -906 -34633 -860 -34599
rect -826 -34633 -780 -34599
rect -746 -34633 -700 -34599
rect -666 -34633 -620 -34599
rect -586 -34633 -540 -34599
rect -506 -34633 -460 -34599
rect -426 -34633 -380 -34599
rect -346 -34633 -300 -34599
rect -266 -34633 -220 -34599
rect -186 -34633 -140 -34599
rect -106 -34633 -60 -34599
rect -26 -34633 20 -34599
rect 54 -34633 100 -34599
rect 134 -34633 180 -34599
rect 214 -34633 260 -34599
rect 294 -34633 340 -34599
rect 374 -34633 420 -34599
rect 454 -34633 500 -34599
rect 534 -34633 580 -34599
rect 614 -34633 660 -34599
rect 694 -34633 740 -34599
rect 774 -34633 820 -34599
rect 854 -34633 900 -34599
rect 934 -34633 980 -34599
rect 1014 -34633 1060 -34599
rect 1094 -34633 1140 -34599
rect 1174 -34633 1220 -34599
rect 1254 -34633 1300 -34599
rect 1334 -34633 1380 -34599
rect 1414 -34633 1460 -34599
rect 1494 -34633 1540 -34599
rect 1574 -34633 1620 -34599
rect 1654 -34633 1700 -34599
rect 1734 -34633 1780 -34599
rect 1814 -34633 1860 -34599
rect 1894 -34633 1940 -34599
rect 1974 -34633 2020 -34599
rect 2054 -34633 2100 -34599
rect 2134 -34633 2180 -34599
rect 2214 -34633 2260 -34599
rect 2294 -34633 2340 -34599
rect 2374 -34633 2420 -34599
rect 2454 -34633 2500 -34599
rect 2534 -34633 2580 -34599
rect 2614 -34633 2660 -34599
rect 2694 -34633 2740 -34599
rect 2774 -34633 2820 -34599
rect 2854 -34633 2900 -34599
rect 2934 -34633 2980 -34599
rect 3014 -34633 3060 -34599
rect 3094 -34633 3140 -34599
rect 3174 -34633 3220 -34599
rect 3254 -34633 3300 -34599
rect 3334 -34633 3380 -34599
rect 3414 -34633 3460 -34599
rect 3494 -34633 3540 -34599
rect 3574 -34633 3620 -34599
rect 3654 -34633 3700 -34599
rect 3734 -34633 3780 -34599
rect 3814 -34633 3860 -34599
rect 3894 -34633 3940 -34599
rect 3974 -34633 4020 -34599
rect 4054 -34633 4100 -34599
rect 4134 -34633 4180 -34599
rect 4214 -34633 4260 -34599
rect 4294 -34633 4340 -34599
rect 4374 -34633 4420 -34599
rect 4454 -34633 4500 -34599
rect 4534 -34633 4580 -34599
rect 4614 -34633 4660 -34599
rect 4694 -34633 4740 -34599
rect 4774 -34633 4820 -34599
rect 4854 -34633 4900 -34599
rect 4934 -34633 4980 -34599
rect 5014 -34633 5060 -34599
rect 5094 -34633 5140 -34599
rect 5174 -34633 5220 -34599
rect 5254 -34633 5300 -34599
rect 5334 -34633 5380 -34599
rect 5414 -34633 5460 -34599
rect 5494 -34633 5540 -34599
rect 5574 -34633 5620 -34599
rect 5654 -34633 5700 -34599
rect 5734 -34633 5780 -34599
rect 5814 -34633 5860 -34599
rect 5894 -34633 5940 -34599
rect 5974 -34633 6020 -34599
rect 6054 -34633 6100 -34599
rect 6134 -34633 6180 -34599
rect 6214 -34633 6260 -34599
rect 6294 -34633 6340 -34599
rect 6374 -34633 6420 -34599
rect 6454 -34633 6500 -34599
rect 6534 -34633 6580 -34599
rect 6614 -34633 6660 -34599
rect 6694 -34633 6740 -34599
rect 6774 -34633 6820 -34599
rect 6854 -34633 6900 -34599
rect 6934 -34633 6980 -34599
rect 7014 -34633 7060 -34599
rect 7094 -34633 7140 -34599
rect 7174 -34633 7220 -34599
rect 7254 -34633 7300 -34599
rect 7334 -34633 7380 -34599
rect 7414 -34633 7460 -34599
rect 7494 -34633 7540 -34599
rect 7574 -34633 7620 -34599
rect 7654 -34633 7700 -34599
rect 7734 -34633 7780 -34599
rect 7814 -34633 7860 -34599
rect 7894 -34633 7940 -34599
rect 7974 -34633 8020 -34599
rect 8054 -34633 8100 -34599
rect 8134 -34633 8180 -34599
rect 8214 -34633 8260 -34599
rect 8294 -34633 8340 -34599
rect 8374 -34633 8420 -34599
rect 8454 -34633 8500 -34599
rect 8534 -34633 8580 -34599
rect 8614 -34633 8660 -34599
rect 8694 -34633 8740 -34599
rect 8774 -34633 8820 -34599
rect 8854 -34633 8900 -34599
rect 8934 -34633 8980 -34599
rect 9014 -34633 9060 -34599
rect 9094 -34633 9140 -34599
rect 9174 -34633 9220 -34599
rect 9254 -34633 9300 -34599
rect 9334 -34633 9380 -34599
rect 9414 -34633 9460 -34599
rect 9494 -34633 9540 -34599
rect 9574 -34633 9620 -34599
rect 9654 -34633 9700 -34599
rect 9734 -34633 9780 -34599
rect 9814 -34633 9860 -34599
rect 9894 -34633 9940 -34599
rect 9974 -34633 10020 -34599
rect 10054 -34633 10100 -34599
rect 10134 -34633 10181 -34599
rect 10215 -34633 10261 -34599
rect 10295 -34633 10341 -34599
rect 10375 -34633 10421 -34599
rect 10455 -34633 10501 -34599
rect 10535 -34633 10581 -34599
rect 10615 -34633 10661 -34599
rect 10695 -34633 10741 -34599
rect 10775 -34633 10821 -34599
rect 10855 -34633 10901 -34599
rect 10935 -34633 10981 -34599
rect 11015 -34633 11061 -34599
rect 11095 -34633 11141 -34599
rect 11175 -34633 11221 -34599
rect 11255 -34633 11301 -34599
rect 11335 -34633 11381 -34599
rect 11415 -34633 11461 -34599
rect 11495 -34633 11541 -34599
rect 11575 -34633 11621 -34599
rect 11655 -34633 11701 -34599
rect 11735 -34633 11781 -34599
rect 11815 -34633 11861 -34599
rect 11895 -34633 11941 -34599
rect 11975 -34633 12021 -34599
rect 12055 -34633 12101 -34599
rect 12135 -34633 12181 -34599
rect 12215 -34633 12261 -34599
rect 12295 -34633 12341 -34599
rect 12375 -34633 12421 -34599
rect 12455 -34633 12501 -34599
rect 12535 -34633 12581 -34599
rect 12615 -34633 12661 -34599
rect 12695 -34633 12741 -34599
rect 12775 -34633 12821 -34599
rect 12855 -34633 12901 -34599
rect 12935 -34633 12981 -34599
rect 13015 -34633 13061 -34599
rect 13095 -34633 13141 -34599
rect 13175 -34633 13221 -34599
rect 13255 -34633 13301 -34599
rect 13335 -34633 13381 -34599
rect 13415 -34633 13461 -34599
rect 13495 -34633 13541 -34599
rect 13575 -34633 13621 -34599
rect 13655 -34633 13701 -34599
rect 13735 -34633 13781 -34599
rect 13815 -34633 13861 -34599
rect 13895 -34633 13941 -34599
rect 13975 -34633 14021 -34599
rect 14055 -34633 14101 -34599
rect 14135 -34633 14181 -34599
rect 14215 -34633 14261 -34599
rect 14295 -34633 14341 -34599
rect 14375 -34633 14421 -34599
rect 14455 -34633 14501 -34599
rect 14535 -34633 14581 -34599
rect 14615 -34633 14661 -34599
rect 14695 -34633 14741 -34599
rect 14775 -34633 14821 -34599
rect 14855 -34633 14901 -34599
rect 14935 -34633 14981 -34599
rect 15015 -34633 15061 -34599
rect 15095 -34633 15141 -34599
rect 15175 -34633 15221 -34599
rect 15255 -34633 15301 -34599
rect 15335 -34633 15381 -34599
rect 15415 -34633 15461 -34599
rect 15495 -34633 15541 -34599
rect 15575 -34633 15621 -34599
rect 15655 -34633 15701 -34599
rect 15735 -34633 15781 -34599
rect 15815 -34633 15861 -34599
rect 15895 -34633 15941 -34599
rect 15975 -34633 16021 -34599
rect 16055 -34633 16101 -34599
rect 16135 -34633 16181 -34599
rect 16215 -34633 16261 -34599
rect 16295 -34633 16341 -34599
rect 16375 -34633 16421 -34599
rect 16455 -34633 16501 -34599
rect 16535 -34633 16581 -34599
rect 16615 -34633 16661 -34599
rect 16695 -34633 16741 -34599
rect 16775 -34633 16821 -34599
rect 16855 -34633 16901 -34599
rect 16935 -34633 16981 -34599
rect 17015 -34633 17061 -34599
rect 17095 -34633 17141 -34599
rect 17175 -34633 17221 -34599
rect 17255 -34633 17301 -34599
rect 17335 -34633 17381 -34599
rect 17415 -34633 17461 -34599
rect 17495 -34633 17541 -34599
rect 17575 -34633 17621 -34599
rect 17655 -34633 17701 -34599
rect 17735 -34633 17781 -34599
rect 17815 -34633 17861 -34599
rect 17895 -34633 17941 -34599
rect 17975 -34633 18021 -34599
rect 18055 -34633 18101 -34599
rect 18135 -34633 18181 -34599
rect 18215 -34633 18261 -34599
rect 18295 -34633 18341 -34599
rect 18375 -34633 18421 -34599
rect 18455 -34633 18501 -34599
rect 18535 -34633 18581 -34599
rect 18615 -34633 18661 -34599
rect 18695 -34633 18741 -34599
rect 18775 -34633 18821 -34599
rect 18855 -34633 18901 -34599
rect 18935 -34633 18981 -34599
rect 19015 -34633 19061 -34599
rect 19095 -34633 19141 -34599
rect 19175 -34633 19221 -34599
rect 19255 -34633 19301 -34599
rect 19335 -34633 19381 -34599
rect 19415 -34633 19461 -34599
rect 19495 -34633 19541 -34599
rect 19575 -34633 19621 -34599
rect 19655 -34633 19701 -34599
rect 19735 -34633 19781 -34599
rect 19815 -34633 19861 -34599
rect 19895 -34633 19941 -34599
rect 19975 -34633 20021 -34599
rect 20055 -34633 20101 -34599
rect 20135 -34633 20181 -34599
rect 20215 -34633 20261 -34599
rect 20295 -34633 20341 -34599
rect 20375 -34633 20421 -34599
rect 20455 -34633 20501 -34599
rect 20535 -34633 20581 -34599
rect 20615 -34633 20661 -34599
rect 20695 -34633 20741 -34599
rect 20775 -34633 20821 -34599
rect 20855 -34633 20901 -34599
rect 20935 -34633 20981 -34599
rect 21015 -34633 21061 -34599
rect 21095 -34633 21141 -34599
rect 21175 -34633 21221 -34599
rect 21255 -34633 21301 -34599
rect 21335 -34633 21381 -34599
rect 21415 -34633 21461 -34599
rect 21495 -34633 21541 -34599
rect 21575 -34633 21621 -34599
rect 21655 -34633 21701 -34599
rect 21735 -34633 21781 -34599
rect 21815 -34633 21861 -34599
rect 21895 -34633 21941 -34599
rect 21975 -34633 22021 -34599
rect 22055 -34633 22101 -34599
rect 22135 -34633 22181 -34599
rect 22215 -34633 22261 -34599
rect 22295 -34633 22341 -34599
rect 22375 -34633 22421 -34599
rect 22455 -34633 22501 -34599
rect 22535 -34633 22581 -34599
rect 22615 -34633 22661 -34599
rect 22695 -34633 22741 -34599
rect 22775 -34633 22821 -34599
rect 22855 -34633 22901 -34599
rect 22935 -34633 22981 -34599
rect 23015 -34633 23061 -34599
rect 23095 -34633 23141 -34599
rect 23175 -34633 23221 -34599
rect 23255 -34633 23301 -34599
rect 23335 -34633 23381 -34599
rect 23415 -34633 23461 -34599
rect 23495 -34633 23541 -34599
rect 23575 -34633 23621 -34599
rect 23655 -34633 23701 -34599
rect 23735 -34633 23781 -34599
rect 23815 -34633 23861 -34599
rect 23895 -34633 23941 -34599
rect 23975 -34633 24021 -34599
rect 24055 -34633 24101 -34599
rect 24135 -34633 24181 -34599
rect 24215 -34633 24261 -34599
rect 24295 -34633 24341 -34599
rect 24375 -34633 24421 -34599
rect 24455 -34633 24501 -34599
rect 24535 -34633 24581 -34599
rect 24615 -34633 24661 -34599
rect 24695 -34633 24741 -34599
rect 24775 -34633 24821 -34599
rect 24855 -34633 24901 -34599
rect 24935 -34633 24981 -34599
rect 25015 -34633 25061 -34599
rect 25095 -34633 25141 -34599
rect 25175 -34633 25221 -34599
rect 25255 -34633 25301 -34599
rect 25335 -34633 25381 -34599
rect 25415 -34633 25461 -34599
rect 25495 -34633 25541 -34599
rect 25575 -34633 25621 -34599
rect 25655 -34633 25701 -34599
rect 25735 -34633 25781 -34599
rect 25815 -34633 25861 -34599
rect 25895 -34633 25941 -34599
rect 25975 -34633 26021 -34599
rect 26055 -34633 26101 -34599
rect 26135 -34633 26181 -34599
rect 26215 -34633 26261 -34599
rect 26295 -34633 26341 -34599
rect 26375 -34633 26421 -34599
rect 26455 -34633 26501 -34599
rect 26535 -34633 26581 -34599
rect 26615 -34633 26661 -34599
rect 26695 -34633 26741 -34599
rect 26775 -34633 26821 -34599
rect 26855 -34633 26901 -34599
rect 26935 -34633 26981 -34599
rect 27015 -34633 27061 -34599
rect 27095 -34633 27141 -34599
rect 27175 -34633 27221 -34599
rect 27255 -34633 27301 -34599
rect 27335 -34633 27381 -34599
rect 27415 -34633 27461 -34599
rect 27495 -34633 27541 -34599
rect 27575 -34633 27621 -34599
rect 27655 -34633 27701 -34599
rect 27735 -34633 27781 -34599
rect 27815 -34633 27861 -34599
rect 27895 -34633 27941 -34599
rect 27975 -34633 28021 -34599
rect 28055 -34633 28101 -34599
rect 28135 -34633 28181 -34599
rect 28215 -34633 28261 -34599
rect 28295 -34633 28341 -34599
rect 28375 -34633 28421 -34599
rect 28455 -34633 28501 -34599
rect 28535 -34633 28581 -34599
rect 28615 -34633 28661 -34599
rect 28695 -34633 28741 -34599
rect 28775 -34633 28821 -34599
rect 28855 -34633 28901 -34599
rect 28935 -34633 28981 -34599
rect 29015 -34633 29061 -34599
rect 29095 -34633 29141 -34599
rect 29175 -34633 29221 -34599
rect 29255 -34633 29301 -34599
rect 29335 -34633 29381 -34599
rect 29415 -34633 29461 -34599
rect 29495 -34633 29541 -34599
rect 29575 -34633 29621 -34599
rect 29655 -34633 29701 -34599
rect 29735 -34633 29781 -34599
rect 29815 -34633 29861 -34599
rect 29895 -34633 29941 -34599
rect 29975 -34633 30021 -34599
rect 30055 -34633 30101 -34599
rect 30135 -34633 30181 -34599
rect 30215 -34633 30261 -34599
rect 30295 -34633 30341 -34599
rect 30375 -34633 30421 -34599
rect 30455 -34633 30501 -34599
rect 30535 -34633 30581 -34599
rect 30615 -34633 30661 -34599
rect 30695 -34633 30741 -34599
rect 30775 -34633 30821 -34599
rect 30855 -34633 30901 -34599
rect 30935 -34633 30981 -34599
rect 31015 -34633 31061 -34599
rect 31095 -34633 31141 -34599
rect 31175 -34633 31221 -34599
rect 31255 -34633 31301 -34599
rect 31335 -34633 31381 -34599
rect 31415 -34633 31461 -34599
rect 31495 -34633 31541 -34599
rect 31575 -34633 31621 -34599
rect 31655 -34633 31701 -34599
rect 31735 -34633 31781 -34599
rect -44482 -34666 31781 -34633
rect -44482 -42425 -43986 -34666
rect -27284 -34710 -27024 -34666
rect -27284 -34762 -27240 -34710
rect -27188 -34762 -27120 -34710
rect -27068 -34762 -27024 -34710
rect -27284 -34830 -27024 -34762
rect -27284 -34882 -27240 -34830
rect -27188 -34882 -27120 -34830
rect -27068 -34882 -27024 -34830
rect -27284 -34926 -27024 -34882
rect 12051 -34711 12311 -34666
rect 12051 -34763 12095 -34711
rect 12147 -34763 12215 -34711
rect 12267 -34763 12311 -34711
rect 12051 -34831 12311 -34763
rect 12051 -34883 12095 -34831
rect 12147 -34883 12215 -34831
rect 12267 -34883 12311 -34831
rect 12051 -34927 12311 -34883
rect -44482 -42458 -624 -42425
rect -44482 -42492 -44422 -42458
rect -44388 -42492 -44342 -42458
rect -44308 -42492 -44262 -42458
rect -44228 -42492 -44182 -42458
rect -44148 -42492 -44102 -42458
rect -44068 -42492 -44022 -42458
rect -43988 -42492 -43942 -42458
rect -43908 -42492 -43862 -42458
rect -43828 -42492 -43782 -42458
rect -43748 -42492 -43702 -42458
rect -43668 -42492 -43622 -42458
rect -43588 -42492 -43542 -42458
rect -43508 -42492 -43462 -42458
rect -43428 -42492 -43382 -42458
rect -43348 -42492 -43302 -42458
rect -43268 -42492 -43222 -42458
rect -43188 -42492 -43142 -42458
rect -43108 -42492 -43062 -42458
rect -43028 -42492 -42982 -42458
rect -42948 -42492 -42902 -42458
rect -42868 -42492 -42822 -42458
rect -42788 -42492 -42742 -42458
rect -42708 -42492 -42662 -42458
rect -42628 -42492 -42582 -42458
rect -42548 -42492 -42502 -42458
rect -42468 -42492 -42422 -42458
rect -42388 -42492 -42342 -42458
rect -42308 -42492 -42262 -42458
rect -42228 -42492 -42182 -42458
rect -42148 -42492 -42102 -42458
rect -42068 -42492 -42022 -42458
rect -41988 -42492 -41942 -42458
rect -41908 -42492 -41862 -42458
rect -41828 -42492 -41782 -42458
rect -41748 -42492 -41702 -42458
rect -41668 -42492 -41622 -42458
rect -41588 -42492 -41542 -42458
rect -41508 -42492 -41462 -42458
rect -41428 -42492 -41382 -42458
rect -41348 -42492 -41302 -42458
rect -41268 -42492 -41222 -42458
rect -41188 -42492 -41142 -42458
rect -41108 -42492 -41062 -42458
rect -41028 -42492 -40982 -42458
rect -40948 -42492 -40902 -42458
rect -40868 -42492 -40822 -42458
rect -40788 -42492 -40742 -42458
rect -40708 -42492 -40662 -42458
rect -40628 -42492 -40582 -42458
rect -40548 -42492 -40502 -42458
rect -40468 -42492 -40422 -42458
rect -40388 -42492 -40342 -42458
rect -40308 -42492 -40262 -42458
rect -40228 -42492 -40182 -42458
rect -40148 -42492 -40102 -42458
rect -40068 -42492 -40022 -42458
rect -39988 -42492 -39942 -42458
rect -39908 -42492 -39862 -42458
rect -39828 -42492 -39782 -42458
rect -39748 -42492 -39702 -42458
rect -39668 -42492 -39622 -42458
rect -39588 -42492 -39542 -42458
rect -39508 -42492 -39462 -42458
rect -39428 -42492 -39382 -42458
rect -39348 -42492 -39302 -42458
rect -39268 -42492 -39222 -42458
rect -39188 -42492 -39142 -42458
rect -39108 -42492 -39062 -42458
rect -39028 -42492 -38982 -42458
rect -38948 -42492 -38902 -42458
rect -38868 -42492 -38822 -42458
rect -38788 -42492 -38742 -42458
rect -38708 -42492 -38662 -42458
rect -38628 -42492 -38582 -42458
rect -38548 -42492 -38502 -42458
rect -38468 -42492 -38422 -42458
rect -38388 -42492 -38342 -42458
rect -38308 -42492 -38262 -42458
rect -38228 -42492 -38182 -42458
rect -38148 -42492 -38102 -42458
rect -38068 -42492 -38022 -42458
rect -37988 -42492 -37942 -42458
rect -37908 -42492 -37862 -42458
rect -37828 -42492 -37782 -42458
rect -37748 -42492 -37702 -42458
rect -37668 -42492 -37622 -42458
rect -37588 -42492 -37542 -42458
rect -37508 -42492 -37462 -42458
rect -37428 -42492 -37382 -42458
rect -37348 -42492 -37302 -42458
rect -37268 -42492 -37222 -42458
rect -37188 -42492 -37142 -42458
rect -37108 -42492 -37062 -42458
rect -37028 -42492 -36982 -42458
rect -36948 -42492 -36902 -42458
rect -36868 -42492 -36822 -42458
rect -36788 -42492 -36742 -42458
rect -36708 -42492 -36662 -42458
rect -36628 -42492 -36582 -42458
rect -36548 -42492 -36502 -42458
rect -36468 -42492 -36422 -42458
rect -36388 -42492 -36342 -42458
rect -36308 -42492 -36262 -42458
rect -36228 -42492 -36182 -42458
rect -36148 -42492 -36102 -42458
rect -36068 -42492 -36022 -42458
rect -35988 -42492 -35942 -42458
rect -35908 -42492 -35862 -42458
rect -35828 -42492 -35782 -42458
rect -35748 -42492 -35702 -42458
rect -35668 -42492 -35622 -42458
rect -35588 -42492 -35542 -42458
rect -35508 -42492 -35462 -42458
rect -35428 -42492 -35382 -42458
rect -35348 -42492 -35302 -42458
rect -35268 -42492 -35222 -42458
rect -35188 -42492 -35142 -42458
rect -35108 -42492 -35062 -42458
rect -35028 -42492 -34982 -42458
rect -34948 -42492 -34902 -42458
rect -34868 -42492 -34822 -42458
rect -34788 -42492 -34742 -42458
rect -34708 -42492 -34662 -42458
rect -34628 -42492 -34582 -42458
rect -34548 -42492 -34502 -42458
rect -34468 -42492 -34422 -42458
rect -34388 -42492 -34342 -42458
rect -34308 -42492 -34262 -42458
rect -34228 -42492 -34182 -42458
rect -34148 -42492 -34102 -42458
rect -34068 -42492 -34022 -42458
rect -33988 -42492 -33942 -42458
rect -33908 -42492 -33862 -42458
rect -33828 -42492 -33782 -42458
rect -33748 -42492 -33702 -42458
rect -33668 -42492 -33622 -42458
rect -33588 -42492 -33542 -42458
rect -33508 -42492 -33462 -42458
rect -33428 -42492 -33382 -42458
rect -33348 -42492 -33302 -42458
rect -33268 -42492 -33222 -42458
rect -33188 -42492 -33142 -42458
rect -33108 -42492 -33062 -42458
rect -33028 -42492 -32982 -42458
rect -32948 -42492 -32902 -42458
rect -32868 -42492 -32822 -42458
rect -32788 -42492 -32742 -42458
rect -32708 -42492 -32662 -42458
rect -32628 -42492 -32582 -42458
rect -32548 -42492 -32502 -42458
rect -32468 -42492 -32422 -42458
rect -32388 -42492 -32342 -42458
rect -32308 -42492 -32262 -42458
rect -32228 -42492 -32182 -42458
rect -32148 -42492 -32102 -42458
rect -32068 -42492 -32022 -42458
rect -31988 -42492 -31942 -42458
rect -31908 -42492 -31862 -42458
rect -31828 -42492 -31782 -42458
rect -31748 -42492 -31702 -42458
rect -31668 -42492 -31622 -42458
rect -31588 -42492 -31542 -42458
rect -31508 -42492 -31461 -42458
rect -31427 -42492 -31381 -42458
rect -31347 -42492 -31301 -42458
rect -31267 -42492 -31221 -42458
rect -31187 -42492 -31141 -42458
rect -31107 -42492 -31061 -42458
rect -31027 -42492 -30981 -42458
rect -30947 -42492 -30901 -42458
rect -30867 -42492 -30821 -42458
rect -30787 -42492 -30741 -42458
rect -30707 -42492 -30661 -42458
rect -30627 -42492 -30581 -42458
rect -30547 -42492 -30501 -42458
rect -30467 -42492 -30421 -42458
rect -30387 -42492 -30341 -42458
rect -30307 -42492 -30261 -42458
rect -30227 -42492 -30181 -42458
rect -30147 -42492 -30101 -42458
rect -30067 -42492 -30021 -42458
rect -29987 -42492 -29941 -42458
rect -29907 -42492 -29861 -42458
rect -29827 -42492 -29781 -42458
rect -29747 -42492 -29701 -42458
rect -29667 -42492 -29621 -42458
rect -29587 -42492 -29541 -42458
rect -29507 -42492 -29461 -42458
rect -29427 -42492 -29381 -42458
rect -29347 -42492 -29301 -42458
rect -29267 -42492 -29221 -42458
rect -29187 -42492 -29141 -42458
rect -29107 -42492 -29061 -42458
rect -29027 -42492 -28981 -42458
rect -28947 -42492 -28901 -42458
rect -28867 -42492 -28821 -42458
rect -28787 -42492 -28741 -42458
rect -28707 -42492 -28661 -42458
rect -28627 -42492 -28581 -42458
rect -28547 -42492 -28501 -42458
rect -28467 -42492 -28421 -42458
rect -28387 -42492 -28341 -42458
rect -28307 -42492 -28261 -42458
rect -28227 -42492 -28181 -42458
rect -28147 -42492 -28101 -42458
rect -28067 -42492 -28021 -42458
rect -27987 -42492 -27941 -42458
rect -27907 -42492 -27861 -42458
rect -27827 -42492 -27781 -42458
rect -27747 -42492 -27701 -42458
rect -27667 -42492 -27621 -42458
rect -27587 -42492 -27541 -42458
rect -27507 -42492 -27461 -42458
rect -27427 -42492 -27381 -42458
rect -27347 -42492 -27301 -42458
rect -27267 -42492 -27221 -42458
rect -27187 -42492 -27141 -42458
rect -27107 -42492 -27061 -42458
rect -27027 -42492 -26981 -42458
rect -26947 -42492 -26901 -42458
rect -26867 -42492 -26821 -42458
rect -26787 -42492 -26741 -42458
rect -26707 -42492 -26661 -42458
rect -26627 -42492 -26581 -42458
rect -26547 -42492 -26501 -42458
rect -26467 -42492 -26421 -42458
rect -26387 -42492 -26341 -42458
rect -26307 -42492 -26261 -42458
rect -26227 -42492 -26181 -42458
rect -26147 -42492 -26101 -42458
rect -26067 -42492 -26021 -42458
rect -25987 -42492 -25941 -42458
rect -25907 -42492 -25861 -42458
rect -25827 -42492 -25781 -42458
rect -25747 -42492 -25701 -42458
rect -25667 -42492 -25621 -42458
rect -25587 -42492 -25541 -42458
rect -25507 -42492 -25461 -42458
rect -25427 -42492 -25381 -42458
rect -25347 -42492 -25301 -42458
rect -25267 -42492 -25221 -42458
rect -25187 -42492 -25141 -42458
rect -25107 -42492 -25061 -42458
rect -25027 -42492 -24981 -42458
rect -24947 -42492 -24901 -42458
rect -24867 -42492 -24821 -42458
rect -24787 -42492 -24741 -42458
rect -24707 -42492 -24661 -42458
rect -24627 -42492 -24581 -42458
rect -24547 -42492 -24501 -42458
rect -24467 -42492 -24421 -42458
rect -24387 -42492 -24341 -42458
rect -24307 -42492 -24261 -42458
rect -24227 -42492 -24181 -42458
rect -24147 -42492 -24101 -42458
rect -24067 -42492 -24021 -42458
rect -23987 -42492 -23941 -42458
rect -23907 -42492 -23861 -42458
rect -23827 -42492 -23781 -42458
rect -23747 -42492 -23701 -42458
rect -23667 -42492 -23621 -42458
rect -23587 -42492 -23541 -42458
rect -23507 -42492 -23461 -42458
rect -23427 -42492 -23381 -42458
rect -23347 -42492 -23301 -42458
rect -23267 -42492 -23221 -42458
rect -23187 -42492 -23141 -42458
rect -23107 -42492 -23061 -42458
rect -23027 -42492 -22981 -42458
rect -22947 -42492 -22901 -42458
rect -22867 -42492 -22821 -42458
rect -22787 -42492 -22741 -42458
rect -22707 -42492 -22661 -42458
rect -22627 -42492 -22581 -42458
rect -22547 -42492 -22501 -42458
rect -22467 -42492 -22421 -42458
rect -22387 -42492 -22341 -42458
rect -22307 -42492 -22261 -42458
rect -22227 -42492 -22181 -42458
rect -22147 -42492 -22101 -42458
rect -22067 -42492 -22021 -42458
rect -21987 -42492 -21941 -42458
rect -21907 -42492 -21861 -42458
rect -21827 -42492 -21781 -42458
rect -21747 -42492 -21701 -42458
rect -21667 -42492 -21621 -42458
rect -21587 -42492 -21541 -42458
rect -21507 -42492 -21461 -42458
rect -21427 -42492 -21381 -42458
rect -21347 -42492 -21301 -42458
rect -21267 -42492 -21221 -42458
rect -21187 -42492 -21141 -42458
rect -21107 -42492 -21061 -42458
rect -21027 -42492 -20981 -42458
rect -20947 -42492 -20901 -42458
rect -20867 -42492 -20821 -42458
rect -20787 -42492 -20741 -42458
rect -20707 -42492 -20661 -42458
rect -20627 -42492 -20581 -42458
rect -20547 -42492 -20501 -42458
rect -20467 -42492 -20421 -42458
rect -20387 -42492 -20341 -42458
rect -20307 -42492 -20261 -42458
rect -20227 -42492 -20181 -42458
rect -20147 -42492 -20101 -42458
rect -20067 -42492 -20021 -42458
rect -19987 -42492 -19941 -42458
rect -19907 -42492 -19861 -42458
rect -19827 -42492 -19781 -42458
rect -19747 -42492 -19701 -42458
rect -19667 -42492 -19621 -42458
rect -19587 -42492 -19541 -42458
rect -19507 -42492 -19461 -42458
rect -19427 -42492 -19381 -42458
rect -19347 -42492 -19301 -42458
rect -19267 -42492 -19221 -42458
rect -19187 -42492 -19141 -42458
rect -19107 -42492 -19061 -42458
rect -19027 -42492 -18981 -42458
rect -18947 -42492 -18901 -42458
rect -18867 -42492 -18821 -42458
rect -18787 -42492 -18741 -42458
rect -18707 -42492 -18661 -42458
rect -18627 -42492 -18581 -42458
rect -18547 -42492 -18500 -42458
rect -18466 -42492 -18420 -42458
rect -18386 -42492 -18340 -42458
rect -18306 -42492 -18260 -42458
rect -18226 -42492 -18180 -42458
rect -18146 -42492 -18100 -42458
rect -18066 -42492 -18020 -42458
rect -17986 -42492 -17940 -42458
rect -17906 -42492 -17860 -42458
rect -17826 -42492 -17780 -42458
rect -17746 -42492 -17700 -42458
rect -17666 -42492 -17620 -42458
rect -17586 -42492 -17540 -42458
rect -17506 -42492 -17460 -42458
rect -17426 -42492 -17380 -42458
rect -17346 -42492 -17300 -42458
rect -17266 -42492 -17220 -42458
rect -17186 -42492 -17140 -42458
rect -17106 -42492 -17060 -42458
rect -17026 -42492 -16980 -42458
rect -16946 -42492 -16900 -42458
rect -16866 -42492 -16820 -42458
rect -16786 -42492 -16740 -42458
rect -16706 -42492 -16660 -42458
rect -16626 -42492 -16580 -42458
rect -16546 -42492 -16500 -42458
rect -16466 -42492 -16420 -42458
rect -16386 -42492 -16340 -42458
rect -16306 -42492 -16260 -42458
rect -16226 -42492 -16180 -42458
rect -16146 -42492 -16100 -42458
rect -16066 -42492 -16020 -42458
rect -15986 -42492 -15940 -42458
rect -15906 -42492 -15860 -42458
rect -15826 -42492 -15780 -42458
rect -15746 -42492 -15700 -42458
rect -15666 -42492 -15620 -42458
rect -15586 -42492 -15540 -42458
rect -15506 -42492 -15460 -42458
rect -15426 -42492 -15380 -42458
rect -15346 -42492 -15300 -42458
rect -15266 -42492 -15220 -42458
rect -15186 -42492 -15140 -42458
rect -15106 -42492 -15060 -42458
rect -15026 -42492 -14980 -42458
rect -14946 -42492 -14900 -42458
rect -14866 -42492 -14820 -42458
rect -14786 -42492 -14740 -42458
rect -14706 -42492 -14660 -42458
rect -14626 -42492 -14580 -42458
rect -14546 -42492 -14500 -42458
rect -14466 -42492 -14420 -42458
rect -14386 -42492 -14340 -42458
rect -14306 -42492 -14260 -42458
rect -14226 -42492 -14180 -42458
rect -14146 -42492 -14100 -42458
rect -14066 -42492 -14020 -42458
rect -13986 -42492 -13940 -42458
rect -13906 -42492 -13860 -42458
rect -13826 -42492 -13780 -42458
rect -13746 -42492 -13700 -42458
rect -13666 -42492 -13620 -42458
rect -13586 -42492 -13540 -42458
rect -13506 -42492 -13460 -42458
rect -13426 -42492 -13380 -42458
rect -13346 -42492 -13300 -42458
rect -13266 -42492 -13220 -42458
rect -13186 -42492 -13140 -42458
rect -13106 -42492 -13060 -42458
rect -13026 -42492 -12980 -42458
rect -12946 -42492 -12900 -42458
rect -12866 -42492 -12820 -42458
rect -12786 -42492 -12740 -42458
rect -12706 -42492 -12660 -42458
rect -12626 -42492 -12580 -42458
rect -12546 -42492 -12500 -42458
rect -12466 -42492 -12420 -42458
rect -12386 -42492 -12340 -42458
rect -12306 -42492 -12260 -42458
rect -12226 -42492 -12180 -42458
rect -12146 -42492 -12100 -42458
rect -12066 -42492 -12020 -42458
rect -11986 -42492 -11940 -42458
rect -11906 -42492 -11860 -42458
rect -11826 -42492 -11780 -42458
rect -11746 -42492 -11700 -42458
rect -11666 -42492 -11620 -42458
rect -11586 -42492 -11540 -42458
rect -11506 -42492 -11460 -42458
rect -11426 -42492 -11380 -42458
rect -11346 -42492 -11300 -42458
rect -11266 -42492 -11220 -42458
rect -11186 -42492 -11140 -42458
rect -11106 -42492 -11060 -42458
rect -11026 -42492 -10980 -42458
rect -10946 -42492 -10900 -42458
rect -10866 -42492 -10820 -42458
rect -10786 -42492 -10740 -42458
rect -10706 -42492 -10660 -42458
rect -10626 -42492 -10580 -42458
rect -10546 -42492 -10500 -42458
rect -10466 -42492 -10420 -42458
rect -10386 -42492 -10340 -42458
rect -10306 -42492 -10260 -42458
rect -10226 -42492 -10180 -42458
rect -10146 -42492 -10100 -42458
rect -10066 -42492 -10020 -42458
rect -9986 -42492 -9940 -42458
rect -9906 -42492 -9859 -42458
rect -9825 -42492 -9779 -42458
rect -9745 -42492 -9699 -42458
rect -9665 -42492 -9619 -42458
rect -9585 -42492 -9539 -42458
rect -9505 -42492 -9459 -42458
rect -9425 -42492 -9379 -42458
rect -9345 -42492 -9299 -42458
rect -9265 -42492 -9219 -42458
rect -9185 -42492 -9139 -42458
rect -9105 -42492 -9059 -42458
rect -9025 -42492 -8979 -42458
rect -8945 -42492 -8899 -42458
rect -8865 -42492 -8819 -42458
rect -8785 -42492 -8739 -42458
rect -8705 -42492 -8659 -42458
rect -8625 -42492 -8579 -42458
rect -8545 -42492 -8499 -42458
rect -8465 -42492 -8419 -42458
rect -8385 -42492 -8339 -42458
rect -8305 -42492 -8259 -42458
rect -8225 -42492 -8179 -42458
rect -8145 -42492 -8099 -42458
rect -8065 -42492 -8019 -42458
rect -7985 -42492 -7939 -42458
rect -7905 -42492 -7859 -42458
rect -7825 -42492 -7779 -42458
rect -7745 -42492 -7699 -42458
rect -7665 -42492 -7619 -42458
rect -7585 -42492 -7539 -42458
rect -7505 -42492 -7459 -42458
rect -7425 -42492 -7379 -42458
rect -7345 -42492 -7299 -42458
rect -7265 -42492 -7219 -42458
rect -7185 -42492 -7139 -42458
rect -7105 -42492 -7059 -42458
rect -7025 -42492 -6979 -42458
rect -6945 -42492 -6899 -42458
rect -6865 -42492 -6819 -42458
rect -6785 -42492 -6739 -42458
rect -6705 -42492 -6659 -42458
rect -6625 -42492 -6579 -42458
rect -6545 -42492 -6499 -42458
rect -6465 -42492 -6419 -42458
rect -6385 -42492 -6339 -42458
rect -6305 -42492 -6259 -42458
rect -6225 -42492 -6179 -42458
rect -6145 -42492 -6099 -42458
rect -6065 -42492 -6019 -42458
rect -5985 -42492 -5939 -42458
rect -5905 -42492 -5859 -42458
rect -5825 -42492 -5779 -42458
rect -5745 -42492 -5699 -42458
rect -5665 -42492 -5619 -42458
rect -5585 -42492 -5539 -42458
rect -5505 -42492 -5459 -42458
rect -5425 -42492 -5379 -42458
rect -5345 -42492 -5299 -42458
rect -5265 -42492 -5219 -42458
rect -5185 -42492 -5139 -42458
rect -5105 -42492 -5059 -42458
rect -5025 -42492 -4979 -42458
rect -4945 -42492 -4899 -42458
rect -4865 -42492 -4819 -42458
rect -4785 -42492 -4739 -42458
rect -4705 -42492 -4659 -42458
rect -4625 -42492 -4579 -42458
rect -4545 -42492 -4499 -42458
rect -4465 -42492 -4419 -42458
rect -4385 -42492 -4339 -42458
rect -4305 -42492 -4259 -42458
rect -4225 -42492 -4140 -42458
rect -4106 -42492 -4060 -42458
rect -4026 -42492 -3980 -42458
rect -3946 -42492 -3900 -42458
rect -3866 -42492 -3820 -42458
rect -3786 -42492 -3740 -42458
rect -3706 -42492 -3660 -42458
rect -3626 -42492 -3580 -42458
rect -3546 -42492 -3500 -42458
rect -3466 -42492 -3420 -42458
rect -3386 -42492 -3340 -42458
rect -3306 -42492 -3260 -42458
rect -3226 -42492 -3180 -42458
rect -3146 -42492 -3100 -42458
rect -3066 -42492 -3020 -42458
rect -2986 -42492 -2940 -42458
rect -2906 -42492 -2860 -42458
rect -2826 -42492 -2780 -42458
rect -2746 -42492 -2700 -42458
rect -2666 -42492 -2620 -42458
rect -2586 -42492 -2540 -42458
rect -2506 -42492 -2460 -42458
rect -2426 -42492 -2380 -42458
rect -2346 -42492 -2300 -42458
rect -2266 -42492 -2220 -42458
rect -2186 -42492 -2140 -42458
rect -2106 -42492 -2060 -42458
rect -2026 -42492 -1980 -42458
rect -1946 -42492 -1900 -42458
rect -1866 -42492 -1820 -42458
rect -1786 -42492 -1740 -42458
rect -1706 -42492 -1660 -42458
rect -1626 -42492 -1580 -42458
rect -1546 -42492 -1500 -42458
rect -1466 -42492 -1420 -42458
rect -1386 -42492 -1340 -42458
rect -1306 -42492 -1260 -42458
rect -1226 -42492 -1180 -42458
rect -1146 -42492 -1100 -42458
rect -1066 -42492 -1020 -42458
rect -986 -42492 -940 -42458
rect -906 -42492 -860 -42458
rect -826 -42492 -780 -42458
rect -746 -42492 -700 -42458
rect -666 -42492 -624 -42458
rect -44482 -42525 -624 -42492
rect -44482 -46942 -43986 -42525
rect -7849 -42710 -7799 -42696
rect -7849 -42744 -7841 -42710
rect -7807 -42744 -7799 -42710
rect -7849 -42782 -7799 -42744
rect -7849 -42816 -7841 -42782
rect -7807 -42816 -7799 -42782
rect -7849 -42854 -7799 -42816
rect -7849 -42888 -7841 -42854
rect -7807 -42888 -7799 -42854
rect -7849 -42926 -7799 -42888
rect -7849 -42960 -7841 -42926
rect -7807 -42960 -7799 -42926
rect -7849 -42998 -7799 -42960
rect -8155 -43041 -8075 -43030
rect -8155 -43100 -8145 -43041
rect -8086 -43100 -8075 -43041
rect -8155 -43110 -8075 -43100
rect -7849 -43032 -7841 -42998
rect -7807 -43032 -7799 -42998
rect -7849 -43070 -7799 -43032
rect -7849 -43104 -7841 -43070
rect -7807 -43104 -7799 -43070
rect -7849 -43117 -7799 -43104
rect -7531 -42710 -7163 -42696
rect -7531 -42744 -7523 -42710
rect -7489 -42744 -7205 -42710
rect -7171 -42744 -7163 -42710
rect -7531 -42782 -7163 -42744
rect -7531 -42816 -7523 -42782
rect -7489 -42816 -7205 -42782
rect -7171 -42816 -7163 -42782
rect -7531 -42854 -7163 -42816
rect -7531 -42888 -7523 -42854
rect -7489 -42888 -7205 -42854
rect -7171 -42888 -7163 -42854
rect -7531 -42926 -7163 -42888
rect -7531 -42960 -7523 -42926
rect -7489 -42960 -7205 -42926
rect -7171 -42960 -7163 -42926
rect -7531 -42976 -7163 -42960
rect -7531 -42998 -7481 -42976
rect -7531 -43032 -7523 -42998
rect -7489 -43032 -7481 -42998
rect -7531 -43070 -7481 -43032
rect -7531 -43104 -7523 -43070
rect -7489 -43104 -7481 -43070
rect -7531 -43117 -7481 -43104
rect -7213 -42998 -7163 -42976
rect -7213 -43032 -7205 -42998
rect -7171 -43032 -7163 -42998
rect -7213 -43070 -7163 -43032
rect -7213 -43104 -7205 -43070
rect -7171 -43104 -7163 -43070
rect -7213 -43117 -7163 -43104
rect -6895 -42710 -6845 -42696
rect -6895 -42744 -6887 -42710
rect -6853 -42744 -6845 -42710
rect -6895 -42782 -6845 -42744
rect -6895 -42816 -6887 -42782
rect -6853 -42816 -6845 -42782
rect -6895 -42854 -6845 -42816
rect -6895 -42888 -6887 -42854
rect -6853 -42888 -6845 -42854
rect -6895 -42926 -6845 -42888
rect -6895 -42960 -6887 -42926
rect -6853 -42960 -6845 -42926
rect -6895 -42998 -6845 -42960
rect -6895 -43032 -6887 -42998
rect -6853 -43032 -6845 -42998
rect -6895 -43070 -6845 -43032
rect -6895 -43104 -6887 -43070
rect -6853 -43104 -6845 -43070
rect -6895 -43117 -6845 -43104
rect -2304 -42711 -2254 -42697
rect -2304 -42745 -2296 -42711
rect -2262 -42745 -2254 -42711
rect -2304 -42783 -2254 -42745
rect -2304 -42817 -2296 -42783
rect -2262 -42817 -2254 -42783
rect -2304 -42855 -2254 -42817
rect -2304 -42889 -2296 -42855
rect -2262 -42889 -2254 -42855
rect -2304 -42927 -2254 -42889
rect -2304 -42961 -2296 -42927
rect -2262 -42961 -2254 -42927
rect -2304 -42999 -2254 -42961
rect -2304 -43033 -2296 -42999
rect -2262 -43033 -2254 -42999
rect -2304 -43071 -2254 -43033
rect -2304 -43105 -2296 -43071
rect -2262 -43105 -2254 -43071
rect -2304 -43118 -2254 -43105
rect -1986 -42711 -1618 -42697
rect -1986 -42745 -1978 -42711
rect -1944 -42745 -1660 -42711
rect -1626 -42745 -1618 -42711
rect -1986 -42783 -1618 -42745
rect -1986 -42817 -1978 -42783
rect -1944 -42817 -1660 -42783
rect -1626 -42817 -1618 -42783
rect -1986 -42855 -1618 -42817
rect -1986 -42889 -1978 -42855
rect -1944 -42889 -1660 -42855
rect -1626 -42889 -1618 -42855
rect -1986 -42927 -1618 -42889
rect -1986 -42961 -1978 -42927
rect -1944 -42961 -1660 -42927
rect -1626 -42961 -1618 -42927
rect -1986 -42977 -1618 -42961
rect -1986 -42999 -1936 -42977
rect -1986 -43033 -1978 -42999
rect -1944 -43033 -1936 -42999
rect -1986 -43071 -1936 -43033
rect -1986 -43105 -1978 -43071
rect -1944 -43105 -1936 -43071
rect -1986 -43118 -1936 -43105
rect -1668 -42999 -1618 -42977
rect -1668 -43033 -1660 -42999
rect -1626 -43033 -1618 -42999
rect -1668 -43071 -1618 -43033
rect -1668 -43105 -1660 -43071
rect -1626 -43105 -1618 -43071
rect -1668 -43118 -1618 -43105
rect -1350 -42711 -1300 -42697
rect -1350 -42745 -1342 -42711
rect -1308 -42745 -1300 -42711
rect -1350 -42783 -1300 -42745
rect -1350 -42817 -1342 -42783
rect -1308 -42817 -1300 -42783
rect -1350 -42855 -1300 -42817
rect -1350 -42889 -1342 -42855
rect -1308 -42889 -1300 -42855
rect -1350 -42927 -1300 -42889
rect -1350 -42961 -1342 -42927
rect -1308 -42961 -1300 -42927
rect -1350 -42999 -1300 -42961
rect -1350 -43033 -1342 -42999
rect -1308 -43033 -1300 -42999
rect -1350 -43071 -1300 -43033
rect -1350 -43105 -1342 -43071
rect -1308 -43105 -1300 -43071
rect -1350 -43118 -1300 -43105
rect -2549 -43150 -2469 -43138
rect -8788 -43224 -8528 -43181
rect -8788 -43278 -8746 -43224
rect -8691 -43278 -8625 -43224
rect -8570 -43278 -8528 -43224
rect -3203 -43223 -2943 -43180
rect -2549 -43206 -2536 -43150
rect -2483 -43206 -2469 -43150
rect -2549 -43218 -2469 -43206
rect -8788 -43343 -8528 -43278
rect -8788 -43397 -8745 -43343
rect -8690 -43344 -8528 -43343
rect -8690 -43397 -8625 -43344
rect -8788 -43398 -8625 -43397
rect -8570 -43398 -8528 -43344
rect -8788 -43441 -8528 -43398
rect -7849 -43279 -7799 -43265
rect -7849 -43313 -7841 -43279
rect -7807 -43313 -7799 -43279
rect -7849 -43351 -7799 -43313
rect -7849 -43385 -7841 -43351
rect -7807 -43385 -7799 -43351
rect -7849 -43406 -7799 -43385
rect -7531 -43279 -7481 -43265
rect -7531 -43313 -7523 -43279
rect -7489 -43313 -7481 -43279
rect -7531 -43351 -7481 -43313
rect -7531 -43385 -7523 -43351
rect -7489 -43385 -7481 -43351
rect -7531 -43406 -7481 -43385
rect -7849 -43423 -7481 -43406
rect -7849 -43457 -7841 -43423
rect -7807 -43457 -7523 -43423
rect -7489 -43457 -7481 -43423
rect -7849 -43495 -7481 -43457
rect -7849 -43529 -7841 -43495
rect -7807 -43529 -7523 -43495
rect -7489 -43529 -7481 -43495
rect -7849 -43567 -7481 -43529
rect -7849 -43601 -7841 -43567
rect -7807 -43601 -7523 -43567
rect -7489 -43601 -7481 -43567
rect -8701 -43640 -8621 -43630
rect -8701 -43700 -8691 -43640
rect -8631 -43700 -8621 -43640
rect -7849 -43639 -7481 -43601
rect -7849 -43673 -7841 -43639
rect -7807 -43673 -7523 -43639
rect -7489 -43673 -7481 -43639
rect -7849 -43686 -7481 -43673
rect -7213 -43279 -7163 -43265
rect -7213 -43313 -7205 -43279
rect -7171 -43313 -7163 -43279
rect -7213 -43351 -7163 -43313
rect -7213 -43385 -7205 -43351
rect -7171 -43385 -7163 -43351
rect -7213 -43406 -7163 -43385
rect -6895 -43279 -6845 -43265
rect -6895 -43313 -6887 -43279
rect -6853 -43313 -6845 -43279
rect -6895 -43351 -6845 -43313
rect -6895 -43385 -6887 -43351
rect -6853 -43385 -6845 -43351
rect -6895 -43406 -6845 -43385
rect -7213 -43423 -6845 -43406
rect -7213 -43457 -7205 -43423
rect -7171 -43457 -6887 -43423
rect -6853 -43457 -6845 -43423
rect -3203 -43277 -3160 -43223
rect -3106 -43277 -3040 -43223
rect -2986 -43277 -2943 -43223
rect -3203 -43342 -2943 -43277
rect -3203 -43343 -3041 -43342
rect -3203 -43397 -3161 -43343
rect -3107 -43396 -3041 -43343
rect -2987 -43396 -2943 -43342
rect -3107 -43397 -2943 -43396
rect -3203 -43440 -2943 -43397
rect -2304 -43280 -2254 -43266
rect -2304 -43314 -2296 -43280
rect -2262 -43314 -2254 -43280
rect -2304 -43352 -2254 -43314
rect -2304 -43386 -2296 -43352
rect -2262 -43386 -2254 -43352
rect -2304 -43407 -2254 -43386
rect -1986 -43280 -1936 -43266
rect -1986 -43314 -1978 -43280
rect -1944 -43314 -1936 -43280
rect -1986 -43352 -1936 -43314
rect -1986 -43386 -1978 -43352
rect -1944 -43386 -1936 -43352
rect -1986 -43407 -1936 -43386
rect -2304 -43424 -1936 -43407
rect -7213 -43495 -6845 -43457
rect -7213 -43529 -7205 -43495
rect -7171 -43529 -6887 -43495
rect -6853 -43529 -6845 -43495
rect -7213 -43567 -6845 -43529
rect -7213 -43601 -7205 -43567
rect -7171 -43601 -6887 -43567
rect -6853 -43601 -6845 -43567
rect -7213 -43639 -6845 -43601
rect -2304 -43458 -2296 -43424
rect -2262 -43458 -1978 -43424
rect -1944 -43458 -1936 -43424
rect -2304 -43496 -1936 -43458
rect -2304 -43530 -2296 -43496
rect -2262 -43530 -1978 -43496
rect -1944 -43530 -1936 -43496
rect -2304 -43568 -1936 -43530
rect -2304 -43602 -2296 -43568
rect -2262 -43602 -1978 -43568
rect -1944 -43602 -1936 -43568
rect -7213 -43673 -7205 -43639
rect -7171 -43673 -6887 -43639
rect -6853 -43673 -6845 -43639
rect -7213 -43686 -6845 -43673
rect -3116 -43639 -3036 -43629
rect -8701 -43710 -8621 -43700
rect -3116 -43699 -3106 -43639
rect -3046 -43699 -3036 -43639
rect -2304 -43640 -1936 -43602
rect -2304 -43674 -2296 -43640
rect -2262 -43674 -1978 -43640
rect -1944 -43674 -1936 -43640
rect -2304 -43687 -1936 -43674
rect -1668 -43280 -1618 -43266
rect -1668 -43314 -1660 -43280
rect -1626 -43314 -1618 -43280
rect -1668 -43352 -1618 -43314
rect -1668 -43386 -1660 -43352
rect -1626 -43386 -1618 -43352
rect -1668 -43407 -1618 -43386
rect -1350 -43280 -1300 -43266
rect -1350 -43314 -1342 -43280
rect -1308 -43314 -1300 -43280
rect -1350 -43352 -1300 -43314
rect -1350 -43386 -1342 -43352
rect -1308 -43386 -1300 -43352
rect -1350 -43407 -1300 -43386
rect -1668 -43424 -1300 -43407
rect -1668 -43458 -1660 -43424
rect -1626 -43458 -1342 -43424
rect -1308 -43458 -1300 -43424
rect -1668 -43496 -1300 -43458
rect -1668 -43530 -1660 -43496
rect -1626 -43530 -1342 -43496
rect -1308 -43530 -1300 -43496
rect -1668 -43568 -1300 -43530
rect -1668 -43602 -1660 -43568
rect -1626 -43602 -1342 -43568
rect -1308 -43602 -1300 -43568
rect -1668 -43640 -1300 -43602
rect -1668 -43674 -1660 -43640
rect -1626 -43674 -1342 -43640
rect -1308 -43674 -1300 -43640
rect -1668 -43687 -1300 -43674
rect -3116 -43709 -3036 -43699
rect -10430 -43753 -10170 -43710
rect -10430 -43809 -10388 -43753
rect -10333 -43757 -10267 -43753
rect -10333 -43807 -10268 -43757
rect -10212 -43807 -10170 -43753
rect -10336 -43809 -10268 -43807
rect -10216 -43809 -10170 -43807
rect -10430 -43813 -10170 -43809
rect -10430 -43829 -5254 -43813
rect -10430 -43863 -5304 -43829
rect -5270 -43863 -5254 -43829
rect -10430 -43872 -5254 -43863
rect -10430 -43877 -10387 -43872
rect -10332 -43873 -5254 -43872
rect -10332 -43877 -10267 -43873
rect -10430 -43929 -10388 -43877
rect -10332 -43926 -10268 -43877
rect -10212 -43879 -5254 -43873
rect -10336 -43929 -10268 -43926
rect -10212 -43927 -10170 -43879
rect -10216 -43929 -10170 -43927
rect -10430 -43970 -10170 -43929
rect -10430 -44989 -10170 -44948
rect -10430 -44991 -10387 -44989
rect -10335 -44991 -10267 -44989
rect -10215 -44991 -10170 -44989
rect -10430 -45047 -10388 -44991
rect -10333 -44995 -10267 -44991
rect -10333 -45045 -10268 -44995
rect -10212 -45043 -10170 -44991
rect -10212 -45045 -7860 -45043
rect -10336 -45047 -10268 -45045
rect -10216 -45047 -7860 -45045
rect -10430 -45059 -7860 -45047
rect -10430 -45093 -7910 -45059
rect -7876 -45093 -7860 -45059
rect -10430 -45109 -7860 -45093
rect -6859 -45081 -6599 -45040
rect -6859 -45083 -6816 -45081
rect -6764 -45083 -6696 -45081
rect -6644 -45083 -6599 -45081
rect -10430 -45115 -10387 -45109
rect -10335 -45110 -10267 -45109
rect -10332 -45115 -10267 -45110
rect -10215 -45111 -10170 -45109
rect -10430 -45167 -10388 -45115
rect -10332 -45164 -10268 -45115
rect -10336 -45167 -10268 -45164
rect -10212 -45165 -10170 -45111
rect -10216 -45167 -10170 -45165
rect -10430 -45208 -10170 -45167
rect -6859 -45139 -6817 -45083
rect -6762 -45087 -6696 -45083
rect -6762 -45137 -6697 -45087
rect -6641 -45137 -6599 -45083
rect -6764 -45139 -6697 -45137
rect -6859 -45140 -6816 -45139
rect -6764 -45140 -6696 -45139
rect -6644 -45140 -6599 -45137
rect -6859 -45201 -6599 -45140
rect -6859 -45207 -6816 -45201
rect -6764 -45202 -6696 -45201
rect -6761 -45207 -6696 -45202
rect -6644 -45203 -6599 -45201
rect -6859 -45259 -6817 -45207
rect -6761 -45256 -6697 -45207
rect -6641 -45243 -6599 -45203
rect -5232 -45080 -4972 -45043
rect -5232 -45081 -5074 -45080
rect -5232 -45146 -5195 -45081
rect -5129 -45145 -5074 -45081
rect -5008 -45145 -4972 -45080
rect -5129 -45146 -4972 -45145
rect -5232 -45200 -4972 -45146
rect -6764 -45259 -6697 -45256
rect -6641 -45257 -6598 -45243
rect -6859 -45260 -6816 -45259
rect -6764 -45260 -6696 -45259
rect -6644 -45260 -6598 -45257
rect -6859 -45300 -6598 -45260
rect -6858 -45303 -6598 -45300
rect -5232 -45265 -5194 -45200
rect -5128 -45265 -5074 -45200
rect -5008 -45265 -4972 -45200
rect -5232 -45303 -4972 -45265
rect -2292 -45403 -2086 -45402
rect -11742 -45436 -2086 -45403
rect -11742 -45470 -11699 -45436
rect -11665 -45470 -11619 -45436
rect -11585 -45470 -11539 -45436
rect -11505 -45470 -11459 -45436
rect -11425 -45470 -11379 -45436
rect -11345 -45470 -11299 -45436
rect -11265 -45470 -11219 -45436
rect -11185 -45470 -11139 -45436
rect -11105 -45470 -11059 -45436
rect -11025 -45470 -10979 -45436
rect -10945 -45470 -10899 -45436
rect -10865 -45470 -10819 -45436
rect -10785 -45470 -10739 -45436
rect -10705 -45470 -10659 -45436
rect -10625 -45470 -10579 -45436
rect -10545 -45470 -10499 -45436
rect -10465 -45470 -10419 -45436
rect -10385 -45470 -10339 -45436
rect -10305 -45470 -10259 -45436
rect -10225 -45470 -10179 -45436
rect -10145 -45470 -10099 -45436
rect -10065 -45470 -10019 -45436
rect -9985 -45470 -9939 -45436
rect -9905 -45470 -9859 -45436
rect -9825 -45470 -9779 -45436
rect -9745 -45470 -9699 -45436
rect -9665 -45470 -9619 -45436
rect -9585 -45470 -9539 -45436
rect -9505 -45470 -9459 -45436
rect -9425 -45470 -9379 -45436
rect -9345 -45470 -9299 -45436
rect -9265 -45470 -9219 -45436
rect -9185 -45470 -9139 -45436
rect -9105 -45470 -9059 -45436
rect -9025 -45470 -8979 -45436
rect -8945 -45470 -8899 -45436
rect -8865 -45470 -8819 -45436
rect -8785 -45470 -8739 -45436
rect -8705 -45470 -8659 -45436
rect -8625 -45470 -8579 -45436
rect -8545 -45470 -8499 -45436
rect -8465 -45470 -8419 -45436
rect -8385 -45470 -8339 -45436
rect -8305 -45470 -8259 -45436
rect -8225 -45470 -8179 -45436
rect -8145 -45470 -8099 -45436
rect -8065 -45470 -8019 -45436
rect -7985 -45470 -7939 -45436
rect -7905 -45470 -7859 -45436
rect -7825 -45470 -7779 -45436
rect -7745 -45470 -7699 -45436
rect -7665 -45470 -7619 -45436
rect -7585 -45470 -7539 -45436
rect -7505 -45470 -7459 -45436
rect -7425 -45470 -7379 -45436
rect -7345 -45470 -7299 -45436
rect -7265 -45470 -7219 -45436
rect -7185 -45470 -7139 -45436
rect -7105 -45470 -7059 -45436
rect -7025 -45470 -6979 -45436
rect -6945 -45470 -6899 -45436
rect -6865 -45470 -6819 -45436
rect -6785 -45470 -6739 -45436
rect -6705 -45470 -6659 -45436
rect -6625 -45470 -6579 -45436
rect -6545 -45470 -6499 -45436
rect -6465 -45470 -6419 -45436
rect -6385 -45470 -6339 -45436
rect -6305 -45470 -6259 -45436
rect -6225 -45470 -6179 -45436
rect -6145 -45470 -6099 -45436
rect -6065 -45470 -6019 -45436
rect -5985 -45470 -5939 -45436
rect -5905 -45470 -5859 -45436
rect -5825 -45470 -5779 -45436
rect -5745 -45470 -5699 -45436
rect -5665 -45470 -5619 -45436
rect -5585 -45470 -5539 -45436
rect -5505 -45470 -5459 -45436
rect -5425 -45470 -5379 -45436
rect -5345 -45470 -5299 -45436
rect -5265 -45470 -5219 -45436
rect -5185 -45470 -5139 -45436
rect -5105 -45470 -5059 -45436
rect -5025 -45470 -4979 -45436
rect -4945 -45470 -4899 -45436
rect -4865 -45470 -4819 -45436
rect -4785 -45470 -4739 -45436
rect -4705 -45470 -4659 -45436
rect -4625 -45470 -4579 -45436
rect -4545 -45470 -4499 -45436
rect -4465 -45470 -4419 -45436
rect -4385 -45470 -4339 -45436
rect -4305 -45470 -4259 -45436
rect -4225 -45470 -4179 -45436
rect -4145 -45470 -4099 -45436
rect -4065 -45470 -4019 -45436
rect -3985 -45470 -3939 -45436
rect -3905 -45470 -3859 -45436
rect -3825 -45470 -3779 -45436
rect -3745 -45470 -3699 -45436
rect -3665 -45470 -3619 -45436
rect -3585 -45470 -3539 -45436
rect -3505 -45470 -3459 -45436
rect -3425 -45470 -3379 -45436
rect -3345 -45470 -3299 -45436
rect -3265 -45470 -3219 -45436
rect -3185 -45470 -3139 -45436
rect -3105 -45470 -3059 -45436
rect -3025 -45470 -2979 -45436
rect -2945 -45470 -2899 -45436
rect -2865 -45470 -2819 -45436
rect -2785 -45470 -2739 -45436
rect -2705 -45470 -2659 -45436
rect -2625 -45470 -2579 -45436
rect -2545 -45470 -2499 -45436
rect -2465 -45470 -2419 -45436
rect -2385 -45470 -2339 -45436
rect -2305 -45470 -2259 -45436
rect -2225 -45470 -2179 -45436
rect -2145 -45470 -2086 -45436
rect -11742 -45503 -2086 -45470
rect -6855 -45942 -6595 -45905
rect -6855 -46007 -6817 -45942
rect -6751 -45943 -6595 -45942
rect -6751 -46007 -6698 -45943
rect -6855 -46008 -6698 -46007
rect -6632 -46008 -6595 -45943
rect -6855 -46063 -6595 -46008
rect -6855 -46064 -6698 -46063
rect -6855 -46129 -6818 -46064
rect -6752 -46128 -6698 -46064
rect -6632 -46128 -6595 -46063
rect -6752 -46129 -6595 -46128
rect -6855 -46165 -6595 -46129
rect -5229 -45943 -4969 -45905
rect -5229 -46008 -5192 -45943
rect -5126 -46008 -5073 -45943
rect -5007 -46008 -4969 -45943
rect -5229 -46062 -4969 -46008
rect -5229 -46063 -5072 -46062
rect -5229 -46128 -5192 -46063
rect -5126 -46127 -5072 -46063
rect -5006 -46127 -4969 -46062
rect -5126 -46128 -4969 -46127
rect -5229 -46165 -4969 -46128
rect -44482 -46975 -4170 -46942
rect -44482 -47009 -44435 -46975
rect -44401 -47009 -44355 -46975
rect -44321 -47009 -44275 -46975
rect -44241 -47009 -44195 -46975
rect -44161 -47009 -44115 -46975
rect -44081 -47009 -44035 -46975
rect -44001 -47009 -43955 -46975
rect -43921 -47009 -43875 -46975
rect -43841 -47009 -43795 -46975
rect -43761 -47009 -43715 -46975
rect -43681 -47009 -43635 -46975
rect -43601 -47009 -43555 -46975
rect -43521 -47009 -43475 -46975
rect -43441 -47009 -43395 -46975
rect -43361 -47009 -43315 -46975
rect -43281 -47009 -43235 -46975
rect -43201 -47009 -43155 -46975
rect -43121 -47009 -43075 -46975
rect -43041 -47009 -42995 -46975
rect -42961 -47009 -42915 -46975
rect -42881 -47009 -42835 -46975
rect -42801 -47009 -42755 -46975
rect -42721 -47009 -42675 -46975
rect -42641 -47009 -42595 -46975
rect -42561 -47009 -42515 -46975
rect -42481 -47009 -42435 -46975
rect -42401 -47009 -42355 -46975
rect -42321 -47009 -42275 -46975
rect -42241 -47009 -42195 -46975
rect -42161 -47009 -42115 -46975
rect -42081 -47009 -42035 -46975
rect -42001 -47009 -41955 -46975
rect -41921 -47009 -41875 -46975
rect -41841 -47009 -41795 -46975
rect -41761 -47009 -41715 -46975
rect -41681 -47009 -41635 -46975
rect -41601 -47009 -41555 -46975
rect -41521 -47009 -41475 -46975
rect -41441 -47009 -41395 -46975
rect -41361 -47009 -41315 -46975
rect -41281 -47009 -41235 -46975
rect -41201 -47009 -41155 -46975
rect -41121 -47009 -41075 -46975
rect -41041 -47009 -40995 -46975
rect -40961 -47009 -40915 -46975
rect -40881 -47009 -40835 -46975
rect -40801 -47009 -40755 -46975
rect -40721 -47009 -40675 -46975
rect -40641 -47009 -40595 -46975
rect -40561 -47009 -40515 -46975
rect -40481 -47009 -40435 -46975
rect -40401 -47009 -40355 -46975
rect -40321 -47009 -40275 -46975
rect -40241 -47009 -40195 -46975
rect -40161 -47009 -40115 -46975
rect -40081 -47009 -40035 -46975
rect -40001 -47009 -39955 -46975
rect -39921 -47009 -39875 -46975
rect -39841 -47009 -39795 -46975
rect -39761 -47009 -39715 -46975
rect -39681 -47009 -39635 -46975
rect -39601 -47009 -39555 -46975
rect -39521 -47009 -39475 -46975
rect -39441 -47009 -39395 -46975
rect -39361 -47009 -39315 -46975
rect -39281 -47009 -39235 -46975
rect -39201 -47009 -39155 -46975
rect -39121 -47009 -39075 -46975
rect -39041 -47009 -38995 -46975
rect -38961 -47009 -38915 -46975
rect -38881 -47009 -38835 -46975
rect -38801 -47009 -38755 -46975
rect -38721 -47009 -38675 -46975
rect -38641 -47009 -38595 -46975
rect -38561 -47009 -38515 -46975
rect -38481 -47009 -38435 -46975
rect -38401 -47009 -38355 -46975
rect -38321 -47009 -38275 -46975
rect -38241 -47009 -38195 -46975
rect -38161 -47009 -38115 -46975
rect -38081 -47009 -38035 -46975
rect -38001 -47009 -37955 -46975
rect -37921 -47009 -37875 -46975
rect -37841 -47009 -37795 -46975
rect -37761 -47009 -37715 -46975
rect -37681 -47009 -37635 -46975
rect -37601 -47009 -37555 -46975
rect -37521 -47009 -37475 -46975
rect -37441 -47009 -37395 -46975
rect -37361 -47009 -37315 -46975
rect -37281 -47009 -37235 -46975
rect -37201 -47009 -37155 -46975
rect -37121 -47009 -37075 -46975
rect -37041 -47009 -36995 -46975
rect -36961 -47009 -36915 -46975
rect -36881 -47009 -36835 -46975
rect -36801 -47009 -36755 -46975
rect -36721 -47009 -36675 -46975
rect -36641 -47009 -36595 -46975
rect -36561 -47009 -36515 -46975
rect -36481 -47009 -36435 -46975
rect -36401 -47009 -36355 -46975
rect -36321 -47009 -36275 -46975
rect -36241 -47009 -36195 -46975
rect -36161 -47009 -36115 -46975
rect -36081 -47009 -36035 -46975
rect -36001 -47009 -35955 -46975
rect -35921 -47009 -35875 -46975
rect -35841 -47009 -35795 -46975
rect -35761 -47009 -35715 -46975
rect -35681 -47009 -35635 -46975
rect -35601 -47009 -35555 -46975
rect -35521 -47009 -35475 -46975
rect -35441 -47009 -35395 -46975
rect -35361 -47009 -35315 -46975
rect -35281 -47009 -35235 -46975
rect -35201 -47009 -35155 -46975
rect -35121 -47009 -35075 -46975
rect -35041 -47009 -34995 -46975
rect -34961 -47009 -34915 -46975
rect -34881 -47009 -34835 -46975
rect -34801 -47009 -34755 -46975
rect -34721 -47009 -34675 -46975
rect -34641 -47009 -34595 -46975
rect -34561 -47009 -34515 -46975
rect -34481 -47009 -34435 -46975
rect -34401 -47009 -34355 -46975
rect -34321 -47009 -34275 -46975
rect -34241 -47009 -34195 -46975
rect -34161 -47009 -34115 -46975
rect -34081 -47009 -34035 -46975
rect -34001 -47009 -33955 -46975
rect -33921 -47009 -33875 -46975
rect -33841 -47009 -33795 -46975
rect -33761 -47009 -33715 -46975
rect -33681 -47009 -33635 -46975
rect -33601 -47009 -33555 -46975
rect -33521 -47009 -33475 -46975
rect -33441 -47009 -33395 -46975
rect -33361 -47009 -33315 -46975
rect -33281 -47009 -33235 -46975
rect -33201 -47009 -33155 -46975
rect -33121 -47009 -33075 -46975
rect -33041 -47009 -32995 -46975
rect -32961 -47009 -32915 -46975
rect -32881 -47009 -32835 -46975
rect -32801 -47009 -32755 -46975
rect -32721 -47009 -32675 -46975
rect -32641 -47009 -32595 -46975
rect -32561 -47009 -32515 -46975
rect -32481 -47009 -32435 -46975
rect -32401 -47009 -32355 -46975
rect -32321 -47009 -32275 -46975
rect -32241 -47009 -32195 -46975
rect -32161 -47009 -32115 -46975
rect -32081 -47009 -32035 -46975
rect -32001 -47009 -31955 -46975
rect -31921 -47009 -31875 -46975
rect -31841 -47009 -31795 -46975
rect -31761 -47009 -31715 -46975
rect -31681 -47009 -31635 -46975
rect -31601 -47009 -31555 -46975
rect -31521 -47009 -31475 -46975
rect -31441 -47009 -31395 -46975
rect -31361 -47009 -31315 -46975
rect -31281 -47009 -31235 -46975
rect -31201 -47009 -31155 -46975
rect -31121 -47009 -31075 -46975
rect -31041 -47009 -30995 -46975
rect -30961 -47009 -30915 -46975
rect -30881 -47009 -30835 -46975
rect -30801 -47009 -30755 -46975
rect -30721 -47009 -30675 -46975
rect -30641 -47009 -30595 -46975
rect -30561 -47009 -30515 -46975
rect -30481 -47009 -30435 -46975
rect -30401 -47009 -30355 -46975
rect -30321 -47009 -30275 -46975
rect -30241 -47009 -30195 -46975
rect -30161 -47009 -30115 -46975
rect -30081 -47009 -30035 -46975
rect -30001 -47009 -29955 -46975
rect -29921 -47009 -29875 -46975
rect -29841 -47009 -29795 -46975
rect -29761 -47009 -29715 -46975
rect -29681 -47009 -29635 -46975
rect -29601 -47009 -29555 -46975
rect -29521 -47009 -29475 -46975
rect -29441 -47009 -29395 -46975
rect -29361 -47009 -29315 -46975
rect -29281 -47009 -29235 -46975
rect -29201 -47009 -29155 -46975
rect -29121 -47009 -29075 -46975
rect -29041 -47009 -28995 -46975
rect -28961 -47009 -28915 -46975
rect -28881 -47009 -28835 -46975
rect -28801 -47009 -28755 -46975
rect -28721 -47009 -28675 -46975
rect -28641 -47009 -28595 -46975
rect -28561 -47009 -28514 -46975
rect -28480 -47009 -28434 -46975
rect -28400 -47009 -28354 -46975
rect -28320 -47009 -28274 -46975
rect -28240 -47009 -28194 -46975
rect -28160 -47009 -28114 -46975
rect -28080 -47009 -28034 -46975
rect -28000 -47009 -27954 -46975
rect -27920 -47009 -27874 -46975
rect -27840 -47009 -27794 -46975
rect -27760 -47009 -27714 -46975
rect -27680 -47009 -27634 -46975
rect -27600 -47009 -27554 -46975
rect -27520 -47009 -27474 -46975
rect -27440 -47009 -27394 -46975
rect -27360 -47009 -27314 -46975
rect -27280 -47009 -27234 -46975
rect -27200 -47009 -27154 -46975
rect -27120 -47009 -27074 -46975
rect -27040 -47009 -26994 -46975
rect -26960 -47009 -26914 -46975
rect -26880 -47009 -26834 -46975
rect -26800 -47009 -26754 -46975
rect -26720 -47009 -26674 -46975
rect -26640 -47009 -26594 -46975
rect -26560 -47009 -26514 -46975
rect -26480 -47009 -26434 -46975
rect -26400 -47009 -26354 -46975
rect -26320 -47009 -26274 -46975
rect -26240 -47009 -26194 -46975
rect -26160 -47009 -26114 -46975
rect -26080 -47009 -26034 -46975
rect -26000 -47009 -25954 -46975
rect -25920 -47009 -25874 -46975
rect -25840 -47009 -25794 -46975
rect -25760 -47009 -25714 -46975
rect -25680 -47009 -25634 -46975
rect -25600 -47009 -25554 -46975
rect -25520 -47009 -25474 -46975
rect -25440 -47009 -25394 -46975
rect -25360 -47009 -25314 -46975
rect -25280 -47009 -25234 -46975
rect -25200 -47009 -25154 -46975
rect -25120 -47009 -25074 -46975
rect -25040 -47009 -24994 -46975
rect -24960 -47009 -24914 -46975
rect -24880 -47009 -24834 -46975
rect -24800 -47009 -24754 -46975
rect -24720 -47009 -24674 -46975
rect -24640 -47009 -24594 -46975
rect -24560 -47009 -24514 -46975
rect -24480 -47009 -24434 -46975
rect -24400 -47009 -24354 -46975
rect -24320 -47009 -24274 -46975
rect -24240 -47009 -24194 -46975
rect -24160 -47009 -24114 -46975
rect -24080 -47009 -24034 -46975
rect -24000 -47009 -23954 -46975
rect -23920 -47009 -23874 -46975
rect -23840 -47009 -23794 -46975
rect -23760 -47009 -23714 -46975
rect -23680 -47009 -23634 -46975
rect -23600 -47009 -23554 -46975
rect -23520 -47009 -23474 -46975
rect -23440 -47009 -23394 -46975
rect -23360 -47009 -23314 -46975
rect -23280 -47009 -23234 -46975
rect -23200 -47009 -23154 -46975
rect -23120 -47009 -23074 -46975
rect -23040 -47009 -22994 -46975
rect -22960 -47009 -22914 -46975
rect -22880 -47009 -22834 -46975
rect -22800 -47009 -22754 -46975
rect -22720 -47009 -22674 -46975
rect -22640 -47009 -22594 -46975
rect -22560 -47009 -22514 -46975
rect -22480 -47009 -22434 -46975
rect -22400 -47009 -22354 -46975
rect -22320 -47009 -22274 -46975
rect -22240 -47009 -22194 -46975
rect -22160 -47009 -22114 -46975
rect -22080 -47009 -22034 -46975
rect -22000 -47009 -21954 -46975
rect -21920 -47009 -21874 -46975
rect -21840 -47009 -21794 -46975
rect -21760 -47009 -21714 -46975
rect -21680 -47009 -21634 -46975
rect -21600 -47009 -21554 -46975
rect -21520 -47009 -21474 -46975
rect -21440 -47009 -21394 -46975
rect -21360 -47009 -21314 -46975
rect -21280 -47009 -21234 -46975
rect -21200 -47009 -21154 -46975
rect -21120 -47009 -21074 -46975
rect -21040 -47009 -20994 -46975
rect -20960 -47009 -20914 -46975
rect -20880 -47009 -20834 -46975
rect -20800 -47009 -20754 -46975
rect -20720 -47009 -20674 -46975
rect -20640 -47009 -20594 -46975
rect -20560 -47009 -20514 -46975
rect -20480 -47009 -20434 -46975
rect -20400 -47009 -20354 -46975
rect -20320 -47009 -20274 -46975
rect -20240 -47009 -20194 -46975
rect -20160 -47009 -20114 -46975
rect -20080 -47009 -20034 -46975
rect -20000 -47009 -19954 -46975
rect -19920 -47009 -19874 -46975
rect -19840 -47009 -19794 -46975
rect -19760 -47009 -19714 -46975
rect -19680 -47009 -19634 -46975
rect -19600 -47009 -19554 -46975
rect -19520 -47009 -19474 -46975
rect -19440 -47009 -19394 -46975
rect -19360 -47009 -19314 -46975
rect -19280 -47009 -19234 -46975
rect -19200 -47009 -19154 -46975
rect -19120 -47009 -19074 -46975
rect -19040 -47009 -18994 -46975
rect -18960 -47009 -18914 -46975
rect -18880 -47009 -18834 -46975
rect -18800 -47009 -18754 -46975
rect -18720 -47009 -18674 -46975
rect -18640 -47009 -18594 -46975
rect -18560 -47009 -18514 -46975
rect -18480 -47009 -18434 -46975
rect -18400 -47009 -18354 -46975
rect -18320 -47009 -18274 -46975
rect -18240 -47009 -18194 -46975
rect -18160 -47009 -18114 -46975
rect -18080 -47009 -18034 -46975
rect -18000 -47009 -17954 -46975
rect -17920 -47009 -17874 -46975
rect -17840 -47009 -17794 -46975
rect -17760 -47009 -17714 -46975
rect -17680 -47009 -17634 -46975
rect -17600 -47009 -17554 -46975
rect -17520 -47009 -17474 -46975
rect -17440 -47009 -17394 -46975
rect -17360 -47009 -17314 -46975
rect -17280 -47009 -17234 -46975
rect -17200 -47009 -17154 -46975
rect -17120 -47009 -17074 -46975
rect -17040 -47009 -16994 -46975
rect -16960 -47009 -16914 -46975
rect -16880 -47009 -16834 -46975
rect -16800 -47009 -16754 -46975
rect -16720 -47009 -16674 -46975
rect -16640 -47009 -16594 -46975
rect -16560 -47009 -16514 -46975
rect -16480 -47009 -16434 -46975
rect -16400 -47009 -16354 -46975
rect -16320 -47009 -16274 -46975
rect -16240 -47009 -16194 -46975
rect -16160 -47009 -16114 -46975
rect -16080 -47009 -16034 -46975
rect -16000 -47009 -15954 -46975
rect -15920 -47009 -15874 -46975
rect -15840 -47009 -15794 -46975
rect -15760 -47009 -15714 -46975
rect -15680 -47009 -15634 -46975
rect -15600 -47009 -15553 -46975
rect -15519 -47009 -15473 -46975
rect -15439 -47009 -15393 -46975
rect -15359 -47009 -15313 -46975
rect -15279 -47009 -15233 -46975
rect -15199 -47009 -15153 -46975
rect -15119 -47009 -15073 -46975
rect -15039 -47009 -14993 -46975
rect -14959 -47009 -14913 -46975
rect -14879 -47009 -14833 -46975
rect -14799 -47009 -14753 -46975
rect -14719 -47009 -14673 -46975
rect -14639 -47009 -14593 -46975
rect -14559 -47009 -14513 -46975
rect -14479 -47009 -14433 -46975
rect -14399 -47009 -14353 -46975
rect -14319 -47009 -14273 -46975
rect -14239 -47009 -14193 -46975
rect -14159 -47009 -14113 -46975
rect -14079 -47009 -14033 -46975
rect -13999 -47009 -13953 -46975
rect -13919 -47009 -13873 -46975
rect -13839 -47009 -13793 -46975
rect -13759 -47009 -13713 -46975
rect -13679 -47009 -13633 -46975
rect -13599 -47009 -13553 -46975
rect -13519 -47009 -13473 -46975
rect -13439 -47009 -13393 -46975
rect -13359 -47009 -13313 -46975
rect -13279 -47009 -13233 -46975
rect -13199 -47009 -13153 -46975
rect -13119 -47009 -13073 -46975
rect -13039 -47009 -12993 -46975
rect -12959 -47009 -12913 -46975
rect -12879 -47009 -12833 -46975
rect -12799 -47009 -12753 -46975
rect -12719 -47009 -12673 -46975
rect -12639 -47009 -12593 -46975
rect -12559 -47009 -12513 -46975
rect -12479 -47009 -12433 -46975
rect -12399 -47009 -12353 -46975
rect -12319 -47009 -12273 -46975
rect -12239 -47009 -12193 -46975
rect -12159 -47009 -12113 -46975
rect -12079 -47009 -12033 -46975
rect -11999 -47009 -11953 -46975
rect -11919 -47009 -11873 -46975
rect -11839 -47009 -11793 -46975
rect -11759 -47009 -11713 -46975
rect -11679 -47009 -11633 -46975
rect -11599 -47009 -11553 -46975
rect -11519 -47009 -11473 -46975
rect -11439 -47009 -11393 -46975
rect -11359 -47009 -11313 -46975
rect -11279 -47009 -11233 -46975
rect -11199 -47009 -11153 -46975
rect -11119 -47009 -11073 -46975
rect -11039 -47009 -10993 -46975
rect -10959 -47009 -10913 -46975
rect -10879 -47009 -10833 -46975
rect -10799 -47009 -10753 -46975
rect -10719 -47009 -10673 -46975
rect -10639 -47009 -10593 -46975
rect -10559 -47009 -10513 -46975
rect -10479 -47009 -10433 -46975
rect -10399 -47009 -10353 -46975
rect -10319 -47009 -10273 -46975
rect -10239 -47009 -10193 -46975
rect -10159 -47009 -10113 -46975
rect -10079 -47009 -10033 -46975
rect -9999 -47009 -9953 -46975
rect -9919 -47009 -9873 -46975
rect -9839 -47009 -9793 -46975
rect -9759 -47009 -9713 -46975
rect -9679 -47009 -9633 -46975
rect -9599 -47009 -9553 -46975
rect -9519 -47009 -9473 -46975
rect -9439 -47009 -9393 -46975
rect -9359 -47009 -9313 -46975
rect -9279 -47009 -9233 -46975
rect -9199 -47009 -9153 -46975
rect -9119 -47009 -9073 -46975
rect -9039 -47009 -8993 -46975
rect -8959 -47009 -8913 -46975
rect -8879 -47009 -8833 -46975
rect -8799 -47009 -8753 -46975
rect -8719 -47009 -8673 -46975
rect -8639 -47009 -8593 -46975
rect -8559 -47009 -8513 -46975
rect -8479 -47009 -8433 -46975
rect -8399 -47009 -8353 -46975
rect -8319 -47009 -8273 -46975
rect -8239 -47009 -8193 -46975
rect -8159 -47009 -8113 -46975
rect -8079 -47009 -8033 -46975
rect -7999 -47009 -7953 -46975
rect -7919 -47009 -7873 -46975
rect -7839 -47009 -7793 -46975
rect -7759 -47009 -7713 -46975
rect -7679 -47009 -7633 -46975
rect -7599 -47009 -7553 -46975
rect -7519 -47009 -7473 -46975
rect -7439 -47009 -7393 -46975
rect -7359 -47009 -7313 -46975
rect -7279 -47009 -7233 -46975
rect -7199 -47009 -7153 -46975
rect -7119 -47009 -7073 -46975
rect -7039 -47009 -6993 -46975
rect -6959 -47009 -6913 -46975
rect -6879 -47009 -6841 -46975
rect -6807 -47009 -6769 -46975
rect -6735 -47009 -6697 -46975
rect -6663 -47009 -6625 -46975
rect -6591 -47009 -6553 -46975
rect -6519 -47009 -6481 -46975
rect -6447 -47009 -6409 -46975
rect -6375 -47009 -6337 -46975
rect -6303 -47009 -6265 -46975
rect -6231 -47009 -6193 -46975
rect -6159 -47009 -6121 -46975
rect -6087 -47009 -6049 -46975
rect -6015 -47009 -5977 -46975
rect -5943 -47009 -5905 -46975
rect -5871 -47009 -5833 -46975
rect -5799 -47009 -5761 -46975
rect -5727 -47009 -5689 -46975
rect -5655 -47009 -5617 -46975
rect -5583 -47009 -5545 -46975
rect -5511 -47009 -5473 -46975
rect -5439 -47009 -5401 -46975
rect -5367 -47009 -5329 -46975
rect -5295 -47009 -5257 -46975
rect -5223 -47009 -5185 -46975
rect -5151 -47009 -5113 -46975
rect -5079 -47009 -5041 -46975
rect -5007 -47009 -4969 -46975
rect -4935 -47009 -4889 -46975
rect -4855 -47009 -4809 -46975
rect -4775 -47009 -4729 -46975
rect -4695 -47009 -4649 -46975
rect -4615 -47009 -4569 -46975
rect -4535 -47009 -4489 -46975
rect -4455 -47009 -4409 -46975
rect -4375 -47009 -4329 -46975
rect -4295 -47009 -4249 -46975
rect -4215 -47009 -4170 -46975
rect -44482 -47042 -4170 -47009
rect -4956 -47111 -4876 -47096
rect -4956 -47163 -4942 -47111
rect -4890 -47163 -4876 -47111
rect -4956 -47176 -4876 -47163
rect -6801 -47801 -6721 -47792
rect -6801 -47835 -6778 -47801
rect -6744 -47835 -6721 -47801
rect -6801 -47844 -6721 -47835
rect -6801 -48213 -6721 -48204
rect -6801 -48247 -6778 -48213
rect -6744 -48247 -6721 -48213
rect -6801 -48256 -6721 -48247
rect -2292 -48312 -2086 -45503
rect -10124 -48345 -2086 -48312
rect -10124 -48379 -10087 -48345
rect -10053 -48379 -10007 -48345
rect -9973 -48379 -9927 -48345
rect -9893 -48379 -9847 -48345
rect -9813 -48379 -9767 -48345
rect -9733 -48379 -9687 -48345
rect -9653 -48379 -9607 -48345
rect -9573 -48379 -9527 -48345
rect -9493 -48379 -9447 -48345
rect -9413 -48379 -9367 -48345
rect -9333 -48379 -9287 -48345
rect -9253 -48379 -9207 -48345
rect -9173 -48379 -9127 -48345
rect -9093 -48379 -9047 -48345
rect -9013 -48379 -8967 -48345
rect -8933 -48379 -8887 -48345
rect -8853 -48379 -8807 -48345
rect -8773 -48379 -8727 -48345
rect -8693 -48379 -8647 -48345
rect -8613 -48379 -8567 -48345
rect -8533 -48379 -8487 -48345
rect -8453 -48379 -8407 -48345
rect -8373 -48379 -8327 -48345
rect -8293 -48379 -8247 -48345
rect -8213 -48379 -8167 -48345
rect -8133 -48379 -8087 -48345
rect -8053 -48379 -8007 -48345
rect -7973 -48379 -7927 -48345
rect -7893 -48379 -7847 -48345
rect -7813 -48379 -7767 -48345
rect -7733 -48379 -7687 -48345
rect -7653 -48379 -7607 -48345
rect -7573 -48379 -7527 -48345
rect -7493 -48379 -7447 -48345
rect -7413 -48379 -7367 -48345
rect -7333 -48379 -7287 -48345
rect -7253 -48379 -7207 -48345
rect -7173 -48379 -7127 -48345
rect -7093 -48379 -7047 -48345
rect -7013 -48379 -6967 -48345
rect -6933 -48379 -6887 -48345
rect -6853 -48379 -6807 -48345
rect -6773 -48379 -6727 -48345
rect -6693 -48379 -6647 -48345
rect -6613 -48379 -6567 -48345
rect -6533 -48379 -6487 -48345
rect -6453 -48379 -6407 -48345
rect -6373 -48379 -6327 -48345
rect -6293 -48379 -6247 -48345
rect -6213 -48379 -6167 -48345
rect -6133 -48379 -6087 -48345
rect -6053 -48379 -6007 -48345
rect -5973 -48379 -5927 -48345
rect -5893 -48379 -5847 -48345
rect -5813 -48379 -5767 -48345
rect -5733 -48379 -5687 -48345
rect -5653 -48379 -5607 -48345
rect -5573 -48379 -5527 -48345
rect -5493 -48379 -5447 -48345
rect -5413 -48379 -5367 -48345
rect -5333 -48379 -5287 -48345
rect -5253 -48379 -5207 -48345
rect -5173 -48379 -5127 -48345
rect -5093 -48379 -5047 -48345
rect -5013 -48379 -4967 -48345
rect -4933 -48379 -4887 -48345
rect -4853 -48379 -4807 -48345
rect -4773 -48379 -4727 -48345
rect -4693 -48379 -4647 -48345
rect -4613 -48379 -4567 -48345
rect -4533 -48379 -4487 -48345
rect -4453 -48379 -4407 -48345
rect -4373 -48379 -4327 -48345
rect -4293 -48379 -4247 -48345
rect -4213 -48379 -4167 -48345
rect -4133 -48379 -4087 -48345
rect -4053 -48379 -4007 -48345
rect -3973 -48379 -3927 -48345
rect -3893 -48379 -3847 -48345
rect -3813 -48379 -3767 -48345
rect -3733 -48379 -3687 -48345
rect -3653 -48379 -3607 -48345
rect -3573 -48379 -3527 -48345
rect -3493 -48379 -3447 -48345
rect -3413 -48379 -3367 -48345
rect -3333 -48379 -3287 -48345
rect -3253 -48379 -3207 -48345
rect -3173 -48379 -3127 -48345
rect -3093 -48379 -3047 -48345
rect -3013 -48379 -2967 -48345
rect -2933 -48379 -2887 -48345
rect -2853 -48379 -2807 -48345
rect -2773 -48379 -2727 -48345
rect -2693 -48379 -2647 -48345
rect -2613 -48379 -2567 -48345
rect -2533 -48379 -2487 -48345
rect -2453 -48379 -2407 -48345
rect -2373 -48379 -2327 -48345
rect -2293 -48379 -2247 -48345
rect -2213 -48379 -2167 -48345
rect -2133 -48379 -2086 -48345
rect -10124 -48412 -2086 -48379
rect -2292 -48414 -2086 -48412
<< via1 >>
rect -27240 -34719 -27188 -34710
rect -27240 -34753 -27231 -34719
rect -27231 -34753 -27197 -34719
rect -27197 -34753 -27188 -34719
rect -27240 -34762 -27188 -34753
rect -27120 -34719 -27068 -34710
rect -27120 -34753 -27111 -34719
rect -27111 -34753 -27077 -34719
rect -27077 -34753 -27068 -34719
rect -27120 -34762 -27068 -34753
rect -27240 -34839 -27188 -34830
rect -27240 -34873 -27231 -34839
rect -27231 -34873 -27197 -34839
rect -27197 -34873 -27188 -34839
rect -27240 -34882 -27188 -34873
rect -27120 -34839 -27068 -34830
rect -27120 -34873 -27111 -34839
rect -27111 -34873 -27077 -34839
rect -27077 -34873 -27068 -34839
rect -27120 -34882 -27068 -34873
rect 12095 -34720 12147 -34711
rect 12095 -34754 12104 -34720
rect 12104 -34754 12138 -34720
rect 12138 -34754 12147 -34720
rect 12095 -34763 12147 -34754
rect 12215 -34720 12267 -34711
rect 12215 -34754 12224 -34720
rect 12224 -34754 12258 -34720
rect 12258 -34754 12267 -34720
rect 12215 -34763 12267 -34754
rect 12095 -34840 12147 -34831
rect 12095 -34874 12104 -34840
rect 12104 -34874 12138 -34840
rect 12138 -34874 12147 -34840
rect 12095 -34883 12147 -34874
rect 12215 -34840 12267 -34831
rect 12215 -34874 12224 -34840
rect 12224 -34874 12258 -34840
rect 12258 -34874 12267 -34840
rect 12215 -34883 12267 -34874
rect -8145 -43053 -8086 -43041
rect -8145 -43087 -8132 -43053
rect -8132 -43087 -8098 -43053
rect -8098 -43087 -8086 -43053
rect -8145 -43100 -8086 -43087
rect -8746 -43234 -8691 -43224
rect -8746 -43268 -8735 -43234
rect -8735 -43268 -8701 -43234
rect -8701 -43268 -8691 -43234
rect -8746 -43278 -8691 -43268
rect -8625 -43234 -8570 -43224
rect -8625 -43268 -8615 -43234
rect -8615 -43268 -8581 -43234
rect -8581 -43268 -8570 -43234
rect -8625 -43278 -8570 -43268
rect -2536 -43161 -2483 -43150
rect -2536 -43195 -2526 -43161
rect -2526 -43195 -2492 -43161
rect -2492 -43195 -2483 -43161
rect -2536 -43206 -2483 -43195
rect -8745 -43354 -8690 -43343
rect -8745 -43388 -8735 -43354
rect -8735 -43388 -8701 -43354
rect -8701 -43388 -8690 -43354
rect -8745 -43397 -8690 -43388
rect -8625 -43354 -8570 -43344
rect -8625 -43388 -8615 -43354
rect -8615 -43388 -8581 -43354
rect -8581 -43388 -8570 -43354
rect -8625 -43398 -8570 -43388
rect -8691 -43650 -8631 -43640
rect -8691 -43690 -8681 -43650
rect -8681 -43690 -8641 -43650
rect -8641 -43690 -8631 -43650
rect -8691 -43700 -8631 -43690
rect -3160 -43233 -3106 -43223
rect -3160 -43267 -3150 -43233
rect -3150 -43267 -3116 -43233
rect -3116 -43267 -3106 -43233
rect -3160 -43277 -3106 -43267
rect -3040 -43233 -2986 -43223
rect -3040 -43267 -3030 -43233
rect -3030 -43267 -2996 -43233
rect -2996 -43267 -2986 -43233
rect -3040 -43277 -2986 -43267
rect -3161 -43353 -3107 -43343
rect -3161 -43387 -3150 -43353
rect -3150 -43387 -3116 -43353
rect -3116 -43387 -3107 -43353
rect -3161 -43397 -3107 -43387
rect -3041 -43353 -2987 -43342
rect -3041 -43387 -3030 -43353
rect -3030 -43387 -2996 -43353
rect -2996 -43387 -2987 -43353
rect -3041 -43396 -2987 -43387
rect -3106 -43649 -3046 -43639
rect -3106 -43689 -3096 -43649
rect -3096 -43689 -3056 -43649
rect -3056 -43689 -3046 -43649
rect -3106 -43699 -3046 -43689
rect -10388 -43763 -10333 -43753
rect -10267 -43757 -10212 -43753
rect -10388 -43766 -10377 -43763
rect -10377 -43766 -10343 -43763
rect -10388 -43800 -10379 -43766
rect -10379 -43797 -10343 -43766
rect -10343 -43797 -10333 -43763
rect -10379 -43800 -10345 -43797
rect -10345 -43800 -10333 -43797
rect -10388 -43807 -10333 -43800
rect -10268 -43763 -10212 -43757
rect -10268 -43766 -10257 -43763
rect -10257 -43766 -10223 -43763
rect -10268 -43800 -10259 -43766
rect -10259 -43797 -10223 -43766
rect -10223 -43797 -10212 -43763
rect -10259 -43800 -10225 -43797
rect -10225 -43800 -10212 -43797
rect -10268 -43807 -10212 -43800
rect -10388 -43809 -10336 -43807
rect -10268 -43809 -10216 -43807
rect -10387 -43877 -10332 -43872
rect -10267 -43877 -10212 -43873
rect -10388 -43883 -10332 -43877
rect -10388 -43886 -10377 -43883
rect -10377 -43886 -10343 -43883
rect -10388 -43920 -10379 -43886
rect -10379 -43917 -10343 -43886
rect -10343 -43917 -10332 -43883
rect -10379 -43920 -10345 -43917
rect -10345 -43920 -10332 -43917
rect -10388 -43926 -10332 -43920
rect -10268 -43883 -10212 -43877
rect -10268 -43886 -10257 -43883
rect -10257 -43886 -10223 -43883
rect -10268 -43920 -10259 -43886
rect -10259 -43917 -10223 -43886
rect -10223 -43917 -10212 -43883
rect -10259 -43920 -10225 -43917
rect -10225 -43920 -10212 -43917
rect -10388 -43929 -10336 -43926
rect -10268 -43927 -10212 -43920
rect -10268 -43929 -10216 -43927
rect -10387 -44991 -10335 -44989
rect -10267 -44991 -10215 -44989
rect -10388 -44998 -10333 -44991
rect -10267 -44995 -10212 -44991
rect -10388 -45004 -10378 -44998
rect -10378 -45001 -10344 -44998
rect -10344 -45001 -10333 -44998
rect -10378 -45004 -10343 -45001
rect -10388 -45038 -10379 -45004
rect -10379 -45035 -10343 -45004
rect -10343 -45035 -10333 -45001
rect -10379 -45038 -10345 -45035
rect -10345 -45038 -10333 -45035
rect -10388 -45045 -10333 -45038
rect -10268 -44998 -10212 -44995
rect -10268 -45004 -10258 -44998
rect -10258 -45001 -10224 -44998
rect -10224 -45001 -10212 -44998
rect -10258 -45004 -10223 -45001
rect -10268 -45038 -10259 -45004
rect -10259 -45035 -10223 -45004
rect -10223 -45035 -10212 -45001
rect -10259 -45038 -10225 -45035
rect -10225 -45038 -10212 -45035
rect -10268 -45045 -10212 -45038
rect -10388 -45047 -10336 -45045
rect -10268 -45047 -10216 -45045
rect -6816 -45083 -6764 -45081
rect -6696 -45083 -6644 -45081
rect -10387 -45110 -10335 -45109
rect -10387 -45115 -10332 -45110
rect -10267 -45111 -10215 -45109
rect -10267 -45115 -10212 -45111
rect -10388 -45118 -10332 -45115
rect -10388 -45124 -10378 -45118
rect -10378 -45121 -10344 -45118
rect -10344 -45121 -10332 -45118
rect -10378 -45124 -10343 -45121
rect -10388 -45158 -10379 -45124
rect -10379 -45155 -10343 -45124
rect -10343 -45155 -10332 -45121
rect -10379 -45158 -10345 -45155
rect -10345 -45158 -10332 -45155
rect -10388 -45164 -10332 -45158
rect -10268 -45118 -10212 -45115
rect -10268 -45124 -10258 -45118
rect -10258 -45121 -10224 -45118
rect -10224 -45121 -10212 -45118
rect -10258 -45124 -10223 -45121
rect -10268 -45158 -10259 -45124
rect -10259 -45155 -10223 -45124
rect -10223 -45155 -10212 -45121
rect -10259 -45158 -10225 -45155
rect -10225 -45158 -10212 -45155
rect -10388 -45167 -10336 -45164
rect -10268 -45165 -10212 -45158
rect -10268 -45167 -10216 -45165
rect -6817 -45090 -6762 -45083
rect -6696 -45087 -6641 -45083
rect -6817 -45096 -6807 -45090
rect -6807 -45093 -6773 -45090
rect -6773 -45093 -6762 -45090
rect -6807 -45096 -6772 -45093
rect -6817 -45130 -6808 -45096
rect -6808 -45127 -6772 -45096
rect -6772 -45127 -6762 -45093
rect -6808 -45130 -6773 -45127
rect -6817 -45131 -6807 -45130
rect -6807 -45131 -6773 -45130
rect -6773 -45131 -6762 -45127
rect -6817 -45137 -6762 -45131
rect -6697 -45090 -6641 -45087
rect -6697 -45096 -6687 -45090
rect -6687 -45093 -6653 -45090
rect -6653 -45093 -6641 -45090
rect -6687 -45096 -6652 -45093
rect -6697 -45130 -6688 -45096
rect -6688 -45127 -6652 -45096
rect -6652 -45127 -6641 -45093
rect -6688 -45130 -6653 -45127
rect -6697 -45131 -6687 -45130
rect -6687 -45131 -6653 -45130
rect -6653 -45131 -6641 -45127
rect -6697 -45137 -6641 -45131
rect -6817 -45139 -6764 -45137
rect -6697 -45139 -6644 -45137
rect -6816 -45140 -6764 -45139
rect -6696 -45140 -6644 -45139
rect -6816 -45202 -6764 -45201
rect -6816 -45207 -6761 -45202
rect -6696 -45203 -6644 -45201
rect -6696 -45207 -6641 -45203
rect -6817 -45210 -6761 -45207
rect -6817 -45216 -6807 -45210
rect -6807 -45213 -6773 -45210
rect -6773 -45213 -6761 -45210
rect -6807 -45216 -6772 -45213
rect -6817 -45250 -6808 -45216
rect -6808 -45247 -6772 -45216
rect -6772 -45247 -6761 -45213
rect -6808 -45250 -6773 -45247
rect -6817 -45251 -6807 -45250
rect -6807 -45251 -6773 -45250
rect -6773 -45251 -6761 -45247
rect -6817 -45256 -6761 -45251
rect -6697 -45210 -6641 -45207
rect -6697 -45216 -6687 -45210
rect -6687 -45213 -6653 -45210
rect -6653 -45213 -6641 -45210
rect -6687 -45216 -6652 -45213
rect -6697 -45250 -6688 -45216
rect -6688 -45247 -6652 -45216
rect -6652 -45247 -6641 -45213
rect -5195 -45096 -5129 -45081
rect -5195 -45130 -5179 -45096
rect -5179 -45130 -5145 -45096
rect -5145 -45130 -5129 -45096
rect -5195 -45146 -5129 -45130
rect -5074 -45096 -5008 -45080
rect -5074 -45130 -5059 -45096
rect -5059 -45130 -5025 -45096
rect -5025 -45130 -5008 -45096
rect -5074 -45145 -5008 -45130
rect -6688 -45250 -6653 -45247
rect -6697 -45251 -6687 -45250
rect -6687 -45251 -6653 -45250
rect -6653 -45251 -6641 -45247
rect -6817 -45259 -6764 -45256
rect -6697 -45257 -6641 -45251
rect -6697 -45259 -6644 -45257
rect -6816 -45260 -6764 -45259
rect -6696 -45260 -6644 -45259
rect -5194 -45216 -5128 -45200
rect -5194 -45250 -5179 -45216
rect -5179 -45250 -5145 -45216
rect -5145 -45250 -5128 -45216
rect -5194 -45265 -5128 -45250
rect -5074 -45216 -5008 -45200
rect -5074 -45250 -5059 -45216
rect -5059 -45250 -5025 -45216
rect -5025 -45250 -5008 -45216
rect -5074 -45265 -5008 -45250
rect -6817 -45958 -6751 -45942
rect -6817 -45992 -6802 -45958
rect -6802 -45992 -6768 -45958
rect -6768 -45992 -6751 -45958
rect -6817 -46007 -6751 -45992
rect -6698 -45958 -6632 -45943
rect -6698 -45992 -6682 -45958
rect -6682 -45992 -6648 -45958
rect -6648 -45992 -6632 -45958
rect -6698 -46008 -6632 -45992
rect -6818 -46078 -6752 -46064
rect -6818 -46112 -6802 -46078
rect -6802 -46112 -6768 -46078
rect -6768 -46112 -6752 -46078
rect -6818 -46129 -6752 -46112
rect -6698 -46078 -6632 -46063
rect -6698 -46112 -6682 -46078
rect -6682 -46112 -6648 -46078
rect -6648 -46112 -6632 -46078
rect -6698 -46128 -6632 -46112
rect -5192 -45958 -5126 -45943
rect -5192 -45992 -5176 -45958
rect -5176 -45992 -5142 -45958
rect -5142 -45992 -5126 -45958
rect -5192 -46008 -5126 -45992
rect -5073 -45958 -5007 -45943
rect -5073 -45992 -5056 -45958
rect -5056 -45992 -5022 -45958
rect -5022 -45992 -5007 -45958
rect -5073 -46008 -5007 -45992
rect -5192 -46078 -5126 -46063
rect -5192 -46112 -5176 -46078
rect -5176 -46112 -5142 -46078
rect -5142 -46112 -5126 -46078
rect -5192 -46128 -5126 -46112
rect -5072 -46078 -5006 -46062
rect -5072 -46112 -5056 -46078
rect -5056 -46112 -5022 -46078
rect -5022 -46112 -5006 -46078
rect -5072 -46127 -5006 -46112
rect -4942 -47119 -4890 -47111
rect -4942 -47153 -4933 -47119
rect -4933 -47153 -4899 -47119
rect -4899 -47153 -4890 -47119
rect -4942 -47163 -4890 -47153
<< metal2 >>
rect -27284 -34700 -27024 -34666
rect -27284 -34770 -27250 -34700
rect -27180 -34770 -27130 -34700
rect -27060 -34770 -27024 -34700
rect -27284 -34820 -27024 -34770
rect -27284 -34890 -27250 -34820
rect -27180 -34890 -27130 -34820
rect -27060 -34890 -27024 -34820
rect -27284 -34926 -27024 -34890
rect 12051 -34700 12311 -34667
rect 12051 -34770 12090 -34700
rect 12160 -34770 12210 -34700
rect 12280 -34770 12311 -34700
rect 12051 -34820 12311 -34770
rect 12051 -34890 12090 -34820
rect 12160 -34890 12210 -34820
rect 12280 -34890 12311 -34820
rect 12051 -34927 12311 -34890
rect -8155 -43041 -8075 -43030
rect -8155 -43100 -8145 -43041
rect -8086 -43053 -8075 -43041
rect -8086 -43087 -584 -43053
rect -8086 -43100 -8075 -43087
rect -8155 -43110 -8075 -43100
rect -2549 -43150 -2469 -43138
rect -8788 -43220 -8528 -43181
rect -8788 -43290 -8750 -43220
rect -8680 -43290 -8630 -43220
rect -8560 -43290 -8528 -43220
rect -8788 -43340 -8528 -43290
rect -8788 -43410 -8750 -43340
rect -8680 -43410 -8630 -43340
rect -8560 -43410 -8528 -43340
rect -8788 -43441 -8528 -43410
rect -3203 -43220 -2943 -43180
rect -2549 -43206 -2536 -43150
rect -2483 -43161 -2469 -43150
rect -2483 -43195 -584 -43161
rect -2483 -43206 -2469 -43195
rect -2549 -43218 -2469 -43206
rect -3203 -43290 -3170 -43220
rect -3100 -43290 -3050 -43220
rect -2980 -43290 -2943 -43220
rect -3203 -43340 -2943 -43290
rect -3203 -43410 -3170 -43340
rect -3100 -43342 -3040 -43340
rect -3100 -43396 -3041 -43342
rect -3100 -43410 -3040 -43396
rect -2970 -43410 -2943 -43340
rect -3203 -43440 -2943 -43410
rect -8721 -43621 -8601 -43610
rect -10430 -43750 -10170 -43710
rect -8721 -43721 -8711 -43621
rect -8610 -43721 -8601 -43621
rect -8721 -43730 -8601 -43721
rect -3136 -43631 -3016 -43609
rect -3136 -43710 -3113 -43631
rect -3040 -43710 -3016 -43631
rect -3136 -43729 -3016 -43710
rect -10430 -43820 -10400 -43750
rect -10330 -43820 -10280 -43750
rect -10210 -43820 -10170 -43750
rect -10430 -43870 -10170 -43820
rect -10430 -43940 -10400 -43870
rect -10330 -43940 -10270 -43870
rect -10200 -43940 -10170 -43870
rect -10430 -43970 -10170 -43940
rect -10430 -44980 -10170 -44948
rect -10430 -45050 -10400 -44980
rect -10330 -45050 -10270 -44980
rect -10200 -45050 -10170 -44980
rect -10430 -45100 -10170 -45050
rect -10430 -45170 -10400 -45100
rect -10330 -45170 -10270 -45100
rect -10200 -45170 -10170 -45100
rect -10430 -45208 -10170 -45170
rect -6859 -45080 -6599 -45040
rect -6859 -45150 -6830 -45080
rect -6760 -45150 -6710 -45080
rect -6640 -45150 -6599 -45080
rect -6859 -45200 -6599 -45150
rect -6859 -45270 -6830 -45200
rect -6760 -45270 -6700 -45200
rect -6630 -45243 -6599 -45200
rect -5232 -45080 -4972 -45043
rect -5232 -45150 -5200 -45080
rect -5130 -45081 -5080 -45080
rect -5129 -45146 -5080 -45081
rect -5008 -45145 -4972 -45080
rect -5130 -45150 -5080 -45146
rect -5010 -45150 -4972 -45145
rect -5232 -45200 -4972 -45150
rect -6630 -45270 -6598 -45243
rect -6859 -45300 -6598 -45270
rect -6858 -45303 -6598 -45300
rect -5232 -45270 -5200 -45200
rect -5128 -45265 -5074 -45200
rect -5130 -45270 -5070 -45265
rect -5000 -45270 -4972 -45200
rect -5232 -45303 -4972 -45270
rect -6855 -45940 -4876 -45905
rect -6855 -46010 -6820 -45940
rect -6750 -46010 -6700 -45940
rect -6630 -45943 -5190 -45940
rect -5120 -45943 -5070 -45940
rect -6630 -46008 -5192 -45943
rect -5120 -46008 -5073 -45943
rect -6630 -46010 -5190 -46008
rect -5120 -46010 -5070 -46008
rect -5000 -46010 -4876 -45940
rect -6855 -46060 -4876 -46010
rect -6855 -46130 -6820 -46060
rect -6750 -46130 -6700 -46060
rect -6630 -46063 -5190 -46060
rect -5120 -46062 -5070 -46060
rect -6630 -46128 -5192 -46063
rect -5120 -46127 -5072 -46062
rect -6630 -46130 -5190 -46128
rect -5120 -46130 -5070 -46127
rect -5000 -46130 -4876 -46060
rect -6855 -46165 -4876 -46130
rect -4956 -47111 -4876 -46165
rect -4956 -47163 -4942 -47111
rect -4890 -47163 -4876 -47111
rect -4956 -47176 -4876 -47163
<< via2 >>
rect -27250 -34710 -27180 -34700
rect -27250 -34762 -27240 -34710
rect -27240 -34762 -27188 -34710
rect -27188 -34762 -27180 -34710
rect -27250 -34770 -27180 -34762
rect -27130 -34710 -27060 -34700
rect -27130 -34762 -27120 -34710
rect -27120 -34762 -27068 -34710
rect -27068 -34762 -27060 -34710
rect -27130 -34770 -27060 -34762
rect -27250 -34830 -27180 -34820
rect -27250 -34882 -27240 -34830
rect -27240 -34882 -27188 -34830
rect -27188 -34882 -27180 -34830
rect -27250 -34890 -27180 -34882
rect -27130 -34830 -27060 -34820
rect -27130 -34882 -27120 -34830
rect -27120 -34882 -27068 -34830
rect -27068 -34882 -27060 -34830
rect -27130 -34890 -27060 -34882
rect 12090 -34711 12160 -34700
rect 12090 -34763 12095 -34711
rect 12095 -34763 12147 -34711
rect 12147 -34763 12160 -34711
rect 12090 -34770 12160 -34763
rect 12210 -34711 12280 -34700
rect 12210 -34763 12215 -34711
rect 12215 -34763 12267 -34711
rect 12267 -34763 12280 -34711
rect 12210 -34770 12280 -34763
rect 12090 -34831 12160 -34820
rect 12090 -34883 12095 -34831
rect 12095 -34883 12147 -34831
rect 12147 -34883 12160 -34831
rect 12090 -34890 12160 -34883
rect 12210 -34831 12280 -34820
rect 12210 -34883 12215 -34831
rect 12215 -34883 12267 -34831
rect 12267 -34883 12280 -34831
rect 12210 -34890 12280 -34883
rect -8750 -43224 -8680 -43220
rect -8750 -43278 -8746 -43224
rect -8746 -43278 -8691 -43224
rect -8691 -43278 -8680 -43224
rect -8750 -43290 -8680 -43278
rect -8630 -43224 -8560 -43220
rect -8630 -43278 -8625 -43224
rect -8625 -43278 -8570 -43224
rect -8570 -43278 -8560 -43224
rect -8630 -43290 -8560 -43278
rect -8750 -43343 -8680 -43340
rect -8750 -43397 -8745 -43343
rect -8745 -43397 -8690 -43343
rect -8690 -43397 -8680 -43343
rect -8750 -43410 -8680 -43397
rect -8630 -43344 -8560 -43340
rect -8630 -43398 -8625 -43344
rect -8625 -43398 -8570 -43344
rect -8570 -43398 -8560 -43344
rect -8630 -43410 -8560 -43398
rect -3170 -43223 -3100 -43220
rect -3170 -43277 -3160 -43223
rect -3160 -43277 -3106 -43223
rect -3106 -43277 -3100 -43223
rect -3170 -43290 -3100 -43277
rect -3050 -43223 -2980 -43220
rect -3050 -43277 -3040 -43223
rect -3040 -43277 -2986 -43223
rect -2986 -43277 -2980 -43223
rect -3050 -43290 -2980 -43277
rect -3170 -43343 -3100 -43340
rect -3040 -43342 -2970 -43340
rect -3170 -43397 -3161 -43343
rect -3161 -43397 -3107 -43343
rect -3107 -43397 -3100 -43343
rect -3040 -43396 -2987 -43342
rect -2987 -43396 -2970 -43342
rect -3170 -43410 -3100 -43397
rect -3040 -43410 -2970 -43396
rect -8711 -43640 -8610 -43621
rect -8711 -43700 -8691 -43640
rect -8691 -43700 -8631 -43640
rect -8631 -43700 -8610 -43640
rect -8711 -43721 -8610 -43700
rect -3113 -43639 -3040 -43631
rect -3113 -43699 -3106 -43639
rect -3106 -43699 -3046 -43639
rect -3046 -43699 -3040 -43639
rect -3113 -43710 -3040 -43699
rect -10400 -43753 -10330 -43750
rect -10400 -43809 -10388 -43753
rect -10388 -43807 -10333 -43753
rect -10333 -43807 -10330 -43753
rect -10388 -43809 -10336 -43807
rect -10336 -43809 -10330 -43807
rect -10400 -43820 -10330 -43809
rect -10280 -43753 -10210 -43750
rect -10280 -43757 -10267 -43753
rect -10267 -43757 -10212 -43753
rect -10280 -43809 -10268 -43757
rect -10268 -43807 -10212 -43757
rect -10212 -43807 -10210 -43753
rect -10268 -43809 -10216 -43807
rect -10216 -43809 -10210 -43807
rect -10280 -43820 -10210 -43809
rect -10400 -43872 -10330 -43870
rect -10400 -43877 -10387 -43872
rect -10387 -43877 -10332 -43872
rect -10400 -43929 -10388 -43877
rect -10388 -43926 -10332 -43877
rect -10332 -43926 -10330 -43872
rect -10388 -43929 -10336 -43926
rect -10336 -43929 -10330 -43926
rect -10400 -43940 -10330 -43929
rect -10270 -43873 -10200 -43870
rect -10270 -43877 -10267 -43873
rect -10267 -43877 -10212 -43873
rect -10270 -43929 -10268 -43877
rect -10268 -43927 -10212 -43877
rect -10212 -43927 -10200 -43873
rect -10268 -43929 -10216 -43927
rect -10216 -43929 -10200 -43927
rect -10270 -43940 -10200 -43929
rect -10400 -44989 -10330 -44980
rect -10400 -44991 -10387 -44989
rect -10387 -44991 -10335 -44989
rect -10335 -44991 -10330 -44989
rect -10400 -45047 -10388 -44991
rect -10388 -45045 -10333 -44991
rect -10333 -45045 -10330 -44991
rect -10388 -45047 -10336 -45045
rect -10336 -45047 -10330 -45045
rect -10400 -45050 -10330 -45047
rect -10270 -44989 -10200 -44980
rect -10270 -44995 -10267 -44989
rect -10267 -44991 -10215 -44989
rect -10215 -44991 -10200 -44989
rect -10267 -44995 -10212 -44991
rect -10270 -45047 -10268 -44995
rect -10268 -45045 -10212 -44995
rect -10212 -45045 -10200 -44991
rect -10268 -45047 -10216 -45045
rect -10216 -45047 -10200 -45045
rect -10270 -45050 -10200 -45047
rect -10400 -45109 -10330 -45100
rect -10400 -45115 -10387 -45109
rect -10387 -45110 -10335 -45109
rect -10335 -45110 -10330 -45109
rect -10387 -45115 -10332 -45110
rect -10400 -45167 -10388 -45115
rect -10388 -45164 -10332 -45115
rect -10332 -45164 -10330 -45110
rect -10388 -45167 -10336 -45164
rect -10336 -45167 -10330 -45164
rect -10400 -45170 -10330 -45167
rect -10270 -45109 -10200 -45100
rect -10270 -45115 -10267 -45109
rect -10267 -45111 -10215 -45109
rect -10215 -45111 -10200 -45109
rect -10267 -45115 -10212 -45111
rect -10270 -45167 -10268 -45115
rect -10268 -45165 -10212 -45115
rect -10212 -45165 -10200 -45111
rect -10268 -45167 -10216 -45165
rect -10216 -45167 -10200 -45165
rect -10270 -45170 -10200 -45167
rect -6830 -45081 -6760 -45080
rect -6830 -45083 -6816 -45081
rect -6816 -45083 -6764 -45081
rect -6764 -45083 -6760 -45081
rect -6830 -45139 -6817 -45083
rect -6817 -45137 -6762 -45083
rect -6762 -45137 -6760 -45083
rect -6817 -45139 -6764 -45137
rect -6830 -45140 -6816 -45139
rect -6816 -45140 -6764 -45139
rect -6764 -45140 -6760 -45137
rect -6830 -45150 -6760 -45140
rect -6710 -45081 -6640 -45080
rect -6710 -45087 -6696 -45081
rect -6696 -45083 -6644 -45081
rect -6644 -45083 -6640 -45081
rect -6696 -45087 -6641 -45083
rect -6710 -45139 -6697 -45087
rect -6697 -45137 -6641 -45087
rect -6641 -45137 -6640 -45083
rect -6697 -45139 -6644 -45137
rect -6710 -45140 -6696 -45139
rect -6696 -45140 -6644 -45139
rect -6644 -45140 -6640 -45137
rect -6710 -45150 -6640 -45140
rect -6830 -45201 -6760 -45200
rect -6830 -45207 -6816 -45201
rect -6816 -45202 -6764 -45201
rect -6764 -45202 -6760 -45201
rect -6816 -45207 -6761 -45202
rect -6830 -45259 -6817 -45207
rect -6817 -45256 -6761 -45207
rect -6761 -45256 -6760 -45202
rect -6817 -45259 -6764 -45256
rect -6830 -45260 -6816 -45259
rect -6816 -45260 -6764 -45259
rect -6764 -45260 -6760 -45256
rect -6830 -45270 -6760 -45260
rect -6700 -45201 -6630 -45200
rect -6700 -45207 -6696 -45201
rect -6696 -45203 -6644 -45201
rect -6644 -45203 -6630 -45201
rect -6696 -45207 -6641 -45203
rect -6700 -45259 -6697 -45207
rect -6697 -45257 -6641 -45207
rect -6641 -45257 -6630 -45203
rect -5200 -45081 -5130 -45080
rect -5200 -45146 -5195 -45081
rect -5195 -45146 -5130 -45081
rect -5080 -45145 -5074 -45080
rect -5074 -45145 -5010 -45080
rect -5200 -45150 -5130 -45146
rect -5080 -45150 -5010 -45145
rect -6697 -45259 -6644 -45257
rect -6700 -45260 -6696 -45259
rect -6696 -45260 -6644 -45259
rect -6644 -45260 -6630 -45257
rect -6700 -45270 -6630 -45260
rect -5200 -45265 -5194 -45200
rect -5194 -45265 -5130 -45200
rect -5070 -45265 -5008 -45200
rect -5008 -45265 -5000 -45200
rect -5200 -45270 -5130 -45265
rect -5070 -45270 -5000 -45265
rect -6820 -45942 -6750 -45940
rect -6820 -46007 -6817 -45942
rect -6817 -46007 -6751 -45942
rect -6751 -46007 -6750 -45942
rect -6820 -46010 -6750 -46007
rect -6700 -45943 -6630 -45940
rect -5190 -45943 -5120 -45940
rect -5070 -45943 -5000 -45940
rect -6700 -46008 -6698 -45943
rect -6698 -46008 -6632 -45943
rect -6632 -46008 -6630 -45943
rect -5190 -46008 -5126 -45943
rect -5126 -46008 -5120 -45943
rect -5070 -46008 -5007 -45943
rect -5007 -46008 -5000 -45943
rect -6700 -46010 -6630 -46008
rect -5190 -46010 -5120 -46008
rect -5070 -46010 -5000 -46008
rect -6820 -46064 -6750 -46060
rect -6820 -46129 -6818 -46064
rect -6818 -46129 -6752 -46064
rect -6752 -46129 -6750 -46064
rect -6820 -46130 -6750 -46129
rect -6700 -46063 -6630 -46060
rect -5190 -46063 -5120 -46060
rect -5070 -46062 -5000 -46060
rect -6700 -46128 -6698 -46063
rect -6698 -46128 -6632 -46063
rect -6632 -46128 -6630 -46063
rect -5190 -46128 -5126 -46063
rect -5126 -46128 -5120 -46063
rect -5070 -46127 -5006 -46062
rect -5006 -46127 -5000 -46062
rect -6700 -46130 -6630 -46128
rect -5190 -46130 -5120 -46128
rect -5070 -46130 -5000 -46127
<< metal3 >>
rect -27284 -34700 -27024 -34666
rect -27284 -34770 -27250 -34700
rect -27180 -34770 -27130 -34700
rect -27060 -34770 -27024 -34700
rect -27284 -34820 -27024 -34770
rect -27284 -34890 -27250 -34820
rect -27180 -34890 -27130 -34820
rect -27060 -34890 -27024 -34820
rect -27284 -34926 -27024 -34890
rect 12051 -34700 12311 -34667
rect 12051 -34705 12090 -34700
rect 12160 -34705 12210 -34700
rect 12051 -34769 12089 -34705
rect 12160 -34769 12209 -34705
rect 12051 -34770 12090 -34769
rect 12160 -34770 12210 -34769
rect 12280 -34770 12311 -34700
rect 12051 -34820 12311 -34770
rect 12051 -34825 12090 -34820
rect 12160 -34825 12210 -34820
rect 12051 -34889 12089 -34825
rect 12160 -34889 12209 -34825
rect 12051 -34890 12090 -34889
rect 12160 -34890 12210 -34889
rect 12280 -34890 12311 -34820
rect 12051 -34927 12311 -34890
rect -8788 -43219 -8528 -43181
rect -8788 -43290 -8750 -43219
rect -8686 -43220 -8630 -43219
rect -8566 -43220 -8528 -43219
rect -8680 -43290 -8630 -43220
rect -8560 -43290 -8528 -43220
rect -8788 -43339 -8528 -43290
rect -8788 -43410 -8750 -43339
rect -8686 -43340 -8630 -43339
rect -8566 -43340 -8528 -43339
rect -8680 -43410 -8630 -43340
rect -8560 -43410 -8528 -43340
rect -8788 -43441 -8528 -43410
rect -3203 -43218 -2943 -43180
rect -3203 -43220 -3165 -43218
rect -3101 -43220 -3045 -43218
rect -2981 -43220 -2943 -43218
rect -3203 -43290 -3170 -43220
rect -3100 -43290 -3050 -43220
rect -2980 -43290 -2943 -43220
rect -3203 -43338 -2943 -43290
rect -3203 -43340 -3165 -43338
rect -3101 -43340 -3045 -43338
rect -2981 -43340 -2943 -43338
rect -3203 -43410 -3170 -43340
rect -3100 -43402 -3045 -43340
rect -3100 -43410 -3040 -43402
rect -2970 -43410 -2943 -43340
rect -3203 -43440 -2943 -43410
rect -8688 -43473 -8628 -43441
rect -8688 -43590 -8628 -43533
rect -3107 -43472 -3047 -43440
rect -3107 -43589 -3047 -43532
rect -8741 -43621 -8581 -43590
rect -10430 -43748 -10170 -43710
rect -10430 -43750 -10392 -43748
rect -10328 -43750 -10272 -43748
rect -10430 -43820 -10400 -43750
rect -10328 -43812 -10280 -43750
rect -10330 -43820 -10280 -43812
rect -10208 -43812 -10170 -43748
rect -8741 -43721 -8711 -43621
rect -8610 -43721 -8581 -43621
rect -8741 -43750 -8581 -43721
rect -3156 -43631 -2996 -43589
rect -3156 -43710 -3113 -43631
rect -3040 -43710 -2996 -43631
rect -3156 -43749 -2996 -43710
rect -10210 -43820 -10170 -43812
rect -10430 -43868 -10170 -43820
rect -10430 -43870 -10392 -43868
rect -10430 -43940 -10400 -43870
rect -10328 -43871 -10272 -43868
rect -10208 -43870 -10170 -43868
rect -10328 -43932 -10274 -43871
rect -10330 -43935 -10274 -43932
rect -10330 -43940 -10270 -43935
rect -10200 -43940 -10170 -43870
rect -10430 -43970 -10170 -43940
rect -10430 -44980 -10170 -44948
rect -10430 -45050 -10400 -44980
rect -10330 -44983 -10270 -44980
rect -10329 -44986 -10273 -44983
rect -10328 -44989 -10273 -44986
rect -10328 -45050 -10274 -44989
rect -10200 -45050 -10170 -44980
rect -10430 -45053 -10394 -45050
rect -10330 -45053 -10274 -45050
rect -10210 -45053 -10170 -45050
rect -10430 -45100 -10170 -45053
rect -10430 -45170 -10400 -45100
rect -10330 -45103 -10270 -45100
rect -10329 -45106 -10273 -45103
rect -10328 -45109 -10273 -45106
rect -10328 -45170 -10274 -45109
rect -10200 -45170 -10170 -45100
rect -10430 -45173 -10394 -45170
rect -10330 -45173 -10274 -45170
rect -10210 -45173 -10170 -45170
rect -10430 -45208 -10170 -45173
rect -6859 -45075 -6599 -45040
rect -6859 -45080 -6822 -45075
rect -6758 -45078 -6702 -45075
rect -6638 -45078 -6599 -45075
rect -6757 -45080 -6702 -45078
rect -6859 -45150 -6830 -45080
rect -6757 -45142 -6710 -45080
rect -6758 -45146 -6710 -45142
rect -6637 -45142 -6599 -45078
rect -6638 -45146 -6599 -45142
rect -6760 -45150 -6710 -45146
rect -6640 -45150 -6599 -45146
rect -6859 -45195 -6599 -45150
rect -6859 -45200 -6822 -45195
rect -6758 -45198 -6702 -45195
rect -6638 -45198 -6599 -45195
rect -6859 -45270 -6830 -45200
rect -6757 -45201 -6702 -45198
rect -6637 -45200 -6599 -45198
rect -6757 -45262 -6703 -45201
rect -6758 -45265 -6703 -45262
rect -6758 -45266 -6702 -45265
rect -6760 -45270 -6700 -45266
rect -6630 -45270 -6599 -45200
rect -6859 -45300 -6599 -45270
rect -5232 -45080 -4972 -45043
rect -5232 -45150 -5200 -45080
rect -5130 -45150 -5080 -45080
rect -5010 -45150 -4972 -45080
rect -5232 -45200 -4972 -45150
rect -5232 -45270 -5200 -45200
rect -5130 -45201 -5070 -45200
rect -5130 -45265 -5074 -45201
rect -5130 -45270 -5070 -45265
rect -5000 -45270 -4972 -45200
rect -6858 -45303 -6598 -45300
rect -5232 -45303 -4972 -45270
rect -6855 -45940 -6595 -45303
rect -6855 -46010 -6820 -45940
rect -6750 -46010 -6700 -45940
rect -6630 -46010 -6595 -45940
rect -6855 -46060 -6595 -46010
rect -6855 -46130 -6820 -46060
rect -6750 -46130 -6700 -46060
rect -6630 -46130 -6595 -46060
rect -6855 -46165 -6595 -46130
rect -5229 -45940 -4969 -45303
rect -5229 -45943 -5190 -45940
rect -5120 -45943 -5070 -45940
rect -5229 -46007 -5191 -45943
rect -5120 -46007 -5071 -45943
rect -5229 -46010 -5190 -46007
rect -5120 -46010 -5070 -46007
rect -5000 -46010 -4969 -45940
rect -5229 -46060 -4969 -46010
rect -5229 -46063 -5190 -46060
rect -5120 -46063 -5070 -46060
rect -5229 -46127 -5191 -46063
rect -5120 -46127 -5071 -46063
rect -5229 -46130 -5190 -46127
rect -5120 -46130 -5070 -46127
rect -5000 -46130 -4969 -46060
rect -5229 -46165 -4969 -46130
<< rmetal3 >>
rect -8688 -43533 -8628 -43473
rect -3107 -43532 -3047 -43472
<< via3 >>
rect -27246 -34768 -27182 -34704
rect -27126 -34768 -27062 -34704
rect -27246 -34888 -27182 -34824
rect -27126 -34888 -27062 -34824
rect 12089 -34769 12090 -34705
rect 12090 -34769 12153 -34705
rect 12209 -34769 12210 -34705
rect 12210 -34769 12273 -34705
rect 12089 -34889 12090 -34825
rect 12090 -34889 12153 -34825
rect 12209 -34889 12210 -34825
rect 12210 -34889 12273 -34825
rect -8750 -43220 -8686 -43219
rect -8630 -43220 -8566 -43219
rect -8750 -43283 -8686 -43220
rect -8630 -43283 -8566 -43220
rect -8750 -43340 -8686 -43339
rect -8630 -43340 -8566 -43339
rect -8750 -43403 -8686 -43340
rect -8630 -43403 -8566 -43340
rect -3165 -43220 -3101 -43218
rect -3045 -43220 -2981 -43218
rect -3165 -43282 -3101 -43220
rect -3045 -43282 -2981 -43220
rect -3165 -43340 -3101 -43338
rect -3045 -43340 -2981 -43338
rect -3165 -43402 -3101 -43340
rect -3045 -43402 -3040 -43340
rect -3040 -43402 -2981 -43340
rect -10392 -43750 -10328 -43748
rect -10272 -43750 -10208 -43748
rect -10392 -43751 -10330 -43750
rect -10394 -43815 -10330 -43751
rect -10330 -43812 -10328 -43750
rect -10272 -43751 -10210 -43750
rect -10274 -43815 -10210 -43751
rect -10210 -43812 -10208 -43750
rect -10392 -43870 -10328 -43868
rect -10392 -43871 -10330 -43870
rect -10394 -43935 -10330 -43871
rect -10330 -43932 -10328 -43870
rect -10272 -43870 -10208 -43868
rect -10272 -43871 -10270 -43870
rect -10274 -43935 -10270 -43871
rect -10270 -43932 -10208 -43870
rect -10270 -43935 -10210 -43932
rect -10393 -44989 -10330 -44983
rect -10330 -44986 -10329 -44983
rect -10394 -45050 -10330 -44989
rect -10330 -45050 -10328 -44986
rect -10273 -44989 -10270 -44983
rect -10270 -44986 -10209 -44983
rect -10274 -45050 -10270 -44989
rect -10270 -45050 -10208 -44986
rect -10394 -45053 -10330 -45050
rect -10274 -45053 -10210 -45050
rect -10393 -45109 -10330 -45103
rect -10330 -45106 -10329 -45103
rect -10394 -45170 -10330 -45109
rect -10330 -45170 -10328 -45106
rect -10273 -45109 -10270 -45103
rect -10270 -45106 -10209 -45103
rect -10274 -45170 -10270 -45109
rect -10270 -45170 -10208 -45106
rect -10394 -45173 -10330 -45170
rect -10274 -45173 -10210 -45170
rect -6822 -45078 -6758 -45075
rect -6702 -45078 -6638 -45075
rect -6822 -45080 -6757 -45078
rect -6702 -45080 -6637 -45078
rect -6822 -45081 -6760 -45080
rect -6823 -45145 -6760 -45081
rect -6760 -45142 -6757 -45080
rect -6702 -45081 -6640 -45080
rect -6822 -45146 -6760 -45145
rect -6760 -45146 -6758 -45142
rect -6703 -45145 -6640 -45081
rect -6640 -45142 -6637 -45080
rect -6702 -45146 -6640 -45145
rect -6640 -45146 -6638 -45142
rect -6822 -45198 -6758 -45195
rect -6702 -45198 -6638 -45195
rect -6822 -45200 -6757 -45198
rect -6822 -45201 -6760 -45200
rect -6823 -45265 -6760 -45201
rect -6760 -45262 -6757 -45200
rect -6702 -45200 -6637 -45198
rect -6702 -45201 -6700 -45200
rect -6822 -45266 -6760 -45265
rect -6760 -45266 -6758 -45262
rect -6703 -45265 -6700 -45201
rect -6700 -45262 -6637 -45200
rect -6702 -45266 -6700 -45265
rect -6700 -45266 -6638 -45262
rect -5194 -45145 -5130 -45081
rect -5074 -45145 -5010 -45081
rect -5194 -45265 -5130 -45201
rect -5074 -45265 -5070 -45201
rect -5070 -45265 -5010 -45201
rect -6817 -46007 -6753 -45943
rect -6697 -46007 -6633 -45943
rect -6817 -46127 -6753 -46063
rect -6697 -46127 -6633 -46063
rect -5191 -46007 -5190 -45943
rect -5190 -46007 -5127 -45943
rect -5071 -46007 -5070 -45943
rect -5070 -46007 -5007 -45943
rect -5191 -46127 -5190 -46063
rect -5190 -46127 -5127 -46063
rect -5071 -46127 -5070 -46063
rect -5070 -46127 -5007 -46063
<< metal4 >>
rect -44425 -5525 -9225 -5325
rect -44425 -39725 -44225 -5525
rect -43825 -6125 -9825 -5925
rect -43825 -39125 -43625 -6125
rect -43225 -6725 -10425 -6525
rect -43225 -38525 -43025 -6725
rect -42625 -7325 -11025 -7125
rect -42625 -37925 -42425 -7325
rect -42025 -7925 -11625 -7725
rect -42025 -37325 -41825 -7925
rect -41425 -8525 -12225 -8325
rect -41425 -36725 -41225 -8525
rect -40825 -9125 -12825 -8925
rect -40825 -36125 -40625 -9125
rect -40225 -9725 -13425 -9525
rect -40225 -35525 -40025 -9725
rect -39625 -10325 -14025 -10125
rect -39625 -34925 -39425 -10325
rect -27284 -34704 -27024 -34666
rect -27284 -34768 -27246 -34704
rect -27182 -34768 -27126 -34704
rect -27062 -34768 -27024 -34704
rect -27284 -34824 -27024 -34768
rect -27284 -34888 -27246 -34824
rect -27182 -34888 -27126 -34824
rect -27062 -34888 -27024 -34824
rect -27284 -34925 -27024 -34888
rect -39625 -34926 -27024 -34925
rect -39625 -35125 -27025 -34926
rect -14225 -35525 -14025 -10325
rect -40225 -35725 -14025 -35525
rect -13625 -36125 -13425 -9725
rect -40825 -36325 -13425 -36125
rect -13025 -36725 -12825 -9125
rect -41425 -36925 -12825 -36725
rect -12425 -37325 -12225 -8525
rect -42025 -37525 -12225 -37325
rect -11825 -37925 -11625 -7925
rect -42625 -38125 -11625 -37925
rect -11225 -38525 -11025 -7325
rect -43225 -38725 -11025 -38525
rect -10625 -39125 -10425 -6725
rect -43825 -39325 -10425 -39125
rect -10025 -39725 -9825 -6125
rect -44425 -39925 -9825 -39725
rect -9425 -40325 -9225 -5525
rect -5089 -5526 30111 -5326
rect -5089 -39726 -4889 -5526
rect -4489 -6126 29511 -5926
rect -4489 -39126 -4289 -6126
rect -3889 -6726 28911 -6526
rect -3889 -38526 -3689 -6726
rect -3289 -7326 28311 -7126
rect -3289 -37926 -3089 -7326
rect -2689 -7926 27711 -7726
rect -2689 -37326 -2489 -7926
rect -2089 -8526 27111 -8326
rect -2089 -36726 -1889 -8526
rect -1489 -9126 26511 -8926
rect -1489 -36126 -1289 -9126
rect -889 -9726 25911 -9526
rect -889 -35526 -689 -9726
rect -289 -10326 25311 -10126
rect -289 -34926 -89 -10326
rect 12051 -34705 12311 -34667
rect 12051 -34769 12089 -34705
rect 12153 -34769 12209 -34705
rect 12273 -34769 12311 -34705
rect 12051 -34825 12311 -34769
rect 12051 -34889 12089 -34825
rect 12153 -34889 12209 -34825
rect 12273 -34889 12311 -34825
rect 12051 -34926 12311 -34889
rect -289 -35126 12311 -34926
rect 25111 -35526 25311 -10326
rect -889 -35726 25311 -35526
rect 25711 -36126 25911 -9726
rect -1489 -36326 25911 -36126
rect 26311 -36726 26511 -9126
rect -2089 -36926 26511 -36726
rect 26911 -37326 27111 -8526
rect -2689 -37526 27111 -37326
rect 27511 -37926 27711 -7926
rect -3289 -38126 27711 -37926
rect 28111 -38526 28311 -7326
rect -3889 -38726 28311 -38526
rect 28711 -39126 28911 -6726
rect -4489 -39326 28911 -39126
rect 29311 -39726 29511 -6126
rect -5089 -39926 29511 -39726
rect -27247 -40525 -9225 -40325
rect 29911 -40326 30111 -5526
rect -27247 -41605 -27047 -40525
rect -3176 -40526 30111 -40326
rect -27247 -41805 -8553 -41605
rect -8753 -43181 -8553 -41805
rect -3176 -43180 -2976 -40526
rect -8788 -43219 -8528 -43181
rect -8788 -43283 -8750 -43219
rect -8686 -43283 -8630 -43219
rect -8566 -43283 -8528 -43219
rect -8788 -43339 -8528 -43283
rect -8788 -43403 -8750 -43339
rect -8686 -43403 -8630 -43339
rect -8566 -43403 -8528 -43339
rect -8788 -43441 -8528 -43403
rect -3203 -43218 -2943 -43180
rect -3203 -43282 -3165 -43218
rect -3101 -43282 -3045 -43218
rect -2981 -43282 -2943 -43218
rect -3203 -43338 -2943 -43282
rect -3203 -43402 -3165 -43338
rect -3101 -43402 -3045 -43338
rect -2981 -43402 -2943 -43338
rect -3203 -43440 -2943 -43402
rect -10430 -43725 -10170 -43710
rect -10430 -43961 -10420 -43725
rect -10184 -43961 -10170 -43725
rect -10430 -43970 -10170 -43961
rect -10430 -44957 -10170 -44948
rect -10430 -44963 -10419 -44957
rect -10430 -45199 -10420 -44963
rect -10183 -45193 -10170 -44957
rect -10184 -45199 -10170 -45193
rect -10430 -45208 -10170 -45199
rect -6859 -45049 -6599 -45040
rect -6859 -45055 -6848 -45049
rect -6859 -45291 -6849 -45055
rect -6612 -45243 -6599 -45049
rect -5232 -45055 -4972 -45043
rect -6859 -45292 -6848 -45291
rect -6612 -45292 -6598 -45243
rect -6859 -45300 -6598 -45292
rect -6858 -45303 -6598 -45300
rect -5232 -45291 -5220 -45055
rect -4984 -45291 -4972 -45055
rect -5232 -45303 -4972 -45291
rect -6855 -45917 -6595 -45905
rect -6855 -46153 -6843 -45917
rect -6607 -46153 -6595 -45917
rect -6855 -46165 -6595 -46153
rect -5229 -45917 -4969 -45905
rect -5229 -46153 -5217 -45917
rect -4981 -46153 -4969 -45917
rect -5229 -46165 -4969 -46153
<< via4 >>
rect -10420 -43748 -10184 -43725
rect -10420 -43751 -10392 -43748
rect -10392 -43751 -10328 -43748
rect -10328 -43751 -10272 -43748
rect -10272 -43751 -10208 -43748
rect -10420 -43815 -10394 -43751
rect -10394 -43812 -10328 -43751
rect -10328 -43812 -10274 -43751
rect -10274 -43812 -10208 -43751
rect -10208 -43812 -10184 -43748
rect -10394 -43815 -10330 -43812
rect -10330 -43815 -10274 -43812
rect -10274 -43815 -10210 -43812
rect -10210 -43815 -10184 -43812
rect -10420 -43868 -10184 -43815
rect -10420 -43871 -10392 -43868
rect -10392 -43871 -10328 -43868
rect -10328 -43871 -10272 -43868
rect -10272 -43871 -10208 -43868
rect -10420 -43935 -10394 -43871
rect -10394 -43932 -10328 -43871
rect -10328 -43932 -10274 -43871
rect -10274 -43932 -10208 -43871
rect -10208 -43932 -10184 -43868
rect -10394 -43935 -10330 -43932
rect -10330 -43935 -10274 -43932
rect -10274 -43935 -10210 -43932
rect -10210 -43935 -10184 -43932
rect -10420 -43961 -10184 -43935
rect -10419 -44963 -10183 -44957
rect -10420 -44983 -10183 -44963
rect -10420 -44989 -10393 -44983
rect -10393 -44986 -10329 -44983
rect -10329 -44986 -10273 -44983
rect -10273 -44986 -10209 -44983
rect -10209 -44986 -10183 -44983
rect -10393 -44989 -10328 -44986
rect -10328 -44989 -10273 -44986
rect -10273 -44989 -10208 -44986
rect -10420 -45053 -10394 -44989
rect -10394 -45050 -10328 -44989
rect -10328 -45050 -10274 -44989
rect -10274 -45050 -10208 -44989
rect -10208 -45050 -10183 -44986
rect -10394 -45053 -10330 -45050
rect -10330 -45053 -10274 -45050
rect -10274 -45053 -10210 -45050
rect -10210 -45053 -10183 -45050
rect -10420 -45103 -10183 -45053
rect -10420 -45109 -10393 -45103
rect -10393 -45106 -10329 -45103
rect -10329 -45106 -10273 -45103
rect -10273 -45106 -10209 -45103
rect -10209 -45106 -10183 -45103
rect -10393 -45109 -10328 -45106
rect -10328 -45109 -10273 -45106
rect -10273 -45109 -10208 -45106
rect -10420 -45173 -10394 -45109
rect -10394 -45170 -10328 -45109
rect -10328 -45170 -10274 -45109
rect -10274 -45170 -10208 -45109
rect -10208 -45170 -10183 -45106
rect -10394 -45173 -10330 -45170
rect -10330 -45173 -10274 -45170
rect -10274 -45173 -10210 -45170
rect -10210 -45173 -10183 -45170
rect -10420 -45193 -10183 -45173
rect -10420 -45199 -10184 -45193
rect -6848 -45055 -6612 -45049
rect -6849 -45075 -6612 -45055
rect -6849 -45081 -6822 -45075
rect -6822 -45078 -6758 -45075
rect -6758 -45078 -6702 -45075
rect -6702 -45078 -6638 -45075
rect -6638 -45078 -6612 -45075
rect -6822 -45081 -6757 -45078
rect -6757 -45081 -6702 -45078
rect -6702 -45081 -6637 -45078
rect -6849 -45145 -6823 -45081
rect -6823 -45142 -6757 -45081
rect -6757 -45142 -6703 -45081
rect -6703 -45142 -6637 -45081
rect -6637 -45142 -6612 -45078
rect -6823 -45145 -6758 -45142
rect -6758 -45145 -6703 -45142
rect -6703 -45145 -6638 -45142
rect -6849 -45146 -6822 -45145
rect -6822 -45146 -6758 -45145
rect -6758 -45146 -6702 -45145
rect -6702 -45146 -6638 -45145
rect -6638 -45146 -6612 -45142
rect -6849 -45195 -6612 -45146
rect -6849 -45201 -6822 -45195
rect -6822 -45198 -6758 -45195
rect -6758 -45198 -6702 -45195
rect -6702 -45198 -6638 -45195
rect -6638 -45198 -6612 -45195
rect -6822 -45201 -6757 -45198
rect -6757 -45201 -6702 -45198
rect -6702 -45201 -6637 -45198
rect -6849 -45265 -6823 -45201
rect -6823 -45262 -6757 -45201
rect -6757 -45262 -6703 -45201
rect -6703 -45262 -6637 -45201
rect -6637 -45262 -6612 -45198
rect -6823 -45265 -6758 -45262
rect -6758 -45265 -6703 -45262
rect -6703 -45265 -6638 -45262
rect -6849 -45266 -6822 -45265
rect -6822 -45266 -6758 -45265
rect -6758 -45266 -6702 -45265
rect -6702 -45266 -6638 -45265
rect -6638 -45266 -6612 -45262
rect -6849 -45291 -6612 -45266
rect -6848 -45292 -6612 -45291
rect -5220 -45081 -4984 -45055
rect -5220 -45145 -5194 -45081
rect -5194 -45145 -5130 -45081
rect -5130 -45145 -5074 -45081
rect -5074 -45145 -5010 -45081
rect -5010 -45145 -4984 -45081
rect -5220 -45201 -4984 -45145
rect -5220 -45265 -5194 -45201
rect -5194 -45265 -5130 -45201
rect -5130 -45265 -5074 -45201
rect -5074 -45265 -5010 -45201
rect -5010 -45265 -4984 -45201
rect -5220 -45291 -4984 -45265
rect -6843 -45943 -6607 -45917
rect -6843 -46007 -6817 -45943
rect -6817 -46007 -6753 -45943
rect -6753 -46007 -6697 -45943
rect -6697 -46007 -6633 -45943
rect -6633 -46007 -6607 -45943
rect -6843 -46063 -6607 -46007
rect -6843 -46127 -6817 -46063
rect -6817 -46127 -6753 -46063
rect -6753 -46127 -6697 -46063
rect -6697 -46127 -6633 -46063
rect -6633 -46127 -6607 -46063
rect -6843 -46153 -6607 -46127
rect -5217 -45943 -4981 -45917
rect -5217 -46007 -5191 -45943
rect -5191 -46007 -5127 -45943
rect -5127 -46007 -5071 -45943
rect -5071 -46007 -5007 -45943
rect -5007 -46007 -4981 -45943
rect -5217 -46063 -4981 -46007
rect -5217 -46127 -5191 -46063
rect -5191 -46127 -5127 -46063
rect -5127 -46127 -5071 -46063
rect -5071 -46127 -5007 -46063
rect -5007 -46127 -4981 -46063
rect -5217 -46153 -4981 -46127
<< metal5 >>
rect -10511 -43725 -10090 -43630
rect -10511 -43961 -10420 -43725
rect -10184 -43961 -10090 -43725
rect -10511 -44050 -10090 -43961
rect -10511 -44957 -10090 -44868
rect -10511 -44963 -10419 -44957
rect -10511 -45199 -10420 -44963
rect -10183 -45193 -10090 -44957
rect -10184 -45199 -10090 -45193
rect -10511 -45288 -10090 -45199
rect -6939 -45049 -6518 -44963
rect -6939 -45055 -6848 -45049
rect -6939 -45291 -6849 -45055
rect -6939 -45292 -6848 -45291
rect -6612 -45292 -6518 -45049
rect -6939 -45383 -6518 -45292
rect -5313 -45055 -4892 -44963
rect -5313 -45291 -5220 -45055
rect -4984 -45291 -4892 -45055
rect -5313 -45383 -4892 -45291
rect -6936 -45917 -6515 -45825
rect -6936 -46153 -6843 -45917
rect -6607 -46153 -6515 -45917
rect -6936 -46245 -6515 -46153
rect -5310 -45917 -4889 -45825
rect -5310 -46153 -5217 -45917
rect -4981 -46153 -4889 -45917
rect -5310 -46245 -4889 -46153
<< labels >>
flabel metal1 s -10030 -43867 -9979 -43824 2 FreeSans 125000 0 0 0 IN1
port 1 nsew
flabel metal1 s -10030 -45097 -9989 -45058 2 FreeSans 125000 0 0 0 IN2
port 2 nsew
flabel metal1 s -7140 -34634 -6466 -34600 2 FreeSans 125000 0 0 0 VDD
port 4 nsew
flabel metal2 s -1081 -43082 -1056 -43059 2 FreeSans 125000 0 0 0 OUT1
port 5 nsew
flabel metal2 s -1080 -43189 -1053 -43169 2 FreeSans 125000 0 0 0 OUT2
port 6 nsew
rlabel metal1 -2226 -47096 -2142 -46954 7 Ground
port 7 w
<< end >>
