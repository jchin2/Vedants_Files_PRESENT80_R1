* NGSPICE file created from EESPFAL_PRESENT80_R1_flat.ext - technology: sky130A

.subckt EESPFAL_PRESENT80_R1_flat GND x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar x2 x2_bar
+ k2 k2_bar x3 x3_bar k3 k3_bar s0 s0_bar Dis0 Dis1 s2 s2_bar s3_bar s3 s1_bar s1
+ Dis2 Dis3 CLK0 CLK2 CLK3 CLK1
X0 s0.t3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B CLK3.t26 GND.t217 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 CLK0.t33 x3_bar.t0 a_1180_5008# GND.t239 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t6 CLK1.t186 CLK1.t185 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 GND.t241 Dis3.t0 s1_bar.t0 GND.t240 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t6 GND.t65 GND.t64 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 GND.t275 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar GND.t274 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X6 a_6287_n6133# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6137_n6133# GND.t135 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X7 CLK1.t11 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A CLK1.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B CLK1.t74 CLK1.t73 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X9 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t6 a_6476_n1173# GND.t134 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X10 CLK1.t29 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6136_4548# GND.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X11 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B CLK0.t38 CLK0.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 GND.t253 Dis2.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B GND.t252 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X13 GND.t71 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t3 GND.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_6436_4548# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t6 CLK1.t105 GND.t97 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_4916_n1173# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B CLK1.t166 GND.t37 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X16 CLK1.t106 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t7 a_4576_4548# GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X17 CLK1.t21 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B CLK1.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X18 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t6 GND.t141 GND.t140 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t6 GND.t300 GND.t156 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X20 a_4876_4548# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A CLK1.t30 GND.t47 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X21 GND.t255 Dis2.t1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT GND.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X22 CLK1.t66 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t6 a_6287_n6133# GND.t114 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X23 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B CLK1.t28 CLK1.t27 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X24 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A CLK1.t162 CLK1.t161 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X25 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A CLK2.t61 CLK2.t60 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X26 CLK0.t21 x1.t0 a_2740_7368# GND.t213 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X27 CLK2.t87 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t3 GND.t299 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X28 CLK1.t141 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar CLK1.t140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X29 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar CLK2.t57 GND.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X30 CLK2.t59 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar CLK2.t58 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X31 CLK1.t132 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A CLK1.t131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X32 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar CLK1.t90 CLK1.t89 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X33 GND.t287 Dis2.t2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT GND.t286 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X34 s3.t0 Dis3.t1 GND.t356 GND.t355 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X35 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t0 Dis1.t0 GND.t154 GND.t153 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X36 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 GND.t328 GND.t327 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X37 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6476_n493# GND.t134 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X38 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t6 GND.t193 GND.t192 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X39 CLK0.t16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t1 CLK0.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X40 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar Dis1.t1 GND.t20 GND.t19 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X41 CLK1.t31 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B GND.t46 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X42 GND.t288 Dis2.t3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT GND.t174 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X43 GND.t18 Dis1.t2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A GND.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X44 GND.t106 s2_bar.t5 s2.t6 GND.t105 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X45 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t6 CLK0.t18 CLK0.t17 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X46 CLK1.t95 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar CLK1.t94 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X47 s2_bar.t4 s2.t7 GND.t340 GND.t339 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X48 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar CLK1.t56 CLK1.t55 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X49 CLK1.t82 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t7 a_6136_n3993# GND.t41 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X50 a_6137_2408# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t7 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A GND.t335 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X51 a_10206_4548# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT GND.t34 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X52 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar Dis1.t3 GND.t264 GND.t263 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X53 CLK2.t66 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t7 a_10206_4548# GND.t208 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X54 a_4576_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t2 GND.t75 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X55 s3.t5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT CLK3.t25 GND.t283 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X56 CLK1.t39 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t8 a_4576_n3313# GND.t49 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X57 a_10206_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT GND.t6 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X58 CLK1.t40 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t9 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B GND.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X59 GND.t138 Dis1.t4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B GND.t119 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X60 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar CLK2.t2 GND.t9 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X61 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t6 CLK1.t170 CLK1.t169 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X62 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 CLK2.t54 CLK2.t53 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X63 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 GND.t73 GND.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X64 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6436_n3313# GND.t133 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X65 a_6436_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t7 CLK1.t151 GND.t172 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X66 CLK2.t103 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t2 CLK2.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X67 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t8 CLK1.t196 CLK1.t195 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X68 CLK1.t164 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B GND.t219 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X69 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar GND.t296 GND.t260 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X70 a_8456_7368# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B GND.t202 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X71 a_1180_7368# k1_bar.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t5 GND.t179 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X72 CLK3.t16 s3_bar.t5 s3.t3 CLK3.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X73 CLK1.t104 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t4 CLK1.t103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X74 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar Dis2.t4 GND.t236 GND.t223 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X75 CLK3.t6 s1_bar.t5 s1.t3 CLK3.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X76 a_10265_n1173# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT GND.t100 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X77 CLK3.t20 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT s3.t4 GND.t273 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X78 a_4876_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A CLK1.t34 GND.t45 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X79 CLK2.t8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t6 a_10206_n3313# GND.t63 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X80 a_6136_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t0 GND.t218 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X81 CLK0.t40 x1_bar.t0 a_1180_7368# GND.t187 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X82 s1_bar.t3 s1.t7 CLK3.t14 CLK3.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X83 GND.t161 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar GND.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X84 CLK2.t40 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B CLK2.t39 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X85 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t1 Dis1.t5 GND.t338 GND.t308 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X86 CLK1.t7 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar CLK1.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X87 CLK1.t44 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t0 CLK1.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X88 CLK0.t29 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t8 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t1 CLK0.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X89 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A k0.t0 a_3040_8048# GND.t50 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X90 a_4576_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t8 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t0 GND.t180 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X91 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X92 GND.t238 Dis2.t5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t0 GND.t237 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X93 GND.t215 Dis0.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A GND.t168 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X94 a_10476_7368# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar s0_bar.t1 GND.t184 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X95 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t8 CLK0.t25 CLK0.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X96 s3_bar.t2 s3.t7 CLK3.t32 CLK3.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X97 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t7 CLK1.t136 CLK1.t135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X98 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4916_n493# GND.t132 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X99 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A CLK1.t121 CLK1.t77 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X100 CLK2.t23 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar CLK2.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X101 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A CLK1.t78 CLK1.t77 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X102 s2.t3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT CLK3.t11 GND.t166 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X103 GND.t329 Dis1.t6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t5 GND.t91 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X104 GND.t222 Dis1.t7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B GND.t83 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X105 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar CLK1.t158 CLK1.t157 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X106 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t0 k2.t0 a_3040_5688# GND.t101 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X107 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t9 CLK1.t150 GND.t284 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X108 GND.t62 Dis1.t8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B GND.t61 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X109 GND.t120 Dis1.t9 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B GND.t119 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X110 GND.t280 Dis0.t1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t3 GND.t266 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X111 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar GND.t227 GND.t226 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X112 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT CLK2.t70 CLK2.t69 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X113 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t9 CLK1.t122 GND.t40 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X114 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t7 CLK2.t114 CLK2.t113 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X115 CLK1.t108 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t4 CLK1.t107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X116 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT CLK2.t31 CLK2.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X117 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t5 CLK2.t89 CLK2.t88 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X118 GND.t307 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t4 GND.t220 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X119 CLK2.t29 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t3 CLK2.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X120 CLK2.t68 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar CLK2.t67 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X121 CLK2.t81 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 CLK2.t80 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X122 a_3040_5008# x3_bar.t1 CLK0.t34 GND.t57 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X123 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B CLK1.t182 CLK1.t181 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X124 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t9 GND.t182 GND.t181 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X125 CLK2.t112 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t8 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT CLK2.t111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X126 a_1480_5008# x3.t0 CLK0.t9 GND.t55 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X127 s2.t5 s2_bar.t6 CLK3.t24 CLK3.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X128 a_6136_5228# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t8 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t0 GND.t60 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X129 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t1 k3.t0 a_1480_5008# GND.t173 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X130 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t1 Dis1.t10 GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X131 a_7196_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t10 CLK1.t177 GND.t164 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X132 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t10 CLK1.t99 GND.t195 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X133 a_4576_5228# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t9 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t0 GND.t194 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X134 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t10 a_7196_8048# GND.t289 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X135 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar CLK1.t52 CLK1.t8 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X136 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t1 Dis2.t6 GND.t245 GND.t148 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X137 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t7 CLK2.t52 GND.t77 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X138 CLK1.t165 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6176_n1173# GND.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X139 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6436_4548# GND.t128 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X140 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B CLK2.t79 CLK2.t78 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X141 GND.t68 Dis1.t11 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t1 GND.t67 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X142 a_2740_8048# k0_bar.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A GND.t56 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X143 CLK3.t8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t7 a_10377_n6134# GND.t111 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X144 a_4616_n1173# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t11 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t5 GND.t139 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X145 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4876_4548# GND.t127 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X146 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t5 Dis0.t2 GND.t352 GND.t102 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X147 GND.t246 Dis2.t7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A GND.t211 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X148 a_10265_n493# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT GND.t100 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X149 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar Dis2.t8 GND.t144 GND.t143 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X150 CLK1.t26 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar CLK1.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X151 CLK1.t117 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B CLK1.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X152 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t0 Dis2.t9 GND.t146 GND.t145 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X153 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t8 CLK2.t1 GND.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X154 GND.t349 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar GND.t158 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X155 GND.t282 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t3 GND.t274 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X156 a_6137_n6133# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A GND.t306 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X157 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B CLK1.t86 CLK1.t85 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X158 a_6476_n1173# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t10 CLK1.t96 GND.t80 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X159 a_2740_5688# k2_bar.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t5 GND.t178 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X160 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar CLK2.t86 CLK2.t85 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X161 CLK1.t88 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B CLK1.t87 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X162 CLK2.t4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar GND.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X163 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t3 Dis0.t3 GND.t214 GND.t136 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X164 CLK1.t97 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t11 a_4616_n1173# GND.t190 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X165 CLK1.t128 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B CLK1.t127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X166 GND.t165 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t4 GND.t150 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X167 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t6 CLK1.t176 CLK1.t175 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X168 s1.t5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t5 CLK3.t12 GND.t196 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X169 a_6176_1648# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t11 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A GND.t290 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X170 CLK0.t12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t10 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A CLK0.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X171 GND.t298 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar GND.t297 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X172 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar Dis1.t12 GND.t231 GND.t230 sky130_fd_pr__nfet_01v8 ad=3.6e+12p pd=1.68e+07u as=0p ps=0u w=1.5e+06u l=150000u
X173 a_6287_2408# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6137_2408# GND.t44 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X174 s0.t0 Dis3.t2 GND.t110 GND.t109 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X175 CLK1.t45 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t12 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar GND.t76 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X176 GND.t244 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar GND.t243 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X177 GND.t12 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar GND.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X178 CLK1.t100 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t12 a_6287_2408# GND.t201 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X179 GND.t233 s0_bar.t5 s0.t1 GND.t232 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X180 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t11 CLK1.t24 GND.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X181 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A CLK1.t81 GND.t131 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X182 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar GND.t257 GND.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X183 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar CLK1.t115 CLK1.t114 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X184 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t8 CLK2.t14 CLK2.t13 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X185 CLK2.t50 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t5 GND.t225 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X186 CLK1.t178 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t11 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar GND.t336 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X187 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B Dis1.t13 GND.t108 GND.t107 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X188 CLK1.t101 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t13 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B GND.t46 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X189 CLK2.t15 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar GND.t117 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X190 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar GND.t272 GND.t271 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X191 GND.t43 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t2 GND.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X192 CLK2.t71 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t6 a_8456_7368# GND.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X193 CLK1.t149 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t9 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t1 CLK1.t148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X194 a_3040_7368# x1_bar.t1 CLK0.t10 GND.t104 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X195 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 Dis2.t10 GND.t52 GND.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X196 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t12 GND.t171 GND.t170 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X197 GND.t291 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar GND.t185 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X198 CLK1.t35 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6136_n3313# GND.t41 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X199 a_6136_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t14 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t1 GND.t58 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X200 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar CLK2.t65 GND.t270 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X201 CLK2.t27 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT CLK2.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X202 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar CLK1.t9 CLK1.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X203 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t7 CLK1.t172 CLK1.t171 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X204 CLK1.t79 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6136_8048# GND.t130 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X205 a_1480_7368# x1.t1 CLK0.t41 GND.t0 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X206 CLK1.t13 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t0 CLK1.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X207 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar GND.t183 GND.t88 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X208 GND.t54 Dis2.t11 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t0 GND.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X209 CLK3.t1 s1.t8 s1_bar.t2 CLK3.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X210 CLK2.t12 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t9 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT CLK2.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X211 GND.t313 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t5 GND.t268 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X212 a_6436_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t12 CLK1.t137 GND.t265 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X213 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t3 k1.t0 a_1480_7368# GND.t81 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X214 a_4576_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t13 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t1 GND.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X215 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar CLK2.t9 GND.t87 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X216 CLK2.t3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t1 GND.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X217 GND.t79 Dis1.t14 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B GND.t78 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X218 CLK1.t154 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t14 a_4576_8048# GND.t292 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X219 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t7 GND.t249 GND.t162 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X220 CLK3.t27 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar a_10476_7368# GND.t295 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X221 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t6 CLK2.t19 GND.t142 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X222 CLK1.t70 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B CLK1.t69 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X223 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 Dis2.t12 GND.t333 GND.t332 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X224 CLK0.t31 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t4 CLK0.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X225 a_4876_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A CLK1.t80 GND.t35 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X226 GND.t113 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 GND.t112 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X227 a_6436_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t13 CLK1.t91 GND.t172 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X228 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t14 CLK1.t197 GND.t303 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X229 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t12 CLK1.t191 GND.t347 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X230 CLK3.t9 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT s2.t2 GND.t152 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X231 GND.t229 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 GND.t228 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X232 s3.t6 s3_bar.t6 CLK3.t46 CLK3.t45 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X233 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t8 CLK1.t58 CLK1.t57 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X234 s2.t1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t7 CLK3.t28 GND.t310 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X235 GND.t189 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t7 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t5 GND.t188 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X236 s1.t0 Dis3.t3 GND.t326 GND.t325 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X237 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B CLK1.t5 CLK1.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X238 CLK1.t145 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A CLK1.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X239 GND.t118 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar GND.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X240 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar Dis1.t15 GND.t66 GND.t28 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X241 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A CLK1.t36 GND.t40 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X242 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar CLK1.t126 CLK1.t125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X243 CLK2.t84 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A CLK2.t83 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X244 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A CLK0.t14 CLK0.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X245 CLK2.t10 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar GND.t90 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X246 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT CLK2.t36 CLK2.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X247 GND.t92 Dis1.t16 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t1 GND.t91 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X248 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t7 GND.t324 GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X249 GND.t342 Dis3.t4 s3_bar.t0 GND.t341 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X250 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t8 CLK2.t49 GND.t217 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X251 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar Dis2.t13 GND.t334 GND.t145 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X252 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t7 CLK2.t93 CLK2.t92 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X253 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 CLK2.t101 CLK2.t100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X254 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B k3.t1 a_3040_5008# GND.t101 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X255 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar GND.t116 GND.t115 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X256 s0.t5 s0_bar.t6 CLK3.t42 CLK3.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X257 GND.t167 Dis1.t17 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B GND.t61 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X258 GND.t99 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar GND.t98 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X259 GND.t151 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar GND.t150 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X260 GND.t210 Dis3.t5 s2_bar.t0 GND.t209 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X261 GND.t267 Dis0.t4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B GND.t266 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X262 CLK2.t91 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t8 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT CLK2.t90 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X263 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 CLK2.t117 CLK2.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X264 CLK3.t39 s0_bar.t7 s0.t4 CLK3.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X265 CLK3.t19 s2_bar.t7 s2.t4 CLK3.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X266 CLK1.t192 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t13 a_6136_5228# GND.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X267 a_10227_2407# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 s1_bar.t4 GND.t216 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X268 GND.t293 Dis1.t18 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B GND.t252 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X269 CLK2.t34 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t3 CLK2.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X270 GND.t82 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t7 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t3 GND.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X271 s2_bar.t2 s2.t8 CLK3.t22 CLK3.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X272 a_6436_5228# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t14 CLK1.t59 GND.t97 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X273 a_10377_2407# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar a_10227_2407# GND.t204 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X274 CLK1.t23 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t15 a_4576_5228# GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X275 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A CLK1.t17 CLK1.t16 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X276 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t7 GND.t281 GND.t140 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X277 CLK0.t5 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t1 CLK0.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X278 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4876_n3993# GND.t126 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X279 a_4876_5228# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t14 CLK1.t119 GND.t47 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X280 a_6176_n493# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t15 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A GND.t197 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X281 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t15 CLK0.t39 CLK0.t24 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X282 CLK2.t6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t1 CLK2.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X283 CLK2.t77 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar CLK2.t76 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X284 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar Dis1.t19 GND.t96 GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X285 a_4616_n493# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t16 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar GND.t139 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X286 CLK0.t26 x0.t0 a_2740_8048# GND.t213 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X287 GND.t124 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar GND.t123 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X288 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar CLK2.t38 CLK2.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X289 CLK2.t16 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_10265_n493# GND.t122 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X290 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t15 CLK0.t28 CLK0.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X291 CLK1.t189 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t16 a_4616_n493# GND.t190 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X292 a_10227_n6134# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 s3_bar.t4 GND.t121 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X293 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar GND.t203 GND.t192 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X294 CLK1.t22 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t16 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B GND.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X295 CLK1.t84 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar CLK1.t83 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X296 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar Dis1.t20 GND.t29 GND.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X297 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT CLK2.t21 CLK2.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X298 GND.t175 Dis2.t14 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT GND.t174 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X299 CLK0.t32 x2.t0 a_2740_5688# GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X300 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar CLK1.t3 CLK1.t2 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X301 a_6176_n1173# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t17 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t2 GND.t197 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X302 GND.t337 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar GND.t98 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X303 CLK1.t174 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t8 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t3 CLK1.t173 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X304 a_10377_n6134# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar a_10227_n6134# GND.t206 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X305 a_10206_5228# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT GND.t34 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X306 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t9 CLK1.t188 CLK1.t187 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X307 a_6326_1648# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6176_1648# GND.t129 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X308 CLK0.t36 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t2 CLK0.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X309 CLK2.t56 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t8 a_10206_5228# GND.t208 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X310 a_6476_1648# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6326_1648# GND.t39 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X311 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t15 CLK0.t8 CLK0.t7 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X312 a_2740_5008# k3_bar.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B GND.t178 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X313 a_10446_1647# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 s2_bar.t1 GND.t322 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X314 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar GND.t86 GND.t85 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X315 CLK1.t111 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t16 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar GND.t219 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X316 s0_bar.t4 s0.t6 GND.t261 GND.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X317 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t0 Dis0.t5 GND.t137 GND.t136 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X318 CLK1.t190 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t17 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar GND.t343 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X319 GND.t277 Dis1.t21 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A GND.t276 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X320 GND.t321 Dis1.t22 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A GND.t320 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X321 CLK1.t102 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t18 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B GND.t202 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X322 a_1180_8048# k0_bar.t1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t3 GND.t179 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X323 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B CLK1.t167 GND.t305 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X324 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar Dis1.t23 GND.t224 GND.t223 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X325 a_6136_7368# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t18 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B GND.t218 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X326 GND.t14 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B GND.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X327 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar Dis1.t24 GND.t309 GND.t308 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X328 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B CLK1.t63 CLK1.t62 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X329 CLK0.t20 x0_bar.t0 a_1180_8048# GND.t187 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X330 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT CLK2.t75 CLK2.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X331 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A k1.t1 a_3040_7368# GND.t50 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X332 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B GND.t33 GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X333 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar Dis1.t25 GND.t279 GND.t278 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X334 GND.t169 Dis0.t6 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A GND.t168 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X335 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t6 GND.t316 GND.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X336 CLK1.t147 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t8 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t3 CLK1.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X337 a_10476_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A GND.t184 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X338 a_1180_5688# k2_bar.t1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t4 GND.t251 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X339 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT CLK2.t110 CLK2.t109 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X340 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6436_8048# GND.t304 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X341 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t8 CLK1.t50 CLK1.t49 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X342 CLK0.t27 x2_bar.t0 a_1180_5688# GND.t239 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X343 CLK1.t184 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t3 CLK1.t183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X344 CLK1.t61 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar CLK1.t60 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X345 GND.t84 Dis1.t26 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t1 GND.t83 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X346 CLK2.t73 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t4 CLK2.t72 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X347 CLK2.t108 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar CLK2.t107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X348 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4876_8048# GND.t284 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X349 CLK2.t82 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t5 GND.t117 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X350 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar GND.t205 GND.t64 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X351 CLK1.t54 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B CLK1.t53 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X352 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 GND.t248 GND.t247 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X353 CLK1.t72 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar CLK1.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X354 GND.t262 Dis1.t27 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t4 GND.t198 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X355 a_6136_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t17 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t0 GND.t58 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X356 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t16 CLK1.t41 GND.t59 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X357 GND.t177 Dis2.t15 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t0 GND.t176 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X358 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t8 CLK1.t47 CLK1.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X359 GND.t331 s1_bar.t6 s1.t4 GND.t330 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X360 s1.t1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT CLK3.t10 GND.t160 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X361 GND.t350 Dis2.t16 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT GND.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X362 s3.t1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t6 CLK3.t33 GND.t323 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X363 s1_bar.t1 s1.t9 GND.t31 GND.t30 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X364 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar CLK1.t68 CLK1.t67 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X365 CLK1.t160 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar CLK1.t159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X366 CLK3.t40 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT s1.t6 GND.t348 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X367 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B CLK1.t168 GND.t303 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X368 CLK1.t42 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t18 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar GND.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X369 a_6136_4548# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t17 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t0 GND.t60 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X370 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t5 Dis1.t28 GND.t314 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X371 CLK2.t32 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar GND.t164 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X372 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t1 Dis1.t29 GND.t318 GND.t153 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X373 GND.t235 s3_bar.t7 s3.t2 GND.t234 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X374 GND.t285 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t9 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t5 GND.t188 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X375 a_4576_4548# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t18 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t0 GND.t194 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X376 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar GND.t157 GND.t156 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X377 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar CLK1.t19 CLK1.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X378 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t19 CLK1.t98 GND.t195 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X379 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t9 CLK2.t99 GND.t289 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X380 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar CLK1.t143 CLK1.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X381 CLK1.t76 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar CLK1.t75 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X382 CLK2.t55 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar GND.t225 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X383 GND.t351 Dis2.t17 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT GND.t286 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X384 s0_bar.t3 s0.t7 CLK3.t37 CLK3.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X385 GND.t5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar GND.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X386 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar Dis1.t30 GND.t315 GND.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X387 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t7 CLK2.t18 CLK2.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X388 CLK3.t2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t9 a_10377_2407# GND.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X389 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6436_5228# GND.t128 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X390 a_2740_7368# k1_bar.t1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A GND.t56 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X391 CLK2.t51 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t4 GND.t242 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X392 CLK1.t15 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar CLK1.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X393 GND.t191 Dis1.t31 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t1 GND.t67 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X394 GND.t212 Dis3.t6 s0_bar.t0 GND.t211 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X395 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B CLK1.t139 CLK1.t138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X396 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t8 GND.t27 GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X397 s3_bar.t3 s3.t8 GND.t95 GND.t94 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X398 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t4 Dis0.t7 GND.t103 GND.t102 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X399 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 Dis2.t18 GND.t345 GND.t344 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X400 CLK1.t37 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6176_n493# GND.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X401 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4876_5228# GND.t127 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X402 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar CLK1.t130 CLK1.t129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X403 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t1 Dis2.t19 GND.t346 GND.t143 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X404 CLK0.t23 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t19 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A CLK0.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X405 GND.t312 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t8 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 GND.t311 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X406 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar GND.t294 GND.t115 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X407 CLK1.t118 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t19 a_4576_n3993# GND.t49 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X408 a_6476_n493# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t20 CLK1.t48 GND.t80 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X409 a_10206_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT GND.t6 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X410 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar CLK2.t25 CLK2.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X411 GND.t159 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t5 GND.t158 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X412 CLK2.t97 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 CLK2.t96 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X413 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar GND.t8 GND.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X414 a_4916_n493# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A CLK1.t38 GND.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X415 s2.t0 Dis3.t7 GND.t354 GND.t353 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X416 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6436_n3993# GND.t133 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X417 GND.t199 Dis1.t32 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A GND.t198 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X418 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B CLK1.t93 CLK1.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X419 CLK2.t0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t0 GND.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X420 CLK2.t115 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t7 a_10265_n1173# GND.t122 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X421 CLK1.t180 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar CLK1.t179 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X422 a_4876_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t17 CLK1.t112 GND.t45 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X423 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4876_n3313# GND.t126 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X424 CLK2.t106 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t9 a_10206_n3993# GND.t63 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X425 CLK2.t105 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t1 CLK2.t104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X426 CLK1.t1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B CLK1.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X427 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t8 CLK1.t65 CLK1.t64 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X428 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar GND.t250 GND.t226 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X429 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t7 CLK2.t64 CLK2.t63 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X430 CLK1.t120 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar CLK1.t75 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X431 CLK2.t95 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t8 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 CLK2.t94 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X432 CLK3.t30 s3.t9 s3_bar.t1 CLK3.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X433 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar Dis2.t20 GND.t147 GND.t109 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X434 CLK1.t134 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t9 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t3 CLK1.t133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X435 CLK1.t194 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t10 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t5 CLK1.t193 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X436 GND.t259 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar GND.t232 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X437 s1.t2 s1_bar.t7 CLK3.t44 CLK3.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X438 CLK1.t156 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B CLK1.t155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X439 CLK1.t124 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t9 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t3 CLK1.t123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X440 CLK1.t198 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t20 a_6476_1648# GND.t357 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X441 CLK0.t43 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t21 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B CLK0.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X442 a_10596_1647# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar a_10446_1647# GND.t155 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X443 CLK0.t1 x3.t1 a_2740_5008# GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X444 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar Dis1.t33 GND.t200 GND.t107 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X445 GND.t125 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t2 GND.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X446 CLK3.t7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t9 a_10596_1647# GND.t93 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X447 a_3040_8048# x0_bar.t1 CLK0.t19 GND.t104 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X448 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A CLK1.t33 GND.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X449 CLK1.t113 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t18 a_6136_7368# GND.t130 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X450 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t19 GND.t319 GND.t170 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X451 GND.t186 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar GND.t185 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X452 a_1480_8048# x0.t1 CLK0.t0 GND.t0 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X453 GND.t269 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar GND.t268 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X454 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar GND.t89 GND.t88 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X455 GND.t317 Dis1.t34 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar GND.t78 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X456 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t4 k0.t1 a_1480_8048# GND.t81 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X457 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar GND.t163 GND.t162 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X458 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t9 CLK2.t62 GND.t142 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X459 GND.t221 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t19 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t2 GND.t220 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X460 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar CLK2.t48 CLK2.t47 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X461 CLK1.t32 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X462 a_3040_5688# x2_bar.t1 CLK0.t30 GND.t57 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X463 CLK2.t98 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t10 a_10476_8048# GND.t295 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X464 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A CLK0.t3 CLK0.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X465 CLK3.t35 s2.t9 s2_bar.t3 CLK3.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X466 CLK3.t4 s0.t8 s0_bar.t2 CLK3.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X467 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t20 GND.t207 GND.t181 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X468 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t3 Dis1.t35 GND.t25 GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X469 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t20 a_4916_n1173# GND.t132 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X470 CLK1.t153 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t9 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t5 CLK1.t152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X471 a_1480_5688# x2.t1 CLK0.t6 GND.t55 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X472 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar CLK2.t44 CLK2.t43 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X473 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t9 CLK1.t110 CLK1.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X474 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t5 k2.t1 a_1480_5688# GND.t173 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X475 CLK1.t51 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A CLK1.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X476 CLK2.t42 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT CLK2.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X477 CLK2.t46 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT CLK2.t45 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X478 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar Dis2.t21 GND.t149 GND.t148 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X479 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t9 CLK2.t7 GND.t77 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X480 GND.t301 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t9 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t2 GND.t123 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X481 a_1180_5008# k3_bar.t1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t5 GND.t251 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X482 CLK3.t17 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A s0.t2 GND.t90 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X483 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B CLK1.t163 GND.t302 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
R0 CLK3.n414 CLK3.n413 407.048
R1 CLK3.n37 CLK3.n28 407.048
R2 CLK3.n345 CLK3.n344 407.048
R3 CLK3.n400 CLK3.n399 407.048
R4 CLK3.n270 CLK3.n269 407.048
R5 CLK3.n324 CLK3.n323 407.048
R6 CLK3.n199 CLK3.n198 407.048
R7 CLK3.n254 CLK3.n253 407.048
R8 CLK3.n72 CLK3.n3 400
R9 CLK3.n413 CLK3.n3 400
R10 CLK3.n38 CLK3.n37 400
R11 CLK3.n39 CLK3.n38 400
R12 CLK3.n346 CLK3.n345 400
R13 CLK3.n346 CLK3.n108 400
R14 CLK3.n354 CLK3.n108 400
R15 CLK3.n355 CLK3.n354 400
R16 CLK3.n389 CLK3.n388 400
R17 CLK3.n389 CLK3.n83 400
R18 CLK3.n398 CLK3.n83 400
R19 CLK3.n399 CLK3.n398 400
R20 CLK3.n281 CLK3.n280 400
R21 CLK3.n280 CLK3.n147 400
R22 CLK3.n271 CLK3.n147 400
R23 CLK3.n271 CLK3.n270 400
R24 CLK3.n323 CLK3.n322 400
R25 CLK3.n322 CLK3.n122 400
R26 CLK3.n314 CLK3.n122 400
R27 CLK3.n314 CLK3.n313 400
R28 CLK3.n200 CLK3.n199 400
R29 CLK3.n200 CLK3.n187 400
R30 CLK3.n208 CLK3.n187 400
R31 CLK3.n209 CLK3.n208 400
R32 CLK3.n243 CLK3.n242 400
R33 CLK3.n243 CLK3.n162 400
R34 CLK3.n252 CLK3.n162 400
R35 CLK3.n253 CLK3.n252 400
R36 CLK3.n72 CLK3.n71 366.379
R37 CLK3.n39 CLK3.n22 366.379
R38 CLK3.n356 CLK3.n355 366.379
R39 CLK3.n388 CLK3.n387 366.379
R40 CLK3.n282 CLK3.n281 366.379
R41 CLK3.n313 CLK3.n312 366.379
R42 CLK3.n210 CLK3.n209 366.379
R43 CLK3.n242 CLK3.n241 366.379
R44 CLK3.n48 CLK3.n22 131.034
R45 CLK3.n49 CLK3.n48 131.034
R46 CLK3.n51 CLK3.n50 131.034
R47 CLK3.n61 CLK3.n60 131.034
R48 CLK3.n70 CLK3.n10 131.034
R49 CLK3.n71 CLK3.n70 131.034
R50 CLK3.n356 CLK3.n102 131.034
R51 CLK3.n365 CLK3.n102 131.034
R52 CLK3.n368 CLK3.n366 131.034
R53 CLK3.n377 CLK3.n376 131.034
R54 CLK3.n378 CLK3.n90 131.034
R55 CLK3.n387 CLK3.n90 131.034
R56 CLK3.n312 CLK3.n128 131.034
R57 CLK3.n303 CLK3.n128 131.034
R58 CLK3.n302 CLK3.n301 131.034
R59 CLK3.n293 CLK3.n292 131.034
R60 CLK3.n291 CLK3.n141 131.034
R61 CLK3.n282 CLK3.n141 131.034
R62 CLK3.n210 CLK3.n181 131.034
R63 CLK3.n219 CLK3.n181 131.034
R64 CLK3.n222 CLK3.n220 131.034
R65 CLK3.n231 CLK3.n230 131.034
R66 CLK3.n232 CLK3.n169 131.034
R67 CLK3.n241 CLK3.n169 131.034
R68 CLK3.n59 CLK3.t36 122.844
R69 CLK3.t38 CLK3.n59 122.844
R70 CLK3.t13 CLK3.n367 122.844
R71 CLK3.n367 CLK3.t5 122.844
R72 CLK3.n140 CLK3.t21 122.844
R73 CLK3.t18 CLK3.n140 122.844
R74 CLK3.t31 CLK3.n221 122.844
R75 CLK3.n221 CLK3.t15 122.844
R76 CLK3.n51 CLK3.t3 106.465
R77 CLK3.n61 CLK3.t41 106.465
R78 CLK3.n366 CLK3.t0 106.465
R79 CLK3.t43 CLK3.n377 106.465
R80 CLK3.t34 CLK3.n302 106.465
R81 CLK3.n292 CLK3.t23 106.465
R82 CLK3.n220 CLK3.t29 106.465
R83 CLK3.t45 CLK3.n231 106.465
R84 CLK3.n36 CLK3.n29 96
R85 CLK3.n36 CLK3.n27 96
R86 CLK3.n40 CLK3.n27 96
R87 CLK3.n40 CLK3.n23 96
R88 CLK3.n47 CLK3.n23 96
R89 CLK3.n47 CLK3.n21 96
R90 CLK3.n52 CLK3.n21 96
R91 CLK3.n52 CLK3.n16 96
R92 CLK3.n58 CLK3.n16 96
R93 CLK3.n58 CLK3.n15 96
R94 CLK3.n62 CLK3.n15 96
R95 CLK3.n62 CLK3.n11 96
R96 CLK3.n69 CLK3.n11 96
R97 CLK3.n69 CLK3.n9 96
R98 CLK3.n73 CLK3.n9 96
R99 CLK3.n73 CLK3.n4 96
R100 CLK3.n412 CLK3.n4 96
R101 CLK3.n412 CLK3.n2 96
R102 CLK3.n343 CLK3.n113 96
R103 CLK3.n347 CLK3.n113 96
R104 CLK3.n347 CLK3.n109 96
R105 CLK3.n353 CLK3.n109 96
R106 CLK3.n353 CLK3.n107 96
R107 CLK3.n357 CLK3.n107 96
R108 CLK3.n357 CLK3.n103 96
R109 CLK3.n364 CLK3.n103 96
R110 CLK3.n364 CLK3.n101 96
R111 CLK3.n369 CLK3.n101 96
R112 CLK3.n369 CLK3.n96 96
R113 CLK3.n375 CLK3.n96 96
R114 CLK3.n375 CLK3.n95 96
R115 CLK3.n379 CLK3.n95 96
R116 CLK3.n379 CLK3.n91 96
R117 CLK3.n386 CLK3.n91 96
R118 CLK3.n386 CLK3.n89 96
R119 CLK3.n390 CLK3.n89 96
R120 CLK3.n390 CLK3.n84 96
R121 CLK3.n397 CLK3.n84 96
R122 CLK3.n397 CLK3.n82 96
R123 CLK3.n401 CLK3.n82 96
R124 CLK3.n325 CLK3.n121 96
R125 CLK3.n321 CLK3.n121 96
R126 CLK3.n321 CLK3.n123 96
R127 CLK3.n315 CLK3.n123 96
R128 CLK3.n315 CLK3.n127 96
R129 CLK3.n311 CLK3.n127 96
R130 CLK3.n311 CLK3.n129 96
R131 CLK3.n304 CLK3.n129 96
R132 CLK3.n304 CLK3.n133 96
R133 CLK3.n300 CLK3.n133 96
R134 CLK3.n300 CLK3.n134 96
R135 CLK3.n294 CLK3.n134 96
R136 CLK3.n294 CLK3.n139 96
R137 CLK3.n290 CLK3.n139 96
R138 CLK3.n290 CLK3.n142 96
R139 CLK3.n283 CLK3.n142 96
R140 CLK3.n283 CLK3.n146 96
R141 CLK3.n279 CLK3.n146 96
R142 CLK3.n279 CLK3.n148 96
R143 CLK3.n272 CLK3.n148 96
R144 CLK3.n272 CLK3.n153 96
R145 CLK3.n268 CLK3.n153 96
R146 CLK3.n197 CLK3.n192 96
R147 CLK3.n201 CLK3.n192 96
R148 CLK3.n201 CLK3.n188 96
R149 CLK3.n207 CLK3.n188 96
R150 CLK3.n207 CLK3.n186 96
R151 CLK3.n211 CLK3.n186 96
R152 CLK3.n211 CLK3.n182 96
R153 CLK3.n218 CLK3.n182 96
R154 CLK3.n218 CLK3.n180 96
R155 CLK3.n223 CLK3.n180 96
R156 CLK3.n223 CLK3.n175 96
R157 CLK3.n229 CLK3.n175 96
R158 CLK3.n229 CLK3.n174 96
R159 CLK3.n233 CLK3.n174 96
R160 CLK3.n233 CLK3.n170 96
R161 CLK3.n240 CLK3.n170 96
R162 CLK3.n240 CLK3.n168 96
R163 CLK3.n244 CLK3.n168 96
R164 CLK3.n244 CLK3.n163 96
R165 CLK3.n251 CLK3.n163 96
R166 CLK3.n251 CLK3.n161 96
R167 CLK3.n255 CLK3.n161 96
R168 CLK3.n31 CLK3.n28 85.261
R169 CLK3.n400 CLK3.n79 85.261
R170 CLK3.n324 CLK3.n118 85.261
R171 CLK3.n254 CLK3.n158 85.261
R172 CLK3.n415 CLK3.n414 85.261
R173 CLK3.n344 CLK3.n114 85.261
R174 CLK3.n269 CLK3.n154 85.261
R175 CLK3.n198 CLK3.n193 85.261
R176 CLK3.n307 CLK3.t35 44.338
R177 CLK3.n287 CLK3.t24 44.338
R178 CLK3.n44 CLK3.t4 44.338
R179 CLK3.n66 CLK3.t42 44.338
R180 CLK3.n382 CLK3.t44 44.337
R181 CLK3.n361 CLK3.t1 44.337
R182 CLK3.n236 CLK3.t46 44.337
R183 CLK3.n215 CLK3.t30 44.337
R184 CLK3.n407 CLK3.n406 44.163
R185 CLK3.n18 CLK3.t37 39.4
R186 CLK3.n18 CLK3.t39 39.4
R187 CLK3.n98 CLK3.t14 39.4
R188 CLK3.n98 CLK3.t6 39.4
R189 CLK3.n136 CLK3.t22 39.4
R190 CLK3.n136 CLK3.t19 39.4
R191 CLK3.n177 CLK3.t32 39.4
R192 CLK3.n177 CLK3.t16 39.4
R193 CLK3.n264 CLK3.t11 30.776
R194 CLK3.n32 CLK3.t27 30.776
R195 CLK3.n404 CLK3.t10 30.775
R196 CLK3.n258 CLK3.t25 30.775
R197 CLK3.n194 CLK3.t8 30.775
R198 CLK3.t3 CLK3.n49 24.568
R199 CLK3.t41 CLK3.n10 24.568
R200 CLK3.t0 CLK3.n365 24.568
R201 CLK3.n378 CLK3.t43 24.568
R202 CLK3.n303 CLK3.t34 24.568
R203 CLK3.t23 CLK3.n291 24.568
R204 CLK3.t29 CLK3.n219 24.568
R205 CLK3.n232 CLK3.t45 24.568
R206 CLK3.n86 CLK3.t12 24
R207 CLK3.n86 CLK3.t40 24
R208 CLK3.n331 CLK3.t7 24
R209 CLK3.n165 CLK3.t33 24
R210 CLK3.n165 CLK3.t20 24
R211 CLK3.n150 CLK3.t28 24
R212 CLK3.n150 CLK3.t9 24
R213 CLK3.n335 CLK3.t2 24
R214 CLK3.n6 CLK3.t26 24
R215 CLK3.n6 CLK3.t17 24
R216 CLK3.n31 CLK3.n30 12.8
R217 CLK3.n35 CLK3.n30 12.8
R218 CLK3.n35 CLK3.n26 12.8
R219 CLK3.n41 CLK3.n26 12.8
R220 CLK3.n41 CLK3.n24 12.8
R221 CLK3.n46 CLK3.n24 12.8
R222 CLK3.n46 CLK3.n20 12.8
R223 CLK3.n53 CLK3.n20 12.8
R224 CLK3.n53 CLK3.n17 12.8
R225 CLK3.n57 CLK3.n17 12.8
R226 CLK3.n57 CLK3.n14 12.8
R227 CLK3.n63 CLK3.n14 12.8
R228 CLK3.n63 CLK3.n12 12.8
R229 CLK3.n68 CLK3.n12 12.8
R230 CLK3.n68 CLK3.n8 12.8
R231 CLK3.n74 CLK3.n8 12.8
R232 CLK3.n74 CLK3.n5 12.8
R233 CLK3.n411 CLK3.n5 12.8
R234 CLK3.n411 CLK3.n1 12.8
R235 CLK3.n415 CLK3.n1 12.8
R236 CLK3.n342 CLK3.n114 12.8
R237 CLK3.n342 CLK3.n112 12.8
R238 CLK3.n348 CLK3.n112 12.8
R239 CLK3.n348 CLK3.n110 12.8
R240 CLK3.n352 CLK3.n110 12.8
R241 CLK3.n352 CLK3.n106 12.8
R242 CLK3.n358 CLK3.n106 12.8
R243 CLK3.n358 CLK3.n104 12.8
R244 CLK3.n363 CLK3.n104 12.8
R245 CLK3.n363 CLK3.n100 12.8
R246 CLK3.n370 CLK3.n100 12.8
R247 CLK3.n370 CLK3.n97 12.8
R248 CLK3.n374 CLK3.n97 12.8
R249 CLK3.n374 CLK3.n94 12.8
R250 CLK3.n380 CLK3.n94 12.8
R251 CLK3.n380 CLK3.n92 12.8
R252 CLK3.n385 CLK3.n92 12.8
R253 CLK3.n385 CLK3.n88 12.8
R254 CLK3.n391 CLK3.n88 12.8
R255 CLK3.n391 CLK3.n85 12.8
R256 CLK3.n396 CLK3.n85 12.8
R257 CLK3.n396 CLK3.n81 12.8
R258 CLK3.n402 CLK3.n81 12.8
R259 CLK3.n402 CLK3.n79 12.8
R260 CLK3.n330 CLK3.n117 12.8
R261 CLK3.n326 CLK3.n118 12.8
R262 CLK3.n326 CLK3.n120 12.8
R263 CLK3.n320 CLK3.n120 12.8
R264 CLK3.n320 CLK3.n124 12.8
R265 CLK3.n316 CLK3.n124 12.8
R266 CLK3.n316 CLK3.n126 12.8
R267 CLK3.n310 CLK3.n126 12.8
R268 CLK3.n310 CLK3.n130 12.8
R269 CLK3.n305 CLK3.n130 12.8
R270 CLK3.n305 CLK3.n132 12.8
R271 CLK3.n299 CLK3.n132 12.8
R272 CLK3.n299 CLK3.n135 12.8
R273 CLK3.n295 CLK3.n135 12.8
R274 CLK3.n295 CLK3.n138 12.8
R275 CLK3.n289 CLK3.n138 12.8
R276 CLK3.n289 CLK3.n143 12.8
R277 CLK3.n284 CLK3.n143 12.8
R278 CLK3.n284 CLK3.n145 12.8
R279 CLK3.n278 CLK3.n145 12.8
R280 CLK3.n278 CLK3.n149 12.8
R281 CLK3.n273 CLK3.n149 12.8
R282 CLK3.n273 CLK3.n152 12.8
R283 CLK3.n196 CLK3.n193 12.8
R284 CLK3.n196 CLK3.n191 12.8
R285 CLK3.n202 CLK3.n191 12.8
R286 CLK3.n202 CLK3.n189 12.8
R287 CLK3.n206 CLK3.n189 12.8
R288 CLK3.n206 CLK3.n185 12.8
R289 CLK3.n212 CLK3.n185 12.8
R290 CLK3.n212 CLK3.n183 12.8
R291 CLK3.n217 CLK3.n183 12.8
R292 CLK3.n217 CLK3.n179 12.8
R293 CLK3.n224 CLK3.n179 12.8
R294 CLK3.n224 CLK3.n176 12.8
R295 CLK3.n228 CLK3.n176 12.8
R296 CLK3.n228 CLK3.n173 12.8
R297 CLK3.n234 CLK3.n173 12.8
R298 CLK3.n234 CLK3.n171 12.8
R299 CLK3.n239 CLK3.n171 12.8
R300 CLK3.n239 CLK3.n167 12.8
R301 CLK3.n245 CLK3.n167 12.8
R302 CLK3.n245 CLK3.n164 12.8
R303 CLK3.n250 CLK3.n164 12.8
R304 CLK3.n250 CLK3.n160 12.8
R305 CLK3.n256 CLK3.n160 12.8
R306 CLK3.n256 CLK3.n158 12.8
R307 CLK3.n337 CLK3.n336 12.8
R308 CLK3.n155 CLK3.n152 12.32
R309 CLK3.n156 CLK3.n154 10.56
R310 EESPFAL_Sbox_0/CLK3 CLK3.n416 9.779
R311 CLK3.n265 CLK3.n156 9.3
R312 CLK3.n267 CLK3.n266 9.3
R313 CLK3.n412 CLK3.n411 8.855
R314 CLK3.n331 CLK3.n330 8.855
R315 CLK3.n153 CLK3.n152 8.855
R316 CLK3.n197 CLK3.n196 8.855
R317 CLK3.n192 CLK3.n191 8.855
R318 CLK3.n199 CLK3.n192 8.855
R319 CLK3.n202 CLK3.n201 8.855
R320 CLK3.n201 CLK3.n200 8.855
R321 CLK3.n189 CLK3.n188 8.855
R322 CLK3.n188 CLK3.n187 8.855
R323 CLK3.n207 CLK3.n206 8.855
R324 CLK3.n208 CLK3.n207 8.855
R325 CLK3.n186 CLK3.n185 8.855
R326 CLK3.n209 CLK3.n186 8.855
R327 CLK3.n212 CLK3.n211 8.855
R328 CLK3.n211 CLK3.n210 8.855
R329 CLK3.n183 CLK3.n182 8.855
R330 CLK3.n182 CLK3.n181 8.855
R331 CLK3.n218 CLK3.n217 8.855
R332 CLK3.n219 CLK3.n218 8.855
R333 CLK3.n180 CLK3.n179 8.855
R334 CLK3.n220 CLK3.n180 8.855
R335 CLK3.n224 CLK3.n223 8.855
R336 CLK3.n223 CLK3.n222 8.855
R337 CLK3.n176 CLK3.n175 8.855
R338 CLK3.n221 CLK3.n175 8.855
R339 CLK3.n229 CLK3.n228 8.855
R340 CLK3.n230 CLK3.n229 8.855
R341 CLK3.n174 CLK3.n173 8.855
R342 CLK3.n231 CLK3.n174 8.855
R343 CLK3.n234 CLK3.n233 8.855
R344 CLK3.n233 CLK3.n232 8.855
R345 CLK3.n171 CLK3.n170 8.855
R346 CLK3.n170 CLK3.n169 8.855
R347 CLK3.n240 CLK3.n239 8.855
R348 CLK3.n241 CLK3.n240 8.855
R349 CLK3.n168 CLK3.n167 8.855
R350 CLK3.n242 CLK3.n168 8.855
R351 CLK3.n245 CLK3.n244 8.855
R352 CLK3.n244 CLK3.n243 8.855
R353 CLK3.n164 CLK3.n163 8.855
R354 CLK3.n163 CLK3.n162 8.855
R355 CLK3.n251 CLK3.n250 8.855
R356 CLK3.n252 CLK3.n251 8.855
R357 CLK3.n161 CLK3.n160 8.855
R358 CLK3.n253 CLK3.n161 8.855
R359 CLK3.n256 CLK3.n255 8.855
R360 CLK3.n326 CLK3.n325 8.855
R361 CLK3.n121 CLK3.n120 8.855
R362 CLK3.n323 CLK3.n121 8.855
R363 CLK3.n321 CLK3.n320 8.855
R364 CLK3.n322 CLK3.n321 8.855
R365 CLK3.n124 CLK3.n123 8.855
R366 CLK3.n123 CLK3.n122 8.855
R367 CLK3.n316 CLK3.n315 8.855
R368 CLK3.n315 CLK3.n314 8.855
R369 CLK3.n127 CLK3.n126 8.855
R370 CLK3.n313 CLK3.n127 8.855
R371 CLK3.n311 CLK3.n310 8.855
R372 CLK3.n312 CLK3.n311 8.855
R373 CLK3.n130 CLK3.n129 8.855
R374 CLK3.n129 CLK3.n128 8.855
R375 CLK3.n305 CLK3.n304 8.855
R376 CLK3.n304 CLK3.n303 8.855
R377 CLK3.n133 CLK3.n132 8.855
R378 CLK3.n302 CLK3.n133 8.855
R379 CLK3.n300 CLK3.n299 8.855
R380 CLK3.n301 CLK3.n300 8.855
R381 CLK3.n135 CLK3.n134 8.855
R382 CLK3.n140 CLK3.n134 8.855
R383 CLK3.n295 CLK3.n294 8.855
R384 CLK3.n294 CLK3.n293 8.855
R385 CLK3.n139 CLK3.n138 8.855
R386 CLK3.n292 CLK3.n139 8.855
R387 CLK3.n290 CLK3.n289 8.855
R388 CLK3.n291 CLK3.n290 8.855
R389 CLK3.n143 CLK3.n142 8.855
R390 CLK3.n142 CLK3.n141 8.855
R391 CLK3.n284 CLK3.n283 8.855
R392 CLK3.n283 CLK3.n282 8.855
R393 CLK3.n146 CLK3.n145 8.855
R394 CLK3.n281 CLK3.n146 8.855
R395 CLK3.n279 CLK3.n278 8.855
R396 CLK3.n280 CLK3.n279 8.855
R397 CLK3.n149 CLK3.n148 8.855
R398 CLK3.n148 CLK3.n147 8.855
R399 CLK3.n273 CLK3.n272 8.855
R400 CLK3.n272 CLK3.n271 8.855
R401 CLK3.n270 CLK3.n153 8.855
R402 CLK3.n268 CLK3.n267 8.855
R403 CLK3.n336 CLK3.n335 8.855
R404 CLK3.n343 CLK3.n342 8.855
R405 CLK3.n113 CLK3.n112 8.855
R406 CLK3.n345 CLK3.n113 8.855
R407 CLK3.n348 CLK3.n347 8.855
R408 CLK3.n347 CLK3.n346 8.855
R409 CLK3.n110 CLK3.n109 8.855
R410 CLK3.n109 CLK3.n108 8.855
R411 CLK3.n353 CLK3.n352 8.855
R412 CLK3.n354 CLK3.n353 8.855
R413 CLK3.n107 CLK3.n106 8.855
R414 CLK3.n355 CLK3.n107 8.855
R415 CLK3.n358 CLK3.n357 8.855
R416 CLK3.n357 CLK3.n356 8.855
R417 CLK3.n104 CLK3.n103 8.855
R418 CLK3.n103 CLK3.n102 8.855
R419 CLK3.n364 CLK3.n363 8.855
R420 CLK3.n365 CLK3.n364 8.855
R421 CLK3.n101 CLK3.n100 8.855
R422 CLK3.n366 CLK3.n101 8.855
R423 CLK3.n370 CLK3.n369 8.855
R424 CLK3.n369 CLK3.n368 8.855
R425 CLK3.n97 CLK3.n96 8.855
R426 CLK3.n367 CLK3.n96 8.855
R427 CLK3.n375 CLK3.n374 8.855
R428 CLK3.n376 CLK3.n375 8.855
R429 CLK3.n95 CLK3.n94 8.855
R430 CLK3.n377 CLK3.n95 8.855
R431 CLK3.n380 CLK3.n379 8.855
R432 CLK3.n379 CLK3.n378 8.855
R433 CLK3.n92 CLK3.n91 8.855
R434 CLK3.n91 CLK3.n90 8.855
R435 CLK3.n386 CLK3.n385 8.855
R436 CLK3.n387 CLK3.n386 8.855
R437 CLK3.n89 CLK3.n88 8.855
R438 CLK3.n388 CLK3.n89 8.855
R439 CLK3.n391 CLK3.n390 8.855
R440 CLK3.n390 CLK3.n389 8.855
R441 CLK3.n85 CLK3.n84 8.855
R442 CLK3.n84 CLK3.n83 8.855
R443 CLK3.n397 CLK3.n396 8.855
R444 CLK3.n398 CLK3.n397 8.855
R445 CLK3.n82 CLK3.n81 8.855
R446 CLK3.n399 CLK3.n82 8.855
R447 CLK3.n402 CLK3.n401 8.855
R448 CLK3.n30 CLK3.n29 8.855
R449 CLK3.n36 CLK3.n35 8.855
R450 CLK3.n37 CLK3.n36 8.855
R451 CLK3.n27 CLK3.n26 8.855
R452 CLK3.n38 CLK3.n27 8.855
R453 CLK3.n41 CLK3.n40 8.855
R454 CLK3.n40 CLK3.n39 8.855
R455 CLK3.n24 CLK3.n23 8.855
R456 CLK3.n23 CLK3.n22 8.855
R457 CLK3.n47 CLK3.n46 8.855
R458 CLK3.n48 CLK3.n47 8.855
R459 CLK3.n21 CLK3.n20 8.855
R460 CLK3.n49 CLK3.n21 8.855
R461 CLK3.n53 CLK3.n52 8.855
R462 CLK3.n52 CLK3.n51 8.855
R463 CLK3.n17 CLK3.n16 8.855
R464 CLK3.n50 CLK3.n16 8.855
R465 CLK3.n58 CLK3.n57 8.855
R466 CLK3.n59 CLK3.n58 8.855
R467 CLK3.n15 CLK3.n14 8.855
R468 CLK3.n60 CLK3.n15 8.855
R469 CLK3.n63 CLK3.n62 8.855
R470 CLK3.n62 CLK3.n61 8.855
R471 CLK3.n12 CLK3.n11 8.855
R472 CLK3.n11 CLK3.n10 8.855
R473 CLK3.n69 CLK3.n68 8.855
R474 CLK3.n70 CLK3.n69 8.855
R475 CLK3.n9 CLK3.n8 8.855
R476 CLK3.n71 CLK3.n9 8.855
R477 CLK3.n74 CLK3.n73 8.855
R478 CLK3.n73 CLK3.n72 8.855
R479 CLK3.n5 CLK3.n4 8.855
R480 CLK3.n4 CLK3.n3 8.855
R481 CLK3.n413 CLK3.n412 8.855
R482 CLK3.n2 CLK3.n1 8.855
R483 CLK3.n339 CLK3.n115 8.365
R484 CLK3.n50 CLK3.t36 8.189
R485 CLK3.n60 CLK3.t38 8.189
R486 CLK3.n368 CLK3.t13 8.189
R487 CLK3.n376 CLK3.t5 8.189
R488 CLK3.n301 CLK3.t21 8.189
R489 CLK3.n293 CLK3.t18 8.189
R490 CLK3.n222 CLK3.t31 8.189
R491 CLK3.n230 CLK3.t15 8.189
R492 CLK3.n393 CLK3.n86 6.776
R493 CLK3.n247 CLK3.n165 6.776
R494 CLK3.n276 CLK3.n150 6.776
R495 CLK3.n77 CLK3.n6 6.776
R496 CLK3.n333 CLK3.n332 6.754
R497 EESPFAL_Sbox_0/EESPFAL_s3_0/CLK3 CLK3.n259 5.161
R498 CLK3.n406 CLK3.n405 4.966
R499 CLK3.n56 CLK3.n18 4.938
R500 CLK3.n372 CLK3.n98 4.938
R501 CLK3.n297 CLK3.n136 4.938
R502 CLK3.n226 CLK3.n177 4.938
R503 CLK3.n194 CLK3.n193 4.687
R504 CLK3.n328 CLK3.n118 4.687
R505 CLK3.n264 CLK3.n154 4.687
R506 CLK3.n340 CLK3.n114 4.687
R507 CLK3.n32 CLK3.n31 4.675
R508 CLK3.n196 CLK3.n195 4.65
R509 CLK3.n191 CLK3.n190 4.65
R510 CLK3.n203 CLK3.n202 4.65
R511 CLK3.n204 CLK3.n189 4.65
R512 CLK3.n206 CLK3.n205 4.65
R513 CLK3.n185 CLK3.n184 4.65
R514 CLK3.n213 CLK3.n212 4.65
R515 CLK3.n214 CLK3.n183 4.65
R516 CLK3.n217 CLK3.n216 4.65
R517 CLK3.n179 CLK3.n178 4.65
R518 CLK3.n225 CLK3.n224 4.65
R519 CLK3.n226 CLK3.n176 4.65
R520 CLK3.n228 CLK3.n227 4.65
R521 CLK3.n173 CLK3.n172 4.65
R522 CLK3.n235 CLK3.n234 4.65
R523 CLK3.n237 CLK3.n171 4.65
R524 CLK3.n239 CLK3.n238 4.65
R525 CLK3.n167 CLK3.n166 4.65
R526 CLK3.n246 CLK3.n245 4.65
R527 CLK3.n248 CLK3.n164 4.65
R528 CLK3.n250 CLK3.n249 4.65
R529 CLK3.n160 CLK3.n159 4.65
R530 CLK3.n257 CLK3.n256 4.65
R531 CLK3.n152 CLK3.n151 4.65
R532 CLK3.n327 CLK3.n326 4.65
R533 CLK3.n120 CLK3.n119 4.65
R534 CLK3.n320 CLK3.n319 4.65
R535 CLK3.n318 CLK3.n124 4.65
R536 CLK3.n317 CLK3.n316 4.65
R537 CLK3.n126 CLK3.n125 4.65
R538 CLK3.n310 CLK3.n309 4.65
R539 CLK3.n308 CLK3.n130 4.65
R540 CLK3.n306 CLK3.n305 4.65
R541 CLK3.n132 CLK3.n131 4.65
R542 CLK3.n299 CLK3.n298 4.65
R543 CLK3.n297 CLK3.n135 4.65
R544 CLK3.n296 CLK3.n295 4.65
R545 CLK3.n138 CLK3.n137 4.65
R546 CLK3.n289 CLK3.n288 4.65
R547 CLK3.n286 CLK3.n143 4.65
R548 CLK3.n285 CLK3.n284 4.65
R549 CLK3.n145 CLK3.n144 4.65
R550 CLK3.n278 CLK3.n277 4.65
R551 CLK3.n275 CLK3.n149 4.65
R552 CLK3.n274 CLK3.n273 4.65
R553 CLK3.n117 CLK3.n116 4.65
R554 CLK3.n330 CLK3.n329 4.65
R555 CLK3.n338 CLK3.n337 4.65
R556 CLK3.n342 CLK3.n341 4.65
R557 CLK3.n112 CLK3.n111 4.65
R558 CLK3.n349 CLK3.n348 4.65
R559 CLK3.n350 CLK3.n110 4.65
R560 CLK3.n352 CLK3.n351 4.65
R561 CLK3.n106 CLK3.n105 4.65
R562 CLK3.n359 CLK3.n358 4.65
R563 CLK3.n360 CLK3.n104 4.65
R564 CLK3.n363 CLK3.n362 4.65
R565 CLK3.n100 CLK3.n99 4.65
R566 CLK3.n371 CLK3.n370 4.65
R567 CLK3.n372 CLK3.n97 4.65
R568 CLK3.n374 CLK3.n373 4.65
R569 CLK3.n94 CLK3.n93 4.65
R570 CLK3.n381 CLK3.n380 4.65
R571 CLK3.n383 CLK3.n92 4.65
R572 CLK3.n385 CLK3.n384 4.65
R573 CLK3.n88 CLK3.n87 4.65
R574 CLK3.n392 CLK3.n391 4.65
R575 CLK3.n394 CLK3.n85 4.65
R576 CLK3.n396 CLK3.n395 4.65
R577 CLK3.n81 CLK3.n80 4.65
R578 CLK3.n403 CLK3.n402 4.65
R579 CLK3.n411 CLK3.n410 4.65
R580 CLK3.n33 CLK3.n30 4.65
R581 CLK3.n35 CLK3.n34 4.65
R582 CLK3.n26 CLK3.n25 4.65
R583 CLK3.n42 CLK3.n41 4.65
R584 CLK3.n43 CLK3.n24 4.65
R585 CLK3.n46 CLK3.n45 4.65
R586 CLK3.n20 CLK3.n19 4.65
R587 CLK3.n54 CLK3.n53 4.65
R588 CLK3.n55 CLK3.n17 4.65
R589 CLK3.n57 CLK3.n56 4.65
R590 CLK3.n14 CLK3.n13 4.65
R591 CLK3.n64 CLK3.n63 4.65
R592 CLK3.n65 CLK3.n12 4.65
R593 CLK3.n68 CLK3.n67 4.65
R594 CLK3.n8 CLK3.n7 4.65
R595 CLK3.n75 CLK3.n74 4.65
R596 CLK3.n76 CLK3.n5 4.65
R597 CLK3.n416 CLK3.n415 4.65
R598 CLK3.n262 CLK3.n261 4.5
R599 CLK3.n263 CLK3.n262 4.5
R600 CLK3.n263 CLK3.n155 4.5
R601 CLK3.n408 CLK3.n0 4.5
R602 CLK3.n409 CLK3.n408 4.5
R603 CLK3.n260 EESPFAL_Sbox_0/EESPFAL_s2_0/CLK3 4.449
R604 CLK3.n334 CLK3.n333 3.724
R605 CLK3.n332 CLK3.n117 3.715
R606 CLK3.n337 CLK3.n115 3.715
R607 CLK3.n336 CLK3.n334 3.039
R608 CLK3.n259 CLK3.n158 3.038
R609 CLK3.n405 CLK3.n79 3.038
R610 CLK3.n78 CLK3.n1 3.033
R611 CLK3.n332 CLK3.n331 2.57
R612 CLK3.n335 CLK3.n115 2.57
R613 CLK3.n267 CLK3.n156 2.24
R614 CLK3.n329 CLK3.n328 2.203
R615 CLK3.n340 CLK3.n339 2.203
R616 CLK3.n255 CLK3.n254 1.655
R617 CLK3.n325 CLK3.n324 1.655
R618 CLK3.n401 CLK3.n400 1.655
R619 CLK3.n29 CLK3.n28 1.655
R620 CLK3.n344 CLK3.n343 1.655
R621 CLK3.n198 CLK3.n197 1.655
R622 CLK3.n269 CLK3.n268 1.655
R623 CLK3.n414 CLK3.n2 1.655
R624 CLK3.n260 CLK3.n157 1.497
R625 CLK3.n407 CLK3.n78 1.121
R626 EESPFAL_Sbox_0/EESPFAL_s2_0/CLK3 EESPFAL_Sbox_0/EESPFAL_s3_0/CLK3 1.018
R627 CLK3.n267 CLK3.n155 0.48
R628 CLK3.n406 EESPFAL_Sbox_0/EESPFAL_s1_0/CLK3 0.195
R629 CLK3.n329 CLK3.n116 0.125
R630 CLK3.n339 CLK3.n338 0.125
R631 CLK3.n333 CLK3.n116 0.119
R632 CLK3.n338 CLK3.n334 0.119
R633 CLK3.n195 CLK3.n190 0.1
R634 CLK3.n203 CLK3.n190 0.1
R635 CLK3.n204 CLK3.n203 0.1
R636 CLK3.n205 CLK3.n204 0.1
R637 CLK3.n205 CLK3.n184 0.1
R638 CLK3.n213 CLK3.n184 0.1
R639 CLK3.n214 CLK3.n213 0.1
R640 CLK3.n216 CLK3.n178 0.1
R641 CLK3.n225 CLK3.n178 0.1
R642 CLK3.n226 CLK3.n225 0.1
R643 CLK3.n227 CLK3.n172 0.1
R644 CLK3.n235 CLK3.n172 0.1
R645 CLK3.n238 CLK3.n237 0.1
R646 CLK3.n238 CLK3.n166 0.1
R647 CLK3.n246 CLK3.n166 0.1
R648 CLK3.n249 CLK3.n248 0.1
R649 CLK3.n249 CLK3.n159 0.1
R650 CLK3.n257 CLK3.n159 0.1
R651 CLK3.n327 CLK3.n119 0.1
R652 CLK3.n319 CLK3.n119 0.1
R653 CLK3.n319 CLK3.n318 0.1
R654 CLK3.n318 CLK3.n317 0.1
R655 CLK3.n317 CLK3.n125 0.1
R656 CLK3.n309 CLK3.n125 0.1
R657 CLK3.n309 CLK3.n308 0.1
R658 CLK3.n306 CLK3.n131 0.1
R659 CLK3.n298 CLK3.n131 0.1
R660 CLK3.n298 CLK3.n297 0.1
R661 CLK3.n296 CLK3.n137 0.1
R662 CLK3.n288 CLK3.n137 0.1
R663 CLK3.n286 CLK3.n285 0.1
R664 CLK3.n285 CLK3.n144 0.1
R665 CLK3.n277 CLK3.n144 0.1
R666 CLK3.n275 CLK3.n274 0.1
R667 CLK3.n274 CLK3.n151 0.1
R668 CLK3.n341 CLK3.n111 0.1
R669 CLK3.n349 CLK3.n111 0.1
R670 CLK3.n350 CLK3.n349 0.1
R671 CLK3.n351 CLK3.n350 0.1
R672 CLK3.n351 CLK3.n105 0.1
R673 CLK3.n359 CLK3.n105 0.1
R674 CLK3.n360 CLK3.n359 0.1
R675 CLK3.n362 CLK3.n99 0.1
R676 CLK3.n371 CLK3.n99 0.1
R677 CLK3.n372 CLK3.n371 0.1
R678 CLK3.n373 CLK3.n93 0.1
R679 CLK3.n381 CLK3.n93 0.1
R680 CLK3.n384 CLK3.n383 0.1
R681 CLK3.n384 CLK3.n87 0.1
R682 CLK3.n392 CLK3.n87 0.1
R683 CLK3.n395 CLK3.n394 0.1
R684 CLK3.n395 CLK3.n80 0.1
R685 CLK3.n403 CLK3.n80 0.1
R686 CLK3.n34 CLK3.n33 0.1
R687 CLK3.n34 CLK3.n25 0.1
R688 CLK3.n42 CLK3.n25 0.1
R689 CLK3.n43 CLK3.n42 0.1
R690 CLK3.n45 CLK3.n43 0.1
R691 CLK3.n54 CLK3.n19 0.1
R692 CLK3.n55 CLK3.n54 0.1
R693 CLK3.n56 CLK3.n55 0.1
R694 CLK3.n64 CLK3.n13 0.1
R695 CLK3.n65 CLK3.n64 0.1
R696 CLK3.n67 CLK3.n7 0.1
R697 CLK3.n75 CLK3.n7 0.1
R698 CLK3.n76 CLK3.n75 0.1
R699 CLK3.n247 CLK3.n246 0.087
R700 CLK3.n277 CLK3.n276 0.087
R701 CLK3.n393 CLK3.n392 0.087
R702 CLK3.n77 CLK3.n76 0.087
R703 CLK3.n216 CLK3.n215 0.075
R704 CLK3.n227 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/CLK 0.075
R705 CLK3.n236 CLK3.n235 0.075
R706 CLK3.n307 CLK3.n306 0.075
R707 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/CLK CLK3.n296 0.075
R708 CLK3.n288 CLK3.n287 0.075
R709 CLK3.n362 CLK3.n361 0.075
R710 CLK3.n373 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/CLK 0.075
R711 CLK3.n382 CLK3.n381 0.075
R712 CLK3.n33 CLK3.n32 0.075
R713 CLK3.n44 CLK3.n19 0.075
R714 CLK3 CLK3.n13 0.075
R715 CLK3.n66 CLK3.n65 0.075
R716 CLK3.n410 CLK3.n409 0.073
R717 CLK3.n416 CLK3.n0 0.072
R718 CLK3.n261 CLK3.n151 0.063
R719 CLK3.n195 CLK3.n194 0.062
R720 CLK3.n258 CLK3.n257 0.062
R721 CLK3.n328 CLK3.n327 0.062
R722 CLK3.n341 CLK3.n340 0.062
R723 CLK3.n404 CLK3.n403 0.062
R724 EESPFAL_Sbox_0/EESPFAL_s0_0/CLK3 EESPFAL_Sbox_0/CLK3 0.046
R725 CLK3.n265 CLK3.n264 0.045
R726 CLK3.n259 CLK3.n258 0.034
R727 CLK3.n405 CLK3.n404 0.034
R728 CLK3.n78 CLK3.n0 0.027
R729 CLK3.n409 CLK3.n78 0.026
R730 CLK3.n215 CLK3.n214 0.025
R731 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/CLK CLK3.n226 0.025
R732 CLK3.n237 CLK3.n236 0.025
R733 CLK3.n308 CLK3.n307 0.025
R734 CLK3.n297 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/CLK 0.025
R735 CLK3.n287 CLK3.n286 0.025
R736 CLK3.n361 CLK3.n360 0.025
R737 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/CLK CLK3.n372 0.025
R738 CLK3.n383 CLK3.n382 0.025
R739 CLK3.n45 CLK3.n44 0.025
R740 CLK3.n56 CLK3 0.025
R741 CLK3.n67 CLK3.n66 0.025
R742 CLK3.n266 CLK3.n265 0.017
R743 CLK3.n261 CLK3.n157 0.016
R744 CLK3.n263 CLK3.n157 0.016
R745 CLK3.n262 CLK3.n260 0.012
R746 CLK3.n248 CLK3.n247 0.012
R747 CLK3.n276 CLK3.n275 0.012
R748 CLK3.n394 CLK3.n393 0.012
R749 CLK3.n410 CLK3.n77 0.012
R750 CLK3.n408 CLK3.n407 0.01
R751 CLK3.n266 CLK3.n263 0.003
R752 s0.t7 s0.t8 819.4
R753 s0.n2 s0.t7 514.133
R754 s0.n2 s0.t6 305.266
R755 s0.n3 s0.n1 166.734
R756 s0.n4 s0.n3 99.2
R757 s0.n5 s0.n4 99.2
R758 s0.n4 s0.t3 97.937
R759 s0.n5 s0.t2 91.537
R760 s0 s0.n2 79.2
R761 s0.n3 s0.n0 73.937
R762 s0.n3 s0 54.4
R763 s0.n1 s0.t4 39.4
R764 s0.n1 s0.t5 39.4
R765 s0.n0 s0.t1 24
R766 s0.n0 s0.t0 24
R767 EESPFAL_Sbox_0/s0 s0.n5 12.406
R768 EESPFAL_Sbox_0/s0 s0 0.081
R769 s0 EESPFAL_Sbox_0/EESPFAL_s0_0/s0 0.003
R770 GND.n1909 GND.n1908 5407.82
R771 GND.n1590 GND.n1589 4632.06
R772 GND.t209 GND.t322 3300
R773 GND.t353 GND.t310 3300
R774 GND.n1760 GND.t160 2526.31
R775 GND.n1589 GND.t93 2526.31
R776 GND.t322 GND.t155 1500
R777 GND.t339 GND.t209 1500
R778 GND.t105 GND.t339 1500
R779 GND.t310 GND.t152 1500
R780 GND.t152 GND.t166 1500
R781 GND.n1569 GND.t353 1150
R782 GND.n1908 GND.t357 1081.56
R783 GND.n1910 GND.n1909 1042.1
R784 GND.n505 GND.n504 594.594
R785 GND.n573 GND.n572 594.594
R786 GND.n1433 GND.n1432 594.594
R787 GND.n1435 GND.n1433 594.594
R788 GND.n1435 GND.n1434 594.594
R789 GND.n1445 GND.n1444 594.594
R790 GND.n1455 GND.n1314 594.594
R791 GND.n1457 GND.n1456 594.594
R792 GND.n1457 GND.n1308 594.594
R793 GND.n1465 GND.n1308 594.594
R794 GND.n1368 GND.n1367 594.594
R795 GND.n1370 GND.n1369 594.594
R796 GND.n1379 GND.n1378 594.594
R797 GND.n1381 GND.n1379 594.594
R798 GND.n1381 GND.n1380 594.594
R799 GND.n1391 GND.n1390 594.594
R800 GND.n1401 GND.n1343 594.594
R801 GND.n1403 GND.n1402 594.594
R802 GND.n1403 GND.n1337 594.594
R803 GND.n1411 GND.n1337 594.594
R804 GND.n1413 GND.n1412 594.594
R805 GND.n1421 GND.n1331 594.594
R806 GND.n1477 GND.n1476 594.594
R807 GND.n1479 GND.n1478 594.594
R808 GND.n1488 GND.n1487 594.594
R809 GND.n1490 GND.n1488 594.594
R810 GND.n1490 GND.n1489 594.594
R811 GND.n1500 GND.n1499 594.594
R812 GND.n1510 GND.n1286 594.594
R813 GND.n1512 GND.n1511 594.594
R814 GND.n1512 GND.n1280 594.594
R815 GND.n1520 GND.n1280 594.594
R816 GND.n1522 GND.n1521 594.594
R817 GND.n1531 GND.n1274 594.594
R818 GND.n1432 GND.t299 557.432
R819 GND.n1446 GND.t72 557.432
R820 GND.n1446 GND.t112 557.432
R821 GND.t270 GND.n1465 557.432
R822 GND.n1378 GND.t121 557.432
R823 GND.n1392 GND.t94 557.432
R824 GND.n1392 GND.t234 557.432
R825 GND.t323 GND.n1411 557.432
R826 GND.n1487 GND.t306 557.432
R827 GND.n1501 GND.t271 557.432
R828 GND.n1501 GND.t297 557.432
R829 GND.t347 GND.n1520 557.432
R830 GND.n1444 GND.t237 483.108
R831 GND.t51 GND.n1455 483.108
R832 GND.n1370 GND.t206 483.108
R833 GND.n1390 GND.t341 483.108
R834 GND.t355 GND.n1401 483.108
R835 GND.n1413 GND.t273 483.108
R836 GND.n1479 GND.t135 483.108
R837 GND.n1499 GND.t17 483.108
R838 GND.t278 GND.n1510 483.108
R839 GND.n1522 GND.t69 483.108
R840 GND.n1367 GND.t111 408.783
R841 GND.t283 GND.n1421 408.783
R842 GND.n1476 GND.t114 408.783
R843 GND.t59 GND.n1531 408.783
R844 GND.n1569 GND.t105 350
R845 GND.n455 GND.n454 341.085
R846 GND.n456 GND.n357 341.085
R847 GND.n465 GND.n357 341.085
R848 GND.n466 GND.n465 341.085
R849 GND.n468 GND.n467 341.085
R850 GND.n478 GND.n477 341.085
R851 GND.n487 GND.n344 341.085
R852 GND.n488 GND.n487 341.085
R853 GND.n489 GND.n488 341.085
R854 GND.n497 GND.n338 341.085
R855 GND.n401 GND.n400 341.085
R856 GND.n402 GND.n387 341.085
R857 GND.n411 GND.n387 341.085
R858 GND.n412 GND.n411 341.085
R859 GND.n414 GND.n413 341.085
R860 GND.n424 GND.n423 341.085
R861 GND.n433 GND.n374 341.085
R862 GND.n434 GND.n433 341.085
R863 GND.n435 GND.n434 341.085
R864 GND.n443 GND.n368 341.085
R865 GND.n513 GND.n329 341.085
R866 GND.n515 GND.n514 341.085
R867 GND.n524 GND.n323 341.085
R868 GND.n525 GND.n524 341.085
R869 GND.n526 GND.n525 341.085
R870 GND.n537 GND.n317 341.085
R871 GND.n540 GND.n539 341.085
R872 GND.n550 GND.n549 341.085
R873 GND.n552 GND.n550 341.085
R874 GND.n552 GND.n551 341.085
R875 GND.n561 GND.n560 341.085
R876 GND.n563 GND.n562 341.085
R877 GND.n581 GND.n580 341.085
R878 GND.n589 GND.n295 341.085
R879 GND.n591 GND.n590 341.085
R880 GND.n600 GND.n289 341.085
R881 GND.n601 GND.n600 341.085
R882 GND.n602 GND.n601 341.085
R883 GND.n613 GND.n283 341.085
R884 GND.n616 GND.n615 341.085
R885 GND.n626 GND.n625 341.085
R886 GND.n628 GND.n626 341.085
R887 GND.n628 GND.n627 341.085
R888 GND.n637 GND.n636 341.085
R889 GND.n639 GND.n638 341.085
R890 GND.n648 GND.n647 341.085
R891 GND.n1161 GND.n1160 341.085
R892 GND.n1163 GND.n1161 341.085
R893 GND.n1163 GND.n1162 341.085
R894 GND.n1173 GND.n1172 341.085
R895 GND.n1183 GND.n1056 341.085
R896 GND.n1185 GND.n1184 341.085
R897 GND.n1185 GND.n1050 341.085
R898 GND.n1193 GND.n1050 341.085
R899 GND.n1107 GND.n1106 341.085
R900 GND.n1108 GND.n1093 341.085
R901 GND.n1117 GND.n1093 341.085
R902 GND.n1118 GND.n1117 341.085
R903 GND.n1120 GND.n1119 341.085
R904 GND.n1130 GND.n1129 341.085
R905 GND.n1139 GND.n1080 341.085
R906 GND.n1140 GND.n1139 341.085
R907 GND.n1141 GND.n1140 341.085
R908 GND.n1149 GND.n1074 341.085
R909 GND.n1201 GND.n1200 341.085
R910 GND.n1209 GND.n1041 341.085
R911 GND.n1211 GND.n1210 341.085
R912 GND.n1220 GND.n1035 341.085
R913 GND.n1221 GND.n1220 341.085
R914 GND.n1222 GND.n1221 341.085
R915 GND.n1233 GND.n1029 341.085
R916 GND.n1236 GND.n1235 341.085
R917 GND.n1246 GND.n1245 341.085
R918 GND.n1248 GND.n1246 341.085
R919 GND.n1248 GND.n1247 341.085
R920 GND.n1257 GND.n1256 341.085
R921 GND.n1259 GND.n1258 341.085
R922 GND.n1269 GND.n1268 341.085
R923 GND.n504 GND.t304 334.459
R924 GND.t180 GND.n573 334.459
R925 GND.n456 GND.t202 319.767
R926 GND.n476 GND.t88 319.767
R927 GND.t185 GND.n476 319.767
R928 GND.n489 GND.t289 319.767
R929 GND.n402 GND.t184 319.767
R930 GND.n422 GND.t260 319.767
R931 GND.t232 GND.n422 319.767
R932 GND.n435 GND.t217 319.767
R933 GND.t218 GND.n323 319.767
R934 GND.n538 GND.t162 319.767
R935 GND.t268 GND.n538 319.767
R936 GND.n551 GND.t284 319.767
R937 GND.t56 GND.n289 319.767
R938 GND.n614 GND.t170 319.767
R939 GND.t42 GND.n614 319.767
R940 GND.n627 GND.t81 319.767
R941 GND.n1160 GND.t46 319.767
R942 GND.n1174 GND.t115 319.767
R943 GND.n1174 GND.t4 319.767
R944 GND.t303 GND.n1193 319.767
R945 GND.n1108 GND.t6 319.767
R946 GND.n1128 GND.t64 319.767
R947 GND.t274 GND.n1128 319.767
R948 GND.n1141 GND.t77 319.767
R949 GND.t58 GND.n1035 319.767
R950 GND.n1234 GND.t26 319.767
R951 GND.t188 GND.n1234 319.767
R952 GND.n1247 GND.t126 319.767
R953 GND.n454 GND.t36 277.131
R954 GND.n468 GND.t252 277.131
R955 GND.n478 GND.t223 277.131
R956 GND.t164 GND.n497 277.131
R957 GND.n400 GND.t295 277.131
R958 GND.n414 GND.t211 277.131
R959 GND.n424 GND.t109 277.131
R960 GND.t90 GND.n443 277.131
R961 GND.n514 GND.t130 277.131
R962 GND.t83 GND.n317 277.131
R963 GND.n539 GND.t308 277.131
R964 GND.t35 GND.n561 277.131
R965 GND.n590 GND.t213 277.131
R966 GND.t168 GND.n283 277.131
R967 GND.n615 GND.t102 277.131
R968 GND.t0 GND.n637 277.131
R969 GND.n1172 GND.t61 277.131
R970 GND.t19 GND.n1183 277.131
R971 GND.n1106 GND.t63 277.131
R972 GND.n1120 GND.t254 277.131
R973 GND.n1130 GND.t148 277.131
R974 GND.t117 GND.n1149 277.131
R975 GND.n1210 GND.t41 277.131
R976 GND.t91 GND.n1029 277.131
R977 GND.n1235 GND.t153 277.131
R978 GND.t45 GND.n1257 277.131
R979 GND.t304 GND.n503 269.289
R980 GND.n574 GND.t180 269.289
R981 GND.t265 GND.n329 234.496
R982 GND.n562 GND.t292 234.496
R983 GND.t104 GND.n295 234.496
R984 GND.n638 GND.t187 234.496
R985 GND.t172 GND.n1041 234.496
R986 GND.n1258 GND.t49 234.496
R987 GND.n752 GND.n751 231.68
R988 GND.n1422 GND.t283 192.984
R989 GND.n1469 GND.t114 192.984
R990 GND.n1362 GND.t111 192.984
R991 GND.n1532 GND.t59 192.984
R992 GND.n580 GND.t50 191.86
R993 GND.t179 GND.n648 191.86
R994 GND.n1200 GND.t133 191.86
R995 GND.t75 GND.n1269 191.86
R996 GND.n1570 GND.n1569 189.88
R997 GND.n578 GND.n577 183.68
R998 GND.n750 GND.t101 158.378
R999 GND.n651 GND.t251 158.378
R1000 GND.n157 GND.t128 158.378
R1001 GND.n257 GND.t194 158.378
R1002 GND.t50 GND.n579 158.378
R1003 GND.n649 GND.t179 158.378
R1004 GND.t133 GND.n1199 158.378
R1005 GND.n1270 GND.t75 158.378
R1006 GND.n911 GND.t134 158.378
R1007 GND.n1011 GND.t139 158.378
R1008 GND.n453 GND.n363 157.6
R1009 GND.n453 GND.n362 157.6
R1010 GND.n457 GND.n362 157.6
R1011 GND.n457 GND.n358 157.6
R1012 GND.n464 GND.n358 157.6
R1013 GND.n464 GND.n356 157.6
R1014 GND.n469 GND.n356 157.6
R1015 GND.n469 GND.n350 157.6
R1016 GND.n475 GND.n350 157.6
R1017 GND.n475 GND.n349 157.6
R1018 GND.n479 GND.n349 157.6
R1019 GND.n479 GND.n345 157.6
R1020 GND.n486 GND.n345 157.6
R1021 GND.n486 GND.n343 157.6
R1022 GND.n490 GND.n343 157.6
R1023 GND.n490 GND.n339 157.6
R1024 GND.n496 GND.n339 157.6
R1025 GND.n496 GND.n337 157.6
R1026 GND.n399 GND.n393 157.6
R1027 GND.n399 GND.n392 157.6
R1028 GND.n403 GND.n392 157.6
R1029 GND.n403 GND.n388 157.6
R1030 GND.n410 GND.n388 157.6
R1031 GND.n410 GND.n386 157.6
R1032 GND.n415 GND.n386 157.6
R1033 GND.n415 GND.n380 157.6
R1034 GND.n421 GND.n380 157.6
R1035 GND.n421 GND.n379 157.6
R1036 GND.n425 GND.n379 157.6
R1037 GND.n425 GND.n375 157.6
R1038 GND.n432 GND.n375 157.6
R1039 GND.n432 GND.n373 157.6
R1040 GND.n436 GND.n373 157.6
R1041 GND.n436 GND.n369 157.6
R1042 GND.n442 GND.n369 157.6
R1043 GND.n442 GND.n367 157.6
R1044 GND.n503 GND.n334 157.6
R1045 GND.n506 GND.n334 157.6
R1046 GND.n506 GND.n330 157.6
R1047 GND.n512 GND.n330 157.6
R1048 GND.n512 GND.n328 157.6
R1049 GND.n516 GND.n328 157.6
R1050 GND.n516 GND.n324 157.6
R1051 GND.n523 GND.n324 157.6
R1052 GND.n523 GND.n322 157.6
R1053 GND.n527 GND.n322 157.6
R1054 GND.n527 GND.n318 157.6
R1055 GND.n536 GND.n318 157.6
R1056 GND.n536 GND.n316 157.6
R1057 GND.n541 GND.n316 157.6
R1058 GND.n541 GND.n313 157.6
R1059 GND.n548 GND.n313 157.6
R1060 GND.n548 GND.n312 157.6
R1061 GND.n553 GND.n312 157.6
R1062 GND.n553 GND.n308 157.6
R1063 GND.n559 GND.n308 157.6
R1064 GND.n559 GND.n307 157.6
R1065 GND.n564 GND.n307 157.6
R1066 GND.n564 GND.n303 157.6
R1067 GND.n571 GND.n303 157.6
R1068 GND.n571 GND.n302 157.6
R1069 GND.n574 GND.n302 157.6
R1070 GND.n579 GND.n300 157.6
R1071 GND.n582 GND.n300 157.6
R1072 GND.n582 GND.n296 157.6
R1073 GND.n588 GND.n296 157.6
R1074 GND.n588 GND.n294 157.6
R1075 GND.n592 GND.n294 157.6
R1076 GND.n592 GND.n290 157.6
R1077 GND.n599 GND.n290 157.6
R1078 GND.n599 GND.n288 157.6
R1079 GND.n603 GND.n288 157.6
R1080 GND.n603 GND.n284 157.6
R1081 GND.n612 GND.n284 157.6
R1082 GND.n612 GND.n282 157.6
R1083 GND.n617 GND.n282 157.6
R1084 GND.n617 GND.n279 157.6
R1085 GND.n624 GND.n279 157.6
R1086 GND.n624 GND.n278 157.6
R1087 GND.n629 GND.n278 157.6
R1088 GND.n629 GND.n274 157.6
R1089 GND.n635 GND.n274 157.6
R1090 GND.n635 GND.n273 157.6
R1091 GND.n640 GND.n273 157.6
R1092 GND.n640 GND.n268 157.6
R1093 GND.n646 GND.n268 157.6
R1094 GND.n646 GND.n267 157.6
R1095 GND.n649 GND.n267 157.6
R1096 GND.n1431 GND.n1326 157.6
R1097 GND.n1431 GND.n1325 157.6
R1098 GND.n1436 GND.n1325 157.6
R1099 GND.n1436 GND.n1321 157.6
R1100 GND.n1443 GND.n1321 157.6
R1101 GND.n1443 GND.n1320 157.6
R1102 GND.n1447 GND.n1320 157.6
R1103 GND.n1447 GND.n1315 157.6
R1104 GND.n1454 GND.n1315 157.6
R1105 GND.n1454 GND.n1313 157.6
R1106 GND.n1458 GND.n1313 157.6
R1107 GND.n1458 GND.n1309 157.6
R1108 GND.n1464 GND.n1309 157.6
R1109 GND.n1464 GND.n1307 157.6
R1110 GND.n1366 GND.n1360 157.6
R1111 GND.n1366 GND.n1359 157.6
R1112 GND.n1371 GND.n1359 157.6
R1113 GND.n1371 GND.n1355 157.6
R1114 GND.n1377 GND.n1355 157.6
R1115 GND.n1377 GND.n1354 157.6
R1116 GND.n1382 GND.n1354 157.6
R1117 GND.n1382 GND.n1350 157.6
R1118 GND.n1389 GND.n1350 157.6
R1119 GND.n1389 GND.n1349 157.6
R1120 GND.n1393 GND.n1349 157.6
R1121 GND.n1393 GND.n1344 157.6
R1122 GND.n1400 GND.n1344 157.6
R1123 GND.n1400 GND.n1342 157.6
R1124 GND.n1404 GND.n1342 157.6
R1125 GND.n1404 GND.n1338 157.6
R1126 GND.n1410 GND.n1338 157.6
R1127 GND.n1410 GND.n1336 157.6
R1128 GND.n1414 GND.n1336 157.6
R1129 GND.n1414 GND.n1332 157.6
R1130 GND.n1420 GND.n1332 157.6
R1131 GND.n1420 GND.n1330 157.6
R1132 GND.n1475 GND.n1303 157.6
R1133 GND.n1475 GND.n1302 157.6
R1134 GND.n1480 GND.n1302 157.6
R1135 GND.n1480 GND.n1298 157.6
R1136 GND.n1486 GND.n1298 157.6
R1137 GND.n1486 GND.n1297 157.6
R1138 GND.n1491 GND.n1297 157.6
R1139 GND.n1491 GND.n1293 157.6
R1140 GND.n1498 GND.n1293 157.6
R1141 GND.n1498 GND.n1292 157.6
R1142 GND.n1502 GND.n1292 157.6
R1143 GND.n1502 GND.n1287 157.6
R1144 GND.n1509 GND.n1287 157.6
R1145 GND.n1509 GND.n1285 157.6
R1146 GND.n1513 GND.n1285 157.6
R1147 GND.n1513 GND.n1281 157.6
R1148 GND.n1519 GND.n1281 157.6
R1149 GND.n1519 GND.n1279 157.6
R1150 GND.n1523 GND.n1279 157.6
R1151 GND.n1523 GND.n1275 157.6
R1152 GND.n1530 GND.n1275 157.6
R1153 GND.n1530 GND.n1273 157.6
R1154 GND.n1159 GND.n1069 157.6
R1155 GND.n1159 GND.n1068 157.6
R1156 GND.n1164 GND.n1068 157.6
R1157 GND.n1164 GND.n1064 157.6
R1158 GND.n1171 GND.n1064 157.6
R1159 GND.n1171 GND.n1063 157.6
R1160 GND.n1175 GND.n1063 157.6
R1161 GND.n1175 GND.n1057 157.6
R1162 GND.n1182 GND.n1057 157.6
R1163 GND.n1182 GND.n1055 157.6
R1164 GND.n1186 GND.n1055 157.6
R1165 GND.n1186 GND.n1051 157.6
R1166 GND.n1192 GND.n1051 157.6
R1167 GND.n1192 GND.n1049 157.6
R1168 GND.n1105 GND.n1099 157.6
R1169 GND.n1105 GND.n1098 157.6
R1170 GND.n1109 GND.n1098 157.6
R1171 GND.n1109 GND.n1094 157.6
R1172 GND.n1116 GND.n1094 157.6
R1173 GND.n1116 GND.n1092 157.6
R1174 GND.n1121 GND.n1092 157.6
R1175 GND.n1121 GND.n1086 157.6
R1176 GND.n1127 GND.n1086 157.6
R1177 GND.n1127 GND.n1085 157.6
R1178 GND.n1131 GND.n1085 157.6
R1179 GND.n1131 GND.n1081 157.6
R1180 GND.n1138 GND.n1081 157.6
R1181 GND.n1138 GND.n1079 157.6
R1182 GND.n1142 GND.n1079 157.6
R1183 GND.n1142 GND.n1075 157.6
R1184 GND.n1148 GND.n1075 157.6
R1185 GND.n1148 GND.n1073 157.6
R1186 GND.n1199 GND.n1046 157.6
R1187 GND.n1202 GND.n1046 157.6
R1188 GND.n1202 GND.n1042 157.6
R1189 GND.n1208 GND.n1042 157.6
R1190 GND.n1208 GND.n1040 157.6
R1191 GND.n1212 GND.n1040 157.6
R1192 GND.n1212 GND.n1036 157.6
R1193 GND.n1219 GND.n1036 157.6
R1194 GND.n1219 GND.n1034 157.6
R1195 GND.n1223 GND.n1034 157.6
R1196 GND.n1223 GND.n1030 157.6
R1197 GND.n1232 GND.n1030 157.6
R1198 GND.n1232 GND.n1028 157.6
R1199 GND.n1237 GND.n1028 157.6
R1200 GND.n1237 GND.n1025 157.6
R1201 GND.n1244 GND.n1025 157.6
R1202 GND.n1244 GND.n1024 157.6
R1203 GND.n1249 GND.n1024 157.6
R1204 GND.n1249 GND.n1020 157.6
R1205 GND.n1255 GND.n1020 157.6
R1206 GND.n1255 GND.n1019 157.6
R1207 GND.n1260 GND.n1019 157.6
R1208 GND.n1260 GND.n1015 157.6
R1209 GND.n1267 GND.n1015 157.6
R1210 GND.n1267 GND.n1014 157.6
R1211 GND.n1270 GND.n1014 157.6
R1212 GND.n1363 GND.n1362 135.387
R1213 GND.n505 GND.t265 133.857
R1214 GND.n572 GND.t292 133.857
R1215 GND.n1426 GND.n1425 132.648
R1216 GND.n1533 GND.n1532 132.648
R1217 GND.n1467 GND.n1466 132.647
R1218 GND.n1423 GND.n1422 132.647
R1219 GND.n1470 GND.n1469 132.647
R1220 GND.n1809 GND.t53 126.679
R1221 GND.n1844 GND.t344 126.679
R1222 GND.n1563 GND.t176 126.679
R1223 GND.n1865 GND.t332 126.679
R1224 GND.n396 GND.n395 118.662
R1225 GND.n1102 GND.n1101 118.662
R1226 GND.n448 GND.n447 115.922
R1227 GND.n1154 GND.n1153 115.922
R1228 GND.n499 GND.n498 115.922
R1229 GND.n445 GND.n444 115.922
R1230 GND.n1195 GND.n1194 115.922
R1231 GND.n1151 GND.n1150 115.922
R1232 GND.n1434 GND.t237 111.486
R1233 GND.n1456 GND.t51 111.486
R1234 GND.t206 GND.n1368 111.486
R1235 GND.n1380 GND.t341 111.486
R1236 GND.n1402 GND.t355 111.486
R1237 GND.t273 GND.n1331 111.486
R1238 GND.t135 GND.n1477 111.486
R1239 GND.n1489 GND.t17 111.486
R1240 GND.n1511 GND.t278 111.486
R1241 GND.t69 GND.n1274 111.486
R1242 GND.n745 GND.t57 106.589
R1243 GND.n657 GND.t239 106.589
R1244 GND.n164 GND.t97 106.589
R1245 GND.n252 GND.t16 106.589
R1246 GND.n581 GND.t104 106.589
R1247 GND.n647 GND.t187 106.589
R1248 GND.n1201 GND.t172 106.589
R1249 GND.n1268 GND.t49 106.589
R1250 GND.n918 GND.t80 106.589
R1251 GND.n1006 GND.t190 106.589
R1252 GND.n1703 GND.t325 98.214
R1253 GND.n1752 GND.t348 98.214
R1254 GND.n87 GND.t1 70.155
R1255 GND.n498 GND.t164 70.155
R1256 GND.n444 GND.t90 70.155
R1257 GND.n1150 GND.t117 70.155
R1258 GND.n841 GND.t225 70.155
R1259 GND.n15 GND.t208 70.155
R1260 GND.n447 GND.t36 70.155
R1261 GND.n395 GND.t295 70.155
R1262 GND.n1101 GND.t63 70.155
R1263 GND.n769 GND.t122 70.155
R1264 GND.n1917 GND.n1916 67.266
R1265 GND.n737 GND.t32 63.953
R1266 GND.n712 GND.t266 63.953
R1267 GND.n690 GND.t136 63.953
R1268 GND.n665 GND.t55 63.953
R1269 GND.n172 GND.t48 63.953
R1270 GND.n197 GND.t67 63.953
R1271 GND.n219 GND.t22 63.953
R1272 GND.n244 GND.t47 63.953
R1273 GND.n112 GND.t78 63.953
R1274 GND.n134 GND.t107 63.953
R1275 GND.n40 GND.t174 63.953
R1276 GND.n62 GND.t143 63.953
R1277 GND.t252 GND.n466 63.953
R1278 GND.t223 GND.n344 63.953
R1279 GND.t211 GND.n412 63.953
R1280 GND.t109 GND.n374 63.953
R1281 GND.t130 GND.n513 63.953
R1282 GND.n526 GND.t83 63.953
R1283 GND.n549 GND.t308 63.953
R1284 GND.n563 GND.t35 63.953
R1285 GND.t213 GND.n589 63.953
R1286 GND.n602 GND.t168 63.953
R1287 GND.n625 GND.t102 63.953
R1288 GND.n639 GND.t0 63.953
R1289 GND.n1162 GND.t61 63.953
R1290 GND.n1184 GND.t19 63.953
R1291 GND.t254 GND.n1118 63.953
R1292 GND.t148 GND.n1080 63.953
R1293 GND.t41 GND.n1209 63.953
R1294 GND.n1222 GND.t91 63.953
R1295 GND.n1245 GND.t153 63.953
R1296 GND.n1259 GND.t45 63.953
R1297 GND.n866 GND.t119 63.953
R1298 GND.n888 GND.t28 63.953
R1299 GND.n794 GND.t286 63.953
R1300 GND.n816 GND.t145 63.953
R1301 GND.n926 GND.t38 63.953
R1302 GND.n951 GND.t198 63.953
R1303 GND.n973 GND.t24 63.953
R1304 GND.n998 GND.t37 63.953
R1305 GND.n1933 GND.t201 63.309
R1306 GND.n2092 GND.t21 63.309
R1307 GND.n1941 GND.t129 59.352
R1308 GND.n1945 GND.t44 59.352
R1309 GND.n1991 GND.t276 59.352
R1310 GND.n1995 GND.t320 59.352
R1311 GND.n2030 GND.t230 59.352
R1312 GND.n2034 GND.t263 59.352
R1313 GND.n2080 GND.t343 59.352
R1314 GND.n2084 GND.t336 59.352
R1315 GND.n1929 GND.t39 55.395
R1316 GND.n2096 GND.t131 55.395
R1317 GND.n1895 GND.t258 49.588
R1318 GND.n1779 GND.t242 49.588
R1319 EESPFAL_Sbox_0/EESPFAL_s3_0/GND GND.n1533 47.3
R1320 GND.n1761 GND.n1760 45.833
R1321 GND.n1466 GND.t270 44.336
R1322 GND.n1425 GND.t299 44.336
R1323 GND.n1560 GND.t327 42.226
R1324 GND.n1834 GND.t311 42.226
R1325 GND.n1878 GND.t87 42.226
R1326 GND.n1796 GND.t10 42.226
R1327 GND.n1553 GND.t247 42.226
R1328 GND.n1848 GND.t228 42.226
R1329 GND.n1628 GND.t204 39.285
R1330 GND.n1586 GND.t240 39.285
R1331 GND.n1535 GND.n1012 37.93
R1332 GND.t72 GND.n1445 37.162
R1333 GND.t112 GND.n1314 37.162
R1334 GND.n1369 GND.t121 37.162
R1335 GND.t94 GND.n1391 37.162
R1336 GND.t234 GND.n1343 37.162
R1337 GND.n1412 GND.t323 37.162
R1338 GND.n1478 GND.t306 37.162
R1339 GND.t271 GND.n1500 37.162
R1340 GND.t297 GND.n1286 37.162
R1341 GND.n1521 GND.t347 37.162
R1342 GND.n652 EESPFAL_4in_XOR_0/GND 35.195
R1343 GND.n1640 GND.t216 32.738
R1344 GND.n1570 GND.t30 32.738
R1345 GND.n1687 GND.t330 32.738
R1346 GND.n1736 GND.t196 32.738
R1347 EESPFAL_4in_XOR_0/GND GND.n650 31.551
R1348 GND.n1534 GND.n1271 31.53
R1349 GND.n716 GND.t280 29.103
R1350 GND.n689 GND.t214 29.103
R1351 GND.n39 GND.t288 29.103
R1352 GND.n66 GND.t346 29.103
R1353 GND.n111 GND.t79 29.103
R1354 GND.n138 GND.t200 29.103
R1355 GND.n196 GND.t191 29.103
R1356 GND.n223 GND.t23 29.103
R1357 GND.n407 GND.t246 29.103
R1358 GND.n429 GND.t147 29.103
R1359 GND.n461 GND.t293 29.103
R1360 GND.n483 GND.t224 29.103
R1361 GND.n320 GND.t84 29.103
R1362 GND.n545 GND.t338 29.103
R1363 GND.n286 GND.t215 29.103
R1364 GND.n621 GND.t352 29.103
R1365 GND.n1666 GND.t241 29.103
R1366 GND.n1711 GND.t326 29.103
R1367 GND.n1825 GND.t177 29.103
R1368 GND.n1873 GND.t333 29.103
R1369 GND.n1990 GND.t321 29.103
R1370 GND.n2043 GND.t264 29.103
R1371 GND.n1385 GND.t342 29.103
R1372 GND.n1340 GND.t356 29.103
R1373 GND.n1439 GND.t238 29.103
R1374 GND.n1311 GND.t52 29.103
R1375 GND.n1494 GND.t18 29.103
R1376 GND.n1283 GND.t279 29.103
R1377 GND.n1113 GND.t255 29.103
R1378 GND.n1135 GND.t245 29.103
R1379 GND.n1167 GND.t167 29.103
R1380 GND.n1053 GND.t20 29.103
R1381 GND.n1032 GND.t92 29.103
R1382 GND.n1241 GND.t154 29.103
R1383 GND.n793 GND.t351 29.103
R1384 GND.n820 GND.t334 29.103
R1385 GND.n865 GND.t120 29.103
R1386 GND.n892 GND.t29 29.103
R1387 GND.n950 GND.t199 29.103
R1388 GND.n977 GND.t96 29.103
R1389 GND.n716 GND.t267 29.102
R1390 GND.n689 GND.t137 29.102
R1391 GND.n39 GND.t175 29.102
R1392 GND.n66 GND.t144 29.102
R1393 GND.n111 GND.t317 29.102
R1394 GND.n138 GND.t108 29.102
R1395 GND.n196 GND.t68 29.102
R1396 GND.n223 GND.t314 29.102
R1397 GND.n407 GND.t212 29.102
R1398 GND.n429 GND.t110 29.102
R1399 GND.n461 GND.t253 29.102
R1400 GND.n483 GND.t236 29.102
R1401 GND.n320 GND.t222 29.102
R1402 GND.n545 GND.t309 29.102
R1403 GND.n286 GND.t169 29.102
R1404 GND.n621 GND.t103 29.102
R1405 GND.n1690 GND.t354 29.102
R1406 GND.n1648 GND.t210 29.102
R1407 GND.n1852 GND.t345 29.102
R1408 GND.n1804 GND.t54 29.102
R1409 GND.n2038 GND.t231 29.102
R1410 GND.n1985 GND.t277 29.102
R1411 GND.n1113 GND.t350 29.102
R1412 GND.n1135 GND.t149 29.102
R1413 GND.n1167 GND.t62 29.102
R1414 GND.n1053 GND.t315 29.102
R1415 GND.n1032 GND.t329 29.102
R1416 GND.n1241 GND.t318 29.102
R1417 GND.n793 GND.t287 29.102
R1418 GND.n820 GND.t146 29.102
R1419 GND.n865 GND.t138 29.102
R1420 GND.n892 GND.t66 29.102
R1421 GND.n950 GND.t262 29.102
R1422 GND.n977 GND.t25 29.102
R1423 GND.n151 GND.t195 27.519
R1424 GND.n1194 GND.t303 27.519
R1425 GND.n905 GND.t40 27.519
R1426 GND.n95 GND.t219 27.519
R1427 GND.n1153 GND.t46 27.519
R1428 GND.n849 GND.t15 27.519
R1429 GND.n577 GND.n575 26.88
R1430 GND.n752 GND.n258 26.88
R1431 GND.n1612 GND.t74 26.19
R1432 GND.n263 GND.t182 24
R1433 GND.n263 GND.t307 24
R1434 GND.n262 GND.t207 24
R1435 GND.n262 GND.t221 24
R1436 GND.n6 GND.t141 24
R1437 GND.n6 GND.t71 24
R1438 GND.n5 GND.t281 24
R1439 GND.n5 GND.t82 24
R1440 GND.n10 GND.t33 24
R1441 GND.n10 GND.t14 24
R1442 GND.n9 GND.t3 24
R1443 GND.n9 GND.t161 24
R1444 GND.n14 GND.t203 24
R1445 GND.n14 GND.t349 24
R1446 GND.n13 GND.t193 24
R1447 GND.n13 GND.t159 24
R1448 GND.n608 GND.t171 24
R1449 GND.n608 GND.t43 24
R1450 GND.n607 GND.t319 24
R1451 GND.n607 GND.t125 24
R1452 GND.n532 GND.t163 24
R1453 GND.n532 GND.t269 24
R1454 GND.n531 GND.t249 24
R1455 GND.n531 GND.t313 24
R1456 GND.n353 GND.t183 24
R1457 GND.n353 GND.t291 24
R1458 GND.n352 GND.t89 24
R1459 GND.n352 GND.t186 24
R1460 GND.n383 GND.t261 24
R1461 GND.n383 GND.t233 24
R1462 GND.n382 GND.t296 24
R1463 GND.n382 GND.t259 24
R1464 GND.n1552 GND.t86 24
R1465 GND.n1552 GND.t244 24
R1466 GND.n1551 GND.t257 24
R1467 GND.n1551 GND.t12 24
R1468 GND.n1568 GND.t328 24
R1469 GND.n1568 GND.t312 24
R1470 GND.n1559 GND.t248 24
R1471 GND.n1559 GND.t229 24
R1472 GND.n1588 GND.t340 24
R1473 GND.n1588 GND.t106 24
R1474 GND.n1576 GND.t31 24
R1475 GND.n1576 GND.t331 24
R1476 GND.n1289 GND.t272 24
R1477 GND.n1289 GND.t298 24
R1478 GND.n1317 GND.t73 24
R1479 GND.n1317 GND.t113 24
R1480 GND.n1346 GND.t95 24
R1481 GND.n1346 GND.t235 24
R1482 GND.n1228 GND.t324 24
R1483 GND.n1228 GND.t189 24
R1484 GND.n1227 GND.t27 24
R1485 GND.n1227 GND.t285 24
R1486 GND.n1060 GND.t116 24
R1487 GND.n1060 GND.t118 24
R1488 GND.n1059 GND.t294 24
R1489 GND.n1059 GND.t5 24
R1490 GND.n1089 GND.t205 24
R1491 GND.n1089 GND.t275 24
R1492 GND.n1088 GND.t65 24
R1493 GND.n1088 GND.t282 24
R1494 GND.n760 GND.t316 24
R1495 GND.n760 GND.t301 24
R1496 GND.n759 GND.t8 24
R1497 GND.n759 GND.t124 24
R1498 GND.n764 GND.t227 24
R1499 GND.n764 GND.t99 24
R1500 GND.n763 GND.t250 24
R1501 GND.n763 GND.t337 24
R1502 GND.n768 GND.t300 24
R1503 GND.n768 GND.t165 24
R1504 GND.n767 GND.t157 24
R1505 GND.n767 GND.t151 24
R1506 GND.n1536 GND.t76 23.741
R1507 GND.n729 GND.t178 21.317
R1508 GND.n704 GND.t181 21.317
R1509 GND.n699 GND.t220 21.317
R1510 GND.n673 GND.t173 21.317
R1511 GND.n180 GND.t60 21.317
R1512 GND.n205 GND.t140 21.317
R1513 GND.n211 GND.t70 21.317
R1514 GND.n236 GND.t127 21.317
R1515 GND.n120 GND.t2 21.317
R1516 GND.n126 GND.t13 21.317
R1517 GND.n23 GND.t34 21.317
R1518 GND.n48 GND.t192 21.317
R1519 GND.n54 GND.t158 21.317
R1520 GND.n79 GND.t142 21.317
R1521 GND.t202 GND.n455 21.317
R1522 GND.n467 GND.t88 21.317
R1523 GND.n477 GND.t185 21.317
R1524 GND.t289 GND.n338 21.317
R1525 GND.t184 GND.n401 21.317
R1526 GND.n413 GND.t260 21.317
R1527 GND.n423 GND.t232 21.317
R1528 GND.t217 GND.n368 21.317
R1529 GND.n515 GND.t218 21.317
R1530 GND.t162 GND.n537 21.317
R1531 GND.n540 GND.t268 21.317
R1532 GND.n560 GND.t284 21.317
R1533 GND.n591 GND.t56 21.317
R1534 GND.t170 GND.n613 21.317
R1535 GND.n616 GND.t42 21.317
R1536 GND.n636 GND.t81 21.317
R1537 GND.t115 GND.n1173 21.317
R1538 GND.t4 GND.n1056 21.317
R1539 GND.t6 GND.n1107 21.317
R1540 GND.n1119 GND.t64 21.317
R1541 GND.n1129 GND.t274 21.317
R1542 GND.t77 GND.n1074 21.317
R1543 GND.n1211 GND.t58 21.317
R1544 GND.t26 GND.n1233 21.317
R1545 GND.n1236 GND.t188 21.317
R1546 GND.n1256 GND.t126 21.317
R1547 GND.n874 GND.t226 21.317
R1548 GND.n880 GND.t98 21.317
R1549 GND.n777 GND.t100 21.317
R1550 GND.n802 GND.t156 21.317
R1551 GND.n808 GND.t150 21.317
R1552 GND.n833 GND.t9 21.317
R1553 GND.n934 GND.t197 21.317
R1554 GND.n959 GND.t7 21.317
R1555 GND.n965 GND.t123 21.317
R1556 GND.n990 GND.t132 21.317
R1557 GND.n1957 GND.t290 19.784
R1558 GND.n1961 GND.t335 19.784
R1559 GND.n1542 GND.t85 19.784
R1560 GND.n1545 GND.t256 19.784
R1561 GND.n2014 GND.t243 19.784
R1562 GND.n2018 GND.t11 19.784
R1563 GND.n2064 GND.t302 19.784
R1564 GND.n2068 GND.t305 19.784
R1565 GND.n1773 GND.n1772 17.357
R1566 GND.n128 GND.n125 12.8
R1567 GND.n56 GND.n53 12.8
R1568 GND.n448 GND.n364 12.8
R1569 GND.n452 GND.n364 12.8
R1570 GND.n452 GND.n361 12.8
R1571 GND.n458 GND.n361 12.8
R1572 GND.n458 GND.n359 12.8
R1573 GND.n463 GND.n359 12.8
R1574 GND.n463 GND.n355 12.8
R1575 GND.n470 GND.n355 12.8
R1576 GND.n470 GND.n351 12.8
R1577 GND.n474 GND.n351 12.8
R1578 GND.n474 GND.n348 12.8
R1579 GND.n480 GND.n348 12.8
R1580 GND.n480 GND.n346 12.8
R1581 GND.n485 GND.n346 12.8
R1582 GND.n485 GND.n342 12.8
R1583 GND.n491 GND.n342 12.8
R1584 GND.n491 GND.n340 12.8
R1585 GND.n495 GND.n340 12.8
R1586 GND.n495 GND.n336 12.8
R1587 GND.n499 GND.n336 12.8
R1588 GND.n398 GND.n394 12.8
R1589 GND.n398 GND.n391 12.8
R1590 GND.n404 GND.n391 12.8
R1591 GND.n404 GND.n389 12.8
R1592 GND.n409 GND.n389 12.8
R1593 GND.n409 GND.n385 12.8
R1594 GND.n416 GND.n385 12.8
R1595 GND.n416 GND.n381 12.8
R1596 GND.n420 GND.n381 12.8
R1597 GND.n420 GND.n378 12.8
R1598 GND.n426 GND.n378 12.8
R1599 GND.n426 GND.n376 12.8
R1600 GND.n431 GND.n376 12.8
R1601 GND.n431 GND.n372 12.8
R1602 GND.n437 GND.n372 12.8
R1603 GND.n437 GND.n370 12.8
R1604 GND.n441 GND.n370 12.8
R1605 GND.n441 GND.n366 12.8
R1606 GND.n445 GND.n366 12.8
R1607 GND.n502 GND.n333 12.8
R1608 GND.n507 GND.n333 12.8
R1609 GND.n507 GND.n331 12.8
R1610 GND.n511 GND.n331 12.8
R1611 GND.n511 GND.n327 12.8
R1612 GND.n517 GND.n327 12.8
R1613 GND.n517 GND.n325 12.8
R1614 GND.n522 GND.n325 12.8
R1615 GND.n522 GND.n321 12.8
R1616 GND.n528 GND.n321 12.8
R1617 GND.n528 GND.n319 12.8
R1618 GND.n535 GND.n319 12.8
R1619 GND.n535 GND.n315 12.8
R1620 GND.n542 GND.n315 12.8
R1621 GND.n542 GND.n314 12.8
R1622 GND.n547 GND.n314 12.8
R1623 GND.n547 GND.n311 12.8
R1624 GND.n554 GND.n311 12.8
R1625 GND.n554 GND.n309 12.8
R1626 GND.n558 GND.n309 12.8
R1627 GND.n558 GND.n306 12.8
R1628 GND.n565 GND.n306 12.8
R1629 GND.n565 GND.n304 12.8
R1630 GND.n570 GND.n304 12.8
R1631 GND.n570 GND.n569 12.8
R1632 GND.n583 GND.n299 12.8
R1633 GND.n583 GND.n297 12.8
R1634 GND.n587 GND.n297 12.8
R1635 GND.n587 GND.n293 12.8
R1636 GND.n593 GND.n293 12.8
R1637 GND.n593 GND.n291 12.8
R1638 GND.n598 GND.n291 12.8
R1639 GND.n598 GND.n287 12.8
R1640 GND.n604 GND.n287 12.8
R1641 GND.n604 GND.n285 12.8
R1642 GND.n611 GND.n285 12.8
R1643 GND.n611 GND.n281 12.8
R1644 GND.n618 GND.n281 12.8
R1645 GND.n618 GND.n280 12.8
R1646 GND.n623 GND.n280 12.8
R1647 GND.n623 GND.n277 12.8
R1648 GND.n630 GND.n277 12.8
R1649 GND.n630 GND.n275 12.8
R1650 GND.n634 GND.n275 12.8
R1651 GND.n634 GND.n272 12.8
R1652 GND.n641 GND.n272 12.8
R1653 GND.n641 GND.n269 12.8
R1654 GND.n645 GND.n269 12.8
R1655 GND.n645 GND.n270 12.8
R1656 GND.n1426 GND.n1327 12.8
R1657 GND.n1430 GND.n1327 12.8
R1658 GND.n1430 GND.n1324 12.8
R1659 GND.n1437 GND.n1324 12.8
R1660 GND.n1437 GND.n1322 12.8
R1661 GND.n1442 GND.n1322 12.8
R1662 GND.n1442 GND.n1319 12.8
R1663 GND.n1448 GND.n1319 12.8
R1664 GND.n1448 GND.n1316 12.8
R1665 GND.n1453 GND.n1316 12.8
R1666 GND.n1453 GND.n1312 12.8
R1667 GND.n1459 GND.n1312 12.8
R1668 GND.n1459 GND.n1310 12.8
R1669 GND.n1463 GND.n1310 12.8
R1670 GND.n1463 GND.n1306 12.8
R1671 GND.n1467 GND.n1306 12.8
R1672 GND.n1365 GND.n1361 12.8
R1673 GND.n1365 GND.n1358 12.8
R1674 GND.n1372 GND.n1358 12.8
R1675 GND.n1372 GND.n1356 12.8
R1676 GND.n1376 GND.n1356 12.8
R1677 GND.n1376 GND.n1353 12.8
R1678 GND.n1383 GND.n1353 12.8
R1679 GND.n1383 GND.n1351 12.8
R1680 GND.n1388 GND.n1351 12.8
R1681 GND.n1388 GND.n1348 12.8
R1682 GND.n1394 GND.n1348 12.8
R1683 GND.n1394 GND.n1345 12.8
R1684 GND.n1399 GND.n1345 12.8
R1685 GND.n1399 GND.n1341 12.8
R1686 GND.n1405 GND.n1341 12.8
R1687 GND.n1405 GND.n1339 12.8
R1688 GND.n1409 GND.n1339 12.8
R1689 GND.n1409 GND.n1335 12.8
R1690 GND.n1415 GND.n1335 12.8
R1691 GND.n1415 GND.n1333 12.8
R1692 GND.n1419 GND.n1333 12.8
R1693 GND.n1419 GND.n1329 12.8
R1694 GND.n1423 GND.n1329 12.8
R1695 GND.n1470 GND.n1304 12.8
R1696 GND.n1474 GND.n1304 12.8
R1697 GND.n1474 GND.n1301 12.8
R1698 GND.n1481 GND.n1301 12.8
R1699 GND.n1481 GND.n1299 12.8
R1700 GND.n1485 GND.n1299 12.8
R1701 GND.n1485 GND.n1296 12.8
R1702 GND.n1492 GND.n1296 12.8
R1703 GND.n1492 GND.n1294 12.8
R1704 GND.n1497 GND.n1294 12.8
R1705 GND.n1497 GND.n1291 12.8
R1706 GND.n1503 GND.n1291 12.8
R1707 GND.n1503 GND.n1288 12.8
R1708 GND.n1508 GND.n1288 12.8
R1709 GND.n1508 GND.n1284 12.8
R1710 GND.n1514 GND.n1284 12.8
R1711 GND.n1514 GND.n1282 12.8
R1712 GND.n1518 GND.n1282 12.8
R1713 GND.n1518 GND.n1278 12.8
R1714 GND.n1524 GND.n1278 12.8
R1715 GND.n1524 GND.n1276 12.8
R1716 GND.n1529 GND.n1276 12.8
R1717 GND.n1529 GND.n1528 12.8
R1718 GND.n1154 GND.n1070 12.8
R1719 GND.n1158 GND.n1070 12.8
R1720 GND.n1158 GND.n1067 12.8
R1721 GND.n1165 GND.n1067 12.8
R1722 GND.n1165 GND.n1065 12.8
R1723 GND.n1170 GND.n1065 12.8
R1724 GND.n1170 GND.n1062 12.8
R1725 GND.n1176 GND.n1062 12.8
R1726 GND.n1176 GND.n1058 12.8
R1727 GND.n1181 GND.n1058 12.8
R1728 GND.n1181 GND.n1054 12.8
R1729 GND.n1187 GND.n1054 12.8
R1730 GND.n1187 GND.n1052 12.8
R1731 GND.n1191 GND.n1052 12.8
R1732 GND.n1191 GND.n1048 12.8
R1733 GND.n1195 GND.n1048 12.8
R1734 GND.n1104 GND.n1100 12.8
R1735 GND.n1104 GND.n1097 12.8
R1736 GND.n1110 GND.n1097 12.8
R1737 GND.n1110 GND.n1095 12.8
R1738 GND.n1115 GND.n1095 12.8
R1739 GND.n1115 GND.n1091 12.8
R1740 GND.n1122 GND.n1091 12.8
R1741 GND.n1122 GND.n1087 12.8
R1742 GND.n1126 GND.n1087 12.8
R1743 GND.n1126 GND.n1084 12.8
R1744 GND.n1132 GND.n1084 12.8
R1745 GND.n1132 GND.n1082 12.8
R1746 GND.n1137 GND.n1082 12.8
R1747 GND.n1137 GND.n1078 12.8
R1748 GND.n1143 GND.n1078 12.8
R1749 GND.n1143 GND.n1076 12.8
R1750 GND.n1147 GND.n1076 12.8
R1751 GND.n1147 GND.n1072 12.8
R1752 GND.n1151 GND.n1072 12.8
R1753 GND.n1198 GND.n1045 12.8
R1754 GND.n1203 GND.n1045 12.8
R1755 GND.n1203 GND.n1043 12.8
R1756 GND.n1207 GND.n1043 12.8
R1757 GND.n1207 GND.n1039 12.8
R1758 GND.n1213 GND.n1039 12.8
R1759 GND.n1213 GND.n1037 12.8
R1760 GND.n1218 GND.n1037 12.8
R1761 GND.n1218 GND.n1033 12.8
R1762 GND.n1224 GND.n1033 12.8
R1763 GND.n1224 GND.n1031 12.8
R1764 GND.n1231 GND.n1031 12.8
R1765 GND.n1231 GND.n1027 12.8
R1766 GND.n1238 GND.n1027 12.8
R1767 GND.n1238 GND.n1026 12.8
R1768 GND.n1243 GND.n1026 12.8
R1769 GND.n1243 GND.n1023 12.8
R1770 GND.n1250 GND.n1023 12.8
R1771 GND.n1250 GND.n1021 12.8
R1772 GND.n1254 GND.n1021 12.8
R1773 GND.n1254 GND.n1018 12.8
R1774 GND.n1261 GND.n1018 12.8
R1775 GND.n1261 GND.n1016 12.8
R1776 GND.n1266 GND.n1016 12.8
R1777 GND.n1266 GND.n1265 12.8
R1778 GND.n882 GND.n879 12.8
R1779 GND.n810 GND.n807 12.8
R1780 GND.n967 GND.n964 12.8
R1781 GND.n213 GND.n210 12.8
R1782 GND.n702 GND.n701 12.8
R1783 GND.n2111 GND.n2110 12.475
R1784 GND.n17 GND.n16 9.154
R1785 GND.n21 GND.n20 9.154
R1786 GND.n20 GND.n19 9.154
R1787 GND.n25 GND.n24 9.154
R1788 GND.n24 GND.n23 9.154
R1789 GND.n29 GND.n28 9.154
R1790 GND.n28 GND.n27 9.154
R1791 GND.n33 GND.n32 9.154
R1792 GND.n32 GND.n31 9.154
R1793 GND.n37 GND.n36 9.154
R1794 GND.n36 GND.n35 9.154
R1795 GND.n42 GND.n41 9.154
R1796 GND.n41 GND.n40 9.154
R1797 GND.n46 GND.n45 9.154
R1798 GND.n45 GND.n44 9.154
R1799 GND.n50 GND.n49 9.154
R1800 GND.n49 GND.n48 9.154
R1801 GND.n53 GND.n12 9.154
R1802 GND.n12 GND.n11 9.154
R1803 GND.n56 GND.n55 9.154
R1804 GND.n55 GND.n54 9.154
R1805 GND.n60 GND.n59 9.154
R1806 GND.n59 GND.n58 9.154
R1807 GND.n64 GND.n63 9.154
R1808 GND.n63 GND.n62 9.154
R1809 GND.n69 GND.n68 9.154
R1810 GND.n68 GND.n67 9.154
R1811 GND.n73 GND.n72 9.154
R1812 GND.n72 GND.n71 9.154
R1813 GND.n77 GND.n76 9.154
R1814 GND.n76 GND.n75 9.154
R1815 GND.n81 GND.n80 9.154
R1816 GND.n80 GND.n79 9.154
R1817 GND.n85 GND.n84 9.154
R1818 GND.n84 GND.n83 9.154
R1819 GND.n89 GND.n88 9.154
R1820 GND.n97 GND.n96 9.154
R1821 GND.n101 GND.n100 9.154
R1822 GND.n100 GND.n99 9.154
R1823 GND.n105 GND.n104 9.154
R1824 GND.n104 GND.n103 9.154
R1825 GND.n109 GND.n108 9.154
R1826 GND.n108 GND.n107 9.154
R1827 GND.n114 GND.n113 9.154
R1828 GND.n113 GND.n112 9.154
R1829 GND.n118 GND.n117 9.154
R1830 GND.n117 GND.n116 9.154
R1831 GND.n122 GND.n121 9.154
R1832 GND.n121 GND.n120 9.154
R1833 GND.n125 GND.n8 9.154
R1834 GND.n8 GND.n7 9.154
R1835 GND.n128 GND.n127 9.154
R1836 GND.n127 GND.n126 9.154
R1837 GND.n132 GND.n131 9.154
R1838 GND.n131 GND.n130 9.154
R1839 GND.n136 GND.n135 9.154
R1840 GND.n135 GND.n134 9.154
R1841 GND.n141 GND.n140 9.154
R1842 GND.n140 GND.n139 9.154
R1843 GND.n145 GND.n144 9.154
R1844 GND.n144 GND.n143 9.154
R1845 GND.n149 GND.n148 9.154
R1846 GND.n148 GND.n147 9.154
R1847 GND.n153 GND.n152 9.154
R1848 GND.n394 GND.n393 9.154
R1849 GND.n399 GND.n398 9.154
R1850 GND.n400 GND.n399 9.154
R1851 GND.n392 GND.n391 9.154
R1852 GND.n401 GND.n392 9.154
R1853 GND.n404 GND.n403 9.154
R1854 GND.n403 GND.n402 9.154
R1855 GND.n389 GND.n388 9.154
R1856 GND.n388 GND.n387 9.154
R1857 GND.n410 GND.n409 9.154
R1858 GND.n411 GND.n410 9.154
R1859 GND.n386 GND.n385 9.154
R1860 GND.n412 GND.n386 9.154
R1861 GND.n416 GND.n415 9.154
R1862 GND.n415 GND.n414 9.154
R1863 GND.n381 GND.n380 9.154
R1864 GND.n413 GND.n380 9.154
R1865 GND.n421 GND.n420 9.154
R1866 GND.n422 GND.n421 9.154
R1867 GND.n379 GND.n378 9.154
R1868 GND.n423 GND.n379 9.154
R1869 GND.n426 GND.n425 9.154
R1870 GND.n425 GND.n424 9.154
R1871 GND.n376 GND.n375 9.154
R1872 GND.n375 GND.n374 9.154
R1873 GND.n432 GND.n431 9.154
R1874 GND.n433 GND.n432 9.154
R1875 GND.n373 GND.n372 9.154
R1876 GND.n434 GND.n373 9.154
R1877 GND.n437 GND.n436 9.154
R1878 GND.n436 GND.n435 9.154
R1879 GND.n370 GND.n369 9.154
R1880 GND.n369 GND.n368 9.154
R1881 GND.n442 GND.n441 9.154
R1882 GND.n443 GND.n442 9.154
R1883 GND.n367 GND.n366 9.154
R1884 GND.n364 GND.n363 9.154
R1885 GND.n453 GND.n452 9.154
R1886 GND.n454 GND.n453 9.154
R1887 GND.n362 GND.n361 9.154
R1888 GND.n455 GND.n362 9.154
R1889 GND.n458 GND.n457 9.154
R1890 GND.n457 GND.n456 9.154
R1891 GND.n359 GND.n358 9.154
R1892 GND.n358 GND.n357 9.154
R1893 GND.n464 GND.n463 9.154
R1894 GND.n465 GND.n464 9.154
R1895 GND.n356 GND.n355 9.154
R1896 GND.n466 GND.n356 9.154
R1897 GND.n470 GND.n469 9.154
R1898 GND.n469 GND.n468 9.154
R1899 GND.n351 GND.n350 9.154
R1900 GND.n467 GND.n350 9.154
R1901 GND.n475 GND.n474 9.154
R1902 GND.n476 GND.n475 9.154
R1903 GND.n349 GND.n348 9.154
R1904 GND.n477 GND.n349 9.154
R1905 GND.n480 GND.n479 9.154
R1906 GND.n479 GND.n478 9.154
R1907 GND.n346 GND.n345 9.154
R1908 GND.n345 GND.n344 9.154
R1909 GND.n486 GND.n485 9.154
R1910 GND.n487 GND.n486 9.154
R1911 GND.n343 GND.n342 9.154
R1912 GND.n488 GND.n343 9.154
R1913 GND.n491 GND.n490 9.154
R1914 GND.n490 GND.n489 9.154
R1915 GND.n340 GND.n339 9.154
R1916 GND.n339 GND.n338 9.154
R1917 GND.n496 GND.n495 9.154
R1918 GND.n497 GND.n496 9.154
R1919 GND.n337 GND.n336 9.154
R1920 GND.n300 GND.n299 9.154
R1921 GND.n580 GND.n300 9.154
R1922 GND.n575 GND.n574 9.154
R1923 GND.n503 GND.n502 9.154
R1924 GND.n334 GND.n333 9.154
R1925 GND.n504 GND.n334 9.154
R1926 GND.n507 GND.n506 9.154
R1927 GND.n506 GND.n505 9.154
R1928 GND.n331 GND.n330 9.154
R1929 GND.n330 GND.n329 9.154
R1930 GND.n512 GND.n511 9.154
R1931 GND.n513 GND.n512 9.154
R1932 GND.n328 GND.n327 9.154
R1933 GND.n514 GND.n328 9.154
R1934 GND.n517 GND.n516 9.154
R1935 GND.n516 GND.n515 9.154
R1936 GND.n325 GND.n324 9.154
R1937 GND.n324 GND.n323 9.154
R1938 GND.n523 GND.n522 9.154
R1939 GND.n524 GND.n523 9.154
R1940 GND.n322 GND.n321 9.154
R1941 GND.n525 GND.n322 9.154
R1942 GND.n528 GND.n527 9.154
R1943 GND.n527 GND.n526 9.154
R1944 GND.n319 GND.n318 9.154
R1945 GND.n318 GND.n317 9.154
R1946 GND.n536 GND.n535 9.154
R1947 GND.n537 GND.n536 9.154
R1948 GND.n316 GND.n315 9.154
R1949 GND.n538 GND.n316 9.154
R1950 GND.n542 GND.n541 9.154
R1951 GND.n541 GND.n540 9.154
R1952 GND.n314 GND.n313 9.154
R1953 GND.n539 GND.n313 9.154
R1954 GND.n548 GND.n547 9.154
R1955 GND.n549 GND.n548 9.154
R1956 GND.n312 GND.n311 9.154
R1957 GND.n550 GND.n312 9.154
R1958 GND.n554 GND.n553 9.154
R1959 GND.n553 GND.n552 9.154
R1960 GND.n309 GND.n308 9.154
R1961 GND.n551 GND.n308 9.154
R1962 GND.n559 GND.n558 9.154
R1963 GND.n560 GND.n559 9.154
R1964 GND.n307 GND.n306 9.154
R1965 GND.n561 GND.n307 9.154
R1966 GND.n565 GND.n564 9.154
R1967 GND.n564 GND.n563 9.154
R1968 GND.n304 GND.n303 9.154
R1969 GND.n562 GND.n303 9.154
R1970 GND.n571 GND.n570 9.154
R1971 GND.n572 GND.n571 9.154
R1972 GND.n569 GND.n302 9.154
R1973 GND.n573 GND.n302 9.154
R1974 GND.n583 GND.n582 9.154
R1975 GND.n582 GND.n581 9.154
R1976 GND.n297 GND.n296 9.154
R1977 GND.n296 GND.n295 9.154
R1978 GND.n588 GND.n587 9.154
R1979 GND.n589 GND.n588 9.154
R1980 GND.n294 GND.n293 9.154
R1981 GND.n590 GND.n294 9.154
R1982 GND.n593 GND.n592 9.154
R1983 GND.n592 GND.n591 9.154
R1984 GND.n291 GND.n290 9.154
R1985 GND.n290 GND.n289 9.154
R1986 GND.n599 GND.n598 9.154
R1987 GND.n600 GND.n599 9.154
R1988 GND.n288 GND.n287 9.154
R1989 GND.n601 GND.n288 9.154
R1990 GND.n604 GND.n603 9.154
R1991 GND.n603 GND.n602 9.154
R1992 GND.n285 GND.n284 9.154
R1993 GND.n284 GND.n283 9.154
R1994 GND.n612 GND.n611 9.154
R1995 GND.n613 GND.n612 9.154
R1996 GND.n282 GND.n281 9.154
R1997 GND.n614 GND.n282 9.154
R1998 GND.n618 GND.n617 9.154
R1999 GND.n617 GND.n616 9.154
R2000 GND.n280 GND.n279 9.154
R2001 GND.n615 GND.n279 9.154
R2002 GND.n624 GND.n623 9.154
R2003 GND.n625 GND.n624 9.154
R2004 GND.n278 GND.n277 9.154
R2005 GND.n626 GND.n278 9.154
R2006 GND.n630 GND.n629 9.154
R2007 GND.n629 GND.n628 9.154
R2008 GND.n275 GND.n274 9.154
R2009 GND.n627 GND.n274 9.154
R2010 GND.n635 GND.n634 9.154
R2011 GND.n636 GND.n635 9.154
R2012 GND.n273 GND.n272 9.154
R2013 GND.n637 GND.n273 9.154
R2014 GND.n641 GND.n640 9.154
R2015 GND.n640 GND.n639 9.154
R2016 GND.n269 GND.n268 9.154
R2017 GND.n638 GND.n268 9.154
R2018 GND.n646 GND.n645 9.154
R2019 GND.n647 GND.n646 9.154
R2020 GND.n270 GND.n267 9.154
R2021 GND.n648 GND.n267 9.154
R2022 GND.n650 GND.n649 9.154
R2023 GND.n579 GND.n578 9.154
R2024 GND.n1798 GND.n1797 9.154
R2025 GND.n1797 GND.n1796 9.154
R2026 GND.n1567 GND.n1566 9.154
R2027 GND.n1602 GND.n1601 9.154
R2028 GND.n1601 GND.n1600 9.154
R2029 GND.n1592 GND.n1591 9.154
R2030 GND.n1598 GND.n1597 9.154
R2031 GND.n1597 GND.n1596 9.154
R2032 GND.n1610 GND.n1609 9.154
R2033 GND.n1609 GND.n1608 9.154
R2034 GND.n1618 GND.n1617 9.154
R2035 GND.n1617 GND.n1616 9.154
R2036 GND.n1626 GND.n1625 9.154
R2037 GND.n1625 GND.n1624 9.154
R2038 GND.n1634 GND.n1633 9.154
R2039 GND.n1633 GND.n1632 9.154
R2040 GND.n1642 GND.n1641 9.154
R2041 GND.n1641 GND.n1640 9.154
R2042 GND.n1651 GND.n1650 9.154
R2043 GND.n1650 GND.n1649 9.154
R2044 GND.n1659 GND.n1658 9.154
R2045 GND.n1658 GND.n1657 9.154
R2046 GND.n1579 GND.n1578 9.154
R2047 GND.n1578 GND.n1577 9.154
R2048 GND.n1585 GND.n1584 9.154
R2049 GND.n1584 GND.n1583 9.154
R2050 GND.n1672 GND.n1671 9.154
R2051 GND.n1671 GND.n1670 9.154
R2052 GND.n1572 GND.n1571 9.154
R2053 GND.n1571 GND.n1570 9.154
R2054 GND.n1683 GND.n1682 9.154
R2055 GND.n1682 GND.n1681 9.154
R2056 GND.n1689 GND.n1688 9.154
R2057 GND.n1688 GND.n1687 9.154
R2058 GND.n1697 GND.n1696 9.154
R2059 GND.n1696 GND.n1695 9.154
R2060 GND.n1705 GND.n1704 9.154
R2061 GND.n1704 GND.n1703 9.154
R2062 GND.n1714 GND.n1713 9.154
R2063 GND.n1713 GND.n1712 9.154
R2064 GND.n1722 GND.n1721 9.154
R2065 GND.n1721 GND.n1720 9.154
R2066 GND.n1730 GND.n1729 9.154
R2067 GND.n1729 GND.n1728 9.154
R2068 GND.n1738 GND.n1737 9.154
R2069 GND.n1737 GND.n1736 9.154
R2070 GND.n1746 GND.n1745 9.154
R2071 GND.n1745 GND.n1744 9.154
R2072 GND.n1754 GND.n1753 9.154
R2073 GND.n1753 GND.n1752 9.154
R2074 GND.n1763 GND.n1762 9.154
R2075 GND.n1762 GND.n1761 9.154
R2076 GND.n1768 GND.n1767 9.154
R2077 GND.n1606 GND.n1605 9.154
R2078 GND.n1605 GND.n1604 9.154
R2079 GND.n1614 GND.n1613 9.154
R2080 GND.n1613 GND.n1612 9.154
R2081 GND.n1622 GND.n1621 9.154
R2082 GND.n1621 GND.n1620 9.154
R2083 GND.n1630 GND.n1629 9.154
R2084 GND.n1629 GND.n1628 9.154
R2085 GND.n1638 GND.n1637 9.154
R2086 GND.n1637 GND.n1636 9.154
R2087 GND.n1646 GND.n1645 9.154
R2088 GND.n1645 GND.n1644 9.154
R2089 GND.n1655 GND.n1654 9.154
R2090 GND.n1654 GND.n1653 9.154
R2091 GND.n1663 GND.n1662 9.154
R2092 GND.n1662 GND.n1661 9.154
R2093 GND.n1582 GND.n1581 9.154
R2094 GND.n1581 GND.n1580 9.154
R2095 GND.n1669 GND.n1587 9.154
R2096 GND.n1587 GND.n1586 9.154
R2097 GND.n1676 GND.n1675 9.154
R2098 GND.n1675 GND.n1674 9.154
R2099 GND.n1575 GND.n1574 9.154
R2100 GND.n1574 GND.n1573 9.154
R2101 GND.n1686 GND.n1685 9.154
R2102 GND.n1685 GND.n1684 9.154
R2103 GND.n1693 GND.n1692 9.154
R2104 GND.n1692 GND.n1691 9.154
R2105 GND.n1701 GND.n1700 9.154
R2106 GND.n1700 GND.n1699 9.154
R2107 GND.n1709 GND.n1708 9.154
R2108 GND.n1708 GND.n1707 9.154
R2109 GND.n1718 GND.n1717 9.154
R2110 GND.n1717 GND.n1716 9.154
R2111 GND.n1726 GND.n1725 9.154
R2112 GND.n1725 GND.n1724 9.154
R2113 GND.n1734 GND.n1733 9.154
R2114 GND.n1733 GND.n1732 9.154
R2115 GND.n1742 GND.n1741 9.154
R2116 GND.n1741 GND.n1740 9.154
R2117 GND.n1750 GND.n1749 9.154
R2118 GND.n1749 GND.n1748 9.154
R2119 GND.n1758 GND.n1757 9.154
R2120 GND.n1757 GND.n1756 9.154
R2121 GND.n1807 GND.n1806 9.154
R2122 GND.n1806 GND.n1805 9.154
R2123 GND.n1815 GND.n1814 9.154
R2124 GND.n1814 GND.n1813 9.154
R2125 GND.n1823 GND.n1822 9.154
R2126 GND.n1822 GND.n1821 9.154
R2127 GND.n1565 GND.n1564 9.154
R2128 GND.n1564 GND.n1563 9.154
R2129 GND.n1832 GND.n1831 9.154
R2130 GND.n1831 GND.n1830 9.154
R2131 GND.n1555 GND.n1554 9.154
R2132 GND.n1554 GND.n1553 9.154
R2133 GND.n1843 GND.n1842 9.154
R2134 GND.n1842 GND.n1841 9.154
R2135 GND.n1850 GND.n1849 9.154
R2136 GND.n1849 GND.n1848 9.154
R2137 GND.n1859 GND.n1858 9.154
R2138 GND.n1858 GND.n1857 9.154
R2139 GND.n1867 GND.n1866 9.154
R2140 GND.n1866 GND.n1865 9.154
R2141 GND.n1876 GND.n1875 9.154
R2142 GND.n1875 GND.n1874 9.154
R2143 GND.n1884 GND.n1883 9.154
R2144 GND.n1883 GND.n1882 9.154
R2145 GND.n1891 GND.n1890 9.154
R2146 GND.n1890 GND.n1889 9.154
R2147 GND.n1897 GND.n1896 9.154
R2148 GND.n1790 GND.n1789 9.154
R2149 GND.n1781 GND.n1780 9.154
R2150 GND.n1787 GND.n1786 9.154
R2151 GND.n1786 GND.n1785 9.154
R2152 GND.n1794 GND.n1793 9.154
R2153 GND.n1793 GND.n1792 9.154
R2154 GND.n1802 GND.n1801 9.154
R2155 GND.n1801 GND.n1800 9.154
R2156 GND.n1811 GND.n1810 9.154
R2157 GND.n1810 GND.n1809 9.154
R2158 GND.n1819 GND.n1818 9.154
R2159 GND.n1818 GND.n1817 9.154
R2160 GND.n1562 GND.n1561 9.154
R2161 GND.n1561 GND.n1560 9.154
R2162 GND.n1829 GND.n1567 9.154
R2163 GND.n1836 GND.n1835 9.154
R2164 GND.n1835 GND.n1834 9.154
R2165 GND.n1558 GND.n1557 9.154
R2166 GND.n1557 GND.n1556 9.154
R2167 GND.n1846 GND.n1845 9.154
R2168 GND.n1845 GND.n1844 9.154
R2169 GND.n1855 GND.n1854 9.154
R2170 GND.n1854 GND.n1853 9.154
R2171 GND.n1863 GND.n1862 9.154
R2172 GND.n1862 GND.n1861 9.154
R2173 GND.n1871 GND.n1870 9.154
R2174 GND.n1870 GND.n1869 9.154
R2175 GND.n1880 GND.n1879 9.154
R2176 GND.n1879 GND.n1878 9.154
R2177 GND.n1887 GND.n1886 9.154
R2178 GND.n1923 GND.n1922 9.154
R2179 GND.n1922 GND.n1921 9.154
R2180 GND.n1931 GND.n1930 9.154
R2181 GND.n1930 GND.n1929 9.154
R2182 GND.n1939 GND.n1938 9.154
R2183 GND.n1938 GND.n1937 9.154
R2184 GND.n1947 GND.n1946 9.154
R2185 GND.n1946 GND.n1945 9.154
R2186 GND.n1955 GND.n1954 9.154
R2187 GND.n1954 GND.n1953 9.154
R2188 GND.n1963 GND.n1962 9.154
R2189 GND.n1962 GND.n1961 9.154
R2190 GND.n1971 GND.n1970 9.154
R2191 GND.n1970 GND.n1969 9.154
R2192 GND.n1979 GND.n1978 9.154
R2193 GND.n1978 GND.n1977 9.154
R2194 GND.n1988 GND.n1987 9.154
R2195 GND.n1987 GND.n1986 9.154
R2196 GND.n1997 GND.n1996 9.154
R2197 GND.n1996 GND.n1995 9.154
R2198 GND.n2005 GND.n2004 9.154
R2199 GND.n2004 GND.n2003 9.154
R2200 GND.n1547 GND.n1546 9.154
R2201 GND.n1546 GND.n1545 9.154
R2202 GND.n2013 GND.n2012 9.154
R2203 GND.n2012 GND.n2011 9.154
R2204 GND.n2020 GND.n2019 9.154
R2205 GND.n2019 GND.n2018 9.154
R2206 GND.n2028 GND.n2027 9.154
R2207 GND.n2027 GND.n2026 9.154
R2208 GND.n2036 GND.n2035 9.154
R2209 GND.n2035 GND.n2034 9.154
R2210 GND.n2046 GND.n2045 9.154
R2211 GND.n2045 GND.n2044 9.154
R2212 GND.n2054 GND.n2053 9.154
R2213 GND.n2053 GND.n2052 9.154
R2214 GND.n2062 GND.n2061 9.154
R2215 GND.n2061 GND.n2060 9.154
R2216 GND.n2070 GND.n2069 9.154
R2217 GND.n2069 GND.n2068 9.154
R2218 GND.n2078 GND.n2077 9.154
R2219 GND.n2077 GND.n2076 9.154
R2220 GND.n2086 GND.n2085 9.154
R2221 GND.n2085 GND.n2084 9.154
R2222 GND.n2094 GND.n2093 9.154
R2223 GND.n2093 GND.n2092 9.154
R2224 GND.n2102 GND.n2101 9.154
R2225 GND.n2101 GND.n2100 9.154
R2226 GND.n1538 GND.n1537 9.154
R2227 GND.n1537 GND.n1536 9.154
R2228 GND.n1904 GND.n1903 9.154
R2229 GND.n1912 GND.n1911 9.154
R2230 GND.n1911 GND.n1910 9.154
R2231 GND.n1919 GND.n1918 9.154
R2232 GND.n1918 GND.n1917 9.154
R2233 GND.n1927 GND.n1926 9.154
R2234 GND.n1926 GND.n1925 9.154
R2235 GND.n1935 GND.n1934 9.154
R2236 GND.n1934 GND.n1933 9.154
R2237 GND.n1943 GND.n1942 9.154
R2238 GND.n1942 GND.n1941 9.154
R2239 GND.n1951 GND.n1950 9.154
R2240 GND.n1950 GND.n1949 9.154
R2241 GND.n1959 GND.n1958 9.154
R2242 GND.n1958 GND.n1957 9.154
R2243 GND.n1967 GND.n1966 9.154
R2244 GND.n1966 GND.n1965 9.154
R2245 GND.n1975 GND.n1974 9.154
R2246 GND.n1974 GND.n1973 9.154
R2247 GND.n1983 GND.n1982 9.154
R2248 GND.n1982 GND.n1981 9.154
R2249 GND.n1993 GND.n1992 9.154
R2250 GND.n1992 GND.n1991 9.154
R2251 GND.n2001 GND.n2000 9.154
R2252 GND.n2000 GND.n1999 9.154
R2253 GND.n1544 GND.n1543 9.154
R2254 GND.n1543 GND.n1542 9.154
R2255 GND.n1550 GND.n1549 9.154
R2256 GND.n1549 GND.n1548 9.154
R2257 GND.n2016 GND.n2015 9.154
R2258 GND.n2015 GND.n2014 9.154
R2259 GND.n2024 GND.n2023 9.154
R2260 GND.n2023 GND.n2022 9.154
R2261 GND.n2032 GND.n2031 9.154
R2262 GND.n2031 GND.n2030 9.154
R2263 GND.n2041 GND.n2040 9.154
R2264 GND.n2040 GND.n2039 9.154
R2265 GND.n2050 GND.n2049 9.154
R2266 GND.n2049 GND.n2048 9.154
R2267 GND.n2058 GND.n2057 9.154
R2268 GND.n2057 GND.n2056 9.154
R2269 GND.n2066 GND.n2065 9.154
R2270 GND.n2065 GND.n2064 9.154
R2271 GND.n2074 GND.n2073 9.154
R2272 GND.n2073 GND.n2072 9.154
R2273 GND.n2082 GND.n2081 9.154
R2274 GND.n2081 GND.n2080 9.154
R2275 GND.n2090 GND.n2089 9.154
R2276 GND.n2089 GND.n2088 9.154
R2277 GND.n2098 GND.n2097 9.154
R2278 GND.n2097 GND.n2096 9.154
R2279 GND.n2106 GND.n2105 9.154
R2280 GND.n2105 GND.n2104 9.154
R2281 GND.n1541 GND.n1540 9.154
R2282 GND.n1361 GND.n1360 9.154
R2283 GND.n1366 GND.n1365 9.154
R2284 GND.n1367 GND.n1366 9.154
R2285 GND.n1359 GND.n1358 9.154
R2286 GND.n1368 GND.n1359 9.154
R2287 GND.n1372 GND.n1371 9.154
R2288 GND.n1371 GND.n1370 9.154
R2289 GND.n1356 GND.n1355 9.154
R2290 GND.n1369 GND.n1355 9.154
R2291 GND.n1377 GND.n1376 9.154
R2292 GND.n1378 GND.n1377 9.154
R2293 GND.n1354 GND.n1353 9.154
R2294 GND.n1379 GND.n1354 9.154
R2295 GND.n1383 GND.n1382 9.154
R2296 GND.n1382 GND.n1381 9.154
R2297 GND.n1351 GND.n1350 9.154
R2298 GND.n1380 GND.n1350 9.154
R2299 GND.n1389 GND.n1388 9.154
R2300 GND.n1390 GND.n1389 9.154
R2301 GND.n1349 GND.n1348 9.154
R2302 GND.n1391 GND.n1349 9.154
R2303 GND.n1394 GND.n1393 9.154
R2304 GND.n1393 GND.n1392 9.154
R2305 GND.n1345 GND.n1344 9.154
R2306 GND.n1344 GND.n1343 9.154
R2307 GND.n1400 GND.n1399 9.154
R2308 GND.n1401 GND.n1400 9.154
R2309 GND.n1342 GND.n1341 9.154
R2310 GND.n1402 GND.n1342 9.154
R2311 GND.n1405 GND.n1404 9.154
R2312 GND.n1404 GND.n1403 9.154
R2313 GND.n1339 GND.n1338 9.154
R2314 GND.n1338 GND.n1337 9.154
R2315 GND.n1410 GND.n1409 9.154
R2316 GND.n1411 GND.n1410 9.154
R2317 GND.n1336 GND.n1335 9.154
R2318 GND.n1412 GND.n1336 9.154
R2319 GND.n1415 GND.n1414 9.154
R2320 GND.n1414 GND.n1413 9.154
R2321 GND.n1333 GND.n1332 9.154
R2322 GND.n1332 GND.n1331 9.154
R2323 GND.n1420 GND.n1419 9.154
R2324 GND.n1421 GND.n1420 9.154
R2325 GND.n1330 GND.n1329 9.154
R2326 GND.n1327 GND.n1326 9.154
R2327 GND.n1431 GND.n1430 9.154
R2328 GND.n1432 GND.n1431 9.154
R2329 GND.n1325 GND.n1324 9.154
R2330 GND.n1433 GND.n1325 9.154
R2331 GND.n1437 GND.n1436 9.154
R2332 GND.n1436 GND.n1435 9.154
R2333 GND.n1322 GND.n1321 9.154
R2334 GND.n1434 GND.n1321 9.154
R2335 GND.n1443 GND.n1442 9.154
R2336 GND.n1444 GND.n1443 9.154
R2337 GND.n1320 GND.n1319 9.154
R2338 GND.n1445 GND.n1320 9.154
R2339 GND.n1448 GND.n1447 9.154
R2340 GND.n1447 GND.n1446 9.154
R2341 GND.n1316 GND.n1315 9.154
R2342 GND.n1315 GND.n1314 9.154
R2343 GND.n1454 GND.n1453 9.154
R2344 GND.n1455 GND.n1454 9.154
R2345 GND.n1313 GND.n1312 9.154
R2346 GND.n1456 GND.n1313 9.154
R2347 GND.n1459 GND.n1458 9.154
R2348 GND.n1458 GND.n1457 9.154
R2349 GND.n1310 GND.n1309 9.154
R2350 GND.n1309 GND.n1308 9.154
R2351 GND.n1464 GND.n1463 9.154
R2352 GND.n1465 GND.n1464 9.154
R2353 GND.n1307 GND.n1306 9.154
R2354 GND.n1304 GND.n1303 9.154
R2355 GND.n1475 GND.n1474 9.154
R2356 GND.n1476 GND.n1475 9.154
R2357 GND.n1302 GND.n1301 9.154
R2358 GND.n1477 GND.n1302 9.154
R2359 GND.n1481 GND.n1480 9.154
R2360 GND.n1480 GND.n1479 9.154
R2361 GND.n1299 GND.n1298 9.154
R2362 GND.n1478 GND.n1298 9.154
R2363 GND.n1486 GND.n1485 9.154
R2364 GND.n1487 GND.n1486 9.154
R2365 GND.n1297 GND.n1296 9.154
R2366 GND.n1488 GND.n1297 9.154
R2367 GND.n1492 GND.n1491 9.154
R2368 GND.n1491 GND.n1490 9.154
R2369 GND.n1294 GND.n1293 9.154
R2370 GND.n1489 GND.n1293 9.154
R2371 GND.n1498 GND.n1497 9.154
R2372 GND.n1499 GND.n1498 9.154
R2373 GND.n1292 GND.n1291 9.154
R2374 GND.n1500 GND.n1292 9.154
R2375 GND.n1503 GND.n1502 9.154
R2376 GND.n1502 GND.n1501 9.154
R2377 GND.n1288 GND.n1287 9.154
R2378 GND.n1287 GND.n1286 9.154
R2379 GND.n1509 GND.n1508 9.154
R2380 GND.n1510 GND.n1509 9.154
R2381 GND.n1285 GND.n1284 9.154
R2382 GND.n1511 GND.n1285 9.154
R2383 GND.n1514 GND.n1513 9.154
R2384 GND.n1513 GND.n1512 9.154
R2385 GND.n1282 GND.n1281 9.154
R2386 GND.n1281 GND.n1280 9.154
R2387 GND.n1519 GND.n1518 9.154
R2388 GND.n1520 GND.n1519 9.154
R2389 GND.n1279 GND.n1278 9.154
R2390 GND.n1521 GND.n1279 9.154
R2391 GND.n1524 GND.n1523 9.154
R2392 GND.n1523 GND.n1522 9.154
R2393 GND.n1276 GND.n1275 9.154
R2394 GND.n1275 GND.n1274 9.154
R2395 GND.n1530 GND.n1529 9.154
R2396 GND.n1531 GND.n1530 9.154
R2397 GND.n1528 GND.n1273 9.154
R2398 GND.n1100 GND.n1099 9.154
R2399 GND.n1105 GND.n1104 9.154
R2400 GND.n1106 GND.n1105 9.154
R2401 GND.n1098 GND.n1097 9.154
R2402 GND.n1107 GND.n1098 9.154
R2403 GND.n1110 GND.n1109 9.154
R2404 GND.n1109 GND.n1108 9.154
R2405 GND.n1095 GND.n1094 9.154
R2406 GND.n1094 GND.n1093 9.154
R2407 GND.n1116 GND.n1115 9.154
R2408 GND.n1117 GND.n1116 9.154
R2409 GND.n1092 GND.n1091 9.154
R2410 GND.n1118 GND.n1092 9.154
R2411 GND.n1122 GND.n1121 9.154
R2412 GND.n1121 GND.n1120 9.154
R2413 GND.n1087 GND.n1086 9.154
R2414 GND.n1119 GND.n1086 9.154
R2415 GND.n1127 GND.n1126 9.154
R2416 GND.n1128 GND.n1127 9.154
R2417 GND.n1085 GND.n1084 9.154
R2418 GND.n1129 GND.n1085 9.154
R2419 GND.n1132 GND.n1131 9.154
R2420 GND.n1131 GND.n1130 9.154
R2421 GND.n1082 GND.n1081 9.154
R2422 GND.n1081 GND.n1080 9.154
R2423 GND.n1138 GND.n1137 9.154
R2424 GND.n1139 GND.n1138 9.154
R2425 GND.n1079 GND.n1078 9.154
R2426 GND.n1140 GND.n1079 9.154
R2427 GND.n1143 GND.n1142 9.154
R2428 GND.n1142 GND.n1141 9.154
R2429 GND.n1076 GND.n1075 9.154
R2430 GND.n1075 GND.n1074 9.154
R2431 GND.n1148 GND.n1147 9.154
R2432 GND.n1149 GND.n1148 9.154
R2433 GND.n1073 GND.n1072 9.154
R2434 GND.n1070 GND.n1069 9.154
R2435 GND.n1159 GND.n1158 9.154
R2436 GND.n1160 GND.n1159 9.154
R2437 GND.n1068 GND.n1067 9.154
R2438 GND.n1161 GND.n1068 9.154
R2439 GND.n1165 GND.n1164 9.154
R2440 GND.n1164 GND.n1163 9.154
R2441 GND.n1065 GND.n1064 9.154
R2442 GND.n1162 GND.n1064 9.154
R2443 GND.n1171 GND.n1170 9.154
R2444 GND.n1172 GND.n1171 9.154
R2445 GND.n1063 GND.n1062 9.154
R2446 GND.n1173 GND.n1063 9.154
R2447 GND.n1176 GND.n1175 9.154
R2448 GND.n1175 GND.n1174 9.154
R2449 GND.n1058 GND.n1057 9.154
R2450 GND.n1057 GND.n1056 9.154
R2451 GND.n1182 GND.n1181 9.154
R2452 GND.n1183 GND.n1182 9.154
R2453 GND.n1055 GND.n1054 9.154
R2454 GND.n1184 GND.n1055 9.154
R2455 GND.n1187 GND.n1186 9.154
R2456 GND.n1186 GND.n1185 9.154
R2457 GND.n1052 GND.n1051 9.154
R2458 GND.n1051 GND.n1050 9.154
R2459 GND.n1192 GND.n1191 9.154
R2460 GND.n1193 GND.n1192 9.154
R2461 GND.n1049 GND.n1048 9.154
R2462 GND.n1271 GND.n1270 9.154
R2463 GND.n1199 GND.n1198 9.154
R2464 GND.n1046 GND.n1045 9.154
R2465 GND.n1200 GND.n1046 9.154
R2466 GND.n1203 GND.n1202 9.154
R2467 GND.n1202 GND.n1201 9.154
R2468 GND.n1043 GND.n1042 9.154
R2469 GND.n1042 GND.n1041 9.154
R2470 GND.n1208 GND.n1207 9.154
R2471 GND.n1209 GND.n1208 9.154
R2472 GND.n1040 GND.n1039 9.154
R2473 GND.n1210 GND.n1040 9.154
R2474 GND.n1213 GND.n1212 9.154
R2475 GND.n1212 GND.n1211 9.154
R2476 GND.n1037 GND.n1036 9.154
R2477 GND.n1036 GND.n1035 9.154
R2478 GND.n1219 GND.n1218 9.154
R2479 GND.n1220 GND.n1219 9.154
R2480 GND.n1034 GND.n1033 9.154
R2481 GND.n1221 GND.n1034 9.154
R2482 GND.n1224 GND.n1223 9.154
R2483 GND.n1223 GND.n1222 9.154
R2484 GND.n1031 GND.n1030 9.154
R2485 GND.n1030 GND.n1029 9.154
R2486 GND.n1232 GND.n1231 9.154
R2487 GND.n1233 GND.n1232 9.154
R2488 GND.n1028 GND.n1027 9.154
R2489 GND.n1234 GND.n1028 9.154
R2490 GND.n1238 GND.n1237 9.154
R2491 GND.n1237 GND.n1236 9.154
R2492 GND.n1026 GND.n1025 9.154
R2493 GND.n1235 GND.n1025 9.154
R2494 GND.n1244 GND.n1243 9.154
R2495 GND.n1245 GND.n1244 9.154
R2496 GND.n1024 GND.n1023 9.154
R2497 GND.n1246 GND.n1024 9.154
R2498 GND.n1250 GND.n1249 9.154
R2499 GND.n1249 GND.n1248 9.154
R2500 GND.n1021 GND.n1020 9.154
R2501 GND.n1247 GND.n1020 9.154
R2502 GND.n1255 GND.n1254 9.154
R2503 GND.n1256 GND.n1255 9.154
R2504 GND.n1019 GND.n1018 9.154
R2505 GND.n1257 GND.n1019 9.154
R2506 GND.n1261 GND.n1260 9.154
R2507 GND.n1260 GND.n1259 9.154
R2508 GND.n1016 GND.n1015 9.154
R2509 GND.n1258 GND.n1015 9.154
R2510 GND.n1267 GND.n1266 9.154
R2511 GND.n1268 GND.n1267 9.154
R2512 GND.n1265 GND.n1014 9.154
R2513 GND.n1269 GND.n1014 9.154
R2514 GND.n771 GND.n770 9.154
R2515 GND.n775 GND.n774 9.154
R2516 GND.n774 GND.n773 9.154
R2517 GND.n779 GND.n778 9.154
R2518 GND.n778 GND.n777 9.154
R2519 GND.n783 GND.n782 9.154
R2520 GND.n782 GND.n781 9.154
R2521 GND.n787 GND.n786 9.154
R2522 GND.n786 GND.n785 9.154
R2523 GND.n791 GND.n790 9.154
R2524 GND.n790 GND.n789 9.154
R2525 GND.n796 GND.n795 9.154
R2526 GND.n795 GND.n794 9.154
R2527 GND.n800 GND.n799 9.154
R2528 GND.n799 GND.n798 9.154
R2529 GND.n804 GND.n803 9.154
R2530 GND.n803 GND.n802 9.154
R2531 GND.n807 GND.n766 9.154
R2532 GND.n766 GND.n765 9.154
R2533 GND.n810 GND.n809 9.154
R2534 GND.n809 GND.n808 9.154
R2535 GND.n814 GND.n813 9.154
R2536 GND.n813 GND.n812 9.154
R2537 GND.n818 GND.n817 9.154
R2538 GND.n817 GND.n816 9.154
R2539 GND.n823 GND.n822 9.154
R2540 GND.n822 GND.n821 9.154
R2541 GND.n827 GND.n826 9.154
R2542 GND.n826 GND.n825 9.154
R2543 GND.n831 GND.n830 9.154
R2544 GND.n830 GND.n829 9.154
R2545 GND.n835 GND.n834 9.154
R2546 GND.n834 GND.n833 9.154
R2547 GND.n839 GND.n838 9.154
R2548 GND.n838 GND.n837 9.154
R2549 GND.n843 GND.n842 9.154
R2550 GND.n851 GND.n850 9.154
R2551 GND.n855 GND.n854 9.154
R2552 GND.n854 GND.n853 9.154
R2553 GND.n859 GND.n858 9.154
R2554 GND.n858 GND.n857 9.154
R2555 GND.n863 GND.n862 9.154
R2556 GND.n862 GND.n861 9.154
R2557 GND.n868 GND.n867 9.154
R2558 GND.n867 GND.n866 9.154
R2559 GND.n872 GND.n871 9.154
R2560 GND.n871 GND.n870 9.154
R2561 GND.n876 GND.n875 9.154
R2562 GND.n875 GND.n874 9.154
R2563 GND.n879 GND.n762 9.154
R2564 GND.n762 GND.n761 9.154
R2565 GND.n882 GND.n881 9.154
R2566 GND.n881 GND.n880 9.154
R2567 GND.n886 GND.n885 9.154
R2568 GND.n885 GND.n884 9.154
R2569 GND.n890 GND.n889 9.154
R2570 GND.n889 GND.n888 9.154
R2571 GND.n895 GND.n894 9.154
R2572 GND.n894 GND.n893 9.154
R2573 GND.n899 GND.n898 9.154
R2574 GND.n898 GND.n897 9.154
R2575 GND.n903 GND.n902 9.154
R2576 GND.n902 GND.n901 9.154
R2577 GND.n907 GND.n906 9.154
R2578 GND.n1012 GND.n1011 9.154
R2579 GND.n912 GND.n911 9.154
R2580 GND.n916 GND.n915 9.154
R2581 GND.n915 GND.n914 9.154
R2582 GND.n920 GND.n919 9.154
R2583 GND.n919 GND.n918 9.154
R2584 GND.n924 GND.n923 9.154
R2585 GND.n923 GND.n922 9.154
R2586 GND.n928 GND.n927 9.154
R2587 GND.n927 GND.n926 9.154
R2588 GND.n932 GND.n931 9.154
R2589 GND.n931 GND.n930 9.154
R2590 GND.n936 GND.n935 9.154
R2591 GND.n935 GND.n934 9.154
R2592 GND.n940 GND.n939 9.154
R2593 GND.n939 GND.n938 9.154
R2594 GND.n944 GND.n943 9.154
R2595 GND.n943 GND.n942 9.154
R2596 GND.n948 GND.n947 9.154
R2597 GND.n947 GND.n946 9.154
R2598 GND.n953 GND.n952 9.154
R2599 GND.n952 GND.n951 9.154
R2600 GND.n957 GND.n956 9.154
R2601 GND.n956 GND.n955 9.154
R2602 GND.n961 GND.n960 9.154
R2603 GND.n960 GND.n959 9.154
R2604 GND.n964 GND.n758 9.154
R2605 GND.n758 GND.n757 9.154
R2606 GND.n967 GND.n966 9.154
R2607 GND.n966 GND.n965 9.154
R2608 GND.n971 GND.n970 9.154
R2609 GND.n970 GND.n969 9.154
R2610 GND.n975 GND.n974 9.154
R2611 GND.n974 GND.n973 9.154
R2612 GND.n980 GND.n979 9.154
R2613 GND.n979 GND.n978 9.154
R2614 GND.n984 GND.n983 9.154
R2615 GND.n983 GND.n982 9.154
R2616 GND.n988 GND.n987 9.154
R2617 GND.n987 GND.n986 9.154
R2618 GND.n992 GND.n991 9.154
R2619 GND.n991 GND.n990 9.154
R2620 GND.n996 GND.n995 9.154
R2621 GND.n995 GND.n994 9.154
R2622 GND.n1000 GND.n999 9.154
R2623 GND.n999 GND.n998 9.154
R2624 GND.n1004 GND.n1003 9.154
R2625 GND.n1003 GND.n1002 9.154
R2626 GND.n1008 GND.n1007 9.154
R2627 GND.n1007 GND.n1006 9.154
R2628 GND.n756 GND.n755 9.154
R2629 GND.n755 GND.n754 9.154
R2630 GND.n258 GND.n257 9.154
R2631 GND.n162 GND.n161 9.154
R2632 GND.n161 GND.n160 9.154
R2633 GND.n166 GND.n165 9.154
R2634 GND.n165 GND.n164 9.154
R2635 GND.n170 GND.n169 9.154
R2636 GND.n169 GND.n168 9.154
R2637 GND.n174 GND.n173 9.154
R2638 GND.n173 GND.n172 9.154
R2639 GND.n178 GND.n177 9.154
R2640 GND.n177 GND.n176 9.154
R2641 GND.n182 GND.n181 9.154
R2642 GND.n181 GND.n180 9.154
R2643 GND.n186 GND.n185 9.154
R2644 GND.n185 GND.n184 9.154
R2645 GND.n190 GND.n189 9.154
R2646 GND.n189 GND.n188 9.154
R2647 GND.n194 GND.n193 9.154
R2648 GND.n193 GND.n192 9.154
R2649 GND.n199 GND.n198 9.154
R2650 GND.n198 GND.n197 9.154
R2651 GND.n203 GND.n202 9.154
R2652 GND.n202 GND.n201 9.154
R2653 GND.n207 GND.n206 9.154
R2654 GND.n206 GND.n205 9.154
R2655 GND.n210 GND.n4 9.154
R2656 GND.n4 GND.n3 9.154
R2657 GND.n213 GND.n212 9.154
R2658 GND.n212 GND.n211 9.154
R2659 GND.n217 GND.n216 9.154
R2660 GND.n216 GND.n215 9.154
R2661 GND.n221 GND.n220 9.154
R2662 GND.n220 GND.n219 9.154
R2663 GND.n226 GND.n225 9.154
R2664 GND.n225 GND.n224 9.154
R2665 GND.n230 GND.n229 9.154
R2666 GND.n229 GND.n228 9.154
R2667 GND.n234 GND.n233 9.154
R2668 GND.n233 GND.n232 9.154
R2669 GND.n238 GND.n237 9.154
R2670 GND.n237 GND.n236 9.154
R2671 GND.n242 GND.n241 9.154
R2672 GND.n241 GND.n240 9.154
R2673 GND.n246 GND.n245 9.154
R2674 GND.n245 GND.n244 9.154
R2675 GND.n250 GND.n249 9.154
R2676 GND.n249 GND.n248 9.154
R2677 GND.n254 GND.n253 9.154
R2678 GND.n253 GND.n252 9.154
R2679 GND.n2 GND.n1 9.154
R2680 GND.n1 GND.n0 9.154
R2681 GND.n158 GND.n157 9.154
R2682 GND.n652 GND.n651 9.154
R2683 GND.n751 GND.n750 9.154
R2684 GND.n261 GND.n260 9.154
R2685 GND.n260 GND.n259 9.154
R2686 GND.n747 GND.n746 9.154
R2687 GND.n746 GND.n745 9.154
R2688 GND.n743 GND.n742 9.154
R2689 GND.n742 GND.n741 9.154
R2690 GND.n739 GND.n738 9.154
R2691 GND.n738 GND.n737 9.154
R2692 GND.n735 GND.n734 9.154
R2693 GND.n734 GND.n733 9.154
R2694 GND.n731 GND.n730 9.154
R2695 GND.n730 GND.n729 9.154
R2696 GND.n727 GND.n726 9.154
R2697 GND.n726 GND.n725 9.154
R2698 GND.n723 GND.n722 9.154
R2699 GND.n722 GND.n721 9.154
R2700 GND.n719 GND.n718 9.154
R2701 GND.n718 GND.n717 9.154
R2702 GND.n714 GND.n713 9.154
R2703 GND.n713 GND.n712 9.154
R2704 GND.n710 GND.n709 9.154
R2705 GND.n709 GND.n708 9.154
R2706 GND.n706 GND.n705 9.154
R2707 GND.n705 GND.n704 9.154
R2708 GND.n702 GND.n265 9.154
R2709 GND.n265 GND.n264 9.154
R2710 GND.n701 GND.n700 9.154
R2711 GND.n700 GND.n699 9.154
R2712 GND.n696 GND.n695 9.154
R2713 GND.n695 GND.n694 9.154
R2714 GND.n692 GND.n691 9.154
R2715 GND.n691 GND.n690 9.154
R2716 GND.n687 GND.n686 9.154
R2717 GND.n686 GND.n685 9.154
R2718 GND.n683 GND.n682 9.154
R2719 GND.n682 GND.n681 9.154
R2720 GND.n679 GND.n678 9.154
R2721 GND.n678 GND.n677 9.154
R2722 GND.n675 GND.n674 9.154
R2723 GND.n674 GND.n673 9.154
R2724 GND.n671 GND.n670 9.154
R2725 GND.n670 GND.n669 9.154
R2726 GND.n667 GND.n666 9.154
R2727 GND.n666 GND.n665 9.154
R2728 GND.n663 GND.n662 9.154
R2729 GND.n662 GND.n661 9.154
R2730 GND.n659 GND.n658 9.154
R2731 GND.n658 GND.n657 9.154
R2732 GND.n655 GND.n654 9.154
R2733 GND.n654 GND.n653 9.154
R2734 GND.n1591 GND.n1590 8.202
R2735 GND.n703 GND.n263 5.103
R2736 GND.n703 GND.n262 5.103
R2737 GND.n209 GND.n6 5.103
R2738 GND.n209 GND.n5 5.103
R2739 GND.n124 GND.n10 5.103
R2740 GND.n124 GND.n9 5.103
R2741 GND.n52 GND.n14 5.103
R2742 GND.n52 GND.n13 5.103
R2743 GND.n609 GND.n608 5.103
R2744 GND.n609 GND.n607 5.103
R2745 GND.n533 GND.n532 5.103
R2746 GND.n533 GND.n531 5.103
R2747 GND.n473 GND.n353 5.103
R2748 GND.n473 GND.n352 5.103
R2749 GND.n419 GND.n383 5.103
R2750 GND.n419 GND.n382 5.103
R2751 GND.n2009 GND.n1552 5.103
R2752 GND.n2010 GND.n1551 5.103
R2753 GND.n1828 GND.n1568 5.103
R2754 GND.n1840 GND.n1559 5.103
R2755 GND.n1668 GND.n1588 5.103
R2756 GND.n1680 GND.n1576 5.103
R2757 GND.n1504 GND.n1289 5.103
R2758 GND.n1449 GND.n1317 5.103
R2759 GND.n1395 GND.n1346 5.103
R2760 GND.n1229 GND.n1228 5.103
R2761 GND.n1229 GND.n1227 5.103
R2762 GND.n1177 GND.n1060 5.103
R2763 GND.n1177 GND.n1059 5.103
R2764 GND.n1125 GND.n1089 5.103
R2765 GND.n1125 GND.n1088 5.103
R2766 GND.n963 GND.n760 5.103
R2767 GND.n963 GND.n759 5.103
R2768 GND.n878 GND.n764 5.103
R2769 GND.n878 GND.n763 5.103
R2770 GND.n806 GND.n768 5.103
R2771 GND.n806 GND.n767 5.103
R2772 GND.n1585 GND.n1582 4.72
R2773 GND.n1672 GND.n1669 4.72
R2774 GND.n1683 GND.n1575 4.72
R2775 GND.n1689 GND.n1686 4.72
R2776 GND.n22 GND.n21 4.65
R2777 GND.n26 GND.n25 4.65
R2778 GND.n30 GND.n29 4.65
R2779 GND.n34 GND.n33 4.65
R2780 GND.n38 GND.n37 4.65
R2781 GND.n43 GND.n42 4.65
R2782 GND.n47 GND.n46 4.65
R2783 GND.n51 GND.n50 4.65
R2784 GND.n53 GND.n52 4.65
R2785 GND.n57 GND.n56 4.65
R2786 GND.n61 GND.n60 4.65
R2787 GND.n65 GND.n64 4.65
R2788 GND.n70 GND.n69 4.65
R2789 GND.n74 GND.n73 4.65
R2790 GND.n78 GND.n77 4.65
R2791 GND.n82 GND.n81 4.65
R2792 GND.n86 GND.n85 4.65
R2793 GND.n90 GND.n89 4.65
R2794 GND.n92 GND.n91 4.65
R2795 GND.n94 GND.n93 4.65
R2796 GND.n98 GND.n97 4.65
R2797 GND.n102 GND.n101 4.65
R2798 GND.n106 GND.n105 4.65
R2799 GND.n110 GND.n109 4.65
R2800 GND.n115 GND.n114 4.65
R2801 GND.n119 GND.n118 4.65
R2802 GND.n123 GND.n122 4.65
R2803 GND.n125 GND.n124 4.65
R2804 GND.n129 GND.n128 4.65
R2805 GND.n133 GND.n132 4.65
R2806 GND.n137 GND.n136 4.65
R2807 GND.n142 GND.n141 4.65
R2808 GND.n146 GND.n145 4.65
R2809 GND.n150 GND.n149 4.65
R2810 GND.n154 GND.n153 4.65
R2811 GND.n156 GND.n155 4.65
R2812 GND.n398 GND.n397 4.65
R2813 GND.n391 GND.n390 4.65
R2814 GND.n405 GND.n404 4.65
R2815 GND.n406 GND.n389 4.65
R2816 GND.n409 GND.n408 4.65
R2817 GND.n385 GND.n384 4.65
R2818 GND.n417 GND.n416 4.65
R2819 GND.n418 GND.n381 4.65
R2820 GND.n420 GND.n419 4.65
R2821 GND.n378 GND.n377 4.65
R2822 GND.n427 GND.n426 4.65
R2823 GND.n428 GND.n376 4.65
R2824 GND.n431 GND.n430 4.65
R2825 GND.n372 GND.n371 4.65
R2826 GND.n438 GND.n437 4.65
R2827 GND.n439 GND.n370 4.65
R2828 GND.n441 GND.n440 4.65
R2829 GND.n366 GND.n365 4.65
R2830 GND.n446 GND.n445 4.65
R2831 GND.n449 GND.n448 4.65
R2832 GND.n450 GND.n364 4.65
R2833 GND.n452 GND.n451 4.65
R2834 GND.n361 GND.n360 4.65
R2835 GND.n459 GND.n458 4.65
R2836 GND.n460 GND.n359 4.65
R2837 GND.n463 GND.n462 4.65
R2838 GND.n355 GND.n354 4.65
R2839 GND.n471 GND.n470 4.65
R2840 GND.n472 GND.n351 4.65
R2841 GND.n474 GND.n473 4.65
R2842 GND.n348 GND.n347 4.65
R2843 GND.n481 GND.n480 4.65
R2844 GND.n482 GND.n346 4.65
R2845 GND.n485 GND.n484 4.65
R2846 GND.n342 GND.n341 4.65
R2847 GND.n492 GND.n491 4.65
R2848 GND.n493 GND.n340 4.65
R2849 GND.n495 GND.n494 4.65
R2850 GND.n336 GND.n335 4.65
R2851 GND.n500 GND.n499 4.65
R2852 GND.n502 GND.n501 4.65
R2853 GND.n333 GND.n332 4.65
R2854 GND.n508 GND.n507 4.65
R2855 GND.n509 GND.n331 4.65
R2856 GND.n511 GND.n510 4.65
R2857 GND.n327 GND.n326 4.65
R2858 GND.n518 GND.n517 4.65
R2859 GND.n519 GND.n325 4.65
R2860 GND.n522 GND.n521 4.65
R2861 GND.n520 GND.n321 4.65
R2862 GND.n529 GND.n528 4.65
R2863 GND.n530 GND.n319 4.65
R2864 GND.n535 GND.n534 4.65
R2865 GND.n533 GND.n315 4.65
R2866 GND.n543 GND.n542 4.65
R2867 GND.n544 GND.n314 4.65
R2868 GND.n547 GND.n546 4.65
R2869 GND.n311 GND.n310 4.65
R2870 GND.n555 GND.n554 4.65
R2871 GND.n556 GND.n309 4.65
R2872 GND.n558 GND.n557 4.65
R2873 GND.n306 GND.n305 4.65
R2874 GND.n566 GND.n565 4.65
R2875 GND.n567 GND.n304 4.65
R2876 GND.n570 GND.n568 4.65
R2877 GND.n584 GND.n583 4.65
R2878 GND.n585 GND.n297 4.65
R2879 GND.n587 GND.n586 4.65
R2880 GND.n293 GND.n292 4.65
R2881 GND.n594 GND.n593 4.65
R2882 GND.n595 GND.n291 4.65
R2883 GND.n598 GND.n597 4.65
R2884 GND.n596 GND.n287 4.65
R2885 GND.n605 GND.n604 4.65
R2886 GND.n606 GND.n285 4.65
R2887 GND.n611 GND.n610 4.65
R2888 GND.n609 GND.n281 4.65
R2889 GND.n619 GND.n618 4.65
R2890 GND.n620 GND.n280 4.65
R2891 GND.n623 GND.n622 4.65
R2892 GND.n277 GND.n276 4.65
R2893 GND.n631 GND.n630 4.65
R2894 GND.n632 GND.n275 4.65
R2895 GND.n634 GND.n633 4.65
R2896 GND.n272 GND.n271 4.65
R2897 GND.n642 GND.n641 4.65
R2898 GND.n643 GND.n269 4.65
R2899 GND.n645 GND.n644 4.65
R2900 GND.n1595 GND.n1594 4.65
R2901 GND.n1599 GND.n1598 4.65
R2902 GND.n1603 GND.n1602 4.65
R2903 GND.n1611 GND.n1610 4.65
R2904 GND.n1619 GND.n1618 4.65
R2905 GND.n1627 GND.n1626 4.65
R2906 GND.n1635 GND.n1634 4.65
R2907 GND.n1643 GND.n1642 4.65
R2908 GND.n1652 GND.n1651 4.65
R2909 GND.n1660 GND.n1659 4.65
R2910 GND.n1673 GND.n1672 4.65
R2911 GND.n1683 GND.n1680 4.65
R2912 GND.n1690 GND.n1689 4.65
R2913 GND.n1698 GND.n1697 4.65
R2914 GND.n1706 GND.n1705 4.65
R2915 GND.n1715 GND.n1714 4.65
R2916 GND.n1723 GND.n1722 4.65
R2917 GND.n1731 GND.n1730 4.65
R2918 GND.n1739 GND.n1738 4.65
R2919 GND.n1747 GND.n1746 4.65
R2920 GND.n1755 GND.n1754 4.65
R2921 GND.n1764 GND.n1763 4.65
R2922 GND.n1769 GND.n1768 4.65
R2923 GND.n1774 GND.n1773 4.65
R2924 GND.n1607 GND.n1606 4.65
R2925 GND.n1615 GND.n1614 4.65
R2926 GND.n1623 GND.n1622 4.65
R2927 GND.n1631 GND.n1630 4.65
R2928 GND.n1639 GND.n1638 4.65
R2929 GND.n1647 GND.n1646 4.65
R2930 GND.n1656 GND.n1655 4.65
R2931 GND.n1664 GND.n1663 4.65
R2932 GND.n1669 GND.n1668 4.65
R2933 GND.n1677 GND.n1676 4.65
R2934 GND.n1686 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/GND 4.65
R2935 GND.n1694 GND.n1693 4.65
R2936 GND.n1702 GND.n1701 4.65
R2937 GND.n1710 GND.n1709 4.65
R2938 GND.n1719 GND.n1718 4.65
R2939 GND.n1727 GND.n1726 4.65
R2940 GND.n1735 GND.n1734 4.65
R2941 GND.n1743 GND.n1742 4.65
R2942 GND.n1751 GND.n1750 4.65
R2943 GND.n1759 GND.n1758 4.65
R2944 GND.n1766 GND.n1765 4.65
R2945 GND.n1771 GND.n1770 4.65
R2946 GND.n1902 GND.n1901 4.65
R2947 GND.n1799 GND.n1798 4.65
R2948 GND.n1808 GND.n1807 4.65
R2949 GND.n1816 GND.n1815 4.65
R2950 GND.n1824 GND.n1823 4.65
R2951 GND.n1833 GND.n1832 4.65
R2952 GND.n1843 GND.n1840 4.65
R2953 GND.n1851 GND.n1850 4.65
R2954 GND.n1860 GND.n1859 4.65
R2955 GND.n1868 GND.n1867 4.65
R2956 GND.n1877 GND.n1876 4.65
R2957 GND.n1885 GND.n1884 4.65
R2958 GND.n1892 GND.n1891 4.65
R2959 GND.n1898 GND.n1897 4.65
R2960 GND.n1791 GND.n1790 4.65
R2961 GND.n1784 GND.n1783 4.65
R2962 GND.n1778 GND.n1777 4.65
R2963 GND.n1776 GND.n1775 4.65
R2964 GND.n1782 GND.n1781 4.65
R2965 GND.n1788 GND.n1787 4.65
R2966 GND.n1795 GND.n1794 4.65
R2967 GND.n1803 GND.n1802 4.65
R2968 GND.n1812 GND.n1811 4.65
R2969 GND.n1820 GND.n1819 4.65
R2970 GND.n1829 GND.n1828 4.65
R2971 GND.n1837 GND.n1836 4.65
R2972 GND.n1847 GND.n1846 4.65
R2973 GND.n1856 GND.n1855 4.65
R2974 GND.n1864 GND.n1863 4.65
R2975 GND.n1872 GND.n1871 4.65
R2976 GND.n1881 GND.n1880 4.65
R2977 GND.n1888 GND.n1887 4.65
R2978 GND.n1894 GND.n1893 4.65
R2979 GND.n1900 GND.n1899 4.65
R2980 GND.n1915 GND.n1914 4.65
R2981 GND.n1924 GND.n1923 4.65
R2982 GND.n1932 GND.n1931 4.65
R2983 GND.n1940 GND.n1939 4.65
R2984 GND.n1948 GND.n1947 4.65
R2985 GND.n1956 GND.n1955 4.65
R2986 GND.n1964 GND.n1963 4.65
R2987 GND.n1972 GND.n1971 4.65
R2988 GND.n1980 GND.n1979 4.65
R2989 GND.n1989 GND.n1988 4.65
R2990 GND.n1998 GND.n1997 4.65
R2991 GND.n2006 GND.n2005 4.65
R2992 GND.n2013 GND.n2010 4.65
R2993 GND.n2021 GND.n2020 4.65
R2994 GND.n2029 GND.n2028 4.65
R2995 GND.n2037 GND.n2036 4.65
R2996 GND.n2047 GND.n2046 4.65
R2997 GND.n2055 GND.n2054 4.65
R2998 GND.n2063 GND.n2062 4.65
R2999 GND.n2071 GND.n2070 4.65
R3000 GND.n2079 GND.n2078 4.65
R3001 GND.n2087 GND.n2086 4.65
R3002 GND.n2095 GND.n2094 4.65
R3003 GND.n2103 GND.n2102 4.65
R3004 GND.n1907 GND.n1906 4.65
R3005 GND.n1905 GND.n1904 4.65
R3006 GND.n1913 GND.n1912 4.65
R3007 GND.n1920 GND.n1919 4.65
R3008 GND.n1928 GND.n1927 4.65
R3009 GND.n1936 GND.n1935 4.65
R3010 GND.n1944 GND.n1943 4.65
R3011 GND.n1952 GND.n1951 4.65
R3012 GND.n1960 GND.n1959 4.65
R3013 GND.n1968 GND.n1967 4.65
R3014 GND.n1976 GND.n1975 4.65
R3015 GND.n1984 GND.n1983 4.65
R3016 GND.n1994 GND.n1993 4.65
R3017 GND.n2002 GND.n2001 4.65
R3018 GND.n2009 GND.n1550 4.65
R3019 GND.n2017 GND.n2016 4.65
R3020 GND.n2025 GND.n2024 4.65
R3021 GND.n2033 GND.n2032 4.65
R3022 GND.n2042 GND.n2041 4.65
R3023 GND.n2051 GND.n2050 4.65
R3024 GND.n2059 GND.n2058 4.65
R3025 GND.n2067 GND.n2066 4.65
R3026 GND.n2075 GND.n2074 4.65
R3027 GND.n2083 GND.n2082 4.65
R3028 GND.n2091 GND.n2090 4.65
R3029 GND.n2099 GND.n2098 4.65
R3030 GND.n2107 GND.n2106 4.65
R3031 GND.n1365 GND.n1364 4.65
R3032 GND.n1358 GND.n1357 4.65
R3033 GND.n1373 GND.n1372 4.65
R3034 GND.n1374 GND.n1356 4.65
R3035 GND.n1376 GND.n1375 4.65
R3036 GND.n1353 GND.n1352 4.65
R3037 GND.n1384 GND.n1383 4.65
R3038 GND.n1386 GND.n1351 4.65
R3039 GND.n1388 GND.n1387 4.65
R3040 GND.n1348 GND.n1347 4.65
R3041 GND.n1395 GND.n1394 4.65
R3042 GND.n1396 GND.n1345 4.65
R3043 GND.n1399 GND.n1398 4.65
R3044 GND.n1397 GND.n1341 4.65
R3045 GND.n1406 GND.n1405 4.65
R3046 GND.n1407 GND.n1339 4.65
R3047 GND.n1409 GND.n1408 4.65
R3048 GND.n1335 GND.n1334 4.65
R3049 GND.n1416 GND.n1415 4.65
R3050 GND.n1417 GND.n1333 4.65
R3051 GND.n1419 GND.n1418 4.65
R3052 GND.n1329 GND.n1328 4.65
R3053 GND.n1424 GND.n1423 4.65
R3054 GND.n1427 GND.n1426 4.65
R3055 GND.n1428 GND.n1327 4.65
R3056 GND.n1430 GND.n1429 4.65
R3057 GND.n1324 GND.n1323 4.65
R3058 GND.n1438 GND.n1437 4.65
R3059 GND.n1440 GND.n1322 4.65
R3060 GND.n1442 GND.n1441 4.65
R3061 GND.n1319 GND.n1318 4.65
R3062 GND.n1449 GND.n1448 4.65
R3063 GND.n1450 GND.n1316 4.65
R3064 GND.n1453 GND.n1452 4.65
R3065 GND.n1451 GND.n1312 4.65
R3066 GND.n1460 GND.n1459 4.65
R3067 GND.n1461 GND.n1310 4.65
R3068 GND.n1463 GND.n1462 4.65
R3069 GND.n1306 GND.n1305 4.65
R3070 GND.n1468 GND.n1467 4.65
R3071 GND.n1471 GND.n1470 4.65
R3072 GND.n1472 GND.n1304 4.65
R3073 GND.n1474 GND.n1473 4.65
R3074 GND.n1301 GND.n1300 4.65
R3075 GND.n1482 GND.n1481 4.65
R3076 GND.n1483 GND.n1299 4.65
R3077 GND.n1485 GND.n1484 4.65
R3078 GND.n1296 GND.n1295 4.65
R3079 GND.n1493 GND.n1492 4.65
R3080 GND.n1495 GND.n1294 4.65
R3081 GND.n1497 GND.n1496 4.65
R3082 GND.n1291 GND.n1290 4.65
R3083 GND.n1504 GND.n1503 4.65
R3084 GND.n1505 GND.n1288 4.65
R3085 GND.n1508 GND.n1507 4.65
R3086 GND.n1506 GND.n1284 4.65
R3087 GND.n1515 GND.n1514 4.65
R3088 GND.n1516 GND.n1282 4.65
R3089 GND.n1518 GND.n1517 4.65
R3090 GND.n1278 GND.n1277 4.65
R3091 GND.n1525 GND.n1524 4.65
R3092 GND.n1526 GND.n1276 4.65
R3093 GND.n1529 GND.n1527 4.65
R3094 GND.n1104 GND.n1103 4.65
R3095 GND.n1097 GND.n1096 4.65
R3096 GND.n1111 GND.n1110 4.65
R3097 GND.n1112 GND.n1095 4.65
R3098 GND.n1115 GND.n1114 4.65
R3099 GND.n1091 GND.n1090 4.65
R3100 GND.n1123 GND.n1122 4.65
R3101 GND.n1124 GND.n1087 4.65
R3102 GND.n1126 GND.n1125 4.65
R3103 GND.n1084 GND.n1083 4.65
R3104 GND.n1133 GND.n1132 4.65
R3105 GND.n1134 GND.n1082 4.65
R3106 GND.n1137 GND.n1136 4.65
R3107 GND.n1078 GND.n1077 4.65
R3108 GND.n1144 GND.n1143 4.65
R3109 GND.n1145 GND.n1076 4.65
R3110 GND.n1147 GND.n1146 4.65
R3111 GND.n1072 GND.n1071 4.65
R3112 GND.n1152 GND.n1151 4.65
R3113 GND.n1155 GND.n1154 4.65
R3114 GND.n1156 GND.n1070 4.65
R3115 GND.n1158 GND.n1157 4.65
R3116 GND.n1067 GND.n1066 4.65
R3117 GND.n1166 GND.n1165 4.65
R3118 GND.n1168 GND.n1065 4.65
R3119 GND.n1170 GND.n1169 4.65
R3120 GND.n1062 GND.n1061 4.65
R3121 GND.n1177 GND.n1176 4.65
R3122 GND.n1178 GND.n1058 4.65
R3123 GND.n1181 GND.n1180 4.65
R3124 GND.n1179 GND.n1054 4.65
R3125 GND.n1188 GND.n1187 4.65
R3126 GND.n1189 GND.n1052 4.65
R3127 GND.n1191 GND.n1190 4.65
R3128 GND.n1048 GND.n1047 4.65
R3129 GND.n1196 GND.n1195 4.65
R3130 GND.n1198 GND.n1197 4.65
R3131 GND.n1045 GND.n1044 4.65
R3132 GND.n1204 GND.n1203 4.65
R3133 GND.n1205 GND.n1043 4.65
R3134 GND.n1207 GND.n1206 4.65
R3135 GND.n1039 GND.n1038 4.65
R3136 GND.n1214 GND.n1213 4.65
R3137 GND.n1215 GND.n1037 4.65
R3138 GND.n1218 GND.n1217 4.65
R3139 GND.n1216 GND.n1033 4.65
R3140 GND.n1225 GND.n1224 4.65
R3141 GND.n1226 GND.n1031 4.65
R3142 GND.n1231 GND.n1230 4.65
R3143 GND.n1229 GND.n1027 4.65
R3144 GND.n1239 GND.n1238 4.65
R3145 GND.n1240 GND.n1026 4.65
R3146 GND.n1243 GND.n1242 4.65
R3147 GND.n1023 GND.n1022 4.65
R3148 GND.n1251 GND.n1250 4.65
R3149 GND.n1252 GND.n1021 4.65
R3150 GND.n1254 GND.n1253 4.65
R3151 GND.n1018 GND.n1017 4.65
R3152 GND.n1262 GND.n1261 4.65
R3153 GND.n1263 GND.n1016 4.65
R3154 GND.n1266 GND.n1264 4.65
R3155 GND.n776 GND.n775 4.65
R3156 GND.n780 GND.n779 4.65
R3157 GND.n784 GND.n783 4.65
R3158 GND.n788 GND.n787 4.65
R3159 GND.n792 GND.n791 4.65
R3160 GND.n797 GND.n796 4.65
R3161 GND.n801 GND.n800 4.65
R3162 GND.n805 GND.n804 4.65
R3163 GND.n807 GND.n806 4.65
R3164 GND.n811 GND.n810 4.65
R3165 GND.n815 GND.n814 4.65
R3166 GND.n819 GND.n818 4.65
R3167 GND.n824 GND.n823 4.65
R3168 GND.n828 GND.n827 4.65
R3169 GND.n832 GND.n831 4.65
R3170 GND.n836 GND.n835 4.65
R3171 GND.n840 GND.n839 4.65
R3172 GND.n844 GND.n843 4.65
R3173 GND.n846 GND.n845 4.65
R3174 GND.n848 GND.n847 4.65
R3175 GND.n852 GND.n851 4.65
R3176 GND.n856 GND.n855 4.65
R3177 GND.n860 GND.n859 4.65
R3178 GND.n864 GND.n863 4.65
R3179 GND.n869 GND.n868 4.65
R3180 GND.n873 GND.n872 4.65
R3181 GND.n877 GND.n876 4.65
R3182 GND.n879 GND.n878 4.65
R3183 GND.n883 GND.n882 4.65
R3184 GND.n887 GND.n886 4.65
R3185 GND.n891 GND.n890 4.65
R3186 GND.n896 GND.n895 4.65
R3187 GND.n900 GND.n899 4.65
R3188 GND.n904 GND.n903 4.65
R3189 GND.n908 GND.n907 4.65
R3190 GND.n910 GND.n909 4.65
R3191 GND.n913 GND.n912 4.65
R3192 GND.n917 GND.n916 4.65
R3193 GND.n921 GND.n920 4.65
R3194 GND.n925 GND.n924 4.65
R3195 GND.n929 GND.n928 4.65
R3196 GND.n933 GND.n932 4.65
R3197 GND.n937 GND.n936 4.65
R3198 GND.n941 GND.n940 4.65
R3199 GND.n945 GND.n944 4.65
R3200 GND.n949 GND.n948 4.65
R3201 GND.n954 GND.n953 4.65
R3202 GND.n958 GND.n957 4.65
R3203 GND.n962 GND.n961 4.65
R3204 GND.n964 GND.n963 4.65
R3205 GND.n968 GND.n967 4.65
R3206 GND.n972 GND.n971 4.65
R3207 GND.n976 GND.n975 4.65
R3208 GND.n981 GND.n980 4.65
R3209 GND.n985 GND.n984 4.65
R3210 GND.n989 GND.n988 4.65
R3211 GND.n993 GND.n992 4.65
R3212 GND.n997 GND.n996 4.65
R3213 GND.n1001 GND.n1000 4.65
R3214 GND.n1005 GND.n1004 4.65
R3215 GND.n1009 GND.n1008 4.65
R3216 GND.n577 GND.n576 4.65
R3217 GND.n753 GND.n752 4.65
R3218 GND.n163 GND.n162 4.65
R3219 GND.n167 GND.n166 4.65
R3220 GND.n171 GND.n170 4.65
R3221 GND.n175 GND.n174 4.65
R3222 GND.n179 GND.n178 4.65
R3223 GND.n183 GND.n182 4.65
R3224 GND.n187 GND.n186 4.65
R3225 GND.n191 GND.n190 4.65
R3226 GND.n195 GND.n194 4.65
R3227 GND.n200 GND.n199 4.65
R3228 GND.n204 GND.n203 4.65
R3229 GND.n208 GND.n207 4.65
R3230 GND.n210 GND.n209 4.65
R3231 GND.n214 GND.n213 4.65
R3232 GND.n218 GND.n217 4.65
R3233 GND.n222 GND.n221 4.65
R3234 GND.n227 GND.n226 4.65
R3235 GND.n231 GND.n230 4.65
R3236 GND.n235 GND.n234 4.65
R3237 GND.n239 GND.n238 4.65
R3238 GND.n243 GND.n242 4.65
R3239 GND.n247 GND.n246 4.65
R3240 GND.n251 GND.n250 4.65
R3241 GND.n255 GND.n254 4.65
R3242 GND.n159 GND.n158 4.65
R3243 GND.n748 GND.n747 4.65
R3244 GND.n744 GND.n743 4.65
R3245 GND.n740 GND.n739 4.65
R3246 GND.n736 GND.n735 4.65
R3247 GND.n732 GND.n731 4.65
R3248 GND.n728 GND.n727 4.65
R3249 GND.n724 GND.n723 4.65
R3250 GND.n720 GND.n719 4.65
R3251 GND.n715 GND.n714 4.65
R3252 GND.n711 GND.n710 4.65
R3253 GND.n707 GND.n706 4.65
R3254 GND.n703 GND.n702 4.65
R3255 GND.n701 GND.n698 4.65
R3256 GND.n697 GND.n696 4.65
R3257 GND.n693 GND.n692 4.65
R3258 GND.n688 GND.n687 4.65
R3259 GND.n684 GND.n683 4.65
R3260 GND.n680 GND.n679 4.65
R3261 GND.n676 GND.n675 4.65
R3262 GND.n672 GND.n671 4.65
R3263 GND.n668 GND.n667 4.65
R3264 GND.n664 GND.n663 4.65
R3265 GND.n660 GND.n659 4.65
R3266 GND.n2111 GND.n1535 4.467
R3267 EESPFAL_Sbox_0/EESPFAL_s1_0/GND GND.n2111 4.432
R3268 EESPFAL_Sbox_0/EESPFAL_s2_0/GND GND.n1534 4.379
R3269 GND.n753 EESPFAL_Sbox_0/EESPFAL_s0_0/GND 4.37
R3270 GND.n1550 GND.n1547 3.28
R3271 GND.n2016 GND.n2013 3.28
R3272 GND.n1541 GND.n1538 3.28
R3273 GND.n1565 GND.n1562 3.18
R3274 GND.n1829 GND.n1565 3.18
R3275 GND.n1832 GND.n1829 3.18
R3276 GND.n1558 GND.n1555 3.18
R3277 GND.n1843 GND.n1558 3.18
R3278 GND.n1846 GND.n1843 3.18
R3279 GND.n1547 GND.n1544 3.12
R3280 GND.n2013 GND.n1550 3.12
R3281 GND.n16 GND.n15 2.791
R3282 GND.n96 GND.n95 2.791
R3283 GND.n395 GND.n393 2.791
R3284 GND.n447 GND.n363 2.791
R3285 GND.n1101 GND.n1099 2.791
R3286 GND.n1153 GND.n1069 2.791
R3287 GND.n770 GND.n769 2.791
R3288 GND.n850 GND.n849 2.791
R3289 GND.n88 GND.n87 2.791
R3290 GND.n152 GND.n151 2.791
R3291 GND.n444 GND.n367 2.791
R3292 GND.n498 GND.n337 2.791
R3293 GND.n1150 GND.n1073 2.791
R3294 GND.n1194 GND.n1049 2.791
R3295 GND.n842 GND.n841 2.791
R3296 GND.n906 GND.n905 2.791
R3297 GND.n751 GND.n749 2.74
R3298 GND.n575 GND.n301 2.739
R3299 GND.n578 GND.n298 2.739
R3300 GND.n650 GND.n266 2.739
R3301 GND.n1533 GND.n1272 2.739
R3302 GND.n1271 GND.n1013 2.739
R3303 GND.n1012 GND.n1010 2.739
R3304 GND.n258 GND.n256 2.739
R3305 GND.n656 GND.n652 2.739
R3306 GND.n18 GND.n17 2.682
R3307 GND.n396 GND.n394 2.682
R3308 GND.n1363 GND.n1361 2.682
R3309 GND.n1102 GND.n1100 2.682
R3310 GND.n772 GND.n771 2.682
R3311 GND.n749 GND.n261 2.682
R3312 GND.n569 GND.n301 2.682
R3313 GND.n299 GND.n298 2.682
R3314 GND.n270 GND.n266 2.682
R3315 GND.n1528 GND.n1272 2.682
R3316 GND.n1265 GND.n1013 2.682
R3317 GND.n1010 GND.n756 2.682
R3318 GND.n256 GND.n2 2.682
R3319 GND.n656 GND.n655 2.682
R3320 GND.n2110 GND.n2109 1.912
R3321 GND.n2109 GND.n1541 1.889
R3322 GND.n1362 GND.n1360 1.873
R3323 GND.n1425 GND.n1326 1.873
R3324 GND.n1532 GND.n1273 1.873
R3325 GND.n1422 GND.n1330 1.873
R3326 GND.n1466 GND.n1307 1.873
R3327 GND.n1469 GND.n1303 1.873
R3328 GND.n1780 GND.n1779 1.695
R3329 GND.n1896 GND.n1895 1.695
R3330 GND.n1582 GND.n1579 1.68
R3331 GND.n1669 GND.n1585 1.68
R3332 GND.n1575 GND.n1572 1.68
R3333 GND.n1686 GND.n1683 1.68
R3334 GND.n1593 GND.n1592 1.588
R3335 GND.n576 EESPFAL_Sbox_0/GND 1.565
R3336 GND.n2109 GND.n2108 1.417
R3337 GND.n749 GND.n748 1.096
R3338 GND.n22 GND.n18 1.096
R3339 GND.n397 GND.n396 1.096
R3340 GND.n1364 GND.n1363 1.096
R3341 GND.n1103 GND.n1102 1.096
R3342 GND.n776 GND.n772 1.096
R3343 GND.n660 GND.n656 1.095
R3344 GND.n256 GND.n255 1.095
R3345 GND.n568 GND.n301 1.095
R3346 GND.n584 GND.n298 1.095
R3347 GND.n644 GND.n266 1.095
R3348 GND.n1527 GND.n1272 1.095
R3349 GND.n1264 GND.n1013 1.095
R3350 GND.n1010 GND.n1009 1.095
R3351 GND.n1595 GND.n1593 0.813
R3352 GND.n913 GND.n910 0.662
R3353 GND.n159 GND.n156 0.637
R3354 GND.n1197 GND.n1196 0.637
R3355 GND.n501 GND.n500 0.6
R3356 GND.n1471 GND.n1468 0.562
R3357 GND.n94 GND.n92 0.55
R3358 GND.n1427 GND.n1424 0.55
R3359 GND.n1155 GND.n1152 0.55
R3360 GND.n848 GND.n846 0.548
R3361 GND.n449 GND.n446 0.525
R3362 GND.n1905 GND.n1902 0.172
R3363 GND.n1776 GND.n1774 0.165
R3364 GND.n748 GND.n744 0.1
R3365 GND.n744 GND.n740 0.1
R3366 GND.n740 GND.n736 0.1
R3367 GND.n736 GND.n732 0.1
R3368 GND.n732 GND.n728 0.1
R3369 GND.n728 GND.n724 0.1
R3370 GND.n724 GND.n720 0.1
R3371 GND.n715 GND.n711 0.1
R3372 GND.n711 GND.n707 0.1
R3373 GND.n707 GND.n703 0.1
R3374 GND.n698 GND.n697 0.1
R3375 GND.n697 GND.n693 0.1
R3376 GND.n688 GND.n684 0.1
R3377 GND.n684 GND.n680 0.1
R3378 GND.n680 GND.n676 0.1
R3379 GND.n676 GND.n672 0.1
R3380 GND.n672 GND.n668 0.1
R3381 GND.n668 GND.n664 0.1
R3382 GND.n664 GND.n660 0.1
R3383 GND.n26 GND.n22 0.1
R3384 GND.n30 GND.n26 0.1
R3385 GND.n34 GND.n30 0.1
R3386 GND.n38 GND.n34 0.1
R3387 GND.n47 GND.n43 0.1
R3388 GND.n51 GND.n47 0.1
R3389 GND.n52 GND.n51 0.1
R3390 GND.n61 GND.n57 0.1
R3391 GND.n65 GND.n61 0.1
R3392 GND.n74 GND.n70 0.1
R3393 GND.n78 GND.n74 0.1
R3394 GND.n82 GND.n78 0.1
R3395 GND.n86 GND.n82 0.1
R3396 GND.n90 GND.n86 0.1
R3397 GND.n92 GND.n90 0.1
R3398 GND.n98 GND.n94 0.1
R3399 GND.n102 GND.n98 0.1
R3400 GND.n106 GND.n102 0.1
R3401 GND.n110 GND.n106 0.1
R3402 GND.n119 GND.n115 0.1
R3403 GND.n123 GND.n119 0.1
R3404 GND.n124 GND.n123 0.1
R3405 GND.n133 GND.n129 0.1
R3406 GND.n137 GND.n133 0.1
R3407 GND.n146 GND.n142 0.1
R3408 GND.n150 GND.n146 0.1
R3409 GND.n154 GND.n150 0.1
R3410 GND.n156 GND.n154 0.1
R3411 GND.n163 GND.n159 0.1
R3412 GND.n167 GND.n163 0.1
R3413 GND.n171 GND.n167 0.1
R3414 GND.n175 GND.n171 0.1
R3415 GND.n179 GND.n175 0.1
R3416 GND.n183 GND.n179 0.1
R3417 GND.n187 GND.n183 0.1
R3418 GND.n191 GND.n187 0.1
R3419 GND.n195 GND.n191 0.1
R3420 GND.n204 GND.n200 0.1
R3421 GND.n208 GND.n204 0.1
R3422 GND.n209 GND.n208 0.1
R3423 GND.n218 GND.n214 0.1
R3424 GND.n222 GND.n218 0.1
R3425 GND.n231 GND.n227 0.1
R3426 GND.n235 GND.n231 0.1
R3427 GND.n239 GND.n235 0.1
R3428 GND.n243 GND.n239 0.1
R3429 GND.n247 GND.n243 0.1
R3430 GND.n251 GND.n247 0.1
R3431 GND.n255 GND.n251 0.1
R3432 GND.n397 GND.n390 0.1
R3433 GND.n405 GND.n390 0.1
R3434 GND.n406 GND.n405 0.1
R3435 GND.n408 GND.n406 0.1
R3436 GND.n417 GND.n384 0.1
R3437 GND.n418 GND.n417 0.1
R3438 GND.n419 GND.n418 0.1
R3439 GND.n427 GND.n377 0.1
R3440 GND.n428 GND.n427 0.1
R3441 GND.n430 GND.n371 0.1
R3442 GND.n438 GND.n371 0.1
R3443 GND.n439 GND.n438 0.1
R3444 GND.n440 GND.n439 0.1
R3445 GND.n440 GND.n365 0.1
R3446 GND.n446 GND.n365 0.1
R3447 GND.n450 GND.n449 0.1
R3448 GND.n451 GND.n450 0.1
R3449 GND.n451 GND.n360 0.1
R3450 GND.n459 GND.n360 0.1
R3451 GND.n460 GND.n459 0.1
R3452 GND.n462 GND.n460 0.1
R3453 GND.n471 GND.n354 0.1
R3454 GND.n472 GND.n471 0.1
R3455 GND.n473 GND.n472 0.1
R3456 GND.n481 GND.n347 0.1
R3457 GND.n482 GND.n481 0.1
R3458 GND.n484 GND.n341 0.1
R3459 GND.n492 GND.n341 0.1
R3460 GND.n493 GND.n492 0.1
R3461 GND.n494 GND.n493 0.1
R3462 GND.n494 GND.n335 0.1
R3463 GND.n500 GND.n335 0.1
R3464 GND.n501 GND.n332 0.1
R3465 GND.n508 GND.n332 0.1
R3466 GND.n509 GND.n508 0.1
R3467 GND.n510 GND.n509 0.1
R3468 GND.n510 GND.n326 0.1
R3469 GND.n518 GND.n326 0.1
R3470 GND.n519 GND.n518 0.1
R3471 GND.n521 GND.n519 0.1
R3472 GND.n521 GND.n520 0.1
R3473 GND.n530 GND.n529 0.1
R3474 GND.n534 GND.n530 0.1
R3475 GND.n534 GND.n533 0.1
R3476 GND.n544 GND.n543 0.1
R3477 GND.n546 GND.n544 0.1
R3478 GND.n555 GND.n310 0.1
R3479 GND.n556 GND.n555 0.1
R3480 GND.n557 GND.n556 0.1
R3481 GND.n557 GND.n305 0.1
R3482 GND.n566 GND.n305 0.1
R3483 GND.n567 GND.n566 0.1
R3484 GND.n568 GND.n567 0.1
R3485 GND.n585 GND.n584 0.1
R3486 GND.n586 GND.n585 0.1
R3487 GND.n586 GND.n292 0.1
R3488 GND.n594 GND.n292 0.1
R3489 GND.n595 GND.n594 0.1
R3490 GND.n597 GND.n595 0.1
R3491 GND.n597 GND.n596 0.1
R3492 GND.n606 GND.n605 0.1
R3493 GND.n610 GND.n606 0.1
R3494 GND.n610 GND.n609 0.1
R3495 GND.n620 GND.n619 0.1
R3496 GND.n622 GND.n620 0.1
R3497 GND.n631 GND.n276 0.1
R3498 GND.n632 GND.n631 0.1
R3499 GND.n633 GND.n632 0.1
R3500 GND.n633 GND.n271 0.1
R3501 GND.n642 GND.n271 0.1
R3502 GND.n643 GND.n642 0.1
R3503 GND.n644 GND.n643 0.1
R3504 GND.n1364 GND.n1357 0.1
R3505 GND.n1373 GND.n1357 0.1
R3506 GND.n1374 GND.n1373 0.1
R3507 GND.n1375 GND.n1374 0.1
R3508 GND.n1375 GND.n1352 0.1
R3509 GND.n1384 GND.n1352 0.1
R3510 GND.n1387 GND.n1386 0.1
R3511 GND.n1387 GND.n1347 0.1
R3512 GND.n1395 GND.n1347 0.1
R3513 GND.n1398 GND.n1396 0.1
R3514 GND.n1398 GND.n1397 0.1
R3515 GND.n1407 GND.n1406 0.1
R3516 GND.n1408 GND.n1407 0.1
R3517 GND.n1408 GND.n1334 0.1
R3518 GND.n1416 GND.n1334 0.1
R3519 GND.n1417 GND.n1416 0.1
R3520 GND.n1418 GND.n1417 0.1
R3521 GND.n1418 GND.n1328 0.1
R3522 GND.n1424 GND.n1328 0.1
R3523 GND.n1428 GND.n1427 0.1
R3524 GND.n1429 GND.n1428 0.1
R3525 GND.n1429 GND.n1323 0.1
R3526 GND.n1438 GND.n1323 0.1
R3527 GND.n1441 GND.n1440 0.1
R3528 GND.n1441 GND.n1318 0.1
R3529 GND.n1449 GND.n1318 0.1
R3530 GND.n1452 GND.n1450 0.1
R3531 GND.n1452 GND.n1451 0.1
R3532 GND.n1461 GND.n1460 0.1
R3533 GND.n1462 GND.n1461 0.1
R3534 GND.n1462 GND.n1305 0.1
R3535 GND.n1468 GND.n1305 0.1
R3536 GND.n1472 GND.n1471 0.1
R3537 GND.n1473 GND.n1472 0.1
R3538 GND.n1473 GND.n1300 0.1
R3539 GND.n1482 GND.n1300 0.1
R3540 GND.n1483 GND.n1482 0.1
R3541 GND.n1484 GND.n1483 0.1
R3542 GND.n1484 GND.n1295 0.1
R3543 GND.n1493 GND.n1295 0.1
R3544 GND.n1496 GND.n1495 0.1
R3545 GND.n1496 GND.n1290 0.1
R3546 GND.n1504 GND.n1290 0.1
R3547 GND.n1507 GND.n1505 0.1
R3548 GND.n1507 GND.n1506 0.1
R3549 GND.n1516 GND.n1515 0.1
R3550 GND.n1517 GND.n1516 0.1
R3551 GND.n1517 GND.n1277 0.1
R3552 GND.n1525 GND.n1277 0.1
R3553 GND.n1526 GND.n1525 0.1
R3554 GND.n1527 GND.n1526 0.1
R3555 GND.n1103 GND.n1096 0.1
R3556 GND.n1111 GND.n1096 0.1
R3557 GND.n1112 GND.n1111 0.1
R3558 GND.n1114 GND.n1112 0.1
R3559 GND.n1123 GND.n1090 0.1
R3560 GND.n1124 GND.n1123 0.1
R3561 GND.n1125 GND.n1124 0.1
R3562 GND.n1133 GND.n1083 0.1
R3563 GND.n1134 GND.n1133 0.1
R3564 GND.n1136 GND.n1077 0.1
R3565 GND.n1144 GND.n1077 0.1
R3566 GND.n1145 GND.n1144 0.1
R3567 GND.n1146 GND.n1145 0.1
R3568 GND.n1146 GND.n1071 0.1
R3569 GND.n1152 GND.n1071 0.1
R3570 GND.n1156 GND.n1155 0.1
R3571 GND.n1157 GND.n1156 0.1
R3572 GND.n1157 GND.n1066 0.1
R3573 GND.n1166 GND.n1066 0.1
R3574 GND.n1169 GND.n1168 0.1
R3575 GND.n1169 GND.n1061 0.1
R3576 GND.n1177 GND.n1061 0.1
R3577 GND.n1180 GND.n1178 0.1
R3578 GND.n1180 GND.n1179 0.1
R3579 GND.n1189 GND.n1188 0.1
R3580 GND.n1190 GND.n1189 0.1
R3581 GND.n1190 GND.n1047 0.1
R3582 GND.n1196 GND.n1047 0.1
R3583 GND.n1197 GND.n1044 0.1
R3584 GND.n1204 GND.n1044 0.1
R3585 GND.n1205 GND.n1204 0.1
R3586 GND.n1206 GND.n1205 0.1
R3587 GND.n1206 GND.n1038 0.1
R3588 GND.n1214 GND.n1038 0.1
R3589 GND.n1215 GND.n1214 0.1
R3590 GND.n1217 GND.n1215 0.1
R3591 GND.n1217 GND.n1216 0.1
R3592 GND.n1226 GND.n1225 0.1
R3593 GND.n1230 GND.n1226 0.1
R3594 GND.n1230 GND.n1229 0.1
R3595 GND.n1240 GND.n1239 0.1
R3596 GND.n1242 GND.n1240 0.1
R3597 GND.n1251 GND.n1022 0.1
R3598 GND.n1252 GND.n1251 0.1
R3599 GND.n1253 GND.n1252 0.1
R3600 GND.n1253 GND.n1017 0.1
R3601 GND.n1262 GND.n1017 0.1
R3602 GND.n1263 GND.n1262 0.1
R3603 GND.n1264 GND.n1263 0.1
R3604 GND.n780 GND.n776 0.1
R3605 GND.n784 GND.n780 0.1
R3606 GND.n788 GND.n784 0.1
R3607 GND.n792 GND.n788 0.1
R3608 GND.n801 GND.n797 0.1
R3609 GND.n805 GND.n801 0.1
R3610 GND.n806 GND.n805 0.1
R3611 GND.n815 GND.n811 0.1
R3612 GND.n819 GND.n815 0.1
R3613 GND.n828 GND.n824 0.1
R3614 GND.n832 GND.n828 0.1
R3615 GND.n836 GND.n832 0.1
R3616 GND.n840 GND.n836 0.1
R3617 GND.n844 GND.n840 0.1
R3618 GND.n846 GND.n844 0.1
R3619 GND.n852 GND.n848 0.1
R3620 GND.n856 GND.n852 0.1
R3621 GND.n860 GND.n856 0.1
R3622 GND.n864 GND.n860 0.1
R3623 GND.n873 GND.n869 0.1
R3624 GND.n877 GND.n873 0.1
R3625 GND.n878 GND.n877 0.1
R3626 GND.n887 GND.n883 0.1
R3627 GND.n891 GND.n887 0.1
R3628 GND.n900 GND.n896 0.1
R3629 GND.n904 GND.n900 0.1
R3630 GND.n908 GND.n904 0.1
R3631 GND.n910 GND.n908 0.1
R3632 GND.n917 GND.n913 0.1
R3633 GND.n921 GND.n917 0.1
R3634 GND.n925 GND.n921 0.1
R3635 GND.n929 GND.n925 0.1
R3636 GND.n933 GND.n929 0.1
R3637 GND.n937 GND.n933 0.1
R3638 GND.n941 GND.n937 0.1
R3639 GND.n945 GND.n941 0.1
R3640 GND.n949 GND.n945 0.1
R3641 GND.n958 GND.n954 0.1
R3642 GND.n962 GND.n958 0.1
R3643 GND.n963 GND.n962 0.1
R3644 GND.n972 GND.n968 0.1
R3645 GND.n976 GND.n972 0.1
R3646 GND.n985 GND.n981 0.1
R3647 GND.n989 GND.n985 0.1
R3648 GND.n993 GND.n989 0.1
R3649 GND.n997 GND.n993 0.1
R3650 GND.n1001 GND.n997 0.1
R3651 GND.n1005 GND.n1001 0.1
R3652 GND.n1009 GND.n1005 0.1
R3653 GND.n716 GND.n715 0.075
R3654 GND.n698 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_2/GND 0.075
R3655 GND.n693 GND.n689 0.075
R3656 GND.n43 GND.n39 0.075
R3657 GND.n57 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/GND 0.075
R3658 GND.n66 GND.n65 0.075
R3659 GND.n115 GND.n111 0.075
R3660 GND.n129 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/GND 0.075
R3661 GND.n138 GND.n137 0.075
R3662 GND.n200 GND.n196 0.075
R3663 GND.n214 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/GND 0.075
R3664 GND.n223 GND.n222 0.075
R3665 GND.n407 GND.n384 0.075
R3666 GND GND.n377 0.075
R3667 GND.n429 GND.n428 0.075
R3668 GND.n461 GND.n354 0.075
R3669 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/GND GND.n347 0.075
R3670 GND.n483 GND.n482 0.075
R3671 GND.n529 GND.n320 0.075
R3672 GND.n543 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/GND 0.075
R3673 GND.n546 GND.n545 0.075
R3674 GND.n605 GND.n286 0.075
R3675 GND.n619 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_0/GND 0.075
R3676 GND.n622 GND.n621 0.075
R3677 GND.n1386 GND.n1385 0.075
R3678 GND.n1396 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/GND 0.075
R3679 GND.n1397 GND.n1340 0.075
R3680 GND.n1440 GND.n1439 0.075
R3681 GND.n1450 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/GND 0.075
R3682 GND.n1451 GND.n1311 0.075
R3683 GND.n1495 GND.n1494 0.075
R3684 GND.n1505 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/GND 0.075
R3685 GND.n1506 GND.n1283 0.075
R3686 GND.n1113 GND.n1090 0.075
R3687 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/GND GND.n1083 0.075
R3688 GND.n1135 GND.n1134 0.075
R3689 GND.n1168 GND.n1167 0.075
R3690 GND.n1178 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/GND 0.075
R3691 GND.n1179 GND.n1053 0.075
R3692 GND.n1225 GND.n1032 0.075
R3693 GND.n1239 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/GND 0.075
R3694 GND.n1242 GND.n1241 0.075
R3695 GND.n797 GND.n793 0.075
R3696 GND.n811 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/GND 0.075
R3697 GND.n820 GND.n819 0.075
R3698 GND.n869 GND.n865 0.075
R3699 GND.n883 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/GND 0.075
R3700 GND.n892 GND.n891 0.075
R3701 GND.n954 GND.n950 0.075
R3702 GND.n968 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/GND 0.075
R3703 GND.n977 GND.n976 0.075
R3704 GND.n1540 GND.n1539 0.053
R3705 GND.n1603 GND.n1599 0.04
R3706 GND.n1611 GND.n1607 0.04
R3707 GND.n1619 GND.n1615 0.04
R3708 GND.n1627 GND.n1623 0.04
R3709 GND.n1635 GND.n1631 0.04
R3710 GND.n1643 GND.n1639 0.04
R3711 GND.n1660 GND.n1656 0.04
R3712 GND.n1665 GND.n1664 0.04
R3713 GND.n1667 GND.n1666 0.04
R3714 GND.n1678 GND.n1677 0.04
R3715 GND.n1680 GND.n1679 0.04
R3716 GND.n1690 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/GND 0.04
R3717 GND.n1698 GND.n1694 0.04
R3718 GND.n1706 GND.n1702 0.04
R3719 GND.n1723 GND.n1719 0.04
R3720 GND.n1731 GND.n1727 0.04
R3721 GND.n1739 GND.n1735 0.04
R3722 GND.n1747 GND.n1743 0.04
R3723 GND.n1755 GND.n1751 0.04
R3724 GND.n1764 GND.n1759 0.04
R3725 GND.n1769 GND.n1766 0.04
R3726 GND.n1774 GND.n1771 0.04
R3727 GND.n1534 EESPFAL_Sbox_0/EESPFAL_s3_0/GND 0.035
R3728 GND.n576 EESPFAL_Sbox_0/EESPFAL_s0_0/GND 0.035
R3729 EESPFAL_Sbox_0/EESPFAL_s1_0/GND GND.n753 0.035
R3730 GND.n1913 GND.n1907 0.028
R3731 GND.n1920 GND.n1915 0.028
R3732 GND.n1928 GND.n1924 0.028
R3733 GND.n1936 GND.n1932 0.028
R3734 GND.n1944 GND.n1940 0.028
R3735 GND.n1952 GND.n1948 0.028
R3736 GND.n1960 GND.n1956 0.028
R3737 GND.n1968 GND.n1964 0.028
R3738 GND.n1976 GND.n1972 0.028
R3739 GND.n1984 GND.n1980 0.028
R3740 GND.n2002 GND.n1998 0.028
R3741 GND.n2007 GND.n2006 0.028
R3742 GND.n2009 GND.n2008 0.028
R3743 GND.n2025 GND.n2021 0.028
R3744 GND.n2033 GND.n2029 0.028
R3745 GND.n2051 GND.n2047 0.028
R3746 GND.n2059 GND.n2055 0.028
R3747 GND.n2067 GND.n2063 0.028
R3748 GND.n2075 GND.n2071 0.028
R3749 GND.n2083 GND.n2079 0.028
R3750 GND.n2091 GND.n2087 0.028
R3751 GND.n2099 GND.n2095 0.028
R3752 GND.n2107 GND.n2103 0.028
R3753 GND.n1652 GND.n1648 0.027
R3754 GND.n1673 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/GND 0.027
R3755 GND.n1711 GND.n1710 0.027
R3756 GND.n1778 GND.n1776 0.027
R3757 GND.n1782 GND.n1778 0.027
R3758 GND.n1784 GND.n1782 0.027
R3759 GND.n1788 GND.n1784 0.027
R3760 GND.n1791 GND.n1788 0.027
R3761 GND.n1795 GND.n1791 0.027
R3762 GND.n1799 GND.n1795 0.027
R3763 GND.n1803 GND.n1799 0.027
R3764 GND.n1812 GND.n1808 0.027
R3765 GND.n1816 GND.n1812 0.027
R3766 GND.n1820 GND.n1816 0.027
R3767 GND.n1824 GND.n1820 0.027
R3768 GND.n1827 GND.n1826 0.027
R3769 GND.n1828 GND.n1827 0.027
R3770 GND.n1837 GND.n1833 0.027
R3771 GND.n1838 GND.n1837 0.027
R3772 GND.n1839 GND.n1838 0.027
R3773 GND.n1840 GND.n1839 0.027
R3774 GND.n1851 GND.n1847 0.027
R3775 GND.n1860 GND.n1856 0.027
R3776 GND.n1864 GND.n1860 0.027
R3777 GND.n1868 GND.n1864 0.027
R3778 GND.n1872 GND.n1868 0.027
R3779 GND.n1881 GND.n1877 0.027
R3780 GND.n1885 GND.n1881 0.027
R3781 GND.n1888 GND.n1885 0.027
R3782 GND.n1892 GND.n1888 0.027
R3783 GND.n1894 GND.n1892 0.027
R3784 GND.n1898 GND.n1894 0.027
R3785 GND.n1900 GND.n1898 0.027
R3786 GND.n1902 GND.n1900 0.027
R3787 GND.n1907 GND.n1905 0.027
R3788 GND.n1915 GND.n1913 0.027
R3789 GND.n1924 GND.n1920 0.027
R3790 GND.n1932 GND.n1928 0.027
R3791 GND.n1940 GND.n1936 0.027
R3792 GND.n1948 GND.n1944 0.027
R3793 GND.n1956 GND.n1952 0.027
R3794 GND.n1964 GND.n1960 0.027
R3795 GND.n1972 GND.n1968 0.027
R3796 GND.n1980 GND.n1976 0.027
R3797 GND.n1998 GND.n1994 0.027
R3798 GND.n2006 GND.n2002 0.027
R3799 GND.n2008 GND.n2007 0.027
R3800 GND.n2021 GND.n2017 0.027
R3801 GND.n2029 GND.n2025 0.027
R3802 GND.n2037 GND.n2033 0.027
R3803 GND.n2055 GND.n2051 0.027
R3804 GND.n2063 GND.n2059 0.027
R3805 GND.n2071 GND.n2067 0.027
R3806 GND.n2079 GND.n2075 0.027
R3807 GND.n2087 GND.n2083 0.027
R3808 GND.n2095 GND.n2091 0.027
R3809 GND.n2103 GND.n2099 0.027
R3810 GND.n2108 GND.n2107 0.027
R3811 GND.n1535 EESPFAL_Sbox_0/EESPFAL_s2_0/GND 0.026
R3812 GND.n720 GND.n716 0.025
R3813 GND.n703 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_2/GND 0.025
R3814 GND.n689 GND.n688 0.025
R3815 GND.n39 GND.n38 0.025
R3816 GND.n52 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/GND 0.025
R3817 GND.n70 GND.n66 0.025
R3818 GND.n111 GND.n110 0.025
R3819 GND.n124 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/GND 0.025
R3820 GND.n142 GND.n138 0.025
R3821 GND.n196 GND.n195 0.025
R3822 GND.n209 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/GND 0.025
R3823 GND.n227 GND.n223 0.025
R3824 GND.n408 GND.n407 0.025
R3825 GND.n419 GND 0.025
R3826 GND.n430 GND.n429 0.025
R3827 GND.n462 GND.n461 0.025
R3828 GND.n473 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/GND 0.025
R3829 GND.n484 GND.n483 0.025
R3830 GND.n520 GND.n320 0.025
R3831 GND.n533 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/GND 0.025
R3832 GND.n545 GND.n310 0.025
R3833 GND.n596 GND.n286 0.025
R3834 GND.n609 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_0/GND 0.025
R3835 GND.n621 GND.n276 0.025
R3836 GND.n1385 GND.n1384 0.025
R3837 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/GND GND.n1395 0.025
R3838 GND.n1406 GND.n1340 0.025
R3839 GND.n1439 GND.n1438 0.025
R3840 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/GND GND.n1449 0.025
R3841 GND.n1460 GND.n1311 0.025
R3842 GND.n1494 GND.n1493 0.025
R3843 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/GND GND.n1504 0.025
R3844 GND.n1515 GND.n1283 0.025
R3845 GND.n1114 GND.n1113 0.025
R3846 GND.n1125 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/GND 0.025
R3847 GND.n1136 GND.n1135 0.025
R3848 GND.n1167 GND.n1166 0.025
R3849 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/GND GND.n1177 0.025
R3850 GND.n1188 GND.n1053 0.025
R3851 GND.n1216 GND.n1032 0.025
R3852 GND.n1229 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/GND 0.025
R3853 GND.n1241 GND.n1022 0.025
R3854 GND.n793 GND.n792 0.025
R3855 GND.n806 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/GND 0.025
R3856 GND.n824 GND.n820 0.025
R3857 GND.n865 GND.n864 0.025
R3858 GND.n878 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/GND 0.025
R3859 GND.n896 GND.n892 0.025
R3860 GND.n950 GND.n949 0.025
R3861 GND.n963 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/GND 0.025
R3862 GND.n981 GND.n977 0.025
R3863 GND.n1599 GND.n1595 0.014
R3864 GND.n1607 GND.n1603 0.014
R3865 GND.n1615 GND.n1611 0.014
R3866 GND.n1623 GND.n1619 0.014
R3867 GND.n1631 GND.n1627 0.014
R3868 GND.n1639 GND.n1635 0.014
R3869 GND.n1647 GND.n1643 0.014
R3870 GND.n1656 GND.n1652 0.014
R3871 GND.n1664 GND.n1660 0.014
R3872 GND.n1668 GND.n1667 0.014
R3873 GND.n1677 GND.n1673 0.014
R3874 GND.n1679 GND.n1678 0.014
R3875 GND.n1702 GND.n1698 0.014
R3876 GND.n1710 GND.n1706 0.014
R3877 GND.n1719 GND.n1715 0.014
R3878 GND.n1727 GND.n1723 0.014
R3879 GND.n1735 GND.n1731 0.014
R3880 GND.n1743 GND.n1739 0.014
R3881 GND.n1751 GND.n1747 0.014
R3882 GND.n1759 GND.n1755 0.014
R3883 GND.n1766 GND.n1764 0.014
R3884 GND.n1771 GND.n1769 0.014
R3885 GND.n1994 GND.n1990 0.014
R3886 GND.n2017 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/GND 0.014
R3887 GND.n2038 GND.n2037 0.014
R3888 GND.n1648 GND.n1647 0.013
R3889 GND.n1666 GND.n1665 0.013
R3890 GND.n1668 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/GND 0.013
R3891 GND.n1680 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/GND 0.013
R3892 GND.n1694 GND.n1690 0.013
R3893 GND.n1715 GND.n1711 0.013
R3894 GND.n1804 GND.n1803 0.013
R3895 GND.n1808 GND.n1804 0.013
R3896 GND.n1825 GND.n1824 0.013
R3897 GND.n1826 GND.n1825 0.013
R3898 GND.n1828 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/GND 0.013
R3899 GND.n1833 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/GND 0.013
R3900 GND.n1840 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/GND 0.013
R3901 GND.n1847 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/GND 0.013
R3902 GND.n1852 GND.n1851 0.013
R3903 GND.n1856 GND.n1852 0.013
R3904 GND.n1873 GND.n1872 0.013
R3905 GND.n1877 GND.n1873 0.013
R3906 GND.n1985 GND.n1984 0.013
R3907 GND.n1989 GND.n1985 0.013
R3908 GND.n1990 GND.n1989 0.013
R3909 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/GND GND.n2009 0.013
R3910 GND.n2010 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/GND 0.013
R3911 GND.n2010 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/GND 0.013
R3912 GND.n2042 GND.n2038 0.013
R3913 GND.n2043 GND.n2042 0.013
R3914 GND.n2047 GND.n2043 0.013
R3915 x3_bar.n0 x3_bar.t1 1077.04
R3916 x3_bar.n0 x3_bar.t0 1015.9
R3917 x3_bar x3_bar.n0 81.6
R3918 x3_bar EESPFAL_4in_XOR_0/x3_bar 35.84
R3919 CLK0.n93 CLK0.t43 44.338
R3920 CLK0.n64 CLK0.t38 44.338
R3921 CLK0.n209 CLK0.t23 44.338
R3922 CLK0.n180 CLK0.t3 44.338
R3923 CLK0.n337 CLK0.t14 44.337
R3924 CLK0.n280 CLK0.t12 44.337
R3925 CLK0.n209 CLK0.t31 44.337
R3926 CLK0.n180 CLK0.t28 44.337
R3927 CLK0.n0 CLK0.t18 39.4
R3928 CLK0.n0 CLK0.t16 39.4
R3929 CLK0.n25 CLK0.t8 39.4
R3930 CLK0.n25 CLK0.t36 39.4
R3931 CLK0.n140 CLK0.t25 39.4
R3932 CLK0.n140 CLK0.t29 39.4
R3933 CLK0.n139 CLK0.t39 39.4
R3934 CLK0.n139 CLK0.t5 39.4
R3935 CLK0.n281 CLK0.t11 24.568
R3936 CLK0.n338 CLK0.t13 24.568
R3937 CLK0.n89 CLK0.t42 24.568
R3938 CLK0.n65 CLK0.t37 24.568
R3939 CLK0.n297 CLK0.t0 24
R3940 CLK0.n297 CLK0.t20 24
R3941 CLK0.n4 CLK0.t10 24
R3942 CLK0.n4 CLK0.t21 24
R3943 CLK0.n10 CLK0.t34 24
R3944 CLK0.n10 CLK0.t1 24
R3945 CLK0.n26 CLK0.t9 24
R3946 CLK0.n26 CLK0.t33 24
R3947 CLK0.n8 CLK0.t30 24
R3948 CLK0.n8 CLK0.t32 24
R3949 CLK0.n142 CLK0.t6 24
R3950 CLK0.n142 CLK0.t27 24
R3951 CLK0.n141 CLK0.t41 24
R3952 CLK0.n141 CLK0.t40 24
R3953 CLK0.n2 CLK0.t19 24
R3954 CLK0.n2 CLK0.t26 24
R3955 CLK0.n205 CLK0.t22 14.843
R3956 CLK0.n181 CLK0.t2 14.843
R3957 CLK0.n79 CLK0.n76 12.8
R3958 CLK0.n195 CLK0.n192 12.8
R3959 CLK0.n15 CLK0.n14 8.855
R3960 CLK0.n19 CLK0.n18 8.855
R3961 CLK0.n18 CLK0.n17 8.855
R3962 CLK0.n23 CLK0.n22 8.855
R3963 CLK0.n22 CLK0.n21 8.855
R3964 CLK0.n116 CLK0.n115 8.855
R3965 CLK0.n115 CLK0.n114 8.855
R3966 CLK0.n112 CLK0.n111 8.855
R3967 CLK0.n111 CLK0.n110 8.855
R3968 CLK0.n108 CLK0.n107 8.855
R3969 CLK0.n107 CLK0.n106 8.855
R3970 CLK0.n104 CLK0.n103 8.855
R3971 CLK0.n103 CLK0.n102 8.855
R3972 CLK0.n100 CLK0.n99 8.855
R3973 CLK0.n99 CLK0.n98 8.855
R3974 CLK0.n96 CLK0.n95 8.855
R3975 CLK0.n95 CLK0.n94 8.855
R3976 CLK0.n91 CLK0.n90 8.855
R3977 CLK0.n90 CLK0.n89 8.855
R3978 CLK0.n87 CLK0.n86 8.855
R3979 CLK0.n86 CLK0.n85 8.855
R3980 CLK0.n83 CLK0.n82 8.855
R3981 CLK0.n82 CLK0.n81 8.855
R3982 CLK0.n79 CLK0.n78 8.855
R3983 CLK0.n78 CLK0.n77 8.855
R3984 CLK0.n76 CLK0.n75 8.855
R3985 CLK0.n75 CLK0.n74 8.855
R3986 CLK0.n71 CLK0.n70 8.855
R3987 CLK0.n70 CLK0.n69 8.855
R3988 CLK0.n67 CLK0.n66 8.855
R3989 CLK0.n66 CLK0.n65 8.855
R3990 CLK0.n62 CLK0.n61 8.855
R3991 CLK0.n61 CLK0.n60 8.855
R3992 CLK0.n58 CLK0.n57 8.855
R3993 CLK0.n57 CLK0.n56 8.855
R3994 CLK0.n54 CLK0.n53 8.855
R3995 CLK0.n53 CLK0.n52 8.855
R3996 CLK0.n50 CLK0.n49 8.855
R3997 CLK0.n49 CLK0.n48 8.855
R3998 CLK0.n46 CLK0.n45 8.855
R3999 CLK0.n45 CLK0.n44 8.855
R4000 CLK0.n42 CLK0.n41 8.855
R4001 CLK0.n41 CLK0.n40 8.855
R4002 CLK0.n37 CLK0.n36 8.855
R4003 CLK0.n36 CLK0.n35 8.855
R4004 CLK0.n33 CLK0.n32 8.855
R4005 CLK0.n32 CLK0.n31 8.855
R4006 CLK0.n29 CLK0.n28 8.855
R4007 CLK0.n129 CLK0.n128 8.855
R4008 CLK0.n133 CLK0.n132 8.855
R4009 CLK0.n132 CLK0.n131 8.855
R4010 CLK0.n137 CLK0.n136 8.855
R4011 CLK0.n136 CLK0.n135 8.855
R4012 CLK0.n232 CLK0.n231 8.855
R4013 CLK0.n231 CLK0.n230 8.855
R4014 CLK0.n228 CLK0.n227 8.855
R4015 CLK0.n227 CLK0.n226 8.855
R4016 CLK0.n224 CLK0.n223 8.855
R4017 CLK0.n223 CLK0.n222 8.855
R4018 CLK0.n220 CLK0.n219 8.855
R4019 CLK0.n219 CLK0.n218 8.855
R4020 CLK0.n216 CLK0.n215 8.855
R4021 CLK0.n215 CLK0.n214 8.855
R4022 CLK0.n212 CLK0.n211 8.855
R4023 CLK0.n211 CLK0.n210 8.855
R4024 CLK0.n207 CLK0.n206 8.855
R4025 CLK0.n206 CLK0.n205 8.855
R4026 CLK0.n203 CLK0.n202 8.855
R4027 CLK0.n202 CLK0.n201 8.855
R4028 CLK0.n199 CLK0.n198 8.855
R4029 CLK0.n198 CLK0.n197 8.855
R4030 CLK0.n195 CLK0.n194 8.855
R4031 CLK0.n194 CLK0.n193 8.855
R4032 CLK0.n192 CLK0.n191 8.855
R4033 CLK0.n191 CLK0.n190 8.855
R4034 CLK0.n187 CLK0.n186 8.855
R4035 CLK0.n186 CLK0.n185 8.855
R4036 CLK0.n183 CLK0.n182 8.855
R4037 CLK0.n182 CLK0.n181 8.855
R4038 CLK0.n178 CLK0.n177 8.855
R4039 CLK0.n177 CLK0.n176 8.855
R4040 CLK0.n174 CLK0.n173 8.855
R4041 CLK0.n173 CLK0.n172 8.855
R4042 CLK0.n170 CLK0.n169 8.855
R4043 CLK0.n169 CLK0.n168 8.855
R4044 CLK0.n166 CLK0.n165 8.855
R4045 CLK0.n165 CLK0.n164 8.855
R4046 CLK0.n162 CLK0.n161 8.855
R4047 CLK0.n161 CLK0.n160 8.855
R4048 CLK0.n158 CLK0.n157 8.855
R4049 CLK0.n157 CLK0.n156 8.855
R4050 CLK0.n153 CLK0.n152 8.855
R4051 CLK0.n152 CLK0.n151 8.855
R4052 CLK0.n149 CLK0.n148 8.855
R4053 CLK0.n148 CLK0.n147 8.855
R4054 CLK0.n145 CLK0.n144 8.855
R4055 CLK0.n245 CLK0.n244 8.855
R4056 CLK0.n249 CLK0.n248 8.855
R4057 CLK0.n248 CLK0.n247 8.855
R4058 CLK0.n253 CLK0.n252 8.855
R4059 CLK0.n252 CLK0.n251 8.855
R4060 CLK0.n258 CLK0.n257 8.855
R4061 CLK0.n257 CLK0.n256 8.855
R4062 CLK0.n262 CLK0.n261 8.855
R4063 CLK0.n261 CLK0.n260 8.855
R4064 CLK0.n266 CLK0.n265 8.855
R4065 CLK0.n265 CLK0.n264 8.855
R4066 CLK0.n270 CLK0.n269 8.855
R4067 CLK0.n269 CLK0.n268 8.855
R4068 CLK0.n274 CLK0.n273 8.855
R4069 CLK0.n273 CLK0.n272 8.855
R4070 CLK0.n278 CLK0.n277 8.855
R4071 CLK0.n277 CLK0.n276 8.855
R4072 CLK0.n283 CLK0.n282 8.855
R4073 CLK0.n282 CLK0.n281 8.855
R4074 CLK0.n287 CLK0.n286 8.855
R4075 CLK0.n286 CLK0.n285 8.855
R4076 CLK0.n291 CLK0.n290 8.855
R4077 CLK0.n290 CLK0.n289 8.855
R4078 CLK0.n295 CLK0.n294 8.855
R4079 CLK0.n294 CLK0.n293 8.855
R4080 CLK0.n348 CLK0.n347 8.855
R4081 CLK0.n347 CLK0.n346 8.855
R4082 CLK0.n344 CLK0.n343 8.855
R4083 CLK0.n343 CLK0.n342 8.855
R4084 CLK0.n340 CLK0.n339 8.855
R4085 CLK0.n339 CLK0.n338 8.855
R4086 CLK0.n335 CLK0.n334 8.855
R4087 CLK0.n334 CLK0.n333 8.855
R4088 CLK0.n331 CLK0.n330 8.855
R4089 CLK0.n330 CLK0.n329 8.855
R4090 CLK0.n327 CLK0.n326 8.855
R4091 CLK0.n326 CLK0.n325 8.855
R4092 CLK0.n323 CLK0.n322 8.855
R4093 CLK0.n322 CLK0.n321 8.855
R4094 CLK0.n319 CLK0.n318 8.855
R4095 CLK0.n318 CLK0.n317 8.855
R4096 CLK0.n315 CLK0.n314 8.855
R4097 CLK0.n314 CLK0.n313 8.855
R4098 CLK0.n310 CLK0.n309 8.855
R4099 CLK0.n309 CLK0.n308 8.855
R4100 CLK0.n306 CLK0.n305 8.855
R4101 CLK0.n305 CLK0.n304 8.855
R4102 CLK0.n302 CLK0.n301 8.855
R4103 CLK0.n289 CLK0.t17 8.189
R4104 CLK0.n346 CLK0.t15 8.189
R4105 CLK0.n81 CLK0.t7 8.189
R4106 CLK0.n74 CLK0.t35 8.189
R4107 CLK0.n312 CLK0.n297 6.776
R4108 CLK0.n39 CLK0.n26 6.776
R4109 CLK0.n155 CLK0.n142 6.776
R4110 CLK0.n155 CLK0.n141 6.776
R4111 CLK0.n123 CLK0.n9 6.754
R4112 CLK0.n239 CLK0.n3 6.754
R4113 CLK0.n197 CLK0.t24 4.947
R4114 CLK0.n190 CLK0.t4 4.947
R4115 CLK0.n296 CLK0.n0 4.938
R4116 CLK0.n80 CLK0.n25 4.938
R4117 CLK0.n196 CLK0.n139 4.938
R4118 CLK0.n196 CLK0.n140 4.938
R4119 CLK0.n20 CLK0.n19 4.65
R4120 CLK0.n24 CLK0.n23 4.65
R4121 CLK0.n117 CLK0.n116 4.65
R4122 CLK0.n113 CLK0.n112 4.65
R4123 CLK0.n109 CLK0.n108 4.65
R4124 CLK0.n105 CLK0.n104 4.65
R4125 CLK0.n101 CLK0.n100 4.65
R4126 CLK0.n97 CLK0.n96 4.65
R4127 CLK0.n92 CLK0.n91 4.65
R4128 CLK0.n88 CLK0.n87 4.65
R4129 CLK0.n84 CLK0.n83 4.65
R4130 CLK0.n80 CLK0.n79 4.65
R4131 CLK0.n76 CLK0.n73 4.65
R4132 CLK0.n72 CLK0.n71 4.65
R4133 CLK0.n68 CLK0.n67 4.65
R4134 CLK0.n63 CLK0.n62 4.65
R4135 CLK0.n59 CLK0.n58 4.65
R4136 CLK0.n55 CLK0.n54 4.65
R4137 CLK0.n51 CLK0.n50 4.65
R4138 CLK0.n47 CLK0.n46 4.65
R4139 CLK0.n43 CLK0.n42 4.65
R4140 CLK0.n38 CLK0.n37 4.65
R4141 CLK0.n34 CLK0.n33 4.65
R4142 CLK0.n120 CLK0.n12 4.65
R4143 CLK0.n126 CLK0.n7 4.65
R4144 CLK0.n125 CLK0.n124 4.65
R4145 CLK0.n134 CLK0.n133 4.65
R4146 CLK0.n138 CLK0.n137 4.65
R4147 CLK0.n233 CLK0.n232 4.65
R4148 CLK0.n229 CLK0.n228 4.65
R4149 CLK0.n225 CLK0.n224 4.65
R4150 CLK0.n221 CLK0.n220 4.65
R4151 CLK0.n217 CLK0.n216 4.65
R4152 CLK0.n213 CLK0.n212 4.65
R4153 CLK0.n208 CLK0.n207 4.65
R4154 CLK0.n204 CLK0.n203 4.65
R4155 CLK0.n200 CLK0.n199 4.65
R4156 CLK0.n196 CLK0.n195 4.65
R4157 CLK0.n192 CLK0.n189 4.65
R4158 CLK0.n188 CLK0.n187 4.65
R4159 CLK0.n184 CLK0.n183 4.65
R4160 CLK0.n179 CLK0.n178 4.65
R4161 CLK0.n175 CLK0.n174 4.65
R4162 CLK0.n171 CLK0.n170 4.65
R4163 CLK0.n167 CLK0.n166 4.65
R4164 CLK0.n163 CLK0.n162 4.65
R4165 CLK0.n159 CLK0.n158 4.65
R4166 CLK0.n154 CLK0.n153 4.65
R4167 CLK0.n150 CLK0.n149 4.65
R4168 CLK0.n236 CLK0.n6 4.65
R4169 CLK0.n242 CLK0.n1 4.65
R4170 CLK0.n241 CLK0.n240 4.65
R4171 CLK0.n250 CLK0.n249 4.65
R4172 CLK0.n254 CLK0.n253 4.65
R4173 CLK0.n259 CLK0.n258 4.65
R4174 CLK0.n263 CLK0.n262 4.65
R4175 CLK0.n267 CLK0.n266 4.65
R4176 CLK0.n271 CLK0.n270 4.65
R4177 CLK0.n275 CLK0.n274 4.65
R4178 CLK0.n279 CLK0.n278 4.65
R4179 CLK0.n284 CLK0.n283 4.65
R4180 CLK0.n288 CLK0.n287 4.65
R4181 CLK0.n292 CLK0.n291 4.65
R4182 CLK0.n296 CLK0.n295 4.65
R4183 CLK0.n349 CLK0.n348 4.65
R4184 CLK0.n345 CLK0.n344 4.65
R4185 CLK0.n341 CLK0.n340 4.65
R4186 CLK0.n336 CLK0.n335 4.65
R4187 CLK0.n332 CLK0.n331 4.65
R4188 CLK0.n328 CLK0.n327 4.65
R4189 CLK0.n324 CLK0.n323 4.65
R4190 CLK0.n320 CLK0.n319 4.65
R4191 CLK0.n316 CLK0.n315 4.65
R4192 CLK0.n311 CLK0.n310 4.65
R4193 CLK0.n307 CLK0.n306 4.65
R4194 CLK0.n303 CLK0.n302 4.65
R4195 CLK0.n6 CLK0.n5 3.715
R4196 CLK0.n12 CLK0.n11 3.715
R4197 CLK0.n122 CLK0.n121 3.039
R4198 CLK0.n238 CLK0.n237 3.039
R4199 CLK0.n299 CLK0.n298 3.037
R4200 CLK0.n246 CLK0.n245 2.682
R4201 CLK0.n16 CLK0.n15 2.682
R4202 CLK0.n30 CLK0.n29 2.682
R4203 CLK0.n130 CLK0.n129 2.682
R4204 CLK0.n146 CLK0.n145 2.682
R4205 CLK0.n5 CLK0.n4 2.57
R4206 CLK0.n11 CLK0.n10 2.57
R4207 CLK0.n9 CLK0.n8 2.57
R4208 CLK0.n3 CLK0.n2 2.57
R4209 CLK0.n123 CLK0.n122 2.224
R4210 CLK0.n239 CLK0.n238 2.224
R4211 CLK0.n119 CLK0.n118 2.203
R4212 CLK0.n234 CLK0.n126 2.203
R4213 CLK0.n235 CLK0.n234 2.203
R4214 CLK0.n255 CLK0.n242 2.203
R4215 CLK0.n128 CLK0.n127 1.722
R4216 CLK0.n144 CLK0.n143 1.722
R4217 CLK0.n244 CLK0.n243 1.655
R4218 CLK0.n14 CLK0.n13 1.655
R4219 CLK0.n28 CLK0.n27 1.655
R4220 CLK0.n301 CLK0.n300 1.655
R4221 CLK0.n250 CLK0.n246 1.096
R4222 CLK0.n20 CLK0.n16 1.095
R4223 CLK0.n34 CLK0.n30 1.095
R4224 CLK0.n134 CLK0.n130 1.095
R4225 CLK0.n150 CLK0.n146 1.095
R4226 CLK0.n299 EESPFAL_4in_XOR_0/CLK 0.764
R4227 CLK0.n120 CLK0.n119 0.125
R4228 CLK0.n126 CLK0.n125 0.125
R4229 CLK0.n236 CLK0.n235 0.125
R4230 CLK0.n242 CLK0.n241 0.125
R4231 CLK0.n125 CLK0.n123 0.12
R4232 CLK0.n241 CLK0.n239 0.12
R4233 CLK0.n122 CLK0.n120 0.119
R4234 CLK0.n238 CLK0.n236 0.119
R4235 CLK0.n24 CLK0.n20 0.1
R4236 CLK0.n117 CLK0.n113 0.1
R4237 CLK0.n113 CLK0.n109 0.1
R4238 CLK0.n109 CLK0.n105 0.1
R4239 CLK0.n105 CLK0.n101 0.1
R4240 CLK0.n101 CLK0.n97 0.1
R4241 CLK0.n92 CLK0.n88 0.1
R4242 CLK0.n88 CLK0.n84 0.1
R4243 CLK0.n84 CLK0.n80 0.1
R4244 CLK0.n73 CLK0.n72 0.1
R4245 CLK0.n72 CLK0.n68 0.1
R4246 CLK0.n63 CLK0.n59 0.1
R4247 CLK0.n59 CLK0.n55 0.1
R4248 CLK0.n55 CLK0.n51 0.1
R4249 CLK0.n51 CLK0.n47 0.1
R4250 CLK0.n47 CLK0.n43 0.1
R4251 CLK0.n38 CLK0.n34 0.1
R4252 CLK0.n138 CLK0.n134 0.1
R4253 CLK0.n233 CLK0.n229 0.1
R4254 CLK0.n229 CLK0.n225 0.1
R4255 CLK0.n225 CLK0.n221 0.1
R4256 CLK0.n221 CLK0.n217 0.1
R4257 CLK0.n217 CLK0.n213 0.1
R4258 CLK0.n208 CLK0.n204 0.1
R4259 CLK0.n204 CLK0.n200 0.1
R4260 CLK0.n200 CLK0.n196 0.1
R4261 CLK0.n189 CLK0.n188 0.1
R4262 CLK0.n188 CLK0.n184 0.1
R4263 CLK0.n179 CLK0.n175 0.1
R4264 CLK0.n175 CLK0.n171 0.1
R4265 CLK0.n171 CLK0.n167 0.1
R4266 CLK0.n167 CLK0.n163 0.1
R4267 CLK0.n163 CLK0.n159 0.1
R4268 CLK0.n154 CLK0.n150 0.1
R4269 CLK0.n254 CLK0.n250 0.1
R4270 CLK0.n263 CLK0.n259 0.1
R4271 CLK0.n267 CLK0.n263 0.1
R4272 CLK0.n271 CLK0.n267 0.1
R4273 CLK0.n275 CLK0.n271 0.1
R4274 CLK0.n279 CLK0.n275 0.1
R4275 CLK0.n288 CLK0.n284 0.1
R4276 CLK0.n292 CLK0.n288 0.1
R4277 CLK0.n296 CLK0.n292 0.1
R4278 CLK0.n349 CLK0.n345 0.1
R4279 CLK0.n345 CLK0.n341 0.1
R4280 CLK0.n336 CLK0.n332 0.1
R4281 CLK0.n332 CLK0.n328 0.1
R4282 CLK0.n328 CLK0.n324 0.1
R4283 CLK0.n324 CLK0.n320 0.1
R4284 CLK0.n320 CLK0.n316 0.1
R4285 CLK0.n311 CLK0.n307 0.1
R4286 CLK0.n307 CLK0.n303 0.1
R4287 CLK0.n303 CLK0.n299 0.095
R4288 CLK0.n118 CLK0.n117 0.075
R4289 CLK0.n93 CLK0.n92 0.075
R4290 CLK0.n73 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/CLK 0.075
R4291 CLK0.n68 CLK0.n64 0.075
R4292 CLK0.n43 CLK0.n39 0.075
R4293 CLK0.n234 CLK0.n233 0.075
R4294 CLK0.n209 CLK0.n208 0.075
R4295 CLK0.n189 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_1/CLK 0.075
R4296 CLK0.n184 CLK0.n180 0.075
R4297 CLK0.n159 CLK0.n155 0.075
R4298 CLK0.n259 CLK0.n255 0.075
R4299 CLK0.n284 CLK0.n280 0.075
R4300 CLK0 CLK0.n349 0.075
R4301 CLK0.n341 CLK0.n337 0.075
R4302 CLK0.n316 CLK0.n312 0.075
R4303 CLK0.n118 CLK0.n24 0.025
R4304 CLK0.n97 CLK0.n93 0.025
R4305 CLK0.n80 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/CLK 0.025
R4306 CLK0.n64 CLK0.n63 0.025
R4307 CLK0.n39 CLK0.n38 0.025
R4308 CLK0.n234 CLK0.n138 0.025
R4309 CLK0.n213 CLK0.n209 0.025
R4310 CLK0.n196 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_1/CLK 0.025
R4311 CLK0.n180 CLK0.n179 0.025
R4312 CLK0.n155 CLK0.n154 0.025
R4313 CLK0.n255 CLK0.n254 0.025
R4314 CLK0.n280 CLK0.n279 0.025
R4315 CLK0 CLK0.n296 0.025
R4316 CLK0.n337 CLK0.n336 0.025
R4317 CLK0.n312 CLK0.n311 0.025
R4318 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t9 1074.82
R4319 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t6 819.4
R4320 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t8 514.133
R4321 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t7 305.266
R4322 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n6 260.333
R4323 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n5 192
R4324 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n1 166.734
R4325 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n4 105.6
R4326 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t1 97.937
R4327 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t3 97.937
R4328 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n2 76
R4329 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n0 73.937
R4330 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n3 57.6
R4331 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t0 39.4
R4332 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t2 39.4
R4333 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t5 24
R4334 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t4 24
R4335 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT 3.2
R4336 CLK1.n277 CLK1.n276 407.048
R4337 CLK1.n232 CLK1.n223 407.048
R4338 CLK1.n1620 CLK1.n1619 407.048
R4339 CLK1.n1553 CLK1.n1552 407.048
R4340 CLK1.n1547 CLK1.n1546 407.048
R4341 CLK1.n1512 CLK1.n1503 407.048
R4342 CLK1.n1253 CLK1.n1252 407.048
R4343 CLK1.n1197 CLK1.n316 407.048
R4344 CLK1.n387 CLK1.n386 407.048
R4345 CLK1.n352 CLK1.n343 407.048
R4346 CLK1.n475 CLK1.n474 407.048
R4347 CLK1.n440 CLK1.n431 407.048
R4348 CLK1.n999 CLK1.n998 407.048
R4349 CLK1.n484 CLK1.n407 407.048
R4350 CLK1.n988 CLK1.n987 407.048
R4351 CLK1.n921 CLK1.n920 407.048
R4352 CLK1.n915 CLK1.n914 407.048
R4353 CLK1.n880 CLK1.n871 407.048
R4354 CLK1.n621 CLK1.n620 407.048
R4355 CLK1.n565 CLK1.n556 407.048
R4356 CLK1.n803 CLK1.n802 407.048
R4357 CLK1.n736 CLK1.n735 407.048
R4358 CLK1.n730 CLK1.n729 407.048
R4359 CLK1.n695 CLK1.n686 407.048
R4360 CLK1.n1435 CLK1.n1434 407.048
R4361 CLK1.n1368 CLK1.n1367 407.048
R4362 CLK1.n1362 CLK1.n1361 407.048
R4363 CLK1.n1327 CLK1.n1318 407.048
R4364 CLK1.n267 CLK1.n198 400
R4365 CLK1.n276 CLK1.n198 400
R4366 CLK1.n233 CLK1.n232 400
R4367 CLK1.n234 CLK1.n233 400
R4368 CLK1.n1607 CLK1.n1453 400
R4369 CLK1.n1608 CLK1.n1607 400
R4370 CLK1.n1609 CLK1.n1608 400
R4371 CLK1.n1609 CLK1.n1445 400
R4372 CLK1.n1619 CLK1.n1445 400
R4373 CLK1.n1553 CLK1.n1475 400
R4374 CLK1.n1562 CLK1.n1475 400
R4375 CLK1.n1563 CLK1.n1562 400
R4376 CLK1.n1564 CLK1.n1563 400
R4377 CLK1.n1564 CLK1.n1469 400
R4378 CLK1.n1242 CLK1.n1241 400
R4379 CLK1.n1243 CLK1.n1242 400
R4380 CLK1.n1243 CLK1.n285 400
R4381 CLK1.n1252 CLK1.n285 400
R4382 CLK1.n1198 CLK1.n1197 400
R4383 CLK1.n1199 CLK1.n1198 400
R4384 CLK1.n1199 CLK1.n310 400
R4385 CLK1.n1207 CLK1.n310 400
R4386 CLK1.n1010 CLK1.n506 400
R4387 CLK1.n1010 CLK1.n1009 400
R4388 CLK1.n1009 CLK1.n1008 400
R4389 CLK1.n1008 CLK1.n513 400
R4390 CLK1.n999 CLK1.n513 400
R4391 CLK1.n485 CLK1.n484 400
R4392 CLK1.n1050 CLK1.n485 400
R4393 CLK1.n1050 CLK1.n1049 400
R4394 CLK1.n1049 CLK1.n1048 400
R4395 CLK1.n1048 CLK1.n486 400
R4396 CLK1.n975 CLK1.n821 400
R4397 CLK1.n976 CLK1.n975 400
R4398 CLK1.n977 CLK1.n976 400
R4399 CLK1.n977 CLK1.n813 400
R4400 CLK1.n987 CLK1.n813 400
R4401 CLK1.n921 CLK1.n843 400
R4402 CLK1.n930 CLK1.n843 400
R4403 CLK1.n931 CLK1.n930 400
R4404 CLK1.n932 CLK1.n931 400
R4405 CLK1.n932 CLK1.n837 400
R4406 CLK1.n610 CLK1.n609 400
R4407 CLK1.n611 CLK1.n610 400
R4408 CLK1.n611 CLK1.n525 400
R4409 CLK1.n620 CLK1.n525 400
R4410 CLK1.n566 CLK1.n565 400
R4411 CLK1.n567 CLK1.n566 400
R4412 CLK1.n567 CLK1.n550 400
R4413 CLK1.n575 CLK1.n550 400
R4414 CLK1.n790 CLK1.n636 400
R4415 CLK1.n791 CLK1.n790 400
R4416 CLK1.n792 CLK1.n791 400
R4417 CLK1.n792 CLK1.n628 400
R4418 CLK1.n802 CLK1.n628 400
R4419 CLK1.n736 CLK1.n658 400
R4420 CLK1.n745 CLK1.n658 400
R4421 CLK1.n746 CLK1.n745 400
R4422 CLK1.n747 CLK1.n746 400
R4423 CLK1.n747 CLK1.n652 400
R4424 CLK1.n1422 CLK1.n1268 400
R4425 CLK1.n1423 CLK1.n1422 400
R4426 CLK1.n1424 CLK1.n1423 400
R4427 CLK1.n1424 CLK1.n1260 400
R4428 CLK1.n1434 CLK1.n1260 400
R4429 CLK1.n1368 CLK1.n1290 400
R4430 CLK1.n1377 CLK1.n1290 400
R4431 CLK1.n1378 CLK1.n1377 400
R4432 CLK1.n1379 CLK1.n1378 400
R4433 CLK1.n1379 CLK1.n1284 400
R4434 CLK1.n267 CLK1.n266 366.379
R4435 CLK1.n234 CLK1.n217 366.379
R4436 CLK1.n1599 CLK1.n1453 366.379
R4437 CLK1.n1573 CLK1.n1469 366.379
R4438 CLK1.n1546 CLK1.n1485 366.379
R4439 CLK1.n1513 CLK1.n1512 366.379
R4440 CLK1.n1241 CLK1.n292 366.379
R4441 CLK1.n1208 CLK1.n1207 366.379
R4442 CLK1.n386 CLK1.n325 366.379
R4443 CLK1.n353 CLK1.n352 366.379
R4444 CLK1.n474 CLK1.n413 366.379
R4445 CLK1.n441 CLK1.n440 366.379
R4446 CLK1.n1018 CLK1.n506 366.379
R4447 CLK1.n1040 CLK1.n486 366.379
R4448 CLK1.n967 CLK1.n821 366.379
R4449 CLK1.n941 CLK1.n837 366.379
R4450 CLK1.n914 CLK1.n853 366.379
R4451 CLK1.n881 CLK1.n880 366.379
R4452 CLK1.n609 CLK1.n532 366.379
R4453 CLK1.n576 CLK1.n575 366.379
R4454 CLK1.n782 CLK1.n636 366.379
R4455 CLK1.n756 CLK1.n652 366.379
R4456 CLK1.n729 CLK1.n668 366.379
R4457 CLK1.n696 CLK1.n695 366.379
R4458 CLK1.n1414 CLK1.n1268 366.379
R4459 CLK1.n1388 CLK1.n1284 366.379
R4460 CLK1.n1361 CLK1.n1300 366.379
R4461 CLK1.n1328 CLK1.n1327 366.379
R4462 CLK1.n1175 CLK1.n1174 240.502
R4463 CLK1.n1118 CLK1.n1117 240.501
R4464 CLK1.n1130 CLK1.n1103 236.76
R4465 CLK1.n1130 CLK1.n1129 236.76
R4466 CLK1.n1129 CLK1.n1128 236.76
R4467 CLK1.n1128 CLK1.n1104 236.76
R4468 CLK1.n1119 CLK1.n1104 236.76
R4469 CLK1.n1119 CLK1.n1118 236.76
R4470 CLK1.n1174 CLK1.n1173 236.76
R4471 CLK1.n1173 CLK1.n395 236.76
R4472 CLK1.n1164 CLK1.n395 236.76
R4473 CLK1.n1164 CLK1.n1163 236.76
R4474 CLK1.n1163 CLK1.n1162 236.76
R4475 CLK1.n1162 CLK1.n1069 236.76
R4476 CLK1.n1103 CLK1.n1095 215.793
R4477 CLK1.n1074 CLK1.n1069 215.793
R4478 CLK1.n243 CLK1.n217 131.034
R4479 CLK1.n244 CLK1.n243 131.034
R4480 CLK1.n246 CLK1.n245 131.034
R4481 CLK1.n256 CLK1.n255 131.034
R4482 CLK1.n265 CLK1.n205 131.034
R4483 CLK1.n266 CLK1.n265 131.034
R4484 CLK1.n1574 CLK1.n1573 131.034
R4485 CLK1.n1575 CLK1.n1574 131.034
R4486 CLK1.n1585 CLK1.n1463 131.034
R4487 CLK1.n1588 CLK1.n1587 131.034
R4488 CLK1.n1598 CLK1.n1597 131.034
R4489 CLK1.n1599 CLK1.n1598 131.034
R4490 CLK1.n1515 CLK1.n1513 131.034
R4491 CLK1.n1515 CLK1.n1514 131.034
R4492 CLK1.n1525 CLK1.n1524 131.034
R4493 CLK1.n1535 CLK1.n1491 131.034
R4494 CLK1.n1537 CLK1.n1536 131.034
R4495 CLK1.n1537 CLK1.n1485 131.034
R4496 CLK1.n1210 CLK1.n1208 131.034
R4497 CLK1.n1210 CLK1.n1209 131.034
R4498 CLK1.n1220 CLK1.n1219 131.034
R4499 CLK1.n1230 CLK1.n298 131.034
R4500 CLK1.n1232 CLK1.n1231 131.034
R4501 CLK1.n1232 CLK1.n292 131.034
R4502 CLK1.n355 CLK1.n353 131.034
R4503 CLK1.n355 CLK1.n354 131.034
R4504 CLK1.n365 CLK1.n364 131.034
R4505 CLK1.n375 CLK1.n331 131.034
R4506 CLK1.n377 CLK1.n376 131.034
R4507 CLK1.n377 CLK1.n325 131.034
R4508 CLK1.n443 CLK1.n441 131.034
R4509 CLK1.n443 CLK1.n442 131.034
R4510 CLK1.n453 CLK1.n452 131.034
R4511 CLK1.n463 CLK1.n419 131.034
R4512 CLK1.n465 CLK1.n464 131.034
R4513 CLK1.n465 CLK1.n413 131.034
R4514 CLK1.n1040 CLK1.n1039 131.034
R4515 CLK1.n1039 CLK1.n1038 131.034
R4516 CLK1.n1030 CLK1.n499 131.034
R4517 CLK1.n1028 CLK1.n500 131.034
R4518 CLK1.n1020 CLK1.n1019 131.034
R4519 CLK1.n1019 CLK1.n1018 131.034
R4520 CLK1.n942 CLK1.n941 131.034
R4521 CLK1.n943 CLK1.n942 131.034
R4522 CLK1.n953 CLK1.n831 131.034
R4523 CLK1.n956 CLK1.n955 131.034
R4524 CLK1.n966 CLK1.n965 131.034
R4525 CLK1.n967 CLK1.n966 131.034
R4526 CLK1.n883 CLK1.n881 131.034
R4527 CLK1.n883 CLK1.n882 131.034
R4528 CLK1.n893 CLK1.n892 131.034
R4529 CLK1.n903 CLK1.n859 131.034
R4530 CLK1.n905 CLK1.n904 131.034
R4531 CLK1.n905 CLK1.n853 131.034
R4532 CLK1.n578 CLK1.n576 131.034
R4533 CLK1.n578 CLK1.n577 131.034
R4534 CLK1.n588 CLK1.n587 131.034
R4535 CLK1.n598 CLK1.n538 131.034
R4536 CLK1.n600 CLK1.n599 131.034
R4537 CLK1.n600 CLK1.n532 131.034
R4538 CLK1.n757 CLK1.n756 131.034
R4539 CLK1.n758 CLK1.n757 131.034
R4540 CLK1.n768 CLK1.n646 131.034
R4541 CLK1.n771 CLK1.n770 131.034
R4542 CLK1.n781 CLK1.n780 131.034
R4543 CLK1.n782 CLK1.n781 131.034
R4544 CLK1.n698 CLK1.n696 131.034
R4545 CLK1.n698 CLK1.n697 131.034
R4546 CLK1.n708 CLK1.n707 131.034
R4547 CLK1.n718 CLK1.n674 131.034
R4548 CLK1.n720 CLK1.n719 131.034
R4549 CLK1.n720 CLK1.n668 131.034
R4550 CLK1.n1389 CLK1.n1388 131.034
R4551 CLK1.n1390 CLK1.n1389 131.034
R4552 CLK1.n1400 CLK1.n1278 131.034
R4553 CLK1.n1403 CLK1.n1402 131.034
R4554 CLK1.n1413 CLK1.n1412 131.034
R4555 CLK1.n1414 CLK1.n1413 131.034
R4556 CLK1.n1330 CLK1.n1328 131.034
R4557 CLK1.n1330 CLK1.n1329 131.034
R4558 CLK1.n1340 CLK1.n1339 131.034
R4559 CLK1.n1350 CLK1.n1306 131.034
R4560 CLK1.n1352 CLK1.n1351 131.034
R4561 CLK1.n1352 CLK1.n1300 131.034
R4562 CLK1.n254 CLK1.t89 122.844
R4563 CLK1.t140 CLK1.n254 122.844
R4564 CLK1.n1586 CLK1.t109 122.844
R4565 CLK1.t152 CLK1.n1586 122.844
R4566 CLK1.n1526 CLK1.t2 122.844
R4567 CLK1.n1526 CLK1.t83 122.844
R4568 CLK1.n1221 CLK1.t129 122.844
R4569 CLK1.n1221 CLK1.t14 122.844
R4570 CLK1.n366 CLK1.t125 122.844
R4571 CLK1.n366 CLK1.t179 122.844
R4572 CLK1.n454 CLK1.t114 122.844
R4573 CLK1.n454 CLK1.t60 122.844
R4574 CLK1.t64 CLK1.n1029 122.844
R4575 CLK1.n1029 CLK1.t43 122.844
R4576 CLK1.n954 CLK1.t135 122.844
R4577 CLK1.t103 CLK1.n954 122.844
R4578 CLK1.n894 CLK1.t157 122.844
R4579 CLK1.n894 CLK1.t6 122.844
R4580 CLK1.n589 CLK1.t142 122.844
R4581 CLK1.n589 CLK1.t159 122.844
R4582 CLK1.n769 CLK1.t46 122.844
R4583 CLK1.t183 CLK1.n769 122.844
R4584 CLK1.n709 CLK1.t67 122.844
R4585 CLK1.n709 CLK1.t71 122.844
R4586 CLK1.n1401 CLK1.t171 122.844
R4587 CLK1.t148 CLK1.n1401 122.844
R4588 CLK1.n1341 CLK1.t27 122.844
R4589 CLK1.n1341 CLK1.t20 122.844
R4590 CLK1.n246 CLK1.t87 106.465
R4591 CLK1.n256 CLK1.t138 106.465
R4592 CLK1.t107 CLK1.n1463 106.465
R4593 CLK1.n1587 CLK1.t49 106.465
R4594 CLK1.n1524 CLK1.t0 106.465
R4595 CLK1.t85 CLK1.n1535 106.465
R4596 CLK1.n1219 CLK1.t131 106.465
R4597 CLK1.t16 CLK1.n1230 106.465
R4598 CLK1.n364 CLK1.t127 106.465
R4599 CLK1.t181 CLK1.n375 106.465
R4600 CLK1.n452 CLK1.t116 106.465
R4601 CLK1.t62 CLK1.n463 106.465
R4602 CLK1.n499 CLK1.t123 106.465
R4603 CLK1.t169 CLK1.n500 106.465
R4604 CLK1.t133 CLK1.n831 106.465
R4605 CLK1.n955 CLK1.t57 106.465
R4606 CLK1.n892 CLK1.t155 106.465
R4607 CLK1.t4 CLK1.n903 106.465
R4608 CLK1.n587 CLK1.t144 106.465
R4609 CLK1.t161 CLK1.n598 106.465
R4610 CLK1.t12 CLK1.n646 106.465
R4611 CLK1.n770 CLK1.t185 106.465
R4612 CLK1.n707 CLK1.t69 106.465
R4613 CLK1.t73 CLK1.n718 106.465
R4614 CLK1.t146 CLK1.n1278 106.465
R4615 CLK1.n1402 CLK1.t195 106.465
R4616 CLK1.n1339 CLK1.t25 106.465
R4617 CLK1.t18 CLK1.n1350 106.465
R4618 CLK1.n231 CLK1.n224 96
R4619 CLK1.n231 CLK1.n222 96
R4620 CLK1.n235 CLK1.n222 96
R4621 CLK1.n235 CLK1.n218 96
R4622 CLK1.n242 CLK1.n218 96
R4623 CLK1.n242 CLK1.n216 96
R4624 CLK1.n247 CLK1.n216 96
R4625 CLK1.n247 CLK1.n211 96
R4626 CLK1.n253 CLK1.n211 96
R4627 CLK1.n253 CLK1.n210 96
R4628 CLK1.n257 CLK1.n210 96
R4629 CLK1.n257 CLK1.n206 96
R4630 CLK1.n264 CLK1.n206 96
R4631 CLK1.n264 CLK1.n204 96
R4632 CLK1.n268 CLK1.n204 96
R4633 CLK1.n268 CLK1.n199 96
R4634 CLK1.n275 CLK1.n199 96
R4635 CLK1.n275 CLK1.n197 96
R4636 CLK1.n1554 CLK1.n1481 96
R4637 CLK1.n1554 CLK1.n1476 96
R4638 CLK1.n1561 CLK1.n1476 96
R4639 CLK1.n1561 CLK1.n1474 96
R4640 CLK1.n1565 CLK1.n1474 96
R4641 CLK1.n1565 CLK1.n1470 96
R4642 CLK1.n1572 CLK1.n1470 96
R4643 CLK1.n1572 CLK1.n1468 96
R4644 CLK1.n1576 CLK1.n1468 96
R4645 CLK1.n1576 CLK1.n1464 96
R4646 CLK1.n1584 CLK1.n1464 96
R4647 CLK1.n1584 CLK1.n1462 96
R4648 CLK1.n1589 CLK1.n1462 96
R4649 CLK1.n1589 CLK1.n1459 96
R4650 CLK1.n1596 CLK1.n1459 96
R4651 CLK1.n1596 CLK1.n1458 96
R4652 CLK1.n1600 CLK1.n1458 96
R4653 CLK1.n1600 CLK1.n1454 96
R4654 CLK1.n1606 CLK1.n1454 96
R4655 CLK1.n1606 CLK1.n1452 96
R4656 CLK1.n1610 CLK1.n1452 96
R4657 CLK1.n1610 CLK1.n1446 96
R4658 CLK1.n1618 CLK1.n1446 96
R4659 CLK1.n1618 CLK1.n1444 96
R4660 CLK1.n1511 CLK1.n1504 96
R4661 CLK1.n1511 CLK1.n1502 96
R4662 CLK1.n1516 CLK1.n1502 96
R4663 CLK1.n1516 CLK1.n1498 96
R4664 CLK1.n1523 CLK1.n1498 96
R4665 CLK1.n1523 CLK1.n1497 96
R4666 CLK1.n1527 CLK1.n1497 96
R4667 CLK1.n1527 CLK1.n1492 96
R4668 CLK1.n1534 CLK1.n1492 96
R4669 CLK1.n1534 CLK1.n1490 96
R4670 CLK1.n1538 CLK1.n1490 96
R4671 CLK1.n1538 CLK1.n1486 96
R4672 CLK1.n1545 CLK1.n1486 96
R4673 CLK1.n1545 CLK1.n1484 96
R4674 CLK1.n1196 CLK1.n317 96
R4675 CLK1.n1196 CLK1.n315 96
R4676 CLK1.n1200 CLK1.n315 96
R4677 CLK1.n1200 CLK1.n311 96
R4678 CLK1.n1206 CLK1.n311 96
R4679 CLK1.n1206 CLK1.n309 96
R4680 CLK1.n1211 CLK1.n309 96
R4681 CLK1.n1211 CLK1.n305 96
R4682 CLK1.n1218 CLK1.n305 96
R4683 CLK1.n1218 CLK1.n304 96
R4684 CLK1.n1222 CLK1.n304 96
R4685 CLK1.n1222 CLK1.n299 96
R4686 CLK1.n1229 CLK1.n299 96
R4687 CLK1.n1229 CLK1.n297 96
R4688 CLK1.n1233 CLK1.n297 96
R4689 CLK1.n1233 CLK1.n293 96
R4690 CLK1.n1240 CLK1.n293 96
R4691 CLK1.n1240 CLK1.n291 96
R4692 CLK1.n1244 CLK1.n291 96
R4693 CLK1.n1244 CLK1.n286 96
R4694 CLK1.n1251 CLK1.n286 96
R4695 CLK1.n1251 CLK1.n284 96
R4696 CLK1.n351 CLK1.n344 96
R4697 CLK1.n351 CLK1.n342 96
R4698 CLK1.n356 CLK1.n342 96
R4699 CLK1.n356 CLK1.n338 96
R4700 CLK1.n363 CLK1.n338 96
R4701 CLK1.n363 CLK1.n337 96
R4702 CLK1.n367 CLK1.n337 96
R4703 CLK1.n367 CLK1.n332 96
R4704 CLK1.n374 CLK1.n332 96
R4705 CLK1.n374 CLK1.n330 96
R4706 CLK1.n378 CLK1.n330 96
R4707 CLK1.n378 CLK1.n326 96
R4708 CLK1.n385 CLK1.n326 96
R4709 CLK1.n385 CLK1.n324 96
R4710 CLK1.n439 CLK1.n432 96
R4711 CLK1.n439 CLK1.n430 96
R4712 CLK1.n444 CLK1.n430 96
R4713 CLK1.n444 CLK1.n426 96
R4714 CLK1.n451 CLK1.n426 96
R4715 CLK1.n451 CLK1.n425 96
R4716 CLK1.n455 CLK1.n425 96
R4717 CLK1.n455 CLK1.n420 96
R4718 CLK1.n462 CLK1.n420 96
R4719 CLK1.n462 CLK1.n418 96
R4720 CLK1.n466 CLK1.n418 96
R4721 CLK1.n466 CLK1.n414 96
R4722 CLK1.n473 CLK1.n414 96
R4723 CLK1.n473 CLK1.n412 96
R4724 CLK1.n483 CLK1.n408 96
R4725 CLK1.n483 CLK1.n405 96
R4726 CLK1.n1051 CLK1.n405 96
R4727 CLK1.n1051 CLK1.n406 96
R4728 CLK1.n1047 CLK1.n406 96
R4729 CLK1.n1047 CLK1.n487 96
R4730 CLK1.n1041 CLK1.n487 96
R4731 CLK1.n1041 CLK1.n491 96
R4732 CLK1.n1037 CLK1.n491 96
R4733 CLK1.n1037 CLK1.n492 96
R4734 CLK1.n1031 CLK1.n492 96
R4735 CLK1.n1031 CLK1.n498 96
R4736 CLK1.n1027 CLK1.n498 96
R4737 CLK1.n1027 CLK1.n501 96
R4738 CLK1.n1021 CLK1.n501 96
R4739 CLK1.n1021 CLK1.n505 96
R4740 CLK1.n1017 CLK1.n505 96
R4741 CLK1.n1017 CLK1.n507 96
R4742 CLK1.n1011 CLK1.n507 96
R4743 CLK1.n1011 CLK1.n512 96
R4744 CLK1.n1007 CLK1.n512 96
R4745 CLK1.n1007 CLK1.n514 96
R4746 CLK1.n1000 CLK1.n514 96
R4747 CLK1.n1000 CLK1.n519 96
R4748 CLK1.n922 CLK1.n849 96
R4749 CLK1.n922 CLK1.n844 96
R4750 CLK1.n929 CLK1.n844 96
R4751 CLK1.n929 CLK1.n842 96
R4752 CLK1.n933 CLK1.n842 96
R4753 CLK1.n933 CLK1.n838 96
R4754 CLK1.n940 CLK1.n838 96
R4755 CLK1.n940 CLK1.n836 96
R4756 CLK1.n944 CLK1.n836 96
R4757 CLK1.n944 CLK1.n832 96
R4758 CLK1.n952 CLK1.n832 96
R4759 CLK1.n952 CLK1.n830 96
R4760 CLK1.n957 CLK1.n830 96
R4761 CLK1.n957 CLK1.n827 96
R4762 CLK1.n964 CLK1.n827 96
R4763 CLK1.n964 CLK1.n826 96
R4764 CLK1.n968 CLK1.n826 96
R4765 CLK1.n968 CLK1.n822 96
R4766 CLK1.n974 CLK1.n822 96
R4767 CLK1.n974 CLK1.n820 96
R4768 CLK1.n978 CLK1.n820 96
R4769 CLK1.n978 CLK1.n814 96
R4770 CLK1.n986 CLK1.n814 96
R4771 CLK1.n986 CLK1.n812 96
R4772 CLK1.n879 CLK1.n872 96
R4773 CLK1.n879 CLK1.n870 96
R4774 CLK1.n884 CLK1.n870 96
R4775 CLK1.n884 CLK1.n866 96
R4776 CLK1.n891 CLK1.n866 96
R4777 CLK1.n891 CLK1.n865 96
R4778 CLK1.n895 CLK1.n865 96
R4779 CLK1.n895 CLK1.n860 96
R4780 CLK1.n902 CLK1.n860 96
R4781 CLK1.n902 CLK1.n858 96
R4782 CLK1.n906 CLK1.n858 96
R4783 CLK1.n906 CLK1.n854 96
R4784 CLK1.n913 CLK1.n854 96
R4785 CLK1.n913 CLK1.n852 96
R4786 CLK1.n564 CLK1.n557 96
R4787 CLK1.n564 CLK1.n555 96
R4788 CLK1.n568 CLK1.n555 96
R4789 CLK1.n568 CLK1.n551 96
R4790 CLK1.n574 CLK1.n551 96
R4791 CLK1.n574 CLK1.n549 96
R4792 CLK1.n579 CLK1.n549 96
R4793 CLK1.n579 CLK1.n545 96
R4794 CLK1.n586 CLK1.n545 96
R4795 CLK1.n586 CLK1.n544 96
R4796 CLK1.n590 CLK1.n544 96
R4797 CLK1.n590 CLK1.n539 96
R4798 CLK1.n597 CLK1.n539 96
R4799 CLK1.n597 CLK1.n537 96
R4800 CLK1.n601 CLK1.n537 96
R4801 CLK1.n601 CLK1.n533 96
R4802 CLK1.n608 CLK1.n533 96
R4803 CLK1.n608 CLK1.n531 96
R4804 CLK1.n612 CLK1.n531 96
R4805 CLK1.n612 CLK1.n526 96
R4806 CLK1.n619 CLK1.n526 96
R4807 CLK1.n619 CLK1.n524 96
R4808 CLK1.n737 CLK1.n664 96
R4809 CLK1.n737 CLK1.n659 96
R4810 CLK1.n744 CLK1.n659 96
R4811 CLK1.n744 CLK1.n657 96
R4812 CLK1.n748 CLK1.n657 96
R4813 CLK1.n748 CLK1.n653 96
R4814 CLK1.n755 CLK1.n653 96
R4815 CLK1.n755 CLK1.n651 96
R4816 CLK1.n759 CLK1.n651 96
R4817 CLK1.n759 CLK1.n647 96
R4818 CLK1.n767 CLK1.n647 96
R4819 CLK1.n767 CLK1.n645 96
R4820 CLK1.n772 CLK1.n645 96
R4821 CLK1.n772 CLK1.n642 96
R4822 CLK1.n779 CLK1.n642 96
R4823 CLK1.n779 CLK1.n641 96
R4824 CLK1.n783 CLK1.n641 96
R4825 CLK1.n783 CLK1.n637 96
R4826 CLK1.n789 CLK1.n637 96
R4827 CLK1.n789 CLK1.n635 96
R4828 CLK1.n793 CLK1.n635 96
R4829 CLK1.n793 CLK1.n629 96
R4830 CLK1.n801 CLK1.n629 96
R4831 CLK1.n801 CLK1.n627 96
R4832 CLK1.n694 CLK1.n687 96
R4833 CLK1.n694 CLK1.n685 96
R4834 CLK1.n699 CLK1.n685 96
R4835 CLK1.n699 CLK1.n681 96
R4836 CLK1.n706 CLK1.n681 96
R4837 CLK1.n706 CLK1.n680 96
R4838 CLK1.n710 CLK1.n680 96
R4839 CLK1.n710 CLK1.n675 96
R4840 CLK1.n717 CLK1.n675 96
R4841 CLK1.n717 CLK1.n673 96
R4842 CLK1.n721 CLK1.n673 96
R4843 CLK1.n721 CLK1.n669 96
R4844 CLK1.n728 CLK1.n669 96
R4845 CLK1.n728 CLK1.n667 96
R4846 CLK1.n1369 CLK1.n1296 96
R4847 CLK1.n1369 CLK1.n1291 96
R4848 CLK1.n1376 CLK1.n1291 96
R4849 CLK1.n1376 CLK1.n1289 96
R4850 CLK1.n1380 CLK1.n1289 96
R4851 CLK1.n1380 CLK1.n1285 96
R4852 CLK1.n1387 CLK1.n1285 96
R4853 CLK1.n1387 CLK1.n1283 96
R4854 CLK1.n1391 CLK1.n1283 96
R4855 CLK1.n1391 CLK1.n1279 96
R4856 CLK1.n1399 CLK1.n1279 96
R4857 CLK1.n1399 CLK1.n1277 96
R4858 CLK1.n1404 CLK1.n1277 96
R4859 CLK1.n1404 CLK1.n1274 96
R4860 CLK1.n1411 CLK1.n1274 96
R4861 CLK1.n1411 CLK1.n1273 96
R4862 CLK1.n1415 CLK1.n1273 96
R4863 CLK1.n1415 CLK1.n1269 96
R4864 CLK1.n1421 CLK1.n1269 96
R4865 CLK1.n1421 CLK1.n1267 96
R4866 CLK1.n1425 CLK1.n1267 96
R4867 CLK1.n1425 CLK1.n1261 96
R4868 CLK1.n1433 CLK1.n1261 96
R4869 CLK1.n1433 CLK1.n1259 96
R4870 CLK1.n1326 CLK1.n1319 96
R4871 CLK1.n1326 CLK1.n1317 96
R4872 CLK1.n1331 CLK1.n1317 96
R4873 CLK1.n1331 CLK1.n1313 96
R4874 CLK1.n1338 CLK1.n1313 96
R4875 CLK1.n1338 CLK1.n1312 96
R4876 CLK1.n1342 CLK1.n1312 96
R4877 CLK1.n1342 CLK1.n1307 96
R4878 CLK1.n1349 CLK1.n1307 96
R4879 CLK1.n1349 CLK1.n1305 96
R4880 CLK1.n1353 CLK1.n1305 96
R4881 CLK1.n1353 CLK1.n1301 96
R4882 CLK1.n1360 CLK1.n1301 96
R4883 CLK1.n1360 CLK1.n1299 96
R4884 CLK1.n226 CLK1.n223 85.261
R4885 CLK1.n1552 CLK1.n1551 85.261
R4886 CLK1.n1506 CLK1.n1503 85.261
R4887 CLK1.n1191 CLK1.n316 85.261
R4888 CLK1.n478 CLK1.n407 85.261
R4889 CLK1.n920 CLK1.n919 85.261
R4890 CLK1.n874 CLK1.n871 85.261
R4891 CLK1.n559 CLK1.n556 85.261
R4892 CLK1.n735 CLK1.n734 85.261
R4893 CLK1.n689 CLK1.n686 85.261
R4894 CLK1.n1367 CLK1.n1366 85.261
R4895 CLK1.n1321 CLK1.n1318 85.261
R4896 CLK1.n278 CLK1.n277 85.261
R4897 CLK1.n1621 CLK1.n1620 85.261
R4898 CLK1.n1548 CLK1.n1547 85.261
R4899 CLK1.n1254 CLK1.n1253 85.261
R4900 CLK1.n346 CLK1.n343 85.261
R4901 CLK1.n388 CLK1.n387 85.261
R4902 CLK1.n434 CLK1.n431 85.261
R4903 CLK1.n476 CLK1.n475 85.261
R4904 CLK1.n998 CLK1.n997 85.261
R4905 CLK1.n989 CLK1.n988 85.261
R4906 CLK1.n916 CLK1.n915 85.261
R4907 CLK1.n622 CLK1.n621 85.261
R4908 CLK1.n804 CLK1.n803 85.261
R4909 CLK1.n731 CLK1.n730 85.261
R4910 CLK1.n1436 CLK1.n1435 85.261
R4911 CLK1.n1363 CLK1.n1362 85.261
R4912 CLK1.n1075 CLK1.n1074 69.028
R4913 CLK1.n1076 CLK1.n1075 69.028
R4914 CLK1.n1085 CLK1.n1084 69.028
R4915 CLK1.n1092 CLK1.n1087 69.028
R4916 CLK1.n1094 CLK1.n1093 69.028
R4917 CLK1.n1095 CLK1.n1094 69.028
R4918 CLK1.n1086 CLK1.t8 64.713
R4919 CLK1.t75 CLK1.n1086 64.713
R4920 CLK1.n1084 CLK1.t10 56.085
R4921 CLK1.t77 CLK1.n1092 56.085
R4922 CLK1.n239 CLK1.t88 44.338
R4923 CLK1.n261 CLK1.t139 44.338
R4924 CLK1.n1079 CLK1.t51 44.338
R4925 CLK1.n1090 CLK1.t121 44.338
R4926 CLK1.n702 CLK1.t70 44.338
R4927 CLK1.n671 CLK1.t74 44.338
R4928 CLK1.n649 CLK1.t13 44.338
R4929 CLK1.n776 CLK1.t186 44.338
R4930 CLK1.n447 CLK1.t117 44.338
R4931 CLK1.n416 CLK1.t63 44.338
R4932 CLK1.n494 CLK1.t124 44.338
R4933 CLK1.n503 CLK1.t170 44.338
R4934 CLK1.n1334 CLK1.t26 44.338
R4935 CLK1.n1303 CLK1.t19 44.338
R4936 CLK1.n1281 CLK1.t147 44.338
R4937 CLK1.n1408 CLK1.t196 44.338
R4938 CLK1.n155 CLK1.t176 44.337
R4939 CLK1.n128 CLK1.t194 44.337
R4940 CLK1.n61 CLK1.t93 44.337
R4941 CLK1.n34 CLK1.t54 44.337
R4942 CLK1.n1593 CLK1.t50 44.337
R4943 CLK1.n1466 CLK1.t108 44.337
R4944 CLK1.n1488 CLK1.t86 44.337
R4945 CLK1.n1519 CLK1.t1 44.337
R4946 CLK1.n295 CLK1.t17 44.337
R4947 CLK1.n1214 CLK1.t132 44.337
R4948 CLK1.n328 CLK1.t182 44.337
R4949 CLK1.n359 CLK1.t128 44.337
R4950 CLK1.n1079 CLK1.t11 44.337
R4951 CLK1.n1090 CLK1.t78 44.337
R4952 CLK1.n961 CLK1.t58 44.337
R4953 CLK1.n834 CLK1.t134 44.337
R4954 CLK1.n856 CLK1.t5 44.337
R4955 CLK1.n887 CLK1.t156 44.337
R4956 CLK1.n535 CLK1.t162 44.337
R4957 CLK1.n582 CLK1.t145 44.337
R4958 CLK1.n1176 CLK1.n394 39.834
R4959 CLK1.n1172 CLK1.n394 39.834
R4960 CLK1.n1172 CLK1.n396 39.834
R4961 CLK1.n1165 CLK1.n396 39.834
R4962 CLK1.n1165 CLK1.n1068 39.834
R4963 CLK1.n1161 CLK1.n1068 39.834
R4964 CLK1.n1161 CLK1.n1070 39.834
R4965 CLK1.n1155 CLK1.n1070 39.834
R4966 CLK1.n1155 CLK1.n1154 39.834
R4967 CLK1.n1154 CLK1.n1153 39.834
R4968 CLK1.n1153 CLK1.n1077 39.834
R4969 CLK1.n1147 CLK1.n1077 39.834
R4970 CLK1.n1147 CLK1.n1146 39.834
R4971 CLK1.n1146 CLK1.n1145 39.834
R4972 CLK1.n1145 CLK1.n1088 39.834
R4973 CLK1.n1139 CLK1.n1088 39.834
R4974 CLK1.n1139 CLK1.n1138 39.834
R4975 CLK1.n1138 CLK1.n1137 39.834
R4976 CLK1.n1137 CLK1.n1096 39.834
R4977 CLK1.n1131 CLK1.n1096 39.834
R4978 CLK1.n1131 CLK1.n1102 39.834
R4979 CLK1.n1127 CLK1.n1102 39.834
R4980 CLK1.n1127 CLK1.n1105 39.834
R4981 CLK1.n1120 CLK1.n1105 39.834
R4982 CLK1.n1120 CLK1.n1112 39.834
R4983 CLK1.n1116 CLK1.n1112 39.834
R4984 CLK1.n3 CLK1.t188 39.4
R4985 CLK1.n3 CLK1.t174 39.4
R4986 CLK1.n7 CLK1.t56 39.4
R4987 CLK1.n7 CLK1.t95 39.4
R4988 CLK1.n213 CLK1.t90 39.4
R4989 CLK1.n213 CLK1.t141 39.4
R4990 CLK1.n1580 CLK1.t110 39.4
R4991 CLK1.n1580 CLK1.t153 39.4
R4992 CLK1.n1494 CLK1.t3 39.4
R4993 CLK1.n1494 CLK1.t84 39.4
R4994 CLK1.n301 CLK1.t130 39.4
R4995 CLK1.n301 CLK1.t15 39.4
R4996 CLK1.n1081 CLK1.t9 39.4
R4997 CLK1.n1081 CLK1.t76 39.4
R4998 CLK1.n1080 CLK1.t52 39.4
R4999 CLK1.n1080 CLK1.t120 39.4
R5000 CLK1.n334 CLK1.t126 39.4
R5001 CLK1.n334 CLK1.t180 39.4
R5002 CLK1.n495 CLK1.t65 39.4
R5003 CLK1.n495 CLK1.t44 39.4
R5004 CLK1.n422 CLK1.t115 39.4
R5005 CLK1.n422 CLK1.t61 39.4
R5006 CLK1.n948 CLK1.t136 39.4
R5007 CLK1.n948 CLK1.t104 39.4
R5008 CLK1.n862 CLK1.t158 39.4
R5009 CLK1.n862 CLK1.t7 39.4
R5010 CLK1.n541 CLK1.t143 39.4
R5011 CLK1.n541 CLK1.t160 39.4
R5012 CLK1.n763 CLK1.t47 39.4
R5013 CLK1.n763 CLK1.t184 39.4
R5014 CLK1.n677 CLK1.t68 39.4
R5015 CLK1.n677 CLK1.t72 39.4
R5016 CLK1.n1395 CLK1.t172 39.4
R5017 CLK1.n1395 CLK1.t149 39.4
R5018 CLK1.n1309 CLK1.t28 39.4
R5019 CLK1.n1309 CLK1.t21 39.4
R5020 CLK1.n1117 CLK1.n1114 39.262
R5021 CLK1.n1175 CLK1.n392 38.088
R5022 CLK1.n227 CLK1.t113 30.776
R5023 CLK1.n86 CLK1.t177 30.775
R5024 CLK1.n282 CLK1.t81 30.775
R5025 CLK1.n522 CLK1.t41 30.775
R5026 CLK1.n560 CLK1.t66 30.775
R5027 CLK1.n690 CLK1.t31 29.713
R5028 CLK1.n665 CLK1.t197 29.713
R5029 CLK1.n435 CLK1.t40 29.713
R5030 CLK1.n410 CLK1.t36 29.713
R5031 CLK1.n1322 CLK1.t111 29.713
R5032 CLK1.n1297 CLK1.t99 29.713
R5033 CLK1.n1482 CLK1.t98 29.712
R5034 CLK1.n1507 CLK1.t164 29.712
R5035 CLK1.n322 CLK1.t122 29.712
R5036 CLK1.n347 CLK1.t22 29.712
R5037 CLK1.n850 CLK1.t168 29.712
R5038 CLK1.n875 CLK1.t101 29.712
R5039 CLK1.n129 CLK1.t193 24.568
R5040 CLK1.n151 CLK1.t175 24.568
R5041 CLK1.n35 CLK1.t53 24.568
R5042 CLK1.n57 CLK1.t92 24.568
R5043 CLK1.t87 CLK1.n244 24.568
R5044 CLK1.t138 CLK1.n205 24.568
R5045 CLK1.n1575 CLK1.t107 24.568
R5046 CLK1.n1597 CLK1.t49 24.568
R5047 CLK1.n1514 CLK1.t0 24.568
R5048 CLK1.n1536 CLK1.t85 24.568
R5049 CLK1.n1209 CLK1.t131 24.568
R5050 CLK1.n1231 CLK1.t16 24.568
R5051 CLK1.n354 CLK1.t127 24.568
R5052 CLK1.n376 CLK1.t181 24.568
R5053 CLK1.n442 CLK1.t116 24.568
R5054 CLK1.n464 CLK1.t62 24.568
R5055 CLK1.n1038 CLK1.t123 24.568
R5056 CLK1.n1020 CLK1.t169 24.568
R5057 CLK1.n943 CLK1.t133 24.568
R5058 CLK1.n965 CLK1.t57 24.568
R5059 CLK1.n882 CLK1.t155 24.568
R5060 CLK1.n904 CLK1.t4 24.568
R5061 CLK1.n577 CLK1.t144 24.568
R5062 CLK1.n599 CLK1.t161 24.568
R5063 CLK1.n758 CLK1.t12 24.568
R5064 CLK1.n780 CLK1.t185 24.568
R5065 CLK1.n697 CLK1.t69 24.568
R5066 CLK1.n719 CLK1.t73 24.568
R5067 CLK1.n1390 CLK1.t146 24.568
R5068 CLK1.n1412 CLK1.t195 24.568
R5069 CLK1.n1329 CLK1.t25 24.568
R5070 CLK1.n1351 CLK1.t18 24.568
R5071 CLK1.n0 CLK1.t80 24
R5072 CLK1.n0 CLK1.t154 24
R5073 CLK1.n4 CLK1.t137 24
R5074 CLK1.n4 CLK1.t79 24
R5075 CLK1.n8 CLK1.t33 24
R5076 CLK1.n8 CLK1.t102 24
R5077 CLK1.n201 CLK1.t150 24
R5078 CLK1.n201 CLK1.t32 24
R5079 CLK1.n1449 CLK1.t119 24
R5080 CLK1.n1449 CLK1.t23 24
R5081 CLK1.n1478 CLK1.t59 24
R5082 CLK1.n1478 CLK1.t192 24
R5083 CLK1.n288 CLK1.t167 24
R5084 CLK1.n288 CLK1.t178 24
R5085 CLK1.n1182 CLK1.t198 24
R5086 CLK1.n1099 CLK1.t163 24
R5087 CLK1.n1099 CLK1.t190 24
R5088 CLK1.n1109 CLK1.t24 24
R5089 CLK1.n1109 CLK1.t45 24
R5090 CLK1.n1108 CLK1.t38 24
R5091 CLK1.n1108 CLK1.t189 24
R5092 CLK1.n1057 CLK1.t96 24
R5093 CLK1.n1057 CLK1.t165 24
R5094 CLK1.n817 CLK1.t34 24
R5095 CLK1.n817 CLK1.t39 24
R5096 CLK1.n846 CLK1.t91 24
R5097 CLK1.n846 CLK1.t35 24
R5098 CLK1.n528 CLK1.t191 24
R5099 CLK1.n528 CLK1.t42 24
R5100 CLK1.n661 CLK1.t151 24
R5101 CLK1.n661 CLK1.t82 24
R5102 CLK1.n632 CLK1.t112 24
R5103 CLK1.n632 CLK1.t118 24
R5104 CLK1.n516 CLK1.t166 24
R5105 CLK1.n516 CLK1.t97 24
R5106 CLK1.n1061 CLK1.t48 24
R5107 CLK1.n1061 CLK1.t37 24
R5108 CLK1.n1186 CLK1.t100 24
R5109 CLK1.n1293 CLK1.t105 24
R5110 CLK1.n1293 CLK1.t29 24
R5111 CLK1.n1264 CLK1.t30 24
R5112 CLK1.n1264 CLK1.t106 24
R5113 CLK1.t10 CLK1.n1076 12.942
R5114 CLK1.n1093 CLK1.t77 12.942
R5115 CLK1.n145 CLK1.n142 12.8
R5116 CLK1.n51 CLK1.n48 12.8
R5117 CLK1.n226 CLK1.n225 12.8
R5118 CLK1.n230 CLK1.n225 12.8
R5119 CLK1.n230 CLK1.n221 12.8
R5120 CLK1.n236 CLK1.n221 12.8
R5121 CLK1.n236 CLK1.n219 12.8
R5122 CLK1.n241 CLK1.n219 12.8
R5123 CLK1.n241 CLK1.n215 12.8
R5124 CLK1.n248 CLK1.n215 12.8
R5125 CLK1.n248 CLK1.n212 12.8
R5126 CLK1.n252 CLK1.n212 12.8
R5127 CLK1.n252 CLK1.n209 12.8
R5128 CLK1.n258 CLK1.n209 12.8
R5129 CLK1.n258 CLK1.n207 12.8
R5130 CLK1.n263 CLK1.n207 12.8
R5131 CLK1.n263 CLK1.n203 12.8
R5132 CLK1.n269 CLK1.n203 12.8
R5133 CLK1.n269 CLK1.n200 12.8
R5134 CLK1.n274 CLK1.n200 12.8
R5135 CLK1.n274 CLK1.n196 12.8
R5136 CLK1.n278 CLK1.n196 12.8
R5137 CLK1.n1551 CLK1.n1480 12.8
R5138 CLK1.n1555 CLK1.n1480 12.8
R5139 CLK1.n1555 CLK1.n1477 12.8
R5140 CLK1.n1560 CLK1.n1477 12.8
R5141 CLK1.n1560 CLK1.n1473 12.8
R5142 CLK1.n1566 CLK1.n1473 12.8
R5143 CLK1.n1566 CLK1.n1471 12.8
R5144 CLK1.n1571 CLK1.n1471 12.8
R5145 CLK1.n1571 CLK1.n1467 12.8
R5146 CLK1.n1577 CLK1.n1467 12.8
R5147 CLK1.n1577 CLK1.n1465 12.8
R5148 CLK1.n1583 CLK1.n1465 12.8
R5149 CLK1.n1583 CLK1.n1461 12.8
R5150 CLK1.n1590 CLK1.n1461 12.8
R5151 CLK1.n1590 CLK1.n1460 12.8
R5152 CLK1.n1595 CLK1.n1460 12.8
R5153 CLK1.n1595 CLK1.n1457 12.8
R5154 CLK1.n1601 CLK1.n1457 12.8
R5155 CLK1.n1601 CLK1.n1455 12.8
R5156 CLK1.n1605 CLK1.n1455 12.8
R5157 CLK1.n1605 CLK1.n1451 12.8
R5158 CLK1.n1611 CLK1.n1451 12.8
R5159 CLK1.n1611 CLK1.n1447 12.8
R5160 CLK1.n1617 CLK1.n1447 12.8
R5161 CLK1.n1617 CLK1.n1448 12.8
R5162 CLK1.n1506 CLK1.n1505 12.8
R5163 CLK1.n1510 CLK1.n1505 12.8
R5164 CLK1.n1510 CLK1.n1501 12.8
R5165 CLK1.n1517 CLK1.n1501 12.8
R5166 CLK1.n1517 CLK1.n1499 12.8
R5167 CLK1.n1522 CLK1.n1499 12.8
R5168 CLK1.n1522 CLK1.n1496 12.8
R5169 CLK1.n1528 CLK1.n1496 12.8
R5170 CLK1.n1528 CLK1.n1493 12.8
R5171 CLK1.n1533 CLK1.n1493 12.8
R5172 CLK1.n1533 CLK1.n1489 12.8
R5173 CLK1.n1539 CLK1.n1489 12.8
R5174 CLK1.n1539 CLK1.n1487 12.8
R5175 CLK1.n1544 CLK1.n1487 12.8
R5176 CLK1.n1544 CLK1.n1483 12.8
R5177 CLK1.n1548 CLK1.n1483 12.8
R5178 CLK1.n1191 CLK1.n318 12.8
R5179 CLK1.n1195 CLK1.n318 12.8
R5180 CLK1.n1195 CLK1.n314 12.8
R5181 CLK1.n1201 CLK1.n314 12.8
R5182 CLK1.n1201 CLK1.n312 12.8
R5183 CLK1.n1205 CLK1.n312 12.8
R5184 CLK1.n1205 CLK1.n308 12.8
R5185 CLK1.n1212 CLK1.n308 12.8
R5186 CLK1.n1212 CLK1.n306 12.8
R5187 CLK1.n1217 CLK1.n306 12.8
R5188 CLK1.n1217 CLK1.n303 12.8
R5189 CLK1.n1223 CLK1.n303 12.8
R5190 CLK1.n1223 CLK1.n300 12.8
R5191 CLK1.n1228 CLK1.n300 12.8
R5192 CLK1.n1228 CLK1.n296 12.8
R5193 CLK1.n1234 CLK1.n296 12.8
R5194 CLK1.n1234 CLK1.n294 12.8
R5195 CLK1.n1239 CLK1.n294 12.8
R5196 CLK1.n1239 CLK1.n290 12.8
R5197 CLK1.n1245 CLK1.n290 12.8
R5198 CLK1.n1245 CLK1.n287 12.8
R5199 CLK1.n1250 CLK1.n287 12.8
R5200 CLK1.n1250 CLK1.n283 12.8
R5201 CLK1.n1254 CLK1.n283 12.8
R5202 CLK1.n1181 CLK1.n321 12.8
R5203 CLK1.n346 CLK1.n345 12.8
R5204 CLK1.n350 CLK1.n345 12.8
R5205 CLK1.n350 CLK1.n341 12.8
R5206 CLK1.n357 CLK1.n341 12.8
R5207 CLK1.n357 CLK1.n339 12.8
R5208 CLK1.n362 CLK1.n339 12.8
R5209 CLK1.n362 CLK1.n336 12.8
R5210 CLK1.n368 CLK1.n336 12.8
R5211 CLK1.n368 CLK1.n333 12.8
R5212 CLK1.n373 CLK1.n333 12.8
R5213 CLK1.n373 CLK1.n329 12.8
R5214 CLK1.n379 CLK1.n329 12.8
R5215 CLK1.n379 CLK1.n327 12.8
R5216 CLK1.n384 CLK1.n327 12.8
R5217 CLK1.n384 CLK1.n323 12.8
R5218 CLK1.n388 CLK1.n323 12.8
R5219 CLK1.n1058 CLK1.n400 12.8
R5220 CLK1.n434 CLK1.n433 12.8
R5221 CLK1.n438 CLK1.n433 12.8
R5222 CLK1.n438 CLK1.n429 12.8
R5223 CLK1.n445 CLK1.n429 12.8
R5224 CLK1.n445 CLK1.n427 12.8
R5225 CLK1.n450 CLK1.n427 12.8
R5226 CLK1.n450 CLK1.n424 12.8
R5227 CLK1.n456 CLK1.n424 12.8
R5228 CLK1.n456 CLK1.n421 12.8
R5229 CLK1.n461 CLK1.n421 12.8
R5230 CLK1.n461 CLK1.n417 12.8
R5231 CLK1.n467 CLK1.n417 12.8
R5232 CLK1.n467 CLK1.n415 12.8
R5233 CLK1.n472 CLK1.n415 12.8
R5234 CLK1.n472 CLK1.n411 12.8
R5235 CLK1.n476 CLK1.n411 12.8
R5236 CLK1.n478 CLK1.n409 12.8
R5237 CLK1.n482 CLK1.n409 12.8
R5238 CLK1.n482 CLK1.n403 12.8
R5239 CLK1.n1052 CLK1.n403 12.8
R5240 CLK1.n1052 CLK1.n404 12.8
R5241 CLK1.n1046 CLK1.n404 12.8
R5242 CLK1.n1046 CLK1.n488 12.8
R5243 CLK1.n1042 CLK1.n488 12.8
R5244 CLK1.n1042 CLK1.n490 12.8
R5245 CLK1.n1036 CLK1.n490 12.8
R5246 CLK1.n1036 CLK1.n493 12.8
R5247 CLK1.n1032 CLK1.n493 12.8
R5248 CLK1.n1032 CLK1.n497 12.8
R5249 CLK1.n1026 CLK1.n497 12.8
R5250 CLK1.n1026 CLK1.n502 12.8
R5251 CLK1.n1022 CLK1.n502 12.8
R5252 CLK1.n1022 CLK1.n504 12.8
R5253 CLK1.n1016 CLK1.n504 12.8
R5254 CLK1.n1016 CLK1.n508 12.8
R5255 CLK1.n1012 CLK1.n508 12.8
R5256 CLK1.n1012 CLK1.n511 12.8
R5257 CLK1.n1006 CLK1.n511 12.8
R5258 CLK1.n1006 CLK1.n515 12.8
R5259 CLK1.n1001 CLK1.n515 12.8
R5260 CLK1.n1001 CLK1.n518 12.8
R5261 CLK1.n997 CLK1.n518 12.8
R5262 CLK1.n919 CLK1.n848 12.8
R5263 CLK1.n923 CLK1.n848 12.8
R5264 CLK1.n923 CLK1.n845 12.8
R5265 CLK1.n928 CLK1.n845 12.8
R5266 CLK1.n928 CLK1.n841 12.8
R5267 CLK1.n934 CLK1.n841 12.8
R5268 CLK1.n934 CLK1.n839 12.8
R5269 CLK1.n939 CLK1.n839 12.8
R5270 CLK1.n939 CLK1.n835 12.8
R5271 CLK1.n945 CLK1.n835 12.8
R5272 CLK1.n945 CLK1.n833 12.8
R5273 CLK1.n951 CLK1.n833 12.8
R5274 CLK1.n951 CLK1.n829 12.8
R5275 CLK1.n958 CLK1.n829 12.8
R5276 CLK1.n958 CLK1.n828 12.8
R5277 CLK1.n963 CLK1.n828 12.8
R5278 CLK1.n963 CLK1.n825 12.8
R5279 CLK1.n969 CLK1.n825 12.8
R5280 CLK1.n969 CLK1.n823 12.8
R5281 CLK1.n973 CLK1.n823 12.8
R5282 CLK1.n973 CLK1.n819 12.8
R5283 CLK1.n979 CLK1.n819 12.8
R5284 CLK1.n979 CLK1.n815 12.8
R5285 CLK1.n985 CLK1.n815 12.8
R5286 CLK1.n985 CLK1.n816 12.8
R5287 CLK1.n874 CLK1.n873 12.8
R5288 CLK1.n878 CLK1.n873 12.8
R5289 CLK1.n878 CLK1.n869 12.8
R5290 CLK1.n885 CLK1.n869 12.8
R5291 CLK1.n885 CLK1.n867 12.8
R5292 CLK1.n890 CLK1.n867 12.8
R5293 CLK1.n890 CLK1.n864 12.8
R5294 CLK1.n896 CLK1.n864 12.8
R5295 CLK1.n896 CLK1.n861 12.8
R5296 CLK1.n901 CLK1.n861 12.8
R5297 CLK1.n901 CLK1.n857 12.8
R5298 CLK1.n907 CLK1.n857 12.8
R5299 CLK1.n907 CLK1.n855 12.8
R5300 CLK1.n912 CLK1.n855 12.8
R5301 CLK1.n912 CLK1.n851 12.8
R5302 CLK1.n916 CLK1.n851 12.8
R5303 CLK1.n559 CLK1.n558 12.8
R5304 CLK1.n563 CLK1.n558 12.8
R5305 CLK1.n563 CLK1.n554 12.8
R5306 CLK1.n569 CLK1.n554 12.8
R5307 CLK1.n569 CLK1.n552 12.8
R5308 CLK1.n573 CLK1.n552 12.8
R5309 CLK1.n573 CLK1.n548 12.8
R5310 CLK1.n580 CLK1.n548 12.8
R5311 CLK1.n580 CLK1.n546 12.8
R5312 CLK1.n585 CLK1.n546 12.8
R5313 CLK1.n585 CLK1.n543 12.8
R5314 CLK1.n591 CLK1.n543 12.8
R5315 CLK1.n591 CLK1.n540 12.8
R5316 CLK1.n596 CLK1.n540 12.8
R5317 CLK1.n596 CLK1.n536 12.8
R5318 CLK1.n602 CLK1.n536 12.8
R5319 CLK1.n602 CLK1.n534 12.8
R5320 CLK1.n607 CLK1.n534 12.8
R5321 CLK1.n607 CLK1.n530 12.8
R5322 CLK1.n613 CLK1.n530 12.8
R5323 CLK1.n613 CLK1.n527 12.8
R5324 CLK1.n618 CLK1.n527 12.8
R5325 CLK1.n618 CLK1.n523 12.8
R5326 CLK1.n622 CLK1.n523 12.8
R5327 CLK1.n734 CLK1.n663 12.8
R5328 CLK1.n738 CLK1.n663 12.8
R5329 CLK1.n738 CLK1.n660 12.8
R5330 CLK1.n743 CLK1.n660 12.8
R5331 CLK1.n743 CLK1.n656 12.8
R5332 CLK1.n749 CLK1.n656 12.8
R5333 CLK1.n749 CLK1.n654 12.8
R5334 CLK1.n754 CLK1.n654 12.8
R5335 CLK1.n754 CLK1.n650 12.8
R5336 CLK1.n760 CLK1.n650 12.8
R5337 CLK1.n760 CLK1.n648 12.8
R5338 CLK1.n766 CLK1.n648 12.8
R5339 CLK1.n766 CLK1.n644 12.8
R5340 CLK1.n773 CLK1.n644 12.8
R5341 CLK1.n773 CLK1.n643 12.8
R5342 CLK1.n778 CLK1.n643 12.8
R5343 CLK1.n778 CLK1.n640 12.8
R5344 CLK1.n784 CLK1.n640 12.8
R5345 CLK1.n784 CLK1.n638 12.8
R5346 CLK1.n788 CLK1.n638 12.8
R5347 CLK1.n788 CLK1.n634 12.8
R5348 CLK1.n794 CLK1.n634 12.8
R5349 CLK1.n794 CLK1.n630 12.8
R5350 CLK1.n800 CLK1.n630 12.8
R5351 CLK1.n800 CLK1.n631 12.8
R5352 CLK1.n689 CLK1.n688 12.8
R5353 CLK1.n693 CLK1.n688 12.8
R5354 CLK1.n693 CLK1.n684 12.8
R5355 CLK1.n700 CLK1.n684 12.8
R5356 CLK1.n700 CLK1.n682 12.8
R5357 CLK1.n705 CLK1.n682 12.8
R5358 CLK1.n705 CLK1.n679 12.8
R5359 CLK1.n711 CLK1.n679 12.8
R5360 CLK1.n711 CLK1.n676 12.8
R5361 CLK1.n716 CLK1.n676 12.8
R5362 CLK1.n716 CLK1.n672 12.8
R5363 CLK1.n722 CLK1.n672 12.8
R5364 CLK1.n722 CLK1.n670 12.8
R5365 CLK1.n727 CLK1.n670 12.8
R5366 CLK1.n727 CLK1.n666 12.8
R5367 CLK1.n731 CLK1.n666 12.8
R5368 CLK1.n1063 CLK1.n398 12.8
R5369 CLK1.n1188 CLK1.n1187 12.8
R5370 CLK1.n1366 CLK1.n1295 12.8
R5371 CLK1.n1370 CLK1.n1295 12.8
R5372 CLK1.n1370 CLK1.n1292 12.8
R5373 CLK1.n1375 CLK1.n1292 12.8
R5374 CLK1.n1375 CLK1.n1288 12.8
R5375 CLK1.n1381 CLK1.n1288 12.8
R5376 CLK1.n1381 CLK1.n1286 12.8
R5377 CLK1.n1386 CLK1.n1286 12.8
R5378 CLK1.n1386 CLK1.n1282 12.8
R5379 CLK1.n1392 CLK1.n1282 12.8
R5380 CLK1.n1392 CLK1.n1280 12.8
R5381 CLK1.n1398 CLK1.n1280 12.8
R5382 CLK1.n1398 CLK1.n1276 12.8
R5383 CLK1.n1405 CLK1.n1276 12.8
R5384 CLK1.n1405 CLK1.n1275 12.8
R5385 CLK1.n1410 CLK1.n1275 12.8
R5386 CLK1.n1410 CLK1.n1272 12.8
R5387 CLK1.n1416 CLK1.n1272 12.8
R5388 CLK1.n1416 CLK1.n1270 12.8
R5389 CLK1.n1420 CLK1.n1270 12.8
R5390 CLK1.n1420 CLK1.n1266 12.8
R5391 CLK1.n1426 CLK1.n1266 12.8
R5392 CLK1.n1426 CLK1.n1262 12.8
R5393 CLK1.n1432 CLK1.n1262 12.8
R5394 CLK1.n1432 CLK1.n1263 12.8
R5395 CLK1.n1321 CLK1.n1320 12.8
R5396 CLK1.n1325 CLK1.n1320 12.8
R5397 CLK1.n1325 CLK1.n1316 12.8
R5398 CLK1.n1332 CLK1.n1316 12.8
R5399 CLK1.n1332 CLK1.n1314 12.8
R5400 CLK1.n1337 CLK1.n1314 12.8
R5401 CLK1.n1337 CLK1.n1311 12.8
R5402 CLK1.n1343 CLK1.n1311 12.8
R5403 CLK1.n1343 CLK1.n1308 12.8
R5404 CLK1.n1348 CLK1.n1308 12.8
R5405 CLK1.n1348 CLK1.n1304 12.8
R5406 CLK1.n1354 CLK1.n1304 12.8
R5407 CLK1.n1354 CLK1.n1302 12.8
R5408 CLK1.n1359 CLK1.n1302 12.8
R5409 CLK1.n1359 CLK1.n1298 12.8
R5410 CLK1.n1363 CLK1.n1298 12.8
R5411 CLK1.n1448 CLK1.n1443 11.36
R5412 CLK1.n816 CLK1.n811 11.36
R5413 CLK1.n631 CLK1.n626 11.36
R5414 CLK1.n1263 CLK1.n1258 11.36
R5415 CLK1.n1443 CLK1.n1442 9.3
R5416 CLK1.n811 CLK1.n810 9.3
R5417 CLK1.n626 CLK1.n625 9.3
R5418 CLK1.n1258 CLK1.n1257 9.3
R5419 CLK1.n11 CLK1.n10 8.855
R5420 CLK1.n15 CLK1.n14 8.855
R5421 CLK1.n14 CLK1.n13 8.855
R5422 CLK1.n20 CLK1.n19 8.855
R5423 CLK1.n19 CLK1.n18 8.855
R5424 CLK1.n24 CLK1.n23 8.855
R5425 CLK1.n23 CLK1.n22 8.855
R5426 CLK1.n28 CLK1.n27 8.855
R5427 CLK1.n27 CLK1.n26 8.855
R5428 CLK1.n32 CLK1.n31 8.855
R5429 CLK1.n31 CLK1.n30 8.855
R5430 CLK1.n37 CLK1.n36 8.855
R5431 CLK1.n36 CLK1.n35 8.855
R5432 CLK1.n41 CLK1.n40 8.855
R5433 CLK1.n40 CLK1.n39 8.855
R5434 CLK1.n45 CLK1.n44 8.855
R5435 CLK1.n44 CLK1.n43 8.855
R5436 CLK1.n48 CLK1.n6 8.855
R5437 CLK1.n6 CLK1.n5 8.855
R5438 CLK1.n51 CLK1.n50 8.855
R5439 CLK1.n50 CLK1.n49 8.855
R5440 CLK1.n55 CLK1.n54 8.855
R5441 CLK1.n54 CLK1.n53 8.855
R5442 CLK1.n59 CLK1.n58 8.855
R5443 CLK1.n58 CLK1.n57 8.855
R5444 CLK1.n64 CLK1.n63 8.855
R5445 CLK1.n63 CLK1.n62 8.855
R5446 CLK1.n68 CLK1.n67 8.855
R5447 CLK1.n67 CLK1.n66 8.855
R5448 CLK1.n72 CLK1.n71 8.855
R5449 CLK1.n71 CLK1.n70 8.855
R5450 CLK1.n76 CLK1.n75 8.855
R5451 CLK1.n75 CLK1.n74 8.855
R5452 CLK1.n80 CLK1.n79 8.855
R5453 CLK1.n79 CLK1.n78 8.855
R5454 CLK1.n84 CLK1.n83 8.855
R5455 CLK1.n93 CLK1.n92 8.855
R5456 CLK1.n97 CLK1.n96 8.855
R5457 CLK1.n96 CLK1.n95 8.855
R5458 CLK1.n101 CLK1.n100 8.855
R5459 CLK1.n100 CLK1.n99 8.855
R5460 CLK1.n106 CLK1.n105 8.855
R5461 CLK1.n105 CLK1.n104 8.855
R5462 CLK1.n110 CLK1.n109 8.855
R5463 CLK1.n109 CLK1.n108 8.855
R5464 CLK1.n114 CLK1.n113 8.855
R5465 CLK1.n113 CLK1.n112 8.855
R5466 CLK1.n118 CLK1.n117 8.855
R5467 CLK1.n117 CLK1.n116 8.855
R5468 CLK1.n122 CLK1.n121 8.855
R5469 CLK1.n121 CLK1.n120 8.855
R5470 CLK1.n126 CLK1.n125 8.855
R5471 CLK1.n125 CLK1.n124 8.855
R5472 CLK1.n131 CLK1.n130 8.855
R5473 CLK1.n130 CLK1.n129 8.855
R5474 CLK1.n135 CLK1.n134 8.855
R5475 CLK1.n134 CLK1.n133 8.855
R5476 CLK1.n139 CLK1.n138 8.855
R5477 CLK1.n138 CLK1.n137 8.855
R5478 CLK1.n142 CLK1.n2 8.855
R5479 CLK1.n2 CLK1.n1 8.855
R5480 CLK1.n145 CLK1.n144 8.855
R5481 CLK1.n144 CLK1.n143 8.855
R5482 CLK1.n149 CLK1.n148 8.855
R5483 CLK1.n148 CLK1.n147 8.855
R5484 CLK1.n153 CLK1.n152 8.855
R5485 CLK1.n152 CLK1.n151 8.855
R5486 CLK1.n158 CLK1.n157 8.855
R5487 CLK1.n157 CLK1.n156 8.855
R5488 CLK1.n162 CLK1.n161 8.855
R5489 CLK1.n161 CLK1.n160 8.855
R5490 CLK1.n166 CLK1.n165 8.855
R5491 CLK1.n165 CLK1.n164 8.855
R5492 CLK1.n170 CLK1.n169 8.855
R5493 CLK1.n169 CLK1.n168 8.855
R5494 CLK1.n174 CLK1.n173 8.855
R5495 CLK1.n173 CLK1.n172 8.855
R5496 CLK1.n178 CLK1.n177 8.855
R5497 CLK1.n177 CLK1.n176 8.855
R5498 CLK1.n183 CLK1.n182 8.855
R5499 CLK1.n182 CLK1.n181 8.855
R5500 CLK1.n187 CLK1.n186 8.855
R5501 CLK1.n186 CLK1.n185 8.855
R5502 CLK1.n191 CLK1.n190 8.855
R5503 CLK1.n225 CLK1.n224 8.855
R5504 CLK1.n231 CLK1.n230 8.855
R5505 CLK1.n232 CLK1.n231 8.855
R5506 CLK1.n222 CLK1.n221 8.855
R5507 CLK1.n233 CLK1.n222 8.855
R5508 CLK1.n236 CLK1.n235 8.855
R5509 CLK1.n235 CLK1.n234 8.855
R5510 CLK1.n219 CLK1.n218 8.855
R5511 CLK1.n218 CLK1.n217 8.855
R5512 CLK1.n242 CLK1.n241 8.855
R5513 CLK1.n243 CLK1.n242 8.855
R5514 CLK1.n216 CLK1.n215 8.855
R5515 CLK1.n244 CLK1.n216 8.855
R5516 CLK1.n248 CLK1.n247 8.855
R5517 CLK1.n247 CLK1.n246 8.855
R5518 CLK1.n212 CLK1.n211 8.855
R5519 CLK1.n245 CLK1.n211 8.855
R5520 CLK1.n253 CLK1.n252 8.855
R5521 CLK1.n254 CLK1.n253 8.855
R5522 CLK1.n210 CLK1.n209 8.855
R5523 CLK1.n255 CLK1.n210 8.855
R5524 CLK1.n258 CLK1.n257 8.855
R5525 CLK1.n257 CLK1.n256 8.855
R5526 CLK1.n207 CLK1.n206 8.855
R5527 CLK1.n206 CLK1.n205 8.855
R5528 CLK1.n264 CLK1.n263 8.855
R5529 CLK1.n265 CLK1.n264 8.855
R5530 CLK1.n204 CLK1.n203 8.855
R5531 CLK1.n266 CLK1.n204 8.855
R5532 CLK1.n269 CLK1.n268 8.855
R5533 CLK1.n268 CLK1.n267 8.855
R5534 CLK1.n200 CLK1.n199 8.855
R5535 CLK1.n199 CLK1.n198 8.855
R5536 CLK1.n275 CLK1.n274 8.855
R5537 CLK1.n276 CLK1.n275 8.855
R5538 CLK1.n197 CLK1.n196 8.855
R5539 CLK1.n1505 CLK1.n1504 8.855
R5540 CLK1.n1511 CLK1.n1510 8.855
R5541 CLK1.n1512 CLK1.n1511 8.855
R5542 CLK1.n1502 CLK1.n1501 8.855
R5543 CLK1.n1513 CLK1.n1502 8.855
R5544 CLK1.n1517 CLK1.n1516 8.855
R5545 CLK1.n1516 CLK1.n1515 8.855
R5546 CLK1.n1499 CLK1.n1498 8.855
R5547 CLK1.n1514 CLK1.n1498 8.855
R5548 CLK1.n1523 CLK1.n1522 8.855
R5549 CLK1.n1524 CLK1.n1523 8.855
R5550 CLK1.n1497 CLK1.n1496 8.855
R5551 CLK1.n1525 CLK1.n1497 8.855
R5552 CLK1.n1528 CLK1.n1527 8.855
R5553 CLK1.n1527 CLK1.n1526 8.855
R5554 CLK1.n1493 CLK1.n1492 8.855
R5555 CLK1.n1492 CLK1.n1491 8.855
R5556 CLK1.n1534 CLK1.n1533 8.855
R5557 CLK1.n1535 CLK1.n1534 8.855
R5558 CLK1.n1490 CLK1.n1489 8.855
R5559 CLK1.n1536 CLK1.n1490 8.855
R5560 CLK1.n1539 CLK1.n1538 8.855
R5561 CLK1.n1538 CLK1.n1537 8.855
R5562 CLK1.n1487 CLK1.n1486 8.855
R5563 CLK1.n1486 CLK1.n1485 8.855
R5564 CLK1.n1545 CLK1.n1544 8.855
R5565 CLK1.n1546 CLK1.n1545 8.855
R5566 CLK1.n1484 CLK1.n1483 8.855
R5567 CLK1.n1481 CLK1.n1480 8.855
R5568 CLK1.n1555 CLK1.n1554 8.855
R5569 CLK1.n1554 CLK1.n1553 8.855
R5570 CLK1.n1477 CLK1.n1476 8.855
R5571 CLK1.n1476 CLK1.n1475 8.855
R5572 CLK1.n1561 CLK1.n1560 8.855
R5573 CLK1.n1562 CLK1.n1561 8.855
R5574 CLK1.n1474 CLK1.n1473 8.855
R5575 CLK1.n1563 CLK1.n1474 8.855
R5576 CLK1.n1566 CLK1.n1565 8.855
R5577 CLK1.n1565 CLK1.n1564 8.855
R5578 CLK1.n1471 CLK1.n1470 8.855
R5579 CLK1.n1470 CLK1.n1469 8.855
R5580 CLK1.n1572 CLK1.n1571 8.855
R5581 CLK1.n1573 CLK1.n1572 8.855
R5582 CLK1.n1468 CLK1.n1467 8.855
R5583 CLK1.n1574 CLK1.n1468 8.855
R5584 CLK1.n1577 CLK1.n1576 8.855
R5585 CLK1.n1576 CLK1.n1575 8.855
R5586 CLK1.n1465 CLK1.n1464 8.855
R5587 CLK1.n1464 CLK1.n1463 8.855
R5588 CLK1.n1584 CLK1.n1583 8.855
R5589 CLK1.n1585 CLK1.n1584 8.855
R5590 CLK1.n1462 CLK1.n1461 8.855
R5591 CLK1.n1586 CLK1.n1462 8.855
R5592 CLK1.n1590 CLK1.n1589 8.855
R5593 CLK1.n1589 CLK1.n1588 8.855
R5594 CLK1.n1460 CLK1.n1459 8.855
R5595 CLK1.n1587 CLK1.n1459 8.855
R5596 CLK1.n1596 CLK1.n1595 8.855
R5597 CLK1.n1597 CLK1.n1596 8.855
R5598 CLK1.n1458 CLK1.n1457 8.855
R5599 CLK1.n1598 CLK1.n1458 8.855
R5600 CLK1.n1601 CLK1.n1600 8.855
R5601 CLK1.n1600 CLK1.n1599 8.855
R5602 CLK1.n1455 CLK1.n1454 8.855
R5603 CLK1.n1454 CLK1.n1453 8.855
R5604 CLK1.n1606 CLK1.n1605 8.855
R5605 CLK1.n1607 CLK1.n1606 8.855
R5606 CLK1.n1452 CLK1.n1451 8.855
R5607 CLK1.n1608 CLK1.n1452 8.855
R5608 CLK1.n1611 CLK1.n1610 8.855
R5609 CLK1.n1610 CLK1.n1609 8.855
R5610 CLK1.n1447 CLK1.n1446 8.855
R5611 CLK1.n1446 CLK1.n1445 8.855
R5612 CLK1.n1618 CLK1.n1617 8.855
R5613 CLK1.n1619 CLK1.n1618 8.855
R5614 CLK1.n1448 CLK1.n1444 8.855
R5615 CLK1.n1182 CLK1.n1181 8.855
R5616 CLK1.n345 CLK1.n344 8.855
R5617 CLK1.n351 CLK1.n350 8.855
R5618 CLK1.n352 CLK1.n351 8.855
R5619 CLK1.n342 CLK1.n341 8.855
R5620 CLK1.n353 CLK1.n342 8.855
R5621 CLK1.n357 CLK1.n356 8.855
R5622 CLK1.n356 CLK1.n355 8.855
R5623 CLK1.n339 CLK1.n338 8.855
R5624 CLK1.n354 CLK1.n338 8.855
R5625 CLK1.n363 CLK1.n362 8.855
R5626 CLK1.n364 CLK1.n363 8.855
R5627 CLK1.n337 CLK1.n336 8.855
R5628 CLK1.n365 CLK1.n337 8.855
R5629 CLK1.n368 CLK1.n367 8.855
R5630 CLK1.n367 CLK1.n366 8.855
R5631 CLK1.n333 CLK1.n332 8.855
R5632 CLK1.n332 CLK1.n331 8.855
R5633 CLK1.n374 CLK1.n373 8.855
R5634 CLK1.n375 CLK1.n374 8.855
R5635 CLK1.n330 CLK1.n329 8.855
R5636 CLK1.n376 CLK1.n330 8.855
R5637 CLK1.n379 CLK1.n378 8.855
R5638 CLK1.n378 CLK1.n377 8.855
R5639 CLK1.n327 CLK1.n326 8.855
R5640 CLK1.n326 CLK1.n325 8.855
R5641 CLK1.n385 CLK1.n384 8.855
R5642 CLK1.n386 CLK1.n385 8.855
R5643 CLK1.n324 CLK1.n323 8.855
R5644 CLK1.n1058 CLK1.n1057 8.855
R5645 CLK1.n433 CLK1.n432 8.855
R5646 CLK1.n519 CLK1.n518 8.855
R5647 CLK1.n873 CLK1.n872 8.855
R5648 CLK1.n879 CLK1.n878 8.855
R5649 CLK1.n880 CLK1.n879 8.855
R5650 CLK1.n870 CLK1.n869 8.855
R5651 CLK1.n881 CLK1.n870 8.855
R5652 CLK1.n885 CLK1.n884 8.855
R5653 CLK1.n884 CLK1.n883 8.855
R5654 CLK1.n867 CLK1.n866 8.855
R5655 CLK1.n882 CLK1.n866 8.855
R5656 CLK1.n891 CLK1.n890 8.855
R5657 CLK1.n892 CLK1.n891 8.855
R5658 CLK1.n865 CLK1.n864 8.855
R5659 CLK1.n893 CLK1.n865 8.855
R5660 CLK1.n896 CLK1.n895 8.855
R5661 CLK1.n895 CLK1.n894 8.855
R5662 CLK1.n861 CLK1.n860 8.855
R5663 CLK1.n860 CLK1.n859 8.855
R5664 CLK1.n902 CLK1.n901 8.855
R5665 CLK1.n903 CLK1.n902 8.855
R5666 CLK1.n858 CLK1.n857 8.855
R5667 CLK1.n904 CLK1.n858 8.855
R5668 CLK1.n907 CLK1.n906 8.855
R5669 CLK1.n906 CLK1.n905 8.855
R5670 CLK1.n855 CLK1.n854 8.855
R5671 CLK1.n854 CLK1.n853 8.855
R5672 CLK1.n913 CLK1.n912 8.855
R5673 CLK1.n914 CLK1.n913 8.855
R5674 CLK1.n852 CLK1.n851 8.855
R5675 CLK1.n849 CLK1.n848 8.855
R5676 CLK1.n923 CLK1.n922 8.855
R5677 CLK1.n922 CLK1.n921 8.855
R5678 CLK1.n845 CLK1.n844 8.855
R5679 CLK1.n844 CLK1.n843 8.855
R5680 CLK1.n929 CLK1.n928 8.855
R5681 CLK1.n930 CLK1.n929 8.855
R5682 CLK1.n842 CLK1.n841 8.855
R5683 CLK1.n931 CLK1.n842 8.855
R5684 CLK1.n934 CLK1.n933 8.855
R5685 CLK1.n933 CLK1.n932 8.855
R5686 CLK1.n839 CLK1.n838 8.855
R5687 CLK1.n838 CLK1.n837 8.855
R5688 CLK1.n940 CLK1.n939 8.855
R5689 CLK1.n941 CLK1.n940 8.855
R5690 CLK1.n836 CLK1.n835 8.855
R5691 CLK1.n942 CLK1.n836 8.855
R5692 CLK1.n945 CLK1.n944 8.855
R5693 CLK1.n944 CLK1.n943 8.855
R5694 CLK1.n833 CLK1.n832 8.855
R5695 CLK1.n832 CLK1.n831 8.855
R5696 CLK1.n952 CLK1.n951 8.855
R5697 CLK1.n953 CLK1.n952 8.855
R5698 CLK1.n830 CLK1.n829 8.855
R5699 CLK1.n954 CLK1.n830 8.855
R5700 CLK1.n958 CLK1.n957 8.855
R5701 CLK1.n957 CLK1.n956 8.855
R5702 CLK1.n828 CLK1.n827 8.855
R5703 CLK1.n955 CLK1.n827 8.855
R5704 CLK1.n964 CLK1.n963 8.855
R5705 CLK1.n965 CLK1.n964 8.855
R5706 CLK1.n826 CLK1.n825 8.855
R5707 CLK1.n966 CLK1.n826 8.855
R5708 CLK1.n969 CLK1.n968 8.855
R5709 CLK1.n968 CLK1.n967 8.855
R5710 CLK1.n823 CLK1.n822 8.855
R5711 CLK1.n822 CLK1.n821 8.855
R5712 CLK1.n974 CLK1.n973 8.855
R5713 CLK1.n975 CLK1.n974 8.855
R5714 CLK1.n820 CLK1.n819 8.855
R5715 CLK1.n976 CLK1.n820 8.855
R5716 CLK1.n979 CLK1.n978 8.855
R5717 CLK1.n978 CLK1.n977 8.855
R5718 CLK1.n815 CLK1.n814 8.855
R5719 CLK1.n814 CLK1.n813 8.855
R5720 CLK1.n986 CLK1.n985 8.855
R5721 CLK1.n987 CLK1.n986 8.855
R5722 CLK1.n816 CLK1.n812 8.855
R5723 CLK1.n558 CLK1.n557 8.855
R5724 CLK1.n564 CLK1.n563 8.855
R5725 CLK1.n565 CLK1.n564 8.855
R5726 CLK1.n555 CLK1.n554 8.855
R5727 CLK1.n566 CLK1.n555 8.855
R5728 CLK1.n569 CLK1.n568 8.855
R5729 CLK1.n568 CLK1.n567 8.855
R5730 CLK1.n552 CLK1.n551 8.855
R5731 CLK1.n551 CLK1.n550 8.855
R5732 CLK1.n574 CLK1.n573 8.855
R5733 CLK1.n575 CLK1.n574 8.855
R5734 CLK1.n549 CLK1.n548 8.855
R5735 CLK1.n576 CLK1.n549 8.855
R5736 CLK1.n580 CLK1.n579 8.855
R5737 CLK1.n579 CLK1.n578 8.855
R5738 CLK1.n546 CLK1.n545 8.855
R5739 CLK1.n577 CLK1.n545 8.855
R5740 CLK1.n586 CLK1.n585 8.855
R5741 CLK1.n587 CLK1.n586 8.855
R5742 CLK1.n544 CLK1.n543 8.855
R5743 CLK1.n588 CLK1.n544 8.855
R5744 CLK1.n591 CLK1.n590 8.855
R5745 CLK1.n590 CLK1.n589 8.855
R5746 CLK1.n540 CLK1.n539 8.855
R5747 CLK1.n539 CLK1.n538 8.855
R5748 CLK1.n597 CLK1.n596 8.855
R5749 CLK1.n598 CLK1.n597 8.855
R5750 CLK1.n537 CLK1.n536 8.855
R5751 CLK1.n599 CLK1.n537 8.855
R5752 CLK1.n602 CLK1.n601 8.855
R5753 CLK1.n601 CLK1.n600 8.855
R5754 CLK1.n534 CLK1.n533 8.855
R5755 CLK1.n533 CLK1.n532 8.855
R5756 CLK1.n608 CLK1.n607 8.855
R5757 CLK1.n609 CLK1.n608 8.855
R5758 CLK1.n531 CLK1.n530 8.855
R5759 CLK1.n610 CLK1.n531 8.855
R5760 CLK1.n613 CLK1.n612 8.855
R5761 CLK1.n612 CLK1.n611 8.855
R5762 CLK1.n527 CLK1.n526 8.855
R5763 CLK1.n526 CLK1.n525 8.855
R5764 CLK1.n619 CLK1.n618 8.855
R5765 CLK1.n620 CLK1.n619 8.855
R5766 CLK1.n524 CLK1.n523 8.855
R5767 CLK1.n688 CLK1.n687 8.855
R5768 CLK1.n694 CLK1.n693 8.855
R5769 CLK1.n695 CLK1.n694 8.855
R5770 CLK1.n685 CLK1.n684 8.855
R5771 CLK1.n696 CLK1.n685 8.855
R5772 CLK1.n700 CLK1.n699 8.855
R5773 CLK1.n699 CLK1.n698 8.855
R5774 CLK1.n682 CLK1.n681 8.855
R5775 CLK1.n697 CLK1.n681 8.855
R5776 CLK1.n706 CLK1.n705 8.855
R5777 CLK1.n707 CLK1.n706 8.855
R5778 CLK1.n680 CLK1.n679 8.855
R5779 CLK1.n708 CLK1.n680 8.855
R5780 CLK1.n711 CLK1.n710 8.855
R5781 CLK1.n710 CLK1.n709 8.855
R5782 CLK1.n676 CLK1.n675 8.855
R5783 CLK1.n675 CLK1.n674 8.855
R5784 CLK1.n717 CLK1.n716 8.855
R5785 CLK1.n718 CLK1.n717 8.855
R5786 CLK1.n673 CLK1.n672 8.855
R5787 CLK1.n719 CLK1.n673 8.855
R5788 CLK1.n722 CLK1.n721 8.855
R5789 CLK1.n721 CLK1.n720 8.855
R5790 CLK1.n670 CLK1.n669 8.855
R5791 CLK1.n669 CLK1.n668 8.855
R5792 CLK1.n728 CLK1.n727 8.855
R5793 CLK1.n729 CLK1.n728 8.855
R5794 CLK1.n667 CLK1.n666 8.855
R5795 CLK1.n664 CLK1.n663 8.855
R5796 CLK1.n738 CLK1.n737 8.855
R5797 CLK1.n737 CLK1.n736 8.855
R5798 CLK1.n660 CLK1.n659 8.855
R5799 CLK1.n659 CLK1.n658 8.855
R5800 CLK1.n744 CLK1.n743 8.855
R5801 CLK1.n745 CLK1.n744 8.855
R5802 CLK1.n657 CLK1.n656 8.855
R5803 CLK1.n746 CLK1.n657 8.855
R5804 CLK1.n749 CLK1.n748 8.855
R5805 CLK1.n748 CLK1.n747 8.855
R5806 CLK1.n654 CLK1.n653 8.855
R5807 CLK1.n653 CLK1.n652 8.855
R5808 CLK1.n755 CLK1.n754 8.855
R5809 CLK1.n756 CLK1.n755 8.855
R5810 CLK1.n651 CLK1.n650 8.855
R5811 CLK1.n757 CLK1.n651 8.855
R5812 CLK1.n760 CLK1.n759 8.855
R5813 CLK1.n759 CLK1.n758 8.855
R5814 CLK1.n648 CLK1.n647 8.855
R5815 CLK1.n647 CLK1.n646 8.855
R5816 CLK1.n767 CLK1.n766 8.855
R5817 CLK1.n768 CLK1.n767 8.855
R5818 CLK1.n645 CLK1.n644 8.855
R5819 CLK1.n769 CLK1.n645 8.855
R5820 CLK1.n773 CLK1.n772 8.855
R5821 CLK1.n772 CLK1.n771 8.855
R5822 CLK1.n643 CLK1.n642 8.855
R5823 CLK1.n770 CLK1.n642 8.855
R5824 CLK1.n779 CLK1.n778 8.855
R5825 CLK1.n780 CLK1.n779 8.855
R5826 CLK1.n641 CLK1.n640 8.855
R5827 CLK1.n781 CLK1.n641 8.855
R5828 CLK1.n784 CLK1.n783 8.855
R5829 CLK1.n783 CLK1.n782 8.855
R5830 CLK1.n638 CLK1.n637 8.855
R5831 CLK1.n637 CLK1.n636 8.855
R5832 CLK1.n789 CLK1.n788 8.855
R5833 CLK1.n790 CLK1.n789 8.855
R5834 CLK1.n635 CLK1.n634 8.855
R5835 CLK1.n791 CLK1.n635 8.855
R5836 CLK1.n794 CLK1.n793 8.855
R5837 CLK1.n793 CLK1.n792 8.855
R5838 CLK1.n630 CLK1.n629 8.855
R5839 CLK1.n629 CLK1.n628 8.855
R5840 CLK1.n801 CLK1.n800 8.855
R5841 CLK1.n802 CLK1.n801 8.855
R5842 CLK1.n631 CLK1.n627 8.855
R5843 CLK1.n439 CLK1.n438 8.855
R5844 CLK1.n440 CLK1.n439 8.855
R5845 CLK1.n430 CLK1.n429 8.855
R5846 CLK1.n441 CLK1.n430 8.855
R5847 CLK1.n445 CLK1.n444 8.855
R5848 CLK1.n444 CLK1.n443 8.855
R5849 CLK1.n427 CLK1.n426 8.855
R5850 CLK1.n442 CLK1.n426 8.855
R5851 CLK1.n451 CLK1.n450 8.855
R5852 CLK1.n452 CLK1.n451 8.855
R5853 CLK1.n425 CLK1.n424 8.855
R5854 CLK1.n453 CLK1.n425 8.855
R5855 CLK1.n456 CLK1.n455 8.855
R5856 CLK1.n455 CLK1.n454 8.855
R5857 CLK1.n421 CLK1.n420 8.855
R5858 CLK1.n420 CLK1.n419 8.855
R5859 CLK1.n462 CLK1.n461 8.855
R5860 CLK1.n463 CLK1.n462 8.855
R5861 CLK1.n418 CLK1.n417 8.855
R5862 CLK1.n464 CLK1.n418 8.855
R5863 CLK1.n467 CLK1.n466 8.855
R5864 CLK1.n466 CLK1.n465 8.855
R5865 CLK1.n415 CLK1.n414 8.855
R5866 CLK1.n414 CLK1.n413 8.855
R5867 CLK1.n473 CLK1.n472 8.855
R5868 CLK1.n474 CLK1.n473 8.855
R5869 CLK1.n412 CLK1.n411 8.855
R5870 CLK1.n409 CLK1.n408 8.855
R5871 CLK1.n483 CLK1.n482 8.855
R5872 CLK1.n484 CLK1.n483 8.855
R5873 CLK1.n405 CLK1.n403 8.855
R5874 CLK1.n485 CLK1.n405 8.855
R5875 CLK1.n1052 CLK1.n1051 8.855
R5876 CLK1.n1051 CLK1.n1050 8.855
R5877 CLK1.n406 CLK1.n404 8.855
R5878 CLK1.n1049 CLK1.n406 8.855
R5879 CLK1.n1047 CLK1.n1046 8.855
R5880 CLK1.n1048 CLK1.n1047 8.855
R5881 CLK1.n488 CLK1.n487 8.855
R5882 CLK1.n487 CLK1.n486 8.855
R5883 CLK1.n1042 CLK1.n1041 8.855
R5884 CLK1.n1041 CLK1.n1040 8.855
R5885 CLK1.n491 CLK1.n490 8.855
R5886 CLK1.n1039 CLK1.n491 8.855
R5887 CLK1.n1037 CLK1.n1036 8.855
R5888 CLK1.n1038 CLK1.n1037 8.855
R5889 CLK1.n493 CLK1.n492 8.855
R5890 CLK1.n499 CLK1.n492 8.855
R5891 CLK1.n1032 CLK1.n1031 8.855
R5892 CLK1.n1031 CLK1.n1030 8.855
R5893 CLK1.n498 CLK1.n497 8.855
R5894 CLK1.n1029 CLK1.n498 8.855
R5895 CLK1.n1027 CLK1.n1026 8.855
R5896 CLK1.n1028 CLK1.n1027 8.855
R5897 CLK1.n502 CLK1.n501 8.855
R5898 CLK1.n501 CLK1.n500 8.855
R5899 CLK1.n1022 CLK1.n1021 8.855
R5900 CLK1.n1021 CLK1.n1020 8.855
R5901 CLK1.n505 CLK1.n504 8.855
R5902 CLK1.n1019 CLK1.n505 8.855
R5903 CLK1.n1017 CLK1.n1016 8.855
R5904 CLK1.n1018 CLK1.n1017 8.855
R5905 CLK1.n508 CLK1.n507 8.855
R5906 CLK1.n507 CLK1.n506 8.855
R5907 CLK1.n1012 CLK1.n1011 8.855
R5908 CLK1.n1011 CLK1.n1010 8.855
R5909 CLK1.n512 CLK1.n511 8.855
R5910 CLK1.n1009 CLK1.n512 8.855
R5911 CLK1.n1007 CLK1.n1006 8.855
R5912 CLK1.n1008 CLK1.n1007 8.855
R5913 CLK1.n515 CLK1.n514 8.855
R5914 CLK1.n514 CLK1.n513 8.855
R5915 CLK1.n1001 CLK1.n1000 8.855
R5916 CLK1.n1000 CLK1.n999 8.855
R5917 CLK1.n1061 CLK1.n398 8.855
R5918 CLK1.n1187 CLK1.n1186 8.855
R5919 CLK1.n318 CLK1.n317 8.855
R5920 CLK1.n1196 CLK1.n1195 8.855
R5921 CLK1.n1197 CLK1.n1196 8.855
R5922 CLK1.n315 CLK1.n314 8.855
R5923 CLK1.n1198 CLK1.n315 8.855
R5924 CLK1.n1201 CLK1.n1200 8.855
R5925 CLK1.n1200 CLK1.n1199 8.855
R5926 CLK1.n312 CLK1.n311 8.855
R5927 CLK1.n311 CLK1.n310 8.855
R5928 CLK1.n1206 CLK1.n1205 8.855
R5929 CLK1.n1207 CLK1.n1206 8.855
R5930 CLK1.n309 CLK1.n308 8.855
R5931 CLK1.n1208 CLK1.n309 8.855
R5932 CLK1.n1212 CLK1.n1211 8.855
R5933 CLK1.n1211 CLK1.n1210 8.855
R5934 CLK1.n306 CLK1.n305 8.855
R5935 CLK1.n1209 CLK1.n305 8.855
R5936 CLK1.n1218 CLK1.n1217 8.855
R5937 CLK1.n1219 CLK1.n1218 8.855
R5938 CLK1.n304 CLK1.n303 8.855
R5939 CLK1.n1220 CLK1.n304 8.855
R5940 CLK1.n1223 CLK1.n1222 8.855
R5941 CLK1.n1222 CLK1.n1221 8.855
R5942 CLK1.n300 CLK1.n299 8.855
R5943 CLK1.n299 CLK1.n298 8.855
R5944 CLK1.n1229 CLK1.n1228 8.855
R5945 CLK1.n1230 CLK1.n1229 8.855
R5946 CLK1.n297 CLK1.n296 8.855
R5947 CLK1.n1231 CLK1.n297 8.855
R5948 CLK1.n1234 CLK1.n1233 8.855
R5949 CLK1.n1233 CLK1.n1232 8.855
R5950 CLK1.n294 CLK1.n293 8.855
R5951 CLK1.n293 CLK1.n292 8.855
R5952 CLK1.n1240 CLK1.n1239 8.855
R5953 CLK1.n1241 CLK1.n1240 8.855
R5954 CLK1.n291 CLK1.n290 8.855
R5955 CLK1.n1242 CLK1.n291 8.855
R5956 CLK1.n1245 CLK1.n1244 8.855
R5957 CLK1.n1244 CLK1.n1243 8.855
R5958 CLK1.n287 CLK1.n286 8.855
R5959 CLK1.n286 CLK1.n285 8.855
R5960 CLK1.n1251 CLK1.n1250 8.855
R5961 CLK1.n1252 CLK1.n1251 8.855
R5962 CLK1.n284 CLK1.n283 8.855
R5963 CLK1.n1320 CLK1.n1319 8.855
R5964 CLK1.n1326 CLK1.n1325 8.855
R5965 CLK1.n1327 CLK1.n1326 8.855
R5966 CLK1.n1317 CLK1.n1316 8.855
R5967 CLK1.n1328 CLK1.n1317 8.855
R5968 CLK1.n1332 CLK1.n1331 8.855
R5969 CLK1.n1331 CLK1.n1330 8.855
R5970 CLK1.n1314 CLK1.n1313 8.855
R5971 CLK1.n1329 CLK1.n1313 8.855
R5972 CLK1.n1338 CLK1.n1337 8.855
R5973 CLK1.n1339 CLK1.n1338 8.855
R5974 CLK1.n1312 CLK1.n1311 8.855
R5975 CLK1.n1340 CLK1.n1312 8.855
R5976 CLK1.n1343 CLK1.n1342 8.855
R5977 CLK1.n1342 CLK1.n1341 8.855
R5978 CLK1.n1308 CLK1.n1307 8.855
R5979 CLK1.n1307 CLK1.n1306 8.855
R5980 CLK1.n1349 CLK1.n1348 8.855
R5981 CLK1.n1350 CLK1.n1349 8.855
R5982 CLK1.n1305 CLK1.n1304 8.855
R5983 CLK1.n1351 CLK1.n1305 8.855
R5984 CLK1.n1354 CLK1.n1353 8.855
R5985 CLK1.n1353 CLK1.n1352 8.855
R5986 CLK1.n1302 CLK1.n1301 8.855
R5987 CLK1.n1301 CLK1.n1300 8.855
R5988 CLK1.n1360 CLK1.n1359 8.855
R5989 CLK1.n1361 CLK1.n1360 8.855
R5990 CLK1.n1299 CLK1.n1298 8.855
R5991 CLK1.n1296 CLK1.n1295 8.855
R5992 CLK1.n1370 CLK1.n1369 8.855
R5993 CLK1.n1369 CLK1.n1368 8.855
R5994 CLK1.n1292 CLK1.n1291 8.855
R5995 CLK1.n1291 CLK1.n1290 8.855
R5996 CLK1.n1376 CLK1.n1375 8.855
R5997 CLK1.n1377 CLK1.n1376 8.855
R5998 CLK1.n1289 CLK1.n1288 8.855
R5999 CLK1.n1378 CLK1.n1289 8.855
R6000 CLK1.n1381 CLK1.n1380 8.855
R6001 CLK1.n1380 CLK1.n1379 8.855
R6002 CLK1.n1286 CLK1.n1285 8.855
R6003 CLK1.n1285 CLK1.n1284 8.855
R6004 CLK1.n1387 CLK1.n1386 8.855
R6005 CLK1.n1388 CLK1.n1387 8.855
R6006 CLK1.n1283 CLK1.n1282 8.855
R6007 CLK1.n1389 CLK1.n1283 8.855
R6008 CLK1.n1392 CLK1.n1391 8.855
R6009 CLK1.n1391 CLK1.n1390 8.855
R6010 CLK1.n1280 CLK1.n1279 8.855
R6011 CLK1.n1279 CLK1.n1278 8.855
R6012 CLK1.n1399 CLK1.n1398 8.855
R6013 CLK1.n1400 CLK1.n1399 8.855
R6014 CLK1.n1277 CLK1.n1276 8.855
R6015 CLK1.n1401 CLK1.n1277 8.855
R6016 CLK1.n1405 CLK1.n1404 8.855
R6017 CLK1.n1404 CLK1.n1403 8.855
R6018 CLK1.n1275 CLK1.n1274 8.855
R6019 CLK1.n1402 CLK1.n1274 8.855
R6020 CLK1.n1411 CLK1.n1410 8.855
R6021 CLK1.n1412 CLK1.n1411 8.855
R6022 CLK1.n1273 CLK1.n1272 8.855
R6023 CLK1.n1413 CLK1.n1273 8.855
R6024 CLK1.n1416 CLK1.n1415 8.855
R6025 CLK1.n1415 CLK1.n1414 8.855
R6026 CLK1.n1270 CLK1.n1269 8.855
R6027 CLK1.n1269 CLK1.n1268 8.855
R6028 CLK1.n1421 CLK1.n1420 8.855
R6029 CLK1.n1422 CLK1.n1421 8.855
R6030 CLK1.n1267 CLK1.n1266 8.855
R6031 CLK1.n1423 CLK1.n1267 8.855
R6032 CLK1.n1426 CLK1.n1425 8.855
R6033 CLK1.n1425 CLK1.n1424 8.855
R6034 CLK1.n1262 CLK1.n1261 8.855
R6035 CLK1.n1261 CLK1.n1260 8.855
R6036 CLK1.n1433 CLK1.n1432 8.855
R6037 CLK1.n1434 CLK1.n1433 8.855
R6038 CLK1.n1263 CLK1.n1259 8.855
R6039 CLK1.n1056 CLK1.n1055 8.365
R6040 CLK1.n1190 CLK1.n319 8.365
R6041 CLK1.n137 CLK1.t187 8.189
R6042 CLK1.n143 CLK1.t173 8.189
R6043 CLK1.n43 CLK1.t55 8.189
R6044 CLK1.n49 CLK1.t94 8.189
R6045 CLK1.n245 CLK1.t89 8.189
R6046 CLK1.n255 CLK1.t140 8.189
R6047 CLK1.t109 CLK1.n1585 8.189
R6048 CLK1.n1588 CLK1.t152 8.189
R6049 CLK1.t2 CLK1.n1525 8.189
R6050 CLK1.t83 CLK1.n1491 8.189
R6051 CLK1.t129 CLK1.n1220 8.189
R6052 CLK1.t14 CLK1.n298 8.189
R6053 CLK1.t125 CLK1.n365 8.189
R6054 CLK1.t179 CLK1.n331 8.189
R6055 CLK1.t114 CLK1.n453 8.189
R6056 CLK1.t60 CLK1.n419 8.189
R6057 CLK1.n1030 CLK1.t64 8.189
R6058 CLK1.t43 CLK1.n1028 8.189
R6059 CLK1.t135 CLK1.n953 8.189
R6060 CLK1.n956 CLK1.t103 8.189
R6061 CLK1.t157 CLK1.n893 8.189
R6062 CLK1.t6 CLK1.n859 8.189
R6063 CLK1.t142 CLK1.n588 8.189
R6064 CLK1.t159 CLK1.n538 8.189
R6065 CLK1.t46 CLK1.n768 8.189
R6066 CLK1.n771 CLK1.t183 8.189
R6067 CLK1.t67 CLK1.n708 8.189
R6068 CLK1.t71 CLK1.n674 8.189
R6069 CLK1.t171 CLK1.n1400 8.189
R6070 CLK1.n1403 CLK1.t148 8.189
R6071 CLK1.t27 CLK1.n1340 8.189
R6072 CLK1.t20 CLK1.n1306 8.189
R6073 CLK1.n1100 CLK1.n1099 7.776
R6074 CLK1.n1110 CLK1.n1109 7.776
R6075 CLK1.n180 CLK1.n0 6.776
R6076 CLK1.n103 CLK1.n4 6.776
R6077 CLK1.n17 CLK1.n8 6.776
R6078 CLK1.n272 CLK1.n201 6.776
R6079 CLK1.n1613 CLK1.n1449 6.776
R6080 CLK1.n1558 CLK1.n1478 6.776
R6081 CLK1.n289 CLK1.n288 6.776
R6082 CLK1.n1124 CLK1.n1108 6.776
R6083 CLK1.n981 CLK1.n817 6.776
R6084 CLK1.n926 CLK1.n846 6.776
R6085 CLK1.n529 CLK1.n528 6.776
R6086 CLK1.n741 CLK1.n661 6.776
R6087 CLK1.n796 CLK1.n632 6.776
R6088 CLK1.n1004 CLK1.n516 6.776
R6089 CLK1.n1373 CLK1.n1293 6.776
R6090 CLK1.n1428 CLK1.n1264 6.776
R6091 CLK1.n1062 CLK1.n1060 6.754
R6092 CLK1.n1184 CLK1.n1183 6.754
R6093 CLK1.n141 CLK1.n3 4.938
R6094 CLK1.n47 CLK1.n7 4.938
R6095 CLK1.n251 CLK1.n213 4.938
R6096 CLK1.n1581 CLK1.n1580 4.938
R6097 CLK1.n1529 CLK1.n1494 4.938
R6098 CLK1.n1224 CLK1.n301 4.938
R6099 CLK1.n1082 CLK1.n1080 4.938
R6100 CLK1.n1082 CLK1.n1081 4.938
R6101 CLK1.n369 CLK1.n334 4.938
R6102 CLK1.n496 CLK1.n495 4.938
R6103 CLK1.n457 CLK1.n422 4.938
R6104 CLK1.n949 CLK1.n948 4.938
R6105 CLK1.n897 CLK1.n862 4.938
R6106 CLK1.n592 CLK1.n541 4.938
R6107 CLK1.n764 CLK1.n763 4.938
R6108 CLK1.n712 CLK1.n677 4.938
R6109 CLK1.n1396 CLK1.n1395 4.938
R6110 CLK1.n1344 CLK1.n1309 4.938
R6111 CLK1.n560 CLK1.n559 4.687
R6112 CLK1.n1192 CLK1.n1191 4.687
R6113 CLK1.n227 CLK1.n226 4.675
R6114 CLK1.n1507 CLK1.n1506 4.662
R6115 CLK1.n347 CLK1.n346 4.662
R6116 CLK1.n875 CLK1.n874 4.662
R6117 CLK1.n690 CLK1.n689 4.662
R6118 CLK1.n435 CLK1.n434 4.662
R6119 CLK1.n1322 CLK1.n1321 4.662
R6120 CLK1.n16 CLK1.n15 4.65
R6121 CLK1.n21 CLK1.n20 4.65
R6122 CLK1.n25 CLK1.n24 4.65
R6123 CLK1.n29 CLK1.n28 4.65
R6124 CLK1.n33 CLK1.n32 4.65
R6125 CLK1.n38 CLK1.n37 4.65
R6126 CLK1.n42 CLK1.n41 4.65
R6127 CLK1.n46 CLK1.n45 4.65
R6128 CLK1.n48 CLK1.n47 4.65
R6129 CLK1.n52 CLK1.n51 4.65
R6130 CLK1.n56 CLK1.n55 4.65
R6131 CLK1.n60 CLK1.n59 4.65
R6132 CLK1.n65 CLK1.n64 4.65
R6133 CLK1.n69 CLK1.n68 4.65
R6134 CLK1.n73 CLK1.n72 4.65
R6135 CLK1.n77 CLK1.n76 4.65
R6136 CLK1.n81 CLK1.n80 4.65
R6137 CLK1.n85 CLK1.n84 4.65
R6138 CLK1.n88 CLK1.n87 4.65
R6139 CLK1.n90 CLK1.n89 4.65
R6140 CLK1.n94 CLK1.n93 4.65
R6141 CLK1.n98 CLK1.n97 4.65
R6142 CLK1.n102 CLK1.n101 4.65
R6143 CLK1.n107 CLK1.n106 4.65
R6144 CLK1.n111 CLK1.n110 4.65
R6145 CLK1.n115 CLK1.n114 4.65
R6146 CLK1.n119 CLK1.n118 4.65
R6147 CLK1.n123 CLK1.n122 4.65
R6148 CLK1.n127 CLK1.n126 4.65
R6149 CLK1.n132 CLK1.n131 4.65
R6150 CLK1.n136 CLK1.n135 4.65
R6151 CLK1.n140 CLK1.n139 4.65
R6152 CLK1.n142 CLK1.n141 4.65
R6153 CLK1.n146 CLK1.n145 4.65
R6154 CLK1.n150 CLK1.n149 4.65
R6155 CLK1.n154 CLK1.n153 4.65
R6156 CLK1.n159 CLK1.n158 4.65
R6157 CLK1.n163 CLK1.n162 4.65
R6158 CLK1.n167 CLK1.n166 4.65
R6159 CLK1.n171 CLK1.n170 4.65
R6160 CLK1.n175 CLK1.n174 4.65
R6161 CLK1.n179 CLK1.n178 4.65
R6162 CLK1.n184 CLK1.n183 4.65
R6163 CLK1.n188 CLK1.n187 4.65
R6164 CLK1.n192 CLK1.n191 4.65
R6165 CLK1.n194 CLK1.n193 4.65
R6166 CLK1.n228 CLK1.n225 4.65
R6167 CLK1.n230 CLK1.n229 4.65
R6168 CLK1.n221 CLK1.n220 4.65
R6169 CLK1.n237 CLK1.n236 4.65
R6170 CLK1.n238 CLK1.n219 4.65
R6171 CLK1.n241 CLK1.n240 4.65
R6172 CLK1.n215 CLK1.n214 4.65
R6173 CLK1.n249 CLK1.n248 4.65
R6174 CLK1.n250 CLK1.n212 4.65
R6175 CLK1.n252 CLK1.n251 4.65
R6176 CLK1.n209 CLK1.n208 4.65
R6177 CLK1.n259 CLK1.n258 4.65
R6178 CLK1.n260 CLK1.n207 4.65
R6179 CLK1.n263 CLK1.n262 4.65
R6180 CLK1.n203 CLK1.n202 4.65
R6181 CLK1.n270 CLK1.n269 4.65
R6182 CLK1.n271 CLK1.n200 4.65
R6183 CLK1.n274 CLK1.n273 4.65
R6184 CLK1.n196 CLK1.n195 4.65
R6185 CLK1.n279 CLK1.n278 4.65
R6186 CLK1.n1508 CLK1.n1505 4.65
R6187 CLK1.n1510 CLK1.n1509 4.65
R6188 CLK1.n1501 CLK1.n1500 4.65
R6189 CLK1.n1518 CLK1.n1517 4.65
R6190 CLK1.n1520 CLK1.n1499 4.65
R6191 CLK1.n1522 CLK1.n1521 4.65
R6192 CLK1.n1496 CLK1.n1495 4.65
R6193 CLK1.n1529 CLK1.n1528 4.65
R6194 CLK1.n1530 CLK1.n1493 4.65
R6195 CLK1.n1533 CLK1.n1532 4.65
R6196 CLK1.n1531 CLK1.n1489 4.65
R6197 CLK1.n1540 CLK1.n1539 4.65
R6198 CLK1.n1541 CLK1.n1487 4.65
R6199 CLK1.n1544 CLK1.n1543 4.65
R6200 CLK1.n1542 CLK1.n1483 4.65
R6201 CLK1.n1549 CLK1.n1548 4.65
R6202 CLK1.n1551 CLK1.n1550 4.65
R6203 CLK1.n1480 CLK1.n1479 4.65
R6204 CLK1.n1556 CLK1.n1555 4.65
R6205 CLK1.n1557 CLK1.n1477 4.65
R6206 CLK1.n1560 CLK1.n1559 4.65
R6207 CLK1.n1473 CLK1.n1472 4.65
R6208 CLK1.n1567 CLK1.n1566 4.65
R6209 CLK1.n1568 CLK1.n1471 4.65
R6210 CLK1.n1571 CLK1.n1570 4.65
R6211 CLK1.n1569 CLK1.n1467 4.65
R6212 CLK1.n1578 CLK1.n1577 4.65
R6213 CLK1.n1579 CLK1.n1465 4.65
R6214 CLK1.n1583 CLK1.n1582 4.65
R6215 CLK1.n1581 CLK1.n1461 4.65
R6216 CLK1.n1591 CLK1.n1590 4.65
R6217 CLK1.n1592 CLK1.n1460 4.65
R6218 CLK1.n1595 CLK1.n1594 4.65
R6219 CLK1.n1457 CLK1.n1456 4.65
R6220 CLK1.n1602 CLK1.n1601 4.65
R6221 CLK1.n1603 CLK1.n1455 4.65
R6222 CLK1.n1605 CLK1.n1604 4.65
R6223 CLK1.n1451 CLK1.n1450 4.65
R6224 CLK1.n1612 CLK1.n1611 4.65
R6225 CLK1.n1614 CLK1.n1447 4.65
R6226 CLK1.n1617 CLK1.n1616 4.65
R6227 CLK1.n1615 CLK1.n1448 4.65
R6228 CLK1.n389 CLK1.n388 4.65
R6229 CLK1.n348 CLK1.n345 4.65
R6230 CLK1.n350 CLK1.n349 4.65
R6231 CLK1.n341 CLK1.n340 4.65
R6232 CLK1.n358 CLK1.n357 4.65
R6233 CLK1.n360 CLK1.n339 4.65
R6234 CLK1.n362 CLK1.n361 4.65
R6235 CLK1.n336 CLK1.n335 4.65
R6236 CLK1.n369 CLK1.n368 4.65
R6237 CLK1.n370 CLK1.n333 4.65
R6238 CLK1.n373 CLK1.n372 4.65
R6239 CLK1.n371 CLK1.n329 4.65
R6240 CLK1.n380 CLK1.n379 4.65
R6241 CLK1.n381 CLK1.n327 4.65
R6242 CLK1.n384 CLK1.n383 4.65
R6243 CLK1.n382 CLK1.n323 4.65
R6244 CLK1.n876 CLK1.n873 4.65
R6245 CLK1.n878 CLK1.n877 4.65
R6246 CLK1.n869 CLK1.n868 4.65
R6247 CLK1.n886 CLK1.n885 4.65
R6248 CLK1.n888 CLK1.n867 4.65
R6249 CLK1.n890 CLK1.n889 4.65
R6250 CLK1.n864 CLK1.n863 4.65
R6251 CLK1.n897 CLK1.n896 4.65
R6252 CLK1.n898 CLK1.n861 4.65
R6253 CLK1.n901 CLK1.n900 4.65
R6254 CLK1.n899 CLK1.n857 4.65
R6255 CLK1.n908 CLK1.n907 4.65
R6256 CLK1.n909 CLK1.n855 4.65
R6257 CLK1.n912 CLK1.n911 4.65
R6258 CLK1.n910 CLK1.n851 4.65
R6259 CLK1.n917 CLK1.n916 4.65
R6260 CLK1.n919 CLK1.n918 4.65
R6261 CLK1.n848 CLK1.n847 4.65
R6262 CLK1.n924 CLK1.n923 4.65
R6263 CLK1.n925 CLK1.n845 4.65
R6264 CLK1.n928 CLK1.n927 4.65
R6265 CLK1.n841 CLK1.n840 4.65
R6266 CLK1.n935 CLK1.n934 4.65
R6267 CLK1.n936 CLK1.n839 4.65
R6268 CLK1.n939 CLK1.n938 4.65
R6269 CLK1.n937 CLK1.n835 4.65
R6270 CLK1.n946 CLK1.n945 4.65
R6271 CLK1.n947 CLK1.n833 4.65
R6272 CLK1.n951 CLK1.n950 4.65
R6273 CLK1.n949 CLK1.n829 4.65
R6274 CLK1.n959 CLK1.n958 4.65
R6275 CLK1.n960 CLK1.n828 4.65
R6276 CLK1.n963 CLK1.n962 4.65
R6277 CLK1.n825 CLK1.n824 4.65
R6278 CLK1.n970 CLK1.n969 4.65
R6279 CLK1.n971 CLK1.n823 4.65
R6280 CLK1.n973 CLK1.n972 4.65
R6281 CLK1.n819 CLK1.n818 4.65
R6282 CLK1.n980 CLK1.n979 4.65
R6283 CLK1.n982 CLK1.n815 4.65
R6284 CLK1.n985 CLK1.n984 4.65
R6285 CLK1.n983 CLK1.n816 4.65
R6286 CLK1.n561 CLK1.n558 4.65
R6287 CLK1.n563 CLK1.n562 4.65
R6288 CLK1.n554 CLK1.n553 4.65
R6289 CLK1.n570 CLK1.n569 4.65
R6290 CLK1.n571 CLK1.n552 4.65
R6291 CLK1.n573 CLK1.n572 4.65
R6292 CLK1.n548 CLK1.n547 4.65
R6293 CLK1.n581 CLK1.n580 4.65
R6294 CLK1.n583 CLK1.n546 4.65
R6295 CLK1.n585 CLK1.n584 4.65
R6296 CLK1.n543 CLK1.n542 4.65
R6297 CLK1.n592 CLK1.n591 4.65
R6298 CLK1.n593 CLK1.n540 4.65
R6299 CLK1.n596 CLK1.n595 4.65
R6300 CLK1.n594 CLK1.n536 4.65
R6301 CLK1.n603 CLK1.n602 4.65
R6302 CLK1.n604 CLK1.n534 4.65
R6303 CLK1.n607 CLK1.n606 4.65
R6304 CLK1.n605 CLK1.n530 4.65
R6305 CLK1.n614 CLK1.n613 4.65
R6306 CLK1.n615 CLK1.n527 4.65
R6307 CLK1.n618 CLK1.n617 4.65
R6308 CLK1.n616 CLK1.n523 4.65
R6309 CLK1.n623 CLK1.n622 4.65
R6310 CLK1.n691 CLK1.n688 4.65
R6311 CLK1.n693 CLK1.n692 4.65
R6312 CLK1.n684 CLK1.n683 4.65
R6313 CLK1.n701 CLK1.n700 4.65
R6314 CLK1.n703 CLK1.n682 4.65
R6315 CLK1.n705 CLK1.n704 4.65
R6316 CLK1.n679 CLK1.n678 4.65
R6317 CLK1.n712 CLK1.n711 4.65
R6318 CLK1.n713 CLK1.n676 4.65
R6319 CLK1.n716 CLK1.n715 4.65
R6320 CLK1.n714 CLK1.n672 4.65
R6321 CLK1.n723 CLK1.n722 4.65
R6322 CLK1.n724 CLK1.n670 4.65
R6323 CLK1.n727 CLK1.n726 4.65
R6324 CLK1.n725 CLK1.n666 4.65
R6325 CLK1.n732 CLK1.n731 4.65
R6326 CLK1.n734 CLK1.n733 4.65
R6327 CLK1.n663 CLK1.n662 4.65
R6328 CLK1.n739 CLK1.n738 4.65
R6329 CLK1.n740 CLK1.n660 4.65
R6330 CLK1.n743 CLK1.n742 4.65
R6331 CLK1.n656 CLK1.n655 4.65
R6332 CLK1.n750 CLK1.n749 4.65
R6333 CLK1.n751 CLK1.n654 4.65
R6334 CLK1.n754 CLK1.n753 4.65
R6335 CLK1.n752 CLK1.n650 4.65
R6336 CLK1.n761 CLK1.n760 4.65
R6337 CLK1.n762 CLK1.n648 4.65
R6338 CLK1.n766 CLK1.n765 4.65
R6339 CLK1.n764 CLK1.n644 4.65
R6340 CLK1.n774 CLK1.n773 4.65
R6341 CLK1.n775 CLK1.n643 4.65
R6342 CLK1.n778 CLK1.n777 4.65
R6343 CLK1.n640 CLK1.n639 4.65
R6344 CLK1.n785 CLK1.n784 4.65
R6345 CLK1.n786 CLK1.n638 4.65
R6346 CLK1.n788 CLK1.n787 4.65
R6347 CLK1.n634 CLK1.n633 4.65
R6348 CLK1.n795 CLK1.n794 4.65
R6349 CLK1.n797 CLK1.n630 4.65
R6350 CLK1.n800 CLK1.n799 4.65
R6351 CLK1.n798 CLK1.n631 4.65
R6352 CLK1.n518 CLK1.n517 4.65
R6353 CLK1.n477 CLK1.n476 4.65
R6354 CLK1.n436 CLK1.n433 4.65
R6355 CLK1.n438 CLK1.n437 4.65
R6356 CLK1.n429 CLK1.n428 4.65
R6357 CLK1.n446 CLK1.n445 4.65
R6358 CLK1.n448 CLK1.n427 4.65
R6359 CLK1.n450 CLK1.n449 4.65
R6360 CLK1.n424 CLK1.n423 4.65
R6361 CLK1.n457 CLK1.n456 4.65
R6362 CLK1.n458 CLK1.n421 4.65
R6363 CLK1.n461 CLK1.n460 4.65
R6364 CLK1.n459 CLK1.n417 4.65
R6365 CLK1.n468 CLK1.n467 4.65
R6366 CLK1.n469 CLK1.n415 4.65
R6367 CLK1.n472 CLK1.n471 4.65
R6368 CLK1.n470 CLK1.n411 4.65
R6369 CLK1.n479 CLK1.n478 4.65
R6370 CLK1.n480 CLK1.n409 4.65
R6371 CLK1.n482 CLK1.n481 4.65
R6372 CLK1.n403 CLK1.n401 4.65
R6373 CLK1.n1053 CLK1.n1052 4.65
R6374 CLK1.n404 CLK1.n402 4.65
R6375 CLK1.n1046 CLK1.n1045 4.65
R6376 CLK1.n1044 CLK1.n488 4.65
R6377 CLK1.n1043 CLK1.n1042 4.65
R6378 CLK1.n490 CLK1.n489 4.65
R6379 CLK1.n1036 CLK1.n1035 4.65
R6380 CLK1.n1034 CLK1.n493 4.65
R6381 CLK1.n1033 CLK1.n1032 4.65
R6382 CLK1.n497 CLK1.n496 4.65
R6383 CLK1.n1026 CLK1.n1025 4.65
R6384 CLK1.n1024 CLK1.n502 4.65
R6385 CLK1.n1023 CLK1.n1022 4.65
R6386 CLK1.n509 CLK1.n504 4.65
R6387 CLK1.n1016 CLK1.n1015 4.65
R6388 CLK1.n1014 CLK1.n508 4.65
R6389 CLK1.n1013 CLK1.n1012 4.65
R6390 CLK1.n511 CLK1.n510 4.65
R6391 CLK1.n1006 CLK1.n1005 4.65
R6392 CLK1.n1003 CLK1.n515 4.65
R6393 CLK1.n1002 CLK1.n1001 4.65
R6394 CLK1.n400 CLK1.n399 4.65
R6395 CLK1.n1065 CLK1.n398 4.65
R6396 CLK1.n1064 CLK1.n1063 4.65
R6397 CLK1.n321 CLK1.n320 4.65
R6398 CLK1.n1181 CLK1.n1180 4.65
R6399 CLK1.n1189 CLK1.n1188 4.65
R6400 CLK1.n1193 CLK1.n318 4.65
R6401 CLK1.n1195 CLK1.n1194 4.65
R6402 CLK1.n314 CLK1.n313 4.65
R6403 CLK1.n1202 CLK1.n1201 4.65
R6404 CLK1.n1203 CLK1.n312 4.65
R6405 CLK1.n1205 CLK1.n1204 4.65
R6406 CLK1.n308 CLK1.n307 4.65
R6407 CLK1.n1213 CLK1.n1212 4.65
R6408 CLK1.n1215 CLK1.n306 4.65
R6409 CLK1.n1217 CLK1.n1216 4.65
R6410 CLK1.n303 CLK1.n302 4.65
R6411 CLK1.n1224 CLK1.n1223 4.65
R6412 CLK1.n1225 CLK1.n300 4.65
R6413 CLK1.n1228 CLK1.n1227 4.65
R6414 CLK1.n1226 CLK1.n296 4.65
R6415 CLK1.n1235 CLK1.n1234 4.65
R6416 CLK1.n1236 CLK1.n294 4.65
R6417 CLK1.n1239 CLK1.n1238 4.65
R6418 CLK1.n1237 CLK1.n290 4.65
R6419 CLK1.n1246 CLK1.n1245 4.65
R6420 CLK1.n1247 CLK1.n287 4.65
R6421 CLK1.n1250 CLK1.n1249 4.65
R6422 CLK1.n1248 CLK1.n283 4.65
R6423 CLK1.n1255 CLK1.n1254 4.65
R6424 CLK1.n1323 CLK1.n1320 4.65
R6425 CLK1.n1325 CLK1.n1324 4.65
R6426 CLK1.n1316 CLK1.n1315 4.65
R6427 CLK1.n1333 CLK1.n1332 4.65
R6428 CLK1.n1335 CLK1.n1314 4.65
R6429 CLK1.n1337 CLK1.n1336 4.65
R6430 CLK1.n1311 CLK1.n1310 4.65
R6431 CLK1.n1344 CLK1.n1343 4.65
R6432 CLK1.n1345 CLK1.n1308 4.65
R6433 CLK1.n1348 CLK1.n1347 4.65
R6434 CLK1.n1346 CLK1.n1304 4.65
R6435 CLK1.n1355 CLK1.n1354 4.65
R6436 CLK1.n1356 CLK1.n1302 4.65
R6437 CLK1.n1359 CLK1.n1358 4.65
R6438 CLK1.n1357 CLK1.n1298 4.65
R6439 CLK1.n1364 CLK1.n1363 4.65
R6440 CLK1.n1366 CLK1.n1365 4.65
R6441 CLK1.n1295 CLK1.n1294 4.65
R6442 CLK1.n1371 CLK1.n1370 4.65
R6443 CLK1.n1372 CLK1.n1292 4.65
R6444 CLK1.n1375 CLK1.n1374 4.65
R6445 CLK1.n1288 CLK1.n1287 4.65
R6446 CLK1.n1382 CLK1.n1381 4.65
R6447 CLK1.n1383 CLK1.n1286 4.65
R6448 CLK1.n1386 CLK1.n1385 4.65
R6449 CLK1.n1384 CLK1.n1282 4.65
R6450 CLK1.n1393 CLK1.n1392 4.65
R6451 CLK1.n1394 CLK1.n1280 4.65
R6452 CLK1.n1398 CLK1.n1397 4.65
R6453 CLK1.n1396 CLK1.n1276 4.65
R6454 CLK1.n1406 CLK1.n1405 4.65
R6455 CLK1.n1407 CLK1.n1275 4.65
R6456 CLK1.n1410 CLK1.n1409 4.65
R6457 CLK1.n1272 CLK1.n1271 4.65
R6458 CLK1.n1417 CLK1.n1416 4.65
R6459 CLK1.n1418 CLK1.n1270 4.65
R6460 CLK1.n1420 CLK1.n1419 4.65
R6461 CLK1.n1266 CLK1.n1265 4.65
R6462 CLK1.n1427 CLK1.n1426 4.65
R6463 CLK1.n1429 CLK1.n1262 4.65
R6464 CLK1.n1432 CLK1.n1431 4.65
R6465 CLK1.n1430 CLK1.n1263 4.65
R6466 CLK1.n1177 CLK1.n392 4.633
R6467 CLK1.n1177 CLK1.n393 4.633
R6468 CLK1.n1171 CLK1.n393 4.633
R6469 CLK1.n1171 CLK1.n397 4.633
R6470 CLK1.n1166 CLK1.n397 4.633
R6471 CLK1.n1166 CLK1.n1067 4.633
R6472 CLK1.n1160 CLK1.n1067 4.633
R6473 CLK1.n1160 CLK1.n1071 4.633
R6474 CLK1.n1156 CLK1.n1071 4.633
R6475 CLK1.n1156 CLK1.n1073 4.633
R6476 CLK1.n1152 CLK1.n1073 4.633
R6477 CLK1.n1152 CLK1.n1078 4.633
R6478 CLK1.n1148 CLK1.n1078 4.633
R6479 CLK1.n1148 CLK1.n1083 4.633
R6480 CLK1.n1144 CLK1.n1083 4.633
R6481 CLK1.n1144 CLK1.n1089 4.633
R6482 CLK1.n1140 CLK1.n1089 4.633
R6483 CLK1.n1140 CLK1.n1091 4.633
R6484 CLK1.n1136 CLK1.n1091 4.633
R6485 CLK1.n1136 CLK1.n1097 4.633
R6486 CLK1.n1132 CLK1.n1097 4.633
R6487 CLK1.n1132 CLK1.n1101 4.633
R6488 CLK1.n1126 CLK1.n1101 4.633
R6489 CLK1.n1126 CLK1.n1106 4.633
R6490 CLK1.n1121 CLK1.n1106 4.633
R6491 CLK1.n1121 CLK1.n1111 4.633
R6492 CLK1.n1115 CLK1.n1111 4.633
R6493 CLK1.n996 CLK1.n994 4.527
R6494 CLK1.n807 CLK1.n624 4.5
R6495 CLK1.n992 CLK1.n809 4.5
R6496 CLK1.n1439 CLK1.n1256 4.5
R6497 CLK1.n1624 CLK1.n1441 4.5
R6498 CLK1.n1177 CLK1.n1176 4.427
R6499 CLK1.n394 CLK1.n393 4.427
R6500 CLK1.n1174 CLK1.n394 4.427
R6501 CLK1.n1172 CLK1.n1171 4.427
R6502 CLK1.n1173 CLK1.n1172 4.427
R6503 CLK1.n397 CLK1.n396 4.427
R6504 CLK1.n396 CLK1.n395 4.427
R6505 CLK1.n1166 CLK1.n1165 4.427
R6506 CLK1.n1165 CLK1.n1164 4.427
R6507 CLK1.n1068 CLK1.n1067 4.427
R6508 CLK1.n1163 CLK1.n1068 4.427
R6509 CLK1.n1161 CLK1.n1160 4.427
R6510 CLK1.n1162 CLK1.n1161 4.427
R6511 CLK1.n1071 CLK1.n1070 4.427
R6512 CLK1.n1070 CLK1.n1069 4.427
R6513 CLK1.n1156 CLK1.n1155 4.427
R6514 CLK1.n1154 CLK1.n1073 4.427
R6515 CLK1.n1153 CLK1.n1152 4.427
R6516 CLK1.n1078 CLK1.n1077 4.427
R6517 CLK1.n1148 CLK1.n1147 4.427
R6518 CLK1.n1146 CLK1.n1083 4.427
R6519 CLK1.n1145 CLK1.n1144 4.427
R6520 CLK1.n1089 CLK1.n1088 4.427
R6521 CLK1.n1140 CLK1.n1139 4.427
R6522 CLK1.n1138 CLK1.n1091 4.427
R6523 CLK1.n1137 CLK1.n1136 4.427
R6524 CLK1.n1097 CLK1.n1096 4.427
R6525 CLK1.n1103 CLK1.n1096 4.427
R6526 CLK1.n1132 CLK1.n1131 4.427
R6527 CLK1.n1131 CLK1.n1130 4.427
R6528 CLK1.n1102 CLK1.n1101 4.427
R6529 CLK1.n1129 CLK1.n1102 4.427
R6530 CLK1.n1127 CLK1.n1126 4.427
R6531 CLK1.n1128 CLK1.n1127 4.427
R6532 CLK1.n1106 CLK1.n1105 4.427
R6533 CLK1.n1105 CLK1.n1104 4.427
R6534 CLK1.n1121 CLK1.n1120 4.427
R6535 CLK1.n1120 CLK1.n1119 4.427
R6536 CLK1.n1112 CLK1.n1111 4.427
R6537 CLK1.n1118 CLK1.n1112 4.427
R6538 CLK1.n1116 CLK1.n1115 4.427
R6539 CLK1.n1155 CLK1.n1074 4.427
R6540 CLK1.n1154 CLK1.n1075 4.427
R6541 CLK1.n1153 CLK1.n1076 4.427
R6542 CLK1.n1084 CLK1.n1077 4.427
R6543 CLK1.n1147 CLK1.n1085 4.427
R6544 CLK1.n1146 CLK1.n1086 4.427
R6545 CLK1.n1145 CLK1.n1087 4.427
R6546 CLK1.n1092 CLK1.n1088 4.427
R6547 CLK1.n1139 CLK1.n1093 4.427
R6548 CLK1.n1138 CLK1.n1094 4.427
R6549 CLK1.n1137 CLK1.n1095 4.427
R6550 CLK1.t8 CLK1.n1085 4.314
R6551 CLK1.n1087 CLK1.t75 4.314
R6552 CLK1.n1183 CLK1.n321 3.715
R6553 CLK1.n1056 CLK1.n400 3.715
R6554 CLK1.n1063 CLK1.n1062 3.715
R6555 CLK1.n1188 CLK1.n319 3.715
R6556 CLK1.n809 CLK1.n808 3.635
R6557 CLK1.n1441 CLK1.n1440 3.635
R6558 CLK1.n1185 CLK1.n1184 3.635
R6559 EESPFAL_Sbox_0/CLK1 CLK1.n1626 3.578
R6560 CLK1.n1622 CLK1.n1621 3.563
R6561 CLK1.n990 CLK1.n989 3.563
R6562 CLK1.n805 CLK1.n804 3.563
R6563 CLK1.n1437 CLK1.n1436 3.563
R6564 CLK1.n1180 CLK1.n1179 3.203
R6565 CLK1.n624 CLK1.n623 3.067
R6566 CLK1.n1256 CLK1.n1255 3.067
R6567 CLK1.n1059 CLK1.n1058 3.039
R6568 CLK1.n1187 CLK1.n1185 3.038
R6569 CLK1.n997 CLK1.n996 3.033
R6570 CLK1.n1060 CLK1.n1059 2.849
R6571 CLK1.n12 CLK1.n11 2.682
R6572 CLK1.n1626 CLK1.n279 2.625
R6573 CLK1.n1183 CLK1.n1182 2.57
R6574 CLK1.n1057 CLK1.n1056 2.57
R6575 CLK1.n1062 CLK1.n1061 2.57
R6576 CLK1.n1186 CLK1.n319 2.57
R6577 EESPFAL_Sbox_0/EESPFAL_s0_0/CLK1 CLK1.n194 2.35
R6578 CLK1.n1178 CLK1.n1177 2.325
R6579 CLK1.n393 CLK1.n391 2.325
R6580 CLK1.n1171 CLK1.n1170 2.325
R6581 CLK1.n1169 CLK1.n397 2.325
R6582 CLK1.n1167 CLK1.n1166 2.325
R6583 CLK1.n1067 CLK1.n1066 2.325
R6584 CLK1.n1160 CLK1.n1159 2.325
R6585 CLK1.n1158 CLK1.n1071 2.325
R6586 CLK1.n1157 CLK1.n1156 2.325
R6587 CLK1.n1073 CLK1.n1072 2.325
R6588 CLK1.n1152 CLK1.n1151 2.325
R6589 CLK1.n1150 CLK1.n1078 2.325
R6590 CLK1.n1149 CLK1.n1148 2.325
R6591 CLK1.n1083 CLK1.n1082 2.325
R6592 CLK1.n1144 CLK1.n1143 2.325
R6593 CLK1.n1142 CLK1.n1089 2.325
R6594 CLK1.n1141 CLK1.n1140 2.325
R6595 CLK1.n1098 CLK1.n1091 2.325
R6596 CLK1.n1136 CLK1.n1135 2.325
R6597 CLK1.n1134 CLK1.n1097 2.325
R6598 CLK1.n1133 CLK1.n1132 2.325
R6599 CLK1.n1107 CLK1.n1101 2.325
R6600 CLK1.n1126 CLK1.n1125 2.325
R6601 CLK1.n1123 CLK1.n1106 2.325
R6602 CLK1.n1122 CLK1.n1121 2.325
R6603 CLK1.n1113 CLK1.n1111 2.325
R6604 CLK1.n392 CLK1.n390 2.325
R6605 CLK1.n993 CLK1.n992 2.246
R6606 CLK1.n1625 CLK1.n1624 2.246
R6607 CLK1.n991 CLK1.n520 2.246
R6608 CLK1.n1623 CLK1.n280 2.246
R6609 CLK1.n808 CLK1.n807 2.245
R6610 CLK1.n1440 CLK1.n1439 2.245
R6611 CLK1.n806 CLK1.n521 2.245
R6612 CLK1.n1438 CLK1.n281 2.245
R6613 CLK1.n1055 CLK1.n1054 2.203
R6614 CLK1.n1168 CLK1.n1065 2.203
R6615 CLK1.n1192 CLK1.n1190 2.203
R6616 CLK1.n10 CLK1.n9 1.655
R6617 CLK1.n92 CLK1.n91 1.655
R6618 CLK1.n224 CLK1.n223 1.655
R6619 CLK1.n1504 CLK1.n1503 1.655
R6620 CLK1.n1552 CLK1.n1481 1.655
R6621 CLK1.n872 CLK1.n871 1.655
R6622 CLK1.n920 CLK1.n849 1.655
R6623 CLK1.n557 CLK1.n556 1.655
R6624 CLK1.n687 CLK1.n686 1.655
R6625 CLK1.n735 CLK1.n664 1.655
R6626 CLK1.n408 CLK1.n407 1.655
R6627 CLK1.n317 CLK1.n316 1.655
R6628 CLK1.n1319 CLK1.n1318 1.655
R6629 CLK1.n1367 CLK1.n1296 1.655
R6630 CLK1.n83 CLK1.n82 1.655
R6631 CLK1.n190 CLK1.n189 1.655
R6632 CLK1.n277 CLK1.n197 1.655
R6633 CLK1.n1547 CLK1.n1484 1.655
R6634 CLK1.n1620 CLK1.n1444 1.655
R6635 CLK1.n344 CLK1.n343 1.655
R6636 CLK1.n387 CLK1.n324 1.655
R6637 CLK1.n432 CLK1.n431 1.655
R6638 CLK1.n915 CLK1.n852 1.655
R6639 CLK1.n988 CLK1.n812 1.655
R6640 CLK1.n621 CLK1.n524 1.655
R6641 CLK1.n730 CLK1.n667 1.655
R6642 CLK1.n803 CLK1.n627 1.655
R6643 CLK1.n475 CLK1.n412 1.655
R6644 CLK1.n998 CLK1.n519 1.655
R6645 CLK1.n1253 CLK1.n284 1.655
R6646 CLK1.n1362 CLK1.n1299 1.655
R6647 CLK1.n1435 CLK1.n1259 1.655
R6648 CLK1.n1621 CLK1.n1443 1.44
R6649 CLK1.n989 CLK1.n811 1.44
R6650 CLK1.n804 CLK1.n626 1.44
R6651 CLK1.n1436 CLK1.n1258 1.44
R6652 CLK1.n1115 CLK1.n1114 1.156
R6653 CLK1.n16 CLK1.n12 1.096
R6654 CLK1.n995 EESPFAL_Sbox_0/EESPFAL_s2_0/CLK1 0.912
R6655 CLK1.n994 CLK1.n993 0.705
R6656 CLK1.n1626 CLK1.n1625 0.7
R6657 CLK1.n479 CLK1.n477 0.662
R6658 CLK1.n1550 CLK1.n1549 0.637
R6659 CLK1.n918 CLK1.n917 0.637
R6660 CLK1.n733 CLK1.n732 0.637
R6661 CLK1.n1365 CLK1.n1364 0.637
R6662 CLK1.n1114 CLK1.n1113 0.631
R6663 CLK1.n1176 CLK1.n1175 0.619
R6664 CLK1.n1117 CLK1.n1116 0.618
R6665 CLK1.n90 CLK1.n88 0.6
R6666 CLK1.n390 CLK1.n389 0.532
R6667 CLK1.n1055 CLK1.n399 0.125
R6668 CLK1.n1065 CLK1.n1064 0.125
R6669 CLK1.n1180 CLK1.n320 0.125
R6670 CLK1.n1190 CLK1.n1189 0.125
R6671 CLK1.n1064 CLK1.n1060 0.12
R6672 CLK1.n1189 CLK1.n1185 0.119
R6673 CLK1.n1059 CLK1.n399 0.119
R6674 CLK1.n1184 CLK1.n320 0.119
R6675 CLK1.n25 CLK1.n21 0.1
R6676 CLK1.n29 CLK1.n25 0.1
R6677 CLK1.n33 CLK1.n29 0.1
R6678 CLK1.n42 CLK1.n38 0.1
R6679 CLK1.n46 CLK1.n42 0.1
R6680 CLK1.n47 CLK1.n46 0.1
R6681 CLK1.n56 CLK1.n52 0.1
R6682 CLK1.n60 CLK1.n56 0.1
R6683 CLK1.n69 CLK1.n65 0.1
R6684 CLK1.n73 CLK1.n69 0.1
R6685 CLK1.n77 CLK1.n73 0.1
R6686 CLK1.n81 CLK1.n77 0.1
R6687 CLK1.n85 CLK1.n81 0.1
R6688 CLK1.n94 CLK1.n90 0.1
R6689 CLK1.n98 CLK1.n94 0.1
R6690 CLK1.n102 CLK1.n98 0.1
R6691 CLK1.n111 CLK1.n107 0.1
R6692 CLK1.n115 CLK1.n111 0.1
R6693 CLK1.n119 CLK1.n115 0.1
R6694 CLK1.n123 CLK1.n119 0.1
R6695 CLK1.n127 CLK1.n123 0.1
R6696 CLK1.n136 CLK1.n132 0.1
R6697 CLK1.n140 CLK1.n136 0.1
R6698 CLK1.n141 CLK1.n140 0.1
R6699 CLK1.n150 CLK1.n146 0.1
R6700 CLK1.n154 CLK1.n150 0.1
R6701 CLK1.n163 CLK1.n159 0.1
R6702 CLK1.n167 CLK1.n163 0.1
R6703 CLK1.n171 CLK1.n167 0.1
R6704 CLK1.n175 CLK1.n171 0.1
R6705 CLK1.n179 CLK1.n175 0.1
R6706 CLK1.n188 CLK1.n184 0.1
R6707 CLK1.n192 CLK1.n188 0.1
R6708 CLK1.n194 CLK1.n192 0.1
R6709 CLK1.n229 CLK1.n228 0.1
R6710 CLK1.n229 CLK1.n220 0.1
R6711 CLK1.n237 CLK1.n220 0.1
R6712 CLK1.n238 CLK1.n237 0.1
R6713 CLK1.n240 CLK1.n238 0.1
R6714 CLK1.n249 CLK1.n214 0.1
R6715 CLK1.n250 CLK1.n249 0.1
R6716 CLK1.n251 CLK1.n250 0.1
R6717 CLK1.n259 CLK1.n208 0.1
R6718 CLK1.n260 CLK1.n259 0.1
R6719 CLK1.n262 CLK1.n202 0.1
R6720 CLK1.n270 CLK1.n202 0.1
R6721 CLK1.n271 CLK1.n270 0.1
R6722 CLK1.n273 CLK1.n195 0.1
R6723 CLK1.n279 CLK1.n195 0.1
R6724 CLK1.n1509 CLK1.n1508 0.1
R6725 CLK1.n1509 CLK1.n1500 0.1
R6726 CLK1.n1518 CLK1.n1500 0.1
R6727 CLK1.n1521 CLK1.n1520 0.1
R6728 CLK1.n1521 CLK1.n1495 0.1
R6729 CLK1.n1529 CLK1.n1495 0.1
R6730 CLK1.n1532 CLK1.n1530 0.1
R6731 CLK1.n1532 CLK1.n1531 0.1
R6732 CLK1.n1541 CLK1.n1540 0.1
R6733 CLK1.n1543 CLK1.n1541 0.1
R6734 CLK1.n1543 CLK1.n1542 0.1
R6735 CLK1.n1550 CLK1.n1479 0.1
R6736 CLK1.n1556 CLK1.n1479 0.1
R6737 CLK1.n1557 CLK1.n1556 0.1
R6738 CLK1.n1559 CLK1.n1472 0.1
R6739 CLK1.n1567 CLK1.n1472 0.1
R6740 CLK1.n1568 CLK1.n1567 0.1
R6741 CLK1.n1570 CLK1.n1568 0.1
R6742 CLK1.n1570 CLK1.n1569 0.1
R6743 CLK1.n1579 CLK1.n1578 0.1
R6744 CLK1.n1582 CLK1.n1579 0.1
R6745 CLK1.n1582 CLK1.n1581 0.1
R6746 CLK1.n1592 CLK1.n1591 0.1
R6747 CLK1.n1594 CLK1.n1592 0.1
R6748 CLK1.n1602 CLK1.n1456 0.1
R6749 CLK1.n1603 CLK1.n1602 0.1
R6750 CLK1.n1604 CLK1.n1603 0.1
R6751 CLK1.n1604 CLK1.n1450 0.1
R6752 CLK1.n1612 CLK1.n1450 0.1
R6753 CLK1.n1616 CLK1.n1614 0.1
R6754 CLK1.n1616 CLK1.n1615 0.1
R6755 CLK1.n349 CLK1.n348 0.1
R6756 CLK1.n349 CLK1.n340 0.1
R6757 CLK1.n358 CLK1.n340 0.1
R6758 CLK1.n361 CLK1.n360 0.1
R6759 CLK1.n361 CLK1.n335 0.1
R6760 CLK1.n369 CLK1.n335 0.1
R6761 CLK1.n372 CLK1.n370 0.1
R6762 CLK1.n372 CLK1.n371 0.1
R6763 CLK1.n381 CLK1.n380 0.1
R6764 CLK1.n383 CLK1.n381 0.1
R6765 CLK1.n383 CLK1.n382 0.1
R6766 CLK1.n877 CLK1.n876 0.1
R6767 CLK1.n877 CLK1.n868 0.1
R6768 CLK1.n886 CLK1.n868 0.1
R6769 CLK1.n889 CLK1.n888 0.1
R6770 CLK1.n889 CLK1.n863 0.1
R6771 CLK1.n897 CLK1.n863 0.1
R6772 CLK1.n900 CLK1.n898 0.1
R6773 CLK1.n900 CLK1.n899 0.1
R6774 CLK1.n909 CLK1.n908 0.1
R6775 CLK1.n911 CLK1.n909 0.1
R6776 CLK1.n911 CLK1.n910 0.1
R6777 CLK1.n918 CLK1.n847 0.1
R6778 CLK1.n924 CLK1.n847 0.1
R6779 CLK1.n925 CLK1.n924 0.1
R6780 CLK1.n927 CLK1.n840 0.1
R6781 CLK1.n935 CLK1.n840 0.1
R6782 CLK1.n936 CLK1.n935 0.1
R6783 CLK1.n938 CLK1.n936 0.1
R6784 CLK1.n938 CLK1.n937 0.1
R6785 CLK1.n947 CLK1.n946 0.1
R6786 CLK1.n950 CLK1.n947 0.1
R6787 CLK1.n950 CLK1.n949 0.1
R6788 CLK1.n960 CLK1.n959 0.1
R6789 CLK1.n962 CLK1.n960 0.1
R6790 CLK1.n970 CLK1.n824 0.1
R6791 CLK1.n971 CLK1.n970 0.1
R6792 CLK1.n972 CLK1.n971 0.1
R6793 CLK1.n972 CLK1.n818 0.1
R6794 CLK1.n980 CLK1.n818 0.1
R6795 CLK1.n984 CLK1.n982 0.1
R6796 CLK1.n984 CLK1.n983 0.1
R6797 CLK1.n562 CLK1.n561 0.1
R6798 CLK1.n562 CLK1.n553 0.1
R6799 CLK1.n570 CLK1.n553 0.1
R6800 CLK1.n571 CLK1.n570 0.1
R6801 CLK1.n572 CLK1.n571 0.1
R6802 CLK1.n572 CLK1.n547 0.1
R6803 CLK1.n581 CLK1.n547 0.1
R6804 CLK1.n584 CLK1.n583 0.1
R6805 CLK1.n584 CLK1.n542 0.1
R6806 CLK1.n592 CLK1.n542 0.1
R6807 CLK1.n595 CLK1.n593 0.1
R6808 CLK1.n595 CLK1.n594 0.1
R6809 CLK1.n604 CLK1.n603 0.1
R6810 CLK1.n606 CLK1.n604 0.1
R6811 CLK1.n606 CLK1.n605 0.1
R6812 CLK1.n615 CLK1.n614 0.1
R6813 CLK1.n617 CLK1.n615 0.1
R6814 CLK1.n617 CLK1.n616 0.1
R6815 CLK1.n692 CLK1.n691 0.1
R6816 CLK1.n692 CLK1.n683 0.1
R6817 CLK1.n701 CLK1.n683 0.1
R6818 CLK1.n704 CLK1.n703 0.1
R6819 CLK1.n704 CLK1.n678 0.1
R6820 CLK1.n712 CLK1.n678 0.1
R6821 CLK1.n715 CLK1.n713 0.1
R6822 CLK1.n715 CLK1.n714 0.1
R6823 CLK1.n724 CLK1.n723 0.1
R6824 CLK1.n726 CLK1.n724 0.1
R6825 CLK1.n726 CLK1.n725 0.1
R6826 CLK1.n733 CLK1.n662 0.1
R6827 CLK1.n739 CLK1.n662 0.1
R6828 CLK1.n740 CLK1.n739 0.1
R6829 CLK1.n742 CLK1.n655 0.1
R6830 CLK1.n750 CLK1.n655 0.1
R6831 CLK1.n751 CLK1.n750 0.1
R6832 CLK1.n753 CLK1.n751 0.1
R6833 CLK1.n753 CLK1.n752 0.1
R6834 CLK1.n762 CLK1.n761 0.1
R6835 CLK1.n765 CLK1.n762 0.1
R6836 CLK1.n765 CLK1.n764 0.1
R6837 CLK1.n775 CLK1.n774 0.1
R6838 CLK1.n777 CLK1.n775 0.1
R6839 CLK1.n785 CLK1.n639 0.1
R6840 CLK1.n786 CLK1.n785 0.1
R6841 CLK1.n787 CLK1.n786 0.1
R6842 CLK1.n787 CLK1.n633 0.1
R6843 CLK1.n795 CLK1.n633 0.1
R6844 CLK1.n799 CLK1.n797 0.1
R6845 CLK1.n799 CLK1.n798 0.1
R6846 CLK1.n437 CLK1.n436 0.1
R6847 CLK1.n437 CLK1.n428 0.1
R6848 CLK1.n446 CLK1.n428 0.1
R6849 CLK1.n449 CLK1.n448 0.1
R6850 CLK1.n449 CLK1.n423 0.1
R6851 CLK1.n457 CLK1.n423 0.1
R6852 CLK1.n460 CLK1.n458 0.1
R6853 CLK1.n460 CLK1.n459 0.1
R6854 CLK1.n469 CLK1.n468 0.1
R6855 CLK1.n471 CLK1.n469 0.1
R6856 CLK1.n471 CLK1.n470 0.1
R6857 CLK1.n480 CLK1.n479 0.1
R6858 CLK1.n481 CLK1.n480 0.1
R6859 CLK1.n481 CLK1.n401 0.1
R6860 CLK1.n1053 CLK1.n402 0.1
R6861 CLK1.n1045 CLK1.n402 0.1
R6862 CLK1.n1045 CLK1.n1044 0.1
R6863 CLK1.n1044 CLK1.n1043 0.1
R6864 CLK1.n1043 CLK1.n489 0.1
R6865 CLK1.n1035 CLK1.n1034 0.1
R6866 CLK1.n1034 CLK1.n1033 0.1
R6867 CLK1.n1033 CLK1.n496 0.1
R6868 CLK1.n1025 CLK1.n1024 0.1
R6869 CLK1.n1024 CLK1.n1023 0.1
R6870 CLK1.n1015 CLK1.n509 0.1
R6871 CLK1.n1015 CLK1.n1014 0.1
R6872 CLK1.n1014 CLK1.n1013 0.1
R6873 CLK1.n1013 CLK1.n510 0.1
R6874 CLK1.n1005 CLK1.n510 0.1
R6875 CLK1.n1003 CLK1.n1002 0.1
R6876 CLK1.n1002 CLK1.n517 0.1
R6877 CLK1.n1194 CLK1.n1193 0.1
R6878 CLK1.n1194 CLK1.n313 0.1
R6879 CLK1.n1202 CLK1.n313 0.1
R6880 CLK1.n1203 CLK1.n1202 0.1
R6881 CLK1.n1204 CLK1.n1203 0.1
R6882 CLK1.n1204 CLK1.n307 0.1
R6883 CLK1.n1213 CLK1.n307 0.1
R6884 CLK1.n1216 CLK1.n1215 0.1
R6885 CLK1.n1216 CLK1.n302 0.1
R6886 CLK1.n1224 CLK1.n302 0.1
R6887 CLK1.n1227 CLK1.n1225 0.1
R6888 CLK1.n1227 CLK1.n1226 0.1
R6889 CLK1.n1236 CLK1.n1235 0.1
R6890 CLK1.n1238 CLK1.n1236 0.1
R6891 CLK1.n1238 CLK1.n1237 0.1
R6892 CLK1.n1247 CLK1.n1246 0.1
R6893 CLK1.n1249 CLK1.n1247 0.1
R6894 CLK1.n1249 CLK1.n1248 0.1
R6895 CLK1.n1324 CLK1.n1323 0.1
R6896 CLK1.n1324 CLK1.n1315 0.1
R6897 CLK1.n1333 CLK1.n1315 0.1
R6898 CLK1.n1336 CLK1.n1335 0.1
R6899 CLK1.n1336 CLK1.n1310 0.1
R6900 CLK1.n1344 CLK1.n1310 0.1
R6901 CLK1.n1347 CLK1.n1345 0.1
R6902 CLK1.n1347 CLK1.n1346 0.1
R6903 CLK1.n1356 CLK1.n1355 0.1
R6904 CLK1.n1358 CLK1.n1356 0.1
R6905 CLK1.n1358 CLK1.n1357 0.1
R6906 CLK1.n1365 CLK1.n1294 0.1
R6907 CLK1.n1371 CLK1.n1294 0.1
R6908 CLK1.n1372 CLK1.n1371 0.1
R6909 CLK1.n1374 CLK1.n1287 0.1
R6910 CLK1.n1382 CLK1.n1287 0.1
R6911 CLK1.n1383 CLK1.n1382 0.1
R6912 CLK1.n1385 CLK1.n1383 0.1
R6913 CLK1.n1385 CLK1.n1384 0.1
R6914 CLK1.n1394 CLK1.n1393 0.1
R6915 CLK1.n1397 CLK1.n1394 0.1
R6916 CLK1.n1397 CLK1.n1396 0.1
R6917 CLK1.n1407 CLK1.n1406 0.1
R6918 CLK1.n1409 CLK1.n1407 0.1
R6919 CLK1.n1417 CLK1.n1271 0.1
R6920 CLK1.n1418 CLK1.n1417 0.1
R6921 CLK1.n1419 CLK1.n1418 0.1
R6922 CLK1.n1419 CLK1.n1265 0.1
R6923 CLK1.n1427 CLK1.n1265 0.1
R6924 CLK1.n1431 CLK1.n1429 0.1
R6925 CLK1.n1431 CLK1.n1430 0.1
R6926 CLK1.n995 CLK1.n517 0.094
R6927 CLK1.n1615 CLK1.n1442 0.088
R6928 CLK1.n983 CLK1.n810 0.088
R6929 CLK1.n798 CLK1.n625 0.088
R6930 CLK1.n1430 CLK1.n1257 0.088
R6931 CLK1.n21 CLK1.n17 0.087
R6932 CLK1.n272 CLK1.n271 0.087
R6933 CLK1.n1508 CLK1.n1507 0.087
R6934 CLK1.n1542 CLK1.n1482 0.087
R6935 CLK1.n348 CLK1.n347 0.087
R6936 CLK1.n382 CLK1.n322 0.087
R6937 CLK1.n876 CLK1.n875 0.087
R6938 CLK1.n910 CLK1.n850 0.087
R6939 CLK1.n605 CLK1.n529 0.087
R6940 CLK1.n691 CLK1.n690 0.087
R6941 CLK1.n725 CLK1.n665 0.087
R6942 CLK1.n436 CLK1.n435 0.087
R6943 CLK1.n470 CLK1.n410 0.087
R6944 CLK1.n1237 CLK1.n289 0.087
R6945 CLK1.n1323 CLK1.n1322 0.087
R6946 CLK1.n1357 CLK1.n1297 0.087
R6947 CLK1 EESPFAL_Sbox_0/CLK1 0.081
R6948 CLK1.n38 CLK1.n34 0.075
R6949 CLK1.n52 CLK1 0.075
R6950 CLK1.n61 CLK1.n60 0.075
R6951 CLK1.n86 CLK1.n85 0.075
R6952 CLK1.n107 CLK1.n103 0.075
R6953 CLK1.n132 CLK1.n128 0.075
R6954 CLK1.n146 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/CLK 0.075
R6955 CLK1.n155 CLK1.n154 0.075
R6956 CLK1.n180 CLK1.n179 0.075
R6957 CLK1.n228 CLK1.n227 0.075
R6958 CLK1.n239 CLK1.n214 0.075
R6959 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/CLK CLK1.n208 0.075
R6960 CLK1.n261 CLK1.n260 0.075
R6961 CLK1.n1520 CLK1.n1519 0.075
R6962 CLK1.n1530 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/CLK 0.075
R6963 CLK1.n1531 CLK1.n1488 0.075
R6964 CLK1.n1559 CLK1.n1558 0.075
R6965 CLK1.n1578 CLK1.n1466 0.075
R6966 CLK1.n1591 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/CLK 0.075
R6967 CLK1.n1594 CLK1.n1593 0.075
R6968 CLK1.n1613 CLK1.n1612 0.075
R6969 CLK1.n360 CLK1.n359 0.075
R6970 CLK1.n370 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/CLK 0.075
R6971 CLK1.n371 CLK1.n328 0.075
R6972 CLK1.n888 CLK1.n887 0.075
R6973 CLK1.n898 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/CLK 0.075
R6974 CLK1.n899 CLK1.n856 0.075
R6975 CLK1.n927 CLK1.n926 0.075
R6976 CLK1.n946 CLK1.n834 0.075
R6977 CLK1.n959 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/CLK 0.075
R6978 CLK1.n962 CLK1.n961 0.075
R6979 CLK1.n981 CLK1.n980 0.075
R6980 CLK1.n583 CLK1.n582 0.075
R6981 CLK1.n593 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/CLK 0.075
R6982 CLK1.n594 CLK1.n535 0.075
R6983 CLK1.n703 CLK1.n702 0.075
R6984 CLK1.n713 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_1/CLK 0.075
R6985 CLK1.n714 CLK1.n671 0.075
R6986 CLK1.n742 CLK1.n741 0.075
R6987 CLK1.n761 CLK1.n649 0.075
R6988 CLK1.n774 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/CLK 0.075
R6989 CLK1.n777 CLK1.n776 0.075
R6990 CLK1.n796 CLK1.n795 0.075
R6991 CLK1.n448 CLK1.n447 0.075
R6992 CLK1.n458 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/CLK 0.075
R6993 CLK1.n459 CLK1.n416 0.075
R6994 CLK1.n1054 CLK1.n1053 0.075
R6995 CLK1.n1035 CLK1.n494 0.075
R6996 CLK1.n1025 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/CLK 0.075
R6997 CLK1.n1023 CLK1.n503 0.075
R6998 CLK1.n1005 CLK1.n1004 0.075
R6999 CLK1.n1215 CLK1.n1214 0.075
R7000 CLK1.n1225 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/CLK 0.075
R7001 CLK1.n1226 CLK1.n295 0.075
R7002 CLK1.n1335 CLK1.n1334 0.075
R7003 CLK1.n1345 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/CLK 0.075
R7004 CLK1.n1346 CLK1.n1303 0.075
R7005 CLK1.n1374 CLK1.n1373 0.075
R7006 CLK1.n1393 CLK1.n1281 0.075
R7007 CLK1.n1406 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/CLK 0.075
R7008 CLK1.n1409 CLK1.n1408 0.075
R7009 CLK1.n1428 CLK1.n1427 0.075
R7010 CLK1.n561 CLK1.n560 0.062
R7011 CLK1.n616 CLK1.n522 0.062
R7012 CLK1.n1193 CLK1.n1192 0.062
R7013 CLK1.n1248 CLK1.n282 0.062
R7014 CLK1.n1178 CLK1.n391 0.041
R7015 CLK1.n1170 CLK1.n391 0.041
R7016 CLK1.n1170 CLK1.n1169 0.041
R7017 CLK1.n1167 CLK1.n1066 0.041
R7018 CLK1.n1159 CLK1.n1066 0.041
R7019 CLK1.n1159 CLK1.n1158 0.041
R7020 CLK1.n1158 CLK1.n1157 0.041
R7021 CLK1.n1157 CLK1.n1072 0.041
R7022 CLK1.n1151 CLK1.n1150 0.041
R7023 CLK1.n1150 CLK1.n1149 0.041
R7024 CLK1.n1149 CLK1.n1082 0.041
R7025 CLK1.n1143 CLK1.n1142 0.041
R7026 CLK1.n1142 CLK1.n1141 0.041
R7027 CLK1.n1135 CLK1.n1098 0.041
R7028 CLK1.n1135 CLK1.n1134 0.041
R7029 CLK1.n1134 CLK1.n1133 0.041
R7030 CLK1.n1125 CLK1.n1107 0.041
R7031 CLK1.n1123 CLK1.n1122 0.041
R7032 CLK1.n623 CLK1.n522 0.037
R7033 CLK1.n1255 CLK1.n282 0.037
R7034 CLK1.n1133 CLK1.n1100 0.036
R7035 CLK1.n624 CLK1.n521 0.034
R7036 CLK1.n1256 CLK1.n281 0.034
R7037 CLK1.n809 EESPFAL_Sbox_0/EESPFAL_s3_0/CLK1 0.032
R7038 CLK1.n1441 EESPFAL_Sbox_0/EESPFAL_s1_0/CLK1 0.032
R7039 CLK1.n1168 CLK1.n1167 0.031
R7040 CLK1.n1151 CLK1.n1079 0.031
R7041 CLK1.n1143 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/CLK 0.031
R7042 CLK1.n1141 CLK1.n1090 0.031
R7043 CLK1.n1125 CLK1.n1124 0.031
R7044 CLK1.n34 CLK1.n33 0.025
R7045 CLK1.n47 CLK1 0.025
R7046 CLK1.n65 CLK1.n61 0.025
R7047 CLK1.n88 CLK1.n86 0.025
R7048 CLK1.n103 CLK1.n102 0.025
R7049 CLK1.n128 CLK1.n127 0.025
R7050 CLK1.n141 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/CLK 0.025
R7051 CLK1.n159 CLK1.n155 0.025
R7052 CLK1.n184 CLK1.n180 0.025
R7053 CLK1.n240 CLK1.n239 0.025
R7054 CLK1.n251 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/CLK 0.025
R7055 CLK1.n262 CLK1.n261 0.025
R7056 CLK1.n1519 CLK1.n1518 0.025
R7057 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/CLK CLK1.n1529 0.025
R7058 CLK1.n1540 CLK1.n1488 0.025
R7059 CLK1.n1558 CLK1.n1557 0.025
R7060 CLK1.n1569 CLK1.n1466 0.025
R7061 CLK1.n1581 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/CLK 0.025
R7062 CLK1.n1593 CLK1.n1456 0.025
R7063 CLK1.n1614 CLK1.n1613 0.025
R7064 CLK1.n359 CLK1.n358 0.025
R7065 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/CLK CLK1.n369 0.025
R7066 CLK1.n380 CLK1.n328 0.025
R7067 CLK1.n887 CLK1.n886 0.025
R7068 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/CLK CLK1.n897 0.025
R7069 CLK1.n908 CLK1.n856 0.025
R7070 CLK1.n926 CLK1.n925 0.025
R7071 CLK1.n937 CLK1.n834 0.025
R7072 CLK1.n949 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/CLK 0.025
R7073 CLK1.n961 CLK1.n824 0.025
R7074 CLK1.n982 CLK1.n981 0.025
R7075 CLK1.n582 CLK1.n581 0.025
R7076 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/CLK CLK1.n592 0.025
R7077 CLK1.n603 CLK1.n535 0.025
R7078 CLK1.n702 CLK1.n701 0.025
R7079 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_1/CLK CLK1.n712 0.025
R7080 CLK1.n723 CLK1.n671 0.025
R7081 CLK1.n741 CLK1.n740 0.025
R7082 CLK1.n752 CLK1.n649 0.025
R7083 CLK1.n764 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/CLK 0.025
R7084 CLK1.n776 CLK1.n639 0.025
R7085 CLK1.n797 CLK1.n796 0.025
R7086 CLK1.n447 CLK1.n446 0.025
R7087 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/CLK CLK1.n457 0.025
R7088 CLK1.n468 CLK1.n416 0.025
R7089 CLK1.n1054 CLK1.n401 0.025
R7090 CLK1.n494 CLK1.n489 0.025
R7091 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/CLK CLK1.n496 0.025
R7092 CLK1.n509 CLK1.n503 0.025
R7093 CLK1.n1004 CLK1.n1003 0.025
R7094 CLK1.n1122 CLK1.n1110 0.025
R7095 CLK1.n1214 CLK1.n1213 0.025
R7096 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/CLK CLK1.n1224 0.025
R7097 CLK1.n1235 CLK1.n295 0.025
R7098 CLK1.n1334 CLK1.n1333 0.025
R7099 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/CLK CLK1.n1344 0.025
R7100 CLK1.n1355 CLK1.n1303 0.025
R7101 CLK1.n1373 CLK1.n1372 0.025
R7102 CLK1.n1384 CLK1.n1281 0.025
R7103 CLK1.n1396 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/CLK 0.025
R7104 CLK1.n1408 CLK1.n1271 0.025
R7105 CLK1.n1429 CLK1.n1428 0.025
R7106 EESPFAL_Sbox_0/EESPFAL_s2_0/CLK1 CLK1.n994 0.02
R7107 CLK1.n1179 CLK1.n390 0.02
R7108 CLK1.n1179 CLK1.n1178 0.02
R7109 CLK1.n1622 CLK1.n1442 0.018
R7110 CLK1.n990 CLK1.n810 0.018
R7111 CLK1.n805 CLK1.n625 0.018
R7112 CLK1.n1437 CLK1.n1257 0.018
R7113 CLK1.n1625 CLK1.n280 0.016
R7114 CLK1.n993 CLK1.n520 0.016
R7115 CLK1.n808 CLK1.n521 0.016
R7116 CLK1.n1440 CLK1.n281 0.016
R7117 CLK1.n806 CLK1.n805 0.015
R7118 CLK1.n1438 CLK1.n1437 0.015
R7119 CLK1.n1113 CLK1.n1110 0.015
R7120 CLK1.n1623 CLK1.n1622 0.015
R7121 CLK1.n991 CLK1.n990 0.015
R7122 CLK1.n17 CLK1.n16 0.012
R7123 CLK1.n273 CLK1.n272 0.012
R7124 CLK1.n1549 CLK1.n1482 0.012
R7125 CLK1.n389 CLK1.n322 0.012
R7126 CLK1.n917 CLK1.n850 0.012
R7127 CLK1.n614 CLK1.n529 0.012
R7128 CLK1.n732 CLK1.n665 0.012
R7129 CLK1.n477 CLK1.n410 0.012
R7130 CLK1.n1246 CLK1.n289 0.012
R7131 CLK1.n1364 CLK1.n1297 0.012
R7132 CLK1.n807 CLK1.n806 0.011
R7133 CLK1.n1439 CLK1.n1438 0.011
R7134 CLK1.n992 CLK1.n991 0.01
R7135 CLK1.n1624 CLK1.n1623 0.01
R7136 CLK1.n1169 CLK1.n1168 0.01
R7137 CLK1.n1079 CLK1.n1072 0.01
R7138 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/CLK CLK1.n1082 0.01
R7139 CLK1.n1098 CLK1.n1090 0.01
R7140 CLK1.n1124 CLK1.n1123 0.01
R7141 CLK1.n996 CLK1.n995 0.006
R7142 CLK1.n1107 CLK1.n1100 0.005
R7143 EESPFAL_Sbox_0/EESPFAL_s0_0/CLK1 CLK1 0.003
R7144 EESPFAL_Sbox_0/EESPFAL_s3_0/CLK1 CLK1.n520 0.001
R7145 EESPFAL_Sbox_0/EESPFAL_s1_0/CLK1 CLK1.n280 0.001
R7146 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t6 819.4
R7147 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t9 736.033
R7148 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t7 506.1
R7149 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 367.829
R7150 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t8 313.3
R7151 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t2 273.936
R7152 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n3 128.336
R7153 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n1 105.6
R7154 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t0 81.937
R7155 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n0 57.937
R7156 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n4 57.6
R7157 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n2 41.6
R7158 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t3 39.4
R7159 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t4 39.4
R7160 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t5 24
R7161 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t1 24
R7162 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n5 8.764
R7163 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n6 4.65
R7164 Dis3 Dis3.t6 392.5
R7165 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/Dis Dis3.t0 392.5
R7166 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/Dis Dis3.t5 392.5
R7167 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/Dis Dis3.t4 392.5
R7168 Dis3.n0 Dis3.t2 389.3
R7169 Dis3.n5 Dis3.t3 389.3
R7170 Dis3.n3 Dis3.t7 389.3
R7171 Dis3.n1 Dis3.t1 389.3
R7172 EESPFAL_Sbox_0/EESPFAL_s3_0/Dis3 Dis3.n1 297.172
R7173 Dis3.n6 Dis3.n5 285.061
R7174 Dis3.n4 Dis3.n3 284.736
R7175 Dis3.n0 Dis3 112
R7176 Dis3.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/Dis 112
R7177 Dis3.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/Dis 112
R7178 Dis3.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/Dis 112
R7179 Dis3.n7 Dis3.n0 98.399
R7180 Dis3.n4 Dis3.n2 12.126
R7181 EESPFAL_Sbox_0/EESPFAL_s1_0/Dis3 Dis3.n6 12.061
R7182 Dis3.n7 EESPFAL_Sbox_0/EESPFAL_s1_0/Dis3 8.969
R7183 EESPFAL_Sbox_0/Dis3 Dis3.n7 4.743
R7184 EESPFAL_Sbox_0/EESPFAL_s2_0/Dis3 EESPFAL_Sbox_0/EESPFAL_s3_0/Dis3 1.73
R7185 Dis3.n6 Dis3.n4 1.496
R7186 Dis3.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/Dis3 0.043
R7187 EESPFAL_Sbox_0/EESPFAL_s0_0/Dis3 EESPFAL_Sbox_0/Dis3 0.04
R7188 Dis3.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/Dis3 0.031
R7189 s1_bar.t5 s1_bar.t7 819.4
R7190 s1_bar.n4 s1_bar.t6 506.1
R7191 s1_bar.n4 s1_bar.t5 313.3
R7192 EESPFAL_Sbox_0/s1_bar s1_bar 188.523
R7193 s1_bar.n2 s1_bar.t4 181.136
R7194 s1_bar.n3 s1_bar.n0 128.334
R7195 s1_bar.n2 s1_bar.n1 57.937
R7196 s1_bar.n5 s1_bar.n3 57.6
R7197 s1_bar.n3 s1_bar.n2 41.6
R7198 s1_bar.n0 s1_bar.t2 39.4
R7199 s1_bar.n0 s1_bar.t3 39.4
R7200 s1_bar.n1 s1_bar.t0 24
R7201 s1_bar.n1 s1_bar.t1 24
R7202 s1_bar.n5 s1_bar.n4 8.764
R7203 s1_bar s1_bar.n5 4.681
R7204 EESPFAL_Sbox_0/s1_bar EESPFAL_Sbox_0/EESPFAL_s1_0/s1_bar 0.115
R7205 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/A_bar 922.56
R7206 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t9 819.4
R7207 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t7 684.833
R7208 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t6 506.1
R7209 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t8 313.3
R7210 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t5 177.936
R7211 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n0 128.334
R7212 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n2 105.6
R7213 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t0 81.939
R7214 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n1 58.265
R7215 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n4 57.6
R7216 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n3 41.6
R7217 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t4 39.4
R7218 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t2 39.4
R7219 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t3 24
R7220 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t1 24
R7221 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n5 8.764
R7222 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n6 4.65
R7223 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t17 1176.57
R7224 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t14 1176.57
R7225 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t7 1149.49
R7226 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t13 1149.49
R7227 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t18 1074.82
R7228 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t8 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t15 819.4
R7229 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n5 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t6 800.452
R7230 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n5 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t20 787.997
R7231 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t16 778.1
R7232 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t12 696.166
R7233 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t10 687.833
R7234 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t8 514.133
R7235 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/D EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t11 444.545
R7236 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t9 392.5
R7237 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t19 305.266
R7238 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/A 257.673
R7239 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A_bar 213.804
R7240 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/A_bar 195.284
R7241 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n17 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n16 192
R7242 EESPFAL_4in_XOR_0/XOR2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n10 191.68
R7243 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n8 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/D 177.673
R7244 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/B 175.745
R7245 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n5 169.6
R7246 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n11 166.734
R7247 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n10 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/A 164.48
R7248 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/A 161.673
R7249 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n3 128
R7250 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n0 128
R7251 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n15 105.6
R7252 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n17 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t0 97.939
R7253 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t5 97.937
R7254 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n14 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n13 76
R7255 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n12 73.937
R7256 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n14 57.6
R7257 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n9 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/A 39.806
R7258 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n11 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t4 39.4
R7259 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n11 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t2 39.4
R7260 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t3 24
R7261 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t1 24
R7262 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar 21.62
R7263 EESPFAL_4in_XOR_0/XOR2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n17 10.56
R7264 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n10 EESPFAL_Sbox_0/EESPFAL_s1_0/x2 4.65
R7265 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n9 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n8 4.347
R7266 EESPFAL_Sbox_0/EESPFAL_s1_0/x2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n9 3.261
R7267 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n14 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_2/OUT 3.2
R7268 EESPFAL_Sbox_0/EESPFAL_s3_0/x2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n4 3.178
R7269 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n8 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n7 2.32
R7270 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n1 2.178
R7271 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n6 1.901
R7272 EESPFAL_Sbox_0/EESPFAL_s1_0/x2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n2 1.338
R7273 EESPFAL_Sbox_0/EESPFAL_s2_0/x2 EESPFAL_Sbox_0/EESPFAL_s3_0/x2 1.192
R7274 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n1 EESPFAL_Sbox_0/x2 0.886
R7275 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/x2 0.312
R7276 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t6 819.4
R7277 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t8 736.033
R7278 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t7 514.133
R7279 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t9 305.266
R7280 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n5 192
R7281 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n1 166.734
R7282 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n6 160.887
R7283 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n4 105.6
R7284 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t0 97.937
R7285 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t2 97.937
R7286 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n2 76
R7287 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n0 73.937
R7288 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n3 57.6
R7289 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t3 39.4
R7290 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t1 39.4
R7291 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t4 24
R7292 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t5 24
R7293 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT 3.2
R7294 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t12 1271.5
R7295 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t10 1077.04
R7296 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t11 1015.9
R7297 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t21 819.4
R7298 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n5 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t14 810.772
R7299 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t17 810.772
R7300 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t7 810.772
R7301 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t13 778.1
R7302 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n5 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t6 694.566
R7303 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t18 694.566
R7304 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t8 694.566
R7305 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n18 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t9 506.1
R7306 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t20 447.076
R7307 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t16 430.966
R7308 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t19 392.5
R7309 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n18 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t15 313.3
R7310 EESPFAL_4in_XOR_0/XOR3_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n12 298.079
R7311 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n14 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t5 273.936
R7312 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/OUT_bar EESPFAL_4in_XOR_0/XOR3_bar 221.36
R7313 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 178.345
R7314 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n17 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n16 128.336
R7315 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n14 105.6
R7316 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n10 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A 103.753
R7317 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C_bar 102.947
R7318 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n14 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t1 81.937
R7319 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n4 81.6
R7320 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n8 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/A_bar 72.49
R7321 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n9 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/A 68.233
R7322 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n13 57.937
R7323 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n19 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n17 57.6
R7324 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n11 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/B_bar 55.433
R7325 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 55.433
R7326 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/B_bar 52.233
R7327 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n17 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n15 41.6
R7328 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n7 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/A 39.542
R7329 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t2 39.4
R7330 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t3 39.4
R7331 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n5 25.6
R7332 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n3 25.6
R7333 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n0 25.6
R7334 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t4 24
R7335 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t0 24
R7336 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n19 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n18 8.764
R7337 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/OUT_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n19 4.65
R7338 EESPFAL_Sbox_0/EESPFAL_s1_0/x3_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n1 4.058
R7339 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n10 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n9 4.035
R7340 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n9 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n8 3.691
R7341 EESPFAL_Sbox_0/EESPFAL_s3_0/x3_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n6 2.609
R7342 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n11 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n10 1.578
R7343 EESPFAL_Sbox_0/EESPFAL_s2_0/x3_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n7 1.142
R7344 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n2 0.932
R7345 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/x3_bar 0.848
R7346 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n11 0.794
R7347 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n1 EESPFAL_Sbox_0/x3_bar 0.346
R7348 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n7 EESPFAL_Sbox_0/EESPFAL_s3_0/x3_bar 0.242
R7349 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n8 EESPFAL_Sbox_0/EESPFAL_s2_0/x3_bar 0.075
R7350 Dis2.n6 Dis2.n4 532.126
R7351 Dis2.n19 Dis2.t3 504.5
R7352 Dis2.n17 Dis2.t14 504.5
R7353 Dis2.n11 Dis2.t17 504.5
R7354 Dis2.n9 Dis2.t2 504.5
R7355 Dis2.n7 Dis2.t1 504.5
R7356 Dis2.n5 Dis2.t16 504.5
R7357 Dis2.n0 Dis2.t7 504.5
R7358 Dis2.n19 Dis2.t19 389.3
R7359 Dis2.n17 Dis2.t8 389.3
R7360 Dis2.n15 Dis2.t15 389.3
R7361 Dis2.n14 Dis2.t12 389.3
R7362 Dis2.n11 Dis2.t13 389.3
R7363 Dis2.n9 Dis2.t9 389.3
R7364 Dis2.n7 Dis2.t6 389.3
R7365 Dis2.n5 Dis2.t21 389.3
R7366 Dis2.n4 Dis2.t5 389.3
R7367 Dis2.n3 Dis2.t10 389.3
R7368 Dis2.n2 Dis2.t11 389.3
R7369 Dis2.n1 Dis2.t18 389.3
R7370 Dis2.n22 Dis2.t0 389.3
R7371 Dis2.n21 Dis2.t4 389.3
R7372 Dis2.n0 Dis2.t20 389.3
R7373 Dis2.n16 Dis2.n15 273.536
R7374 Dis2.n24 Dis2.n23 265.28
R7375 Dis2.n18 Dis2.n16 258.592
R7376 Dis2.n13 Dis2.n12 243.072
R7377 Dis2.n12 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/Dis 177.536
R7378 Dis2.n20 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/Dis 177.216
R7379 Dis2.n18 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/Dis 177.216
R7380 Dis2.n8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/Dis 177.216
R7381 Dis2.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/Dis 177.216
R7382 Dis2.n10 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/Dis 176.896
R7383 Dis2.n13 Dis2.n2 165.061
R7384 Dis2.n24 Dis2 149.76
R7385 Dis2.n23 Dis2.n22 125.76
R7386 Dis2.n15 Dis2.n14 115.2
R7387 Dis2.n4 Dis2.n3 115.2
R7388 Dis2.n2 Dis2.n1 115.2
R7389 Dis2.n22 Dis2.n21 115.2
R7390 Dis2.n23 EESPFAL_Sbox_0/EESPFAL_s1_0/Dis2 9.259
R7391 EESPFAL_Sbox_0/Dis2 Dis2.n24 6.908
R7392 EESPFAL_Sbox_0/EESPFAL_s2_0/Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/Dis2 5.575
R7393 Dis2.n10 EESPFAL_Sbox_0/EESPFAL_s2_0/Dis2 3.357
R7394 EESPFAL_Sbox_0/EESPFAL_s1_0/Dis2 Dis2.n20 3.284
R7395 EESPFAL_Sbox_0/EESPFAL_s3_0/Dis2 Dis2.n8 3.284
R7396 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/Dis Dis2.n19 3.2
R7397 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/Dis Dis2.n17 3.2
R7398 Dis2.n14 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/Dis 3.2
R7399 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/Dis Dis2.n11 3.2
R7400 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/Dis Dis2.n9 3.2
R7401 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/Dis Dis2.n7 3.2
R7402 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/Dis Dis2.n5 3.2
R7403 Dis2.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/Dis 3.2
R7404 Dis2.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/Dis 3.2
R7405 Dis2.n21 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/Dis 3.2
R7406 Dis2 Dis2.n0 3.2
R7407 Dis2.n16 Dis2.n13 2.039
R7408 Dis2.n12 Dis2.n10 0.627
R7409 Dis2.n8 Dis2.n6 0.623
R7410 Dis2.n20 Dis2.n18 0.623
R7411 EESPFAL_Sbox_0/Dis2 Dis2 0.106
R7412 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/Dis2 0.056
R7413 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t7 1074.82
R7414 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t9 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t8 819.4
R7415 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t9 514.133
R7416 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t6 305.266
R7417 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n6 260.333
R7418 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n5 192
R7419 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n1 166.734
R7420 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n4 105.6
R7421 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t0 97.937
R7422 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t4 97.937
R7423 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n2 76
R7424 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n0 73.937
R7425 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n3 57.6
R7426 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t3 39.4
R7427 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t5 39.4
R7428 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t1 24
R7429 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t2 24
R7430 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT 3.2
R7431 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t7 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t8 819.4
R7432 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t9 736.033
R7433 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t6 506.1
R7434 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t7 313.3
R7435 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t0 273.936
R7436 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 266.318
R7437 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n3 128.336
R7438 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n1 105.6
R7439 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t4 81.937
R7440 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n0 57.937
R7441 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n4 57.6
R7442 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n2 41.6
R7443 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t1 39.4
R7444 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t2 39.4
R7445 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t3 24
R7446 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t5 24
R7447 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n5 8.764
R7448 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n6 4.65
R7449 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t13 1077.04
R7450 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t20 1077.04
R7451 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t6 1077.04
R7452 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t8 1015.9
R7453 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t16 1015.9
R7454 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t7 1015.9
R7455 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t17 912.566
R7456 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t18 881.55
R7457 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t19 819.4
R7458 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t9 778.1
R7459 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t11 604.112
R7460 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n17 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t12 506.1
R7461 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t10 479.166
R7462 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t14 392.5
R7463 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n17 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t15 313.3
R7464 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n11 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/B 293.928
R7465 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t5 273.936
R7466 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n8 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B_bar 249.673
R7467 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_1/OUT_bar EESPFAL_4in_XOR_0/XOR1_bar 220.4
R7468 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/A_bar 218.41
R7469 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/B_bar 214.153
R7470 EESPFAL_Sbox_0/EESPFAL_s3_0/x1_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/A_bar 205.61
R7471 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n9 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/A_bar 198.153
R7472 EESPFAL_4in_XOR_0/XOR1_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n11 187.688
R7473 EESPFAL_Sbox_0/EESPFAL_s3_0/x1_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_1/A_bar 183.517
R7474 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n15 128.336
R7475 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n14 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n13 105.6
R7476 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t3 81.937
R7477 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n4 81.6
R7478 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n2 81.6
R7479 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n1 81.6
R7480 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n14 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n12 57.937
R7481 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n18 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n16 57.6
R7482 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n14 41.6
R7483 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t1 39.4
R7484 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t0 39.4
R7485 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/A 38.977
R7486 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t2 24
R7487 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t4 24
R7488 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar 21.897
R7489 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n18 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n17 8.764
R7490 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n18 4.65
R7491 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/x1_bar 3.014
R7492 EESPFAL_Sbox_0/EESPFAL_s1_0/x1_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n9 2.92
R7493 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n8 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n7 2.551
R7494 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n11 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n10 2.298
R7495 EESPFAL_Sbox_0/EESPFAL_s2_0/x1_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n3 2
R7496 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n3 1.996
R7497 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n9 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n8 1.844
R7498 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n10 EESPFAL_Sbox_0/EESPFAL_s1_0/x1_bar 1.704
R7499 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n6 1.591
R7500 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n10 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n0 1.535
R7501 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/x1_bar 1.299
R7502 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n0 EESPFAL_Sbox_0/x1_bar 1.164
R7503 EESPFAL_Sbox_0/EESPFAL_s2_0/x1_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n5 0.124
R7504 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/A_bar 951.139
R7505 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t8 819.4
R7506 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t9 684.833
R7507 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t6 506.1
R7508 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t7 313.3
R7509 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t5 177.936
R7510 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n0 128.334
R7511 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n1 105.6
R7512 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t1 81.937
R7513 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n2 58.265
R7514 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n4 57.6
R7515 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n3 41.6
R7516 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t3 39.4
R7517 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t2 39.4
R7518 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t4 24
R7519 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t0 24
R7520 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n5 8.764
R7521 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n6 4.65
R7522 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t6 1271.5
R7523 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t7 1077.04
R7524 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t14 1077.04
R7525 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t19 1015.9
R7526 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t15 1015.9
R7527 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t18 833.352
R7528 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t8 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t13 819.4
R7529 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t17 810.772
R7530 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t16 778.1
R7531 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t9 736.033
R7532 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t11 694.566
R7533 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t20 506.1
R7534 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/D_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t12 495.233
R7535 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t10 392.5
R7536 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t8 313.3
R7537 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t4 273.936
R7538 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/A_bar 228.65
R7539 EESPFAL_4in_XOR_0/XOR2_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n10 227.121
R7540 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_2/OUT_bar EESPFAL_4in_XOR_0/XOR2_bar 221.04
R7541 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n9 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/A_bar 181.404
R7542 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A 174.778
R7543 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/B_bar 141.193
R7544 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n8 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/D_bar 141.193
R7545 EESPFAL_Sbox_0/EESPFAL_s1_0/x2_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/A_bar 132.65
R7546 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n14 128.334
R7547 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/A_bar 125.193
R7548 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n12 105.6
R7549 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t5 81.937
R7550 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n4 81.6
R7551 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n2 81.6
R7552 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n11 57.937
R7553 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n17 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n15 57.6
R7554 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n13 41.6
R7555 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/A 39.762
R7556 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n14 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t1 39.4
R7557 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n14 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t0 39.4
R7558 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n3 25.6
R7559 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n11 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t2 24
R7560 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n11 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t3 24
R7561 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B 21.031
R7562 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n17 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n16 8.764
R7563 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n9 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n8 4.827
R7564 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_2/OUT_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n17 4.65
R7565 EESPFAL_Sbox_0/EESPFAL_s3_0/x2_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n5 2.922
R7566 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n6 2.82
R7567 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n0 2.504
R7568 EESPFAL_Sbox_0/EESPFAL_s1_0/x2_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n9 2.061
R7569 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n8 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n7 1.803
R7570 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n10 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n1 1.487
R7571 EESPFAL_Sbox_0/EESPFAL_s2_0/x2_bar EESPFAL_Sbox_0/EESPFAL_s3_0/x2_bar 1.387
R7572 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/x2_bar 0.441
R7573 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n10 EESPFAL_Sbox_0/EESPFAL_s1_0/x2_bar 0.324
R7574 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n0 EESPFAL_Sbox_0/x2_bar 0.086
R7575 CLK2.n311 CLK2.n137 407.048
R7576 CLK2.n357 CLK2.n117 407.048
R7577 CLK2.n251 CLK2.n250 407.048
R7578 CLK2.n292 CLK2.n291 407.048
R7579 CLK2.n207 CLK2.n206 407.048
R7580 CLK2.n240 CLK2.n239 407.048
R7581 CLK2.n319 CLK2.n137 400
R7582 CLK2.n320 CLK2.n319 400
R7583 CLK2.n356 CLK2.n355 400
R7584 CLK2.n357 CLK2.n356 400
R7585 CLK2.n252 CLK2.n168 400
R7586 CLK2.n252 CLK2.n251 400
R7587 CLK2.n291 CLK2.n290 400
R7588 CLK2.n290 CLK2.n148 400
R7589 CLK2.n321 CLK2.n320 366.379
R7590 CLK2.n355 CLK2.n118 366.379
R7591 CLK2.n260 CLK2.n168 366.379
R7592 CLK2.n282 CLK2.n148 366.379
R7593 CLK2.n208 CLK2.n207 366.379
R7594 CLK2.n239 CLK2.n238 366.379
R7595 CLK2.n321 CLK2.n131 131.034
R7596 CLK2.n330 CLK2.n131 131.034
R7597 CLK2.n333 CLK2.n331 131.034
R7598 CLK2.n342 CLK2.n341 131.034
R7599 CLK2.n344 CLK2.n343 131.034
R7600 CLK2.n343 CLK2.n118 131.034
R7601 CLK2.n282 CLK2.n281 131.034
R7602 CLK2.n281 CLK2.n280 131.034
R7603 CLK2.n272 CLK2.n161 131.034
R7604 CLK2.n270 CLK2.n162 131.034
R7605 CLK2.n262 CLK2.n261 131.034
R7606 CLK2.n261 CLK2.n260 131.034
R7607 CLK2.n238 CLK2.n182 131.034
R7608 CLK2.n229 CLK2.n182 131.034
R7609 CLK2.n228 CLK2.n227 131.034
R7610 CLK2.n219 CLK2.n218 131.034
R7611 CLK2.n217 CLK2.n195 131.034
R7612 CLK2.n208 CLK2.n195 131.034
R7613 CLK2.t13 CLK2.n332 122.844
R7614 CLK2.n332 CLK2.t72 122.844
R7615 CLK2.t47 CLK2.n271 122.844
R7616 CLK2.n271 CLK2.t67 122.844
R7617 CLK2.n194 CLK2.t116 122.844
R7618 CLK2.t96 CLK2.n194 122.844
R7619 CLK2.n331 CLK2.t11 106.465
R7620 CLK2.t74 CLK2.n342 106.465
R7621 CLK2.n161 CLK2.t45 106.465
R7622 CLK2.t69 CLK2.n162 106.465
R7623 CLK2.t5 CLK2.n228 106.465
R7624 CLK2.n218 CLK2.t17 106.465
R7625 CLK2.n858 CLK2.n857 104.32
R7626 CLK2.n312 CLK2.n138 96
R7627 CLK2.n318 CLK2.n138 96
R7628 CLK2.n318 CLK2.n136 96
R7629 CLK2.n322 CLK2.n136 96
R7630 CLK2.n322 CLK2.n132 96
R7631 CLK2.n329 CLK2.n132 96
R7632 CLK2.n329 CLK2.n130 96
R7633 CLK2.n334 CLK2.n130 96
R7634 CLK2.n334 CLK2.n125 96
R7635 CLK2.n340 CLK2.n125 96
R7636 CLK2.n340 CLK2.n124 96
R7637 CLK2.n345 CLK2.n124 96
R7638 CLK2.n345 CLK2.n119 96
R7639 CLK2.n353 CLK2.n119 96
R7640 CLK2.n354 CLK2.n353 96
R7641 CLK2.n354 CLK2.n114 96
R7642 CLK2.n358 CLK2.n114 96
R7643 CLK2.n359 CLK2.n358 96
R7644 CLK2.n293 CLK2.n147 96
R7645 CLK2.n289 CLK2.n147 96
R7646 CLK2.n289 CLK2.n149 96
R7647 CLK2.n283 CLK2.n149 96
R7648 CLK2.n283 CLK2.n153 96
R7649 CLK2.n279 CLK2.n153 96
R7650 CLK2.n279 CLK2.n154 96
R7651 CLK2.n273 CLK2.n154 96
R7652 CLK2.n273 CLK2.n160 96
R7653 CLK2.n269 CLK2.n160 96
R7654 CLK2.n269 CLK2.n163 96
R7655 CLK2.n263 CLK2.n163 96
R7656 CLK2.n263 CLK2.n167 96
R7657 CLK2.n259 CLK2.n167 96
R7658 CLK2.n259 CLK2.n169 96
R7659 CLK2.n253 CLK2.n169 96
R7660 CLK2.n253 CLK2.n175 96
R7661 CLK2.n249 CLK2.n175 96
R7662 CLK2.n241 CLK2.n181 96
R7663 CLK2.n237 CLK2.n181 96
R7664 CLK2.n237 CLK2.n183 96
R7665 CLK2.n230 CLK2.n183 96
R7666 CLK2.n230 CLK2.n187 96
R7667 CLK2.n226 CLK2.n187 96
R7668 CLK2.n226 CLK2.n188 96
R7669 CLK2.n220 CLK2.n188 96
R7670 CLK2.n220 CLK2.n193 96
R7671 CLK2.n216 CLK2.n193 96
R7672 CLK2.n216 CLK2.n196 96
R7673 CLK2.n209 CLK2.n196 96
R7674 CLK2.n209 CLK2.n200 96
R7675 CLK2.n205 CLK2.n200 96
R7676 CLK2.n361 CLK2.n117 88
R7677 CLK2.n292 CLK2.n144 85.261
R7678 CLK2.n250 CLK2.n176 85.261
R7679 CLK2.n240 CLK2.n178 85.261
R7680 CLK2.n206 CLK2.n201 85.261
R7681 CLK2.n311 CLK2.n310 85.261
R7682 CLK2.n745 CLK2.t42 44.338
R7683 CLK2.n716 CLK2.t110 44.338
R7684 CLK2.n596 CLK2.t105 44.338
R7685 CLK2.n567 CLK2.t89 44.338
R7686 CLK2.n156 CLK2.t46 44.338
R7687 CLK2.n165 CLK2.t70 44.338
R7688 CLK2.n427 CLK2.t112 44.338
R7689 CLK2.n398 CLK2.t36 44.338
R7690 CLK2.n915 CLK2.t40 44.338
R7691 CLK2.n886 CLK2.t79 44.338
R7692 CLK2.n836 CLK2.t31 44.337
R7693 CLK2.n809 CLK2.t91 44.337
R7694 CLK2.n642 CLK2.t64 44.337
R7695 CLK2.n671 CLK2.t103 44.337
R7696 CLK2.n520 CLK2.t21 44.337
R7697 CLK2.n491 CLK2.t27 44.337
R7698 CLK2.n348 CLK2.t75 44.337
R7699 CLK2.n326 CLK2.t12 44.337
R7700 CLK2.n213 CLK2.t18 44.337
R7701 CLK2.n233 CLK2.t6 44.337
R7702 CLK2.n56 CLK2.t61 44.337
R7703 CLK2.n27 CLK2.t84 44.337
R7704 CLK2.n859 CLK2.t38 39.4
R7705 CLK2.n859 CLK2.t77 39.4
R7706 CLK2.n83 CLK2.t93 39.4
R7707 CLK2.n83 CLK2.t29 39.4
R7708 CLK2.n89 CLK2.t44 39.4
R7709 CLK2.n89 CLK2.t108 39.4
R7710 CLK2.n623 CLK2.t54 39.4
R7711 CLK2.n623 CLK2.t95 39.4
R7712 CLK2.n548 CLK2.t101 39.4
R7713 CLK2.n548 CLK2.t81 39.4
R7714 CLK2.n101 CLK2.t25 39.4
R7715 CLK2.n101 CLK2.t23 39.4
R7716 CLK2.n105 CLK2.t114 39.4
R7717 CLK2.n105 CLK2.t34 39.4
R7718 CLK2.n127 CLK2.t14 39.4
R7719 CLK2.n127 CLK2.t73 39.4
R7720 CLK2.n157 CLK2.t48 39.4
R7721 CLK2.n157 CLK2.t68 39.4
R7722 CLK2.n190 CLK2.t117 39.4
R7723 CLK2.n190 CLK2.t97 39.4
R7724 CLK2.n0 CLK2.t86 39.4
R7725 CLK2.n0 CLK2.t59 39.4
R7726 CLK2.n2 CLK2.t98 30.775
R7727 CLK2.n550 CLK2.t9 29.713
R7728 CLK2.n625 CLK2.t57 29.712
R7729 CLK2.n202 CLK2.t65 29.712
R7730 CLK2.n244 CLK2.t87 29.712
R7731 CLK2.n911 CLK2.t39 24.568
R7732 CLK2.n887 CLK2.t78 24.568
R7733 CLK2.n810 CLK2.t90 24.568
R7734 CLK2.n832 CLK2.t30 24.568
R7735 CLK2.n741 CLK2.t41 24.568
R7736 CLK2.n717 CLK2.t109 24.568
R7737 CLK2.n667 CLK2.t102 24.568
R7738 CLK2.n643 CLK2.t63 24.568
R7739 CLK2.n592 CLK2.t104 24.568
R7740 CLK2.n568 CLK2.t88 24.568
R7741 CLK2.n492 CLK2.t26 24.568
R7742 CLK2.n516 CLK2.t20 24.568
R7743 CLK2.n423 CLK2.t111 24.568
R7744 CLK2.n399 CLK2.t35 24.568
R7745 CLK2.t11 CLK2.n330 24.568
R7746 CLK2.n344 CLK2.t74 24.568
R7747 CLK2.n280 CLK2.t45 24.568
R7748 CLK2.n262 CLK2.t69 24.568
R7749 CLK2.n229 CLK2.t5 24.568
R7750 CLK2.t17 CLK2.n217 24.568
R7751 CLK2.n28 CLK2.t83 24.568
R7752 CLK2.n52 CLK2.t60 24.568
R7753 CLK2.n945 CLK2.t71 24
R7754 CLK2.n80 CLK2.t19 24
R7755 CLK2.n80 CLK2.t0 24
R7756 CLK2.n774 CLK2.t66 24
R7757 CLK2.n90 CLK2.t62 24
R7758 CLK2.n90 CLK2.t4 24
R7759 CLK2.n96 CLK2.t51 24
R7760 CLK2.n100 CLK2.t2 24
R7761 CLK2.n100 CLK2.t55 24
R7762 CLK2.n462 CLK2.t16 24
R7763 CLK2.n456 CLK2.t115 24
R7764 CLK2.n116 CLK2.t52 24
R7765 CLK2.n116 CLK2.t82 24
R7766 CLK2.n299 CLK2.t106 24
R7767 CLK2.n172 CLK2.t7 24
R7768 CLK2.n172 CLK2.t15 24
R7769 CLK2.n303 CLK2.t8 24
R7770 CLK2.n372 CLK2.t1 24
R7771 CLK2.n372 CLK2.t50 24
R7772 CLK2.n93 CLK2.t3 24
R7773 CLK2.n84 CLK2.t56 24
R7774 CLK2.n860 CLK2.t99 24
R7775 CLK2.n860 CLK2.t32 24
R7776 CLK2.n949 CLK2.t49 24
R7777 CLK2.n949 CLK2.t10 24
R7778 CLK2.n731 CLK2.n728 12.8
R7779 CLK2.n657 CLK2.n654 12.8
R7780 CLK2.n582 CLK2.n579 12.8
R7781 CLK2.n510 CLK2.n507 12.8
R7782 CLK2.n413 CLK2.n410 12.8
R7783 CLK2.n313 CLK2.n310 12.8
R7784 CLK2.n313 CLK2.n139 12.8
R7785 CLK2.n317 CLK2.n139 12.8
R7786 CLK2.n317 CLK2.n135 12.8
R7787 CLK2.n323 CLK2.n135 12.8
R7788 CLK2.n323 CLK2.n133 12.8
R7789 CLK2.n328 CLK2.n133 12.8
R7790 CLK2.n328 CLK2.n129 12.8
R7791 CLK2.n335 CLK2.n129 12.8
R7792 CLK2.n335 CLK2.n126 12.8
R7793 CLK2.n339 CLK2.n126 12.8
R7794 CLK2.n339 CLK2.n123 12.8
R7795 CLK2.n346 CLK2.n123 12.8
R7796 CLK2.n346 CLK2.n120 12.8
R7797 CLK2.n352 CLK2.n120 12.8
R7798 CLK2.n365 CLK2.n115 12.8
R7799 CLK2.n360 CLK2.n115 12.8
R7800 CLK2.n298 CLK2.n143 12.8
R7801 CLK2.n294 CLK2.n144 12.8
R7802 CLK2.n294 CLK2.n146 12.8
R7803 CLK2.n288 CLK2.n146 12.8
R7804 CLK2.n288 CLK2.n150 12.8
R7805 CLK2.n284 CLK2.n150 12.8
R7806 CLK2.n284 CLK2.n152 12.8
R7807 CLK2.n278 CLK2.n152 12.8
R7808 CLK2.n278 CLK2.n155 12.8
R7809 CLK2.n274 CLK2.n155 12.8
R7810 CLK2.n274 CLK2.n159 12.8
R7811 CLK2.n268 CLK2.n159 12.8
R7812 CLK2.n268 CLK2.n164 12.8
R7813 CLK2.n264 CLK2.n164 12.8
R7814 CLK2.n264 CLK2.n166 12.8
R7815 CLK2.n258 CLK2.n166 12.8
R7816 CLK2.n258 CLK2.n170 12.8
R7817 CLK2.n254 CLK2.n170 12.8
R7818 CLK2.n254 CLK2.n174 12.8
R7819 CLK2.n248 CLK2.n174 12.8
R7820 CLK2.n248 CLK2.n176 12.8
R7821 CLK2.n242 CLK2.n178 12.8
R7822 CLK2.n242 CLK2.n180 12.8
R7823 CLK2.n236 CLK2.n180 12.8
R7824 CLK2.n236 CLK2.n184 12.8
R7825 CLK2.n231 CLK2.n184 12.8
R7826 CLK2.n231 CLK2.n186 12.8
R7827 CLK2.n225 CLK2.n186 12.8
R7828 CLK2.n225 CLK2.n189 12.8
R7829 CLK2.n221 CLK2.n189 12.8
R7830 CLK2.n221 CLK2.n192 12.8
R7831 CLK2.n215 CLK2.n192 12.8
R7832 CLK2.n215 CLK2.n197 12.8
R7833 CLK2.n210 CLK2.n197 12.8
R7834 CLK2.n210 CLK2.n199 12.8
R7835 CLK2.n204 CLK2.n199 12.8
R7836 CLK2.n204 CLK2.n201 12.8
R7837 CLK2.n305 CLK2.n304 12.8
R7838 CLK2.n826 CLK2.n823 12.8
R7839 CLK2.n901 CLK2.n898 12.8
R7840 CLK2.n46 CLK2.n43 12.8
R7841 CLK2.n366 CLK2.n365 11.84
R7842 CLK2.n352 CLK2.n121 11.04
R7843 CLK2.n350 CLK2.n121 9.3
R7844 CLK2.n113 CLK2.n112 9.3
R7845 CLK2.n768 CLK2.n767 8.855
R7846 CLK2.n686 CLK2.n685 8.855
R7847 CLK2.n612 CLK2.n611 8.855
R7848 CLK2.n469 CLK2.n468 8.855
R7849 CLK2.n108 CLK2.n107 8.855
R7850 CLK2.n358 CLK2.n115 8.855
R7851 CLK2.n358 CLK2.n357 8.855
R7852 CLK2.n313 CLK2.n312 8.855
R7853 CLK2.n299 CLK2.n298 8.855
R7854 CLK2.n294 CLK2.n293 8.855
R7855 CLK2.n242 CLK2.n241 8.855
R7856 CLK2.n181 CLK2.n180 8.855
R7857 CLK2.n239 CLK2.n181 8.855
R7858 CLK2.n237 CLK2.n236 8.855
R7859 CLK2.n238 CLK2.n237 8.855
R7860 CLK2.n184 CLK2.n183 8.855
R7861 CLK2.n183 CLK2.n182 8.855
R7862 CLK2.n231 CLK2.n230 8.855
R7863 CLK2.n230 CLK2.n229 8.855
R7864 CLK2.n187 CLK2.n186 8.855
R7865 CLK2.n228 CLK2.n187 8.855
R7866 CLK2.n226 CLK2.n225 8.855
R7867 CLK2.n227 CLK2.n226 8.855
R7868 CLK2.n189 CLK2.n188 8.855
R7869 CLK2.n194 CLK2.n188 8.855
R7870 CLK2.n221 CLK2.n220 8.855
R7871 CLK2.n220 CLK2.n219 8.855
R7872 CLK2.n193 CLK2.n192 8.855
R7873 CLK2.n218 CLK2.n193 8.855
R7874 CLK2.n216 CLK2.n215 8.855
R7875 CLK2.n217 CLK2.n216 8.855
R7876 CLK2.n197 CLK2.n196 8.855
R7877 CLK2.n196 CLK2.n195 8.855
R7878 CLK2.n210 CLK2.n209 8.855
R7879 CLK2.n209 CLK2.n208 8.855
R7880 CLK2.n200 CLK2.n199 8.855
R7881 CLK2.n207 CLK2.n200 8.855
R7882 CLK2.n205 CLK2.n204 8.855
R7883 CLK2.n147 CLK2.n146 8.855
R7884 CLK2.n291 CLK2.n147 8.855
R7885 CLK2.n289 CLK2.n288 8.855
R7886 CLK2.n290 CLK2.n289 8.855
R7887 CLK2.n150 CLK2.n149 8.855
R7888 CLK2.n149 CLK2.n148 8.855
R7889 CLK2.n284 CLK2.n283 8.855
R7890 CLK2.n283 CLK2.n282 8.855
R7891 CLK2.n153 CLK2.n152 8.855
R7892 CLK2.n281 CLK2.n153 8.855
R7893 CLK2.n279 CLK2.n278 8.855
R7894 CLK2.n280 CLK2.n279 8.855
R7895 CLK2.n155 CLK2.n154 8.855
R7896 CLK2.n161 CLK2.n154 8.855
R7897 CLK2.n274 CLK2.n273 8.855
R7898 CLK2.n273 CLK2.n272 8.855
R7899 CLK2.n160 CLK2.n159 8.855
R7900 CLK2.n271 CLK2.n160 8.855
R7901 CLK2.n269 CLK2.n268 8.855
R7902 CLK2.n270 CLK2.n269 8.855
R7903 CLK2.n164 CLK2.n163 8.855
R7904 CLK2.n163 CLK2.n162 8.855
R7905 CLK2.n264 CLK2.n263 8.855
R7906 CLK2.n263 CLK2.n262 8.855
R7907 CLK2.n167 CLK2.n166 8.855
R7908 CLK2.n261 CLK2.n167 8.855
R7909 CLK2.n259 CLK2.n258 8.855
R7910 CLK2.n260 CLK2.n259 8.855
R7911 CLK2.n170 CLK2.n169 8.855
R7912 CLK2.n169 CLK2.n168 8.855
R7913 CLK2.n254 CLK2.n253 8.855
R7914 CLK2.n253 CLK2.n252 8.855
R7915 CLK2.n175 CLK2.n174 8.855
R7916 CLK2.n251 CLK2.n175 8.855
R7917 CLK2.n249 CLK2.n248 8.855
R7918 CLK2.n304 CLK2.n303 8.855
R7919 CLK2.n360 CLK2.n359 8.855
R7920 CLK2.n139 CLK2.n138 8.855
R7921 CLK2.n138 CLK2.n137 8.855
R7922 CLK2.n318 CLK2.n317 8.855
R7923 CLK2.n319 CLK2.n318 8.855
R7924 CLK2.n136 CLK2.n135 8.855
R7925 CLK2.n320 CLK2.n136 8.855
R7926 CLK2.n323 CLK2.n322 8.855
R7927 CLK2.n322 CLK2.n321 8.855
R7928 CLK2.n133 CLK2.n132 8.855
R7929 CLK2.n132 CLK2.n131 8.855
R7930 CLK2.n329 CLK2.n328 8.855
R7931 CLK2.n330 CLK2.n329 8.855
R7932 CLK2.n130 CLK2.n129 8.855
R7933 CLK2.n331 CLK2.n130 8.855
R7934 CLK2.n335 CLK2.n334 8.855
R7935 CLK2.n334 CLK2.n333 8.855
R7936 CLK2.n126 CLK2.n125 8.855
R7937 CLK2.n332 CLK2.n125 8.855
R7938 CLK2.n340 CLK2.n339 8.855
R7939 CLK2.n341 CLK2.n340 8.855
R7940 CLK2.n124 CLK2.n123 8.855
R7941 CLK2.n342 CLK2.n124 8.855
R7942 CLK2.n346 CLK2.n345 8.855
R7943 CLK2.n345 CLK2.n344 8.855
R7944 CLK2.n120 CLK2.n119 8.855
R7945 CLK2.n343 CLK2.n119 8.855
R7946 CLK2.n353 CLK2.n352 8.855
R7947 CLK2.n353 CLK2.n118 8.855
R7948 CLK2.n354 CLK2.n113 8.855
R7949 CLK2.n355 CLK2.n354 8.855
R7950 CLK2.n365 CLK2.n114 8.855
R7951 CLK2.n356 CLK2.n114 8.855
R7952 CLK2.n450 CLK2.n449 8.855
R7953 CLK2.n446 CLK2.n445 8.855
R7954 CLK2.n445 CLK2.n444 8.855
R7955 CLK2.n442 CLK2.n441 8.855
R7956 CLK2.n441 CLK2.n440 8.855
R7957 CLK2.n438 CLK2.n437 8.855
R7958 CLK2.n437 CLK2.n436 8.855
R7959 CLK2.n434 CLK2.n433 8.855
R7960 CLK2.n433 CLK2.n432 8.855
R7961 CLK2.n430 CLK2.n429 8.855
R7962 CLK2.n429 CLK2.n428 8.855
R7963 CLK2.n425 CLK2.n424 8.855
R7964 CLK2.n424 CLK2.n423 8.855
R7965 CLK2.n421 CLK2.n420 8.855
R7966 CLK2.n420 CLK2.n419 8.855
R7967 CLK2.n417 CLK2.n416 8.855
R7968 CLK2.n416 CLK2.n415 8.855
R7969 CLK2.n413 CLK2.n412 8.855
R7970 CLK2.n412 CLK2.n411 8.855
R7971 CLK2.n410 CLK2.n409 8.855
R7972 CLK2.n409 CLK2.n408 8.855
R7973 CLK2.n405 CLK2.n404 8.855
R7974 CLK2.n404 CLK2.n403 8.855
R7975 CLK2.n401 CLK2.n400 8.855
R7976 CLK2.n400 CLK2.n399 8.855
R7977 CLK2.n396 CLK2.n395 8.855
R7978 CLK2.n395 CLK2.n394 8.855
R7979 CLK2.n392 CLK2.n391 8.855
R7980 CLK2.n391 CLK2.n390 8.855
R7981 CLK2.n107 CLK2.n106 8.855
R7982 CLK2.n385 CLK2.n384 8.855
R7983 CLK2.n384 CLK2.n383 8.855
R7984 CLK2.n379 CLK2.n378 8.855
R7985 CLK2.n378 CLK2.n377 8.855
R7986 CLK2.n375 CLK2.n374 8.855
R7987 CLK2.n473 CLK2.n472 8.855
R7988 CLK2.n472 CLK2.n471 8.855
R7989 CLK2.n477 CLK2.n476 8.855
R7990 CLK2.n476 CLK2.n475 8.855
R7991 CLK2.n481 CLK2.n480 8.855
R7992 CLK2.n480 CLK2.n479 8.855
R7993 CLK2.n485 CLK2.n484 8.855
R7994 CLK2.n484 CLK2.n483 8.855
R7995 CLK2.n489 CLK2.n488 8.855
R7996 CLK2.n488 CLK2.n487 8.855
R7997 CLK2.n494 CLK2.n493 8.855
R7998 CLK2.n493 CLK2.n492 8.855
R7999 CLK2.n498 CLK2.n497 8.855
R8000 CLK2.n497 CLK2.n496 8.855
R8001 CLK2.n502 CLK2.n501 8.855
R8002 CLK2.n501 CLK2.n500 8.855
R8003 CLK2.n507 CLK2.n506 8.855
R8004 CLK2.n506 CLK2.n505 8.855
R8005 CLK2.n510 CLK2.n509 8.855
R8006 CLK2.n509 CLK2.n508 8.855
R8007 CLK2.n514 CLK2.n513 8.855
R8008 CLK2.n513 CLK2.n512 8.855
R8009 CLK2.n518 CLK2.n517 8.855
R8010 CLK2.n517 CLK2.n516 8.855
R8011 CLK2.n523 CLK2.n522 8.855
R8012 CLK2.n522 CLK2.n521 8.855
R8013 CLK2.n527 CLK2.n526 8.855
R8014 CLK2.n526 CLK2.n525 8.855
R8015 CLK2.n531 CLK2.n530 8.855
R8016 CLK2.n530 CLK2.n529 8.855
R8017 CLK2.n535 CLK2.n534 8.855
R8018 CLK2.n534 CLK2.n533 8.855
R8019 CLK2.n540 CLK2.n539 8.855
R8020 CLK2.n539 CLK2.n538 8.855
R8021 CLK2.n544 CLK2.n543 8.855
R8022 CLK2.n607 CLK2.n606 8.855
R8023 CLK2.n606 CLK2.n605 8.855
R8024 CLK2.n603 CLK2.n602 8.855
R8025 CLK2.n602 CLK2.n601 8.855
R8026 CLK2.n599 CLK2.n598 8.855
R8027 CLK2.n598 CLK2.n597 8.855
R8028 CLK2.n594 CLK2.n593 8.855
R8029 CLK2.n593 CLK2.n592 8.855
R8030 CLK2.n590 CLK2.n589 8.855
R8031 CLK2.n589 CLK2.n588 8.855
R8032 CLK2.n586 CLK2.n585 8.855
R8033 CLK2.n585 CLK2.n584 8.855
R8034 CLK2.n582 CLK2.n581 8.855
R8035 CLK2.n581 CLK2.n580 8.855
R8036 CLK2.n579 CLK2.n578 8.855
R8037 CLK2.n578 CLK2.n577 8.855
R8038 CLK2.n574 CLK2.n573 8.855
R8039 CLK2.n573 CLK2.n572 8.855
R8040 CLK2.n570 CLK2.n569 8.855
R8041 CLK2.n569 CLK2.n568 8.855
R8042 CLK2.n565 CLK2.n564 8.855
R8043 CLK2.n564 CLK2.n563 8.855
R8044 CLK2.n561 CLK2.n560 8.855
R8045 CLK2.n560 CLK2.n559 8.855
R8046 CLK2.n557 CLK2.n556 8.855
R8047 CLK2.n556 CLK2.n555 8.855
R8048 CLK2.n553 CLK2.n552 8.855
R8049 CLK2.n682 CLK2.n681 8.855
R8050 CLK2.n681 CLK2.n680 8.855
R8051 CLK2.n678 CLK2.n677 8.855
R8052 CLK2.n677 CLK2.n676 8.855
R8053 CLK2.n674 CLK2.n673 8.855
R8054 CLK2.n673 CLK2.n672 8.855
R8055 CLK2.n669 CLK2.n668 8.855
R8056 CLK2.n668 CLK2.n667 8.855
R8057 CLK2.n665 CLK2.n664 8.855
R8058 CLK2.n664 CLK2.n663 8.855
R8059 CLK2.n661 CLK2.n660 8.855
R8060 CLK2.n660 CLK2.n659 8.855
R8061 CLK2.n657 CLK2.n656 8.855
R8062 CLK2.n656 CLK2.n655 8.855
R8063 CLK2.n654 CLK2.n653 8.855
R8064 CLK2.n653 CLK2.n652 8.855
R8065 CLK2.n649 CLK2.n648 8.855
R8066 CLK2.n648 CLK2.n647 8.855
R8067 CLK2.n645 CLK2.n644 8.855
R8068 CLK2.n644 CLK2.n643 8.855
R8069 CLK2.n640 CLK2.n639 8.855
R8070 CLK2.n639 CLK2.n638 8.855
R8071 CLK2.n636 CLK2.n635 8.855
R8072 CLK2.n635 CLK2.n634 8.855
R8073 CLK2.n632 CLK2.n631 8.855
R8074 CLK2.n631 CLK2.n630 8.855
R8075 CLK2.n628 CLK2.n627 8.855
R8076 CLK2.n764 CLK2.n763 8.855
R8077 CLK2.n763 CLK2.n762 8.855
R8078 CLK2.n760 CLK2.n759 8.855
R8079 CLK2.n759 CLK2.n758 8.855
R8080 CLK2.n756 CLK2.n755 8.855
R8081 CLK2.n755 CLK2.n754 8.855
R8082 CLK2.n752 CLK2.n751 8.855
R8083 CLK2.n751 CLK2.n750 8.855
R8084 CLK2.n748 CLK2.n747 8.855
R8085 CLK2.n747 CLK2.n746 8.855
R8086 CLK2.n743 CLK2.n742 8.855
R8087 CLK2.n742 CLK2.n741 8.855
R8088 CLK2.n739 CLK2.n738 8.855
R8089 CLK2.n738 CLK2.n737 8.855
R8090 CLK2.n735 CLK2.n734 8.855
R8091 CLK2.n734 CLK2.n733 8.855
R8092 CLK2.n731 CLK2.n730 8.855
R8093 CLK2.n730 CLK2.n729 8.855
R8094 CLK2.n728 CLK2.n727 8.855
R8095 CLK2.n727 CLK2.n726 8.855
R8096 CLK2.n723 CLK2.n722 8.855
R8097 CLK2.n722 CLK2.n721 8.855
R8098 CLK2.n719 CLK2.n718 8.855
R8099 CLK2.n718 CLK2.n717 8.855
R8100 CLK2.n714 CLK2.n713 8.855
R8101 CLK2.n713 CLK2.n712 8.855
R8102 CLK2.n710 CLK2.n709 8.855
R8103 CLK2.n709 CLK2.n708 8.855
R8104 CLK2.n706 CLK2.n705 8.855
R8105 CLK2.n705 CLK2.n704 8.855
R8106 CLK2.n702 CLK2.n701 8.855
R8107 CLK2.n701 CLK2.n700 8.855
R8108 CLK2.n697 CLK2.n696 8.855
R8109 CLK2.n696 CLK2.n695 8.855
R8110 CLK2.n693 CLK2.n692 8.855
R8111 CLK2.n787 CLK2.n786 8.855
R8112 CLK2.n791 CLK2.n790 8.855
R8113 CLK2.n790 CLK2.n789 8.855
R8114 CLK2.n795 CLK2.n794 8.855
R8115 CLK2.n794 CLK2.n793 8.855
R8116 CLK2.n799 CLK2.n798 8.855
R8117 CLK2.n798 CLK2.n797 8.855
R8118 CLK2.n803 CLK2.n802 8.855
R8119 CLK2.n802 CLK2.n801 8.855
R8120 CLK2.n807 CLK2.n806 8.855
R8121 CLK2.n806 CLK2.n805 8.855
R8122 CLK2.n812 CLK2.n811 8.855
R8123 CLK2.n811 CLK2.n810 8.855
R8124 CLK2.n816 CLK2.n815 8.855
R8125 CLK2.n815 CLK2.n814 8.855
R8126 CLK2.n820 CLK2.n819 8.855
R8127 CLK2.n819 CLK2.n818 8.855
R8128 CLK2.n823 CLK2.n82 8.855
R8129 CLK2.n82 CLK2.n81 8.855
R8130 CLK2.n826 CLK2.n825 8.855
R8131 CLK2.n825 CLK2.n824 8.855
R8132 CLK2.n830 CLK2.n829 8.855
R8133 CLK2.n829 CLK2.n828 8.855
R8134 CLK2.n834 CLK2.n833 8.855
R8135 CLK2.n833 CLK2.n832 8.855
R8136 CLK2.n839 CLK2.n838 8.855
R8137 CLK2.n838 CLK2.n837 8.855
R8138 CLK2.n843 CLK2.n842 8.855
R8139 CLK2.n842 CLK2.n841 8.855
R8140 CLK2.n847 CLK2.n846 8.855
R8141 CLK2.n846 CLK2.n845 8.855
R8142 CLK2.n851 CLK2.n850 8.855
R8143 CLK2.n850 CLK2.n849 8.855
R8144 CLK2.n77 CLK2.n76 8.855
R8145 CLK2.n76 CLK2.n75 8.855
R8146 CLK2.n856 CLK2.n79 8.855
R8147 CLK2.n938 CLK2.n937 8.855
R8148 CLK2.n934 CLK2.n933 8.855
R8149 CLK2.n933 CLK2.n932 8.855
R8150 CLK2.n930 CLK2.n929 8.855
R8151 CLK2.n929 CLK2.n928 8.855
R8152 CLK2.n926 CLK2.n925 8.855
R8153 CLK2.n925 CLK2.n924 8.855
R8154 CLK2.n922 CLK2.n921 8.855
R8155 CLK2.n921 CLK2.n920 8.855
R8156 CLK2.n918 CLK2.n917 8.855
R8157 CLK2.n917 CLK2.n916 8.855
R8158 CLK2.n913 CLK2.n912 8.855
R8159 CLK2.n912 CLK2.n911 8.855
R8160 CLK2.n909 CLK2.n908 8.855
R8161 CLK2.n908 CLK2.n907 8.855
R8162 CLK2.n905 CLK2.n904 8.855
R8163 CLK2.n904 CLK2.n903 8.855
R8164 CLK2.n901 CLK2.n900 8.855
R8165 CLK2.n900 CLK2.n899 8.855
R8166 CLK2.n898 CLK2.n897 8.855
R8167 CLK2.n897 CLK2.n896 8.855
R8168 CLK2.n893 CLK2.n892 8.855
R8169 CLK2.n892 CLK2.n891 8.855
R8170 CLK2.n889 CLK2.n888 8.855
R8171 CLK2.n888 CLK2.n887 8.855
R8172 CLK2.n884 CLK2.n883 8.855
R8173 CLK2.n883 CLK2.n882 8.855
R8174 CLK2.n880 CLK2.n879 8.855
R8175 CLK2.n879 CLK2.n878 8.855
R8176 CLK2.n876 CLK2.n875 8.855
R8177 CLK2.n875 CLK2.n874 8.855
R8178 CLK2.n872 CLK2.n871 8.855
R8179 CLK2.n871 CLK2.n870 8.855
R8180 CLK2.n867 CLK2.n866 8.855
R8181 CLK2.n866 CLK2.n865 8.855
R8182 CLK2.n863 CLK2.n862 8.855
R8183 CLK2.n5 CLK2.n4 8.855
R8184 CLK2.n9 CLK2.n8 8.855
R8185 CLK2.n8 CLK2.n7 8.855
R8186 CLK2.n13 CLK2.n12 8.855
R8187 CLK2.n12 CLK2.n11 8.855
R8188 CLK2.n17 CLK2.n16 8.855
R8189 CLK2.n16 CLK2.n15 8.855
R8190 CLK2.n21 CLK2.n20 8.855
R8191 CLK2.n20 CLK2.n19 8.855
R8192 CLK2.n25 CLK2.n24 8.855
R8193 CLK2.n24 CLK2.n23 8.855
R8194 CLK2.n30 CLK2.n29 8.855
R8195 CLK2.n29 CLK2.n28 8.855
R8196 CLK2.n34 CLK2.n33 8.855
R8197 CLK2.n33 CLK2.n32 8.855
R8198 CLK2.n38 CLK2.n37 8.855
R8199 CLK2.n37 CLK2.n36 8.855
R8200 CLK2.n43 CLK2.n42 8.855
R8201 CLK2.n42 CLK2.n41 8.855
R8202 CLK2.n46 CLK2.n45 8.855
R8203 CLK2.n45 CLK2.n44 8.855
R8204 CLK2.n50 CLK2.n49 8.855
R8205 CLK2.n49 CLK2.n48 8.855
R8206 CLK2.n54 CLK2.n53 8.855
R8207 CLK2.n53 CLK2.n52 8.855
R8208 CLK2.n59 CLK2.n58 8.855
R8209 CLK2.n58 CLK2.n57 8.855
R8210 CLK2.n63 CLK2.n62 8.855
R8211 CLK2.n62 CLK2.n61 8.855
R8212 CLK2.n67 CLK2.n66 8.855
R8213 CLK2.n66 CLK2.n65 8.855
R8214 CLK2.n71 CLK2.n70 8.855
R8215 CLK2.n70 CLK2.n69 8.855
R8216 CLK2.n962 CLK2.n960 8.855
R8217 CLK2.n960 CLK2.n959 8.855
R8218 CLK2.n956 CLK2.n955 8.855
R8219 CLK2.n464 CLK2.n463 8.365
R8220 CLK2.n307 CLK2.n141 8.365
R8221 CLK2.n622 CLK2.n94 8.365
R8222 CLK2.n780 CLK2.n85 8.365
R8223 CLK2.n947 CLK2.n946 8.365
R8224 CLK2.n903 CLK2.t37 8.189
R8225 CLK2.n896 CLK2.t76 8.189
R8226 CLK2.n818 CLK2.t92 8.189
R8227 CLK2.n824 CLK2.t28 8.189
R8228 CLK2.n733 CLK2.t43 8.189
R8229 CLK2.n726 CLK2.t107 8.189
R8230 CLK2.n659 CLK2.t53 8.189
R8231 CLK2.n652 CLK2.t94 8.189
R8232 CLK2.n584 CLK2.t100 8.189
R8233 CLK2.n577 CLK2.t80 8.189
R8234 CLK2.n500 CLK2.t24 8.189
R8235 CLK2.n508 CLK2.t22 8.189
R8236 CLK2.n415 CLK2.t113 8.189
R8237 CLK2.n408 CLK2.t33 8.189
R8238 CLK2.n333 CLK2.t13 8.189
R8239 CLK2.n341 CLK2.t72 8.189
R8240 CLK2.n272 CLK2.t47 8.189
R8241 CLK2.t67 CLK2.n270 8.189
R8242 CLK2.n227 CLK2.t116 8.189
R8243 CLK2.n219 CLK2.t96 8.189
R8244 CLK2.n36 CLK2.t85 8.189
R8245 CLK2.n44 CLK2.t58 8.189
R8246 CLK2.n948 CLK2.n947 7.422
R8247 CLK2.n853 CLK2.n80 6.776
R8248 CLK2.n699 CLK2.n90 6.776
R8249 CLK2.n537 CLK2.n100 6.776
R8250 CLK2.n363 CLK2.n116 6.776
R8251 CLK2.n173 CLK2.n172 6.776
R8252 CLK2.n381 CLK2.n372 6.776
R8253 CLK2.n869 CLK2.n860 6.776
R8254 CLK2.n618 CLK2.n97 6.755
R8255 CLK2.n301 CLK2.n300 6.754
R8256 CLK2.n776 CLK2.n775 6.754
R8257 CLK2.n458 CLK2.n457 6.754
R8258 CLK2.n857 CLK2.n856 6.72
R8259 CLK2.n857 CLK2.n77 6.08
R8260 CLK2.n902 CLK2.n859 4.938
R8261 CLK2.n822 CLK2.n83 4.938
R8262 CLK2.n732 CLK2.n89 4.938
R8263 CLK2.n658 CLK2.n623 4.938
R8264 CLK2.n583 CLK2.n548 4.938
R8265 CLK2.n504 CLK2.n101 4.938
R8266 CLK2.n414 CLK2.n105 4.938
R8267 CLK2.n337 CLK2.n127 4.938
R8268 CLK2.n158 CLK2.n157 4.938
R8269 CLK2.n223 CLK2.n190 4.938
R8270 CLK2.n40 CLK2.n0 4.938
R8271 CLK2.n296 CLK2.n144 4.675
R8272 CLK2.n452 CLK2.n104 4.675
R8273 CLK2.n466 CLK2.n465 4.675
R8274 CLK2.n770 CLK2.n88 4.675
R8275 CLK2.n940 CLK2.n858 4.675
R8276 CLK2.n2 CLK2.n1 4.675
R8277 CLK2.n202 CLK2.n201 4.662
R8278 CLK2.n614 CLK2.n99 4.662
R8279 CLK2.n550 CLK2.n549 4.662
R8280 CLK2.n625 CLK2.n624 4.662
R8281 CLK2.n243 CLK2.n242 4.65
R8282 CLK2.n180 CLK2.n179 4.65
R8283 CLK2.n236 CLK2.n235 4.65
R8284 CLK2.n234 CLK2.n184 4.65
R8285 CLK2.n232 CLK2.n231 4.65
R8286 CLK2.n186 CLK2.n185 4.65
R8287 CLK2.n225 CLK2.n224 4.65
R8288 CLK2.n223 CLK2.n189 4.65
R8289 CLK2.n222 CLK2.n221 4.65
R8290 CLK2.n192 CLK2.n191 4.65
R8291 CLK2.n215 CLK2.n214 4.65
R8292 CLK2.n212 CLK2.n197 4.65
R8293 CLK2.n211 CLK2.n210 4.65
R8294 CLK2.n199 CLK2.n198 4.65
R8295 CLK2.n204 CLK2.n203 4.65
R8296 CLK2.n245 CLK2.n178 4.65
R8297 CLK2.n246 CLK2.n176 4.65
R8298 CLK2.n295 CLK2.n294 4.65
R8299 CLK2.n146 CLK2.n145 4.65
R8300 CLK2.n288 CLK2.n287 4.65
R8301 CLK2.n286 CLK2.n150 4.65
R8302 CLK2.n285 CLK2.n284 4.65
R8303 CLK2.n152 CLK2.n151 4.65
R8304 CLK2.n278 CLK2.n277 4.65
R8305 CLK2.n276 CLK2.n155 4.65
R8306 CLK2.n275 CLK2.n274 4.65
R8307 CLK2.n159 CLK2.n158 4.65
R8308 CLK2.n268 CLK2.n267 4.65
R8309 CLK2.n266 CLK2.n164 4.65
R8310 CLK2.n265 CLK2.n264 4.65
R8311 CLK2.n171 CLK2.n166 4.65
R8312 CLK2.n258 CLK2.n257 4.65
R8313 CLK2.n256 CLK2.n170 4.65
R8314 CLK2.n255 CLK2.n254 4.65
R8315 CLK2.n177 CLK2.n174 4.65
R8316 CLK2.n248 CLK2.n247 4.65
R8317 CLK2.n143 CLK2.n142 4.65
R8318 CLK2.n298 CLK2.n297 4.65
R8319 CLK2.n306 CLK2.n305 4.65
R8320 CLK2.n314 CLK2.n313 4.65
R8321 CLK2.n362 CLK2.n115 4.65
R8322 CLK2.n315 CLK2.n139 4.65
R8323 CLK2.n317 CLK2.n316 4.65
R8324 CLK2.n135 CLK2.n134 4.65
R8325 CLK2.n324 CLK2.n323 4.65
R8326 CLK2.n325 CLK2.n133 4.65
R8327 CLK2.n328 CLK2.n327 4.65
R8328 CLK2.n129 CLK2.n128 4.65
R8329 CLK2.n336 CLK2.n335 4.65
R8330 CLK2.n337 CLK2.n126 4.65
R8331 CLK2.n339 CLK2.n338 4.65
R8332 CLK2.n123 CLK2.n122 4.65
R8333 CLK2.n347 CLK2.n346 4.65
R8334 CLK2.n349 CLK2.n120 4.65
R8335 CLK2.n352 CLK2.n351 4.65
R8336 CLK2.n365 CLK2.n364 4.65
R8337 CLK2.n389 CLK2.n108 4.65
R8338 CLK2.n451 CLK2.n450 4.65
R8339 CLK2.n447 CLK2.n446 4.65
R8340 CLK2.n443 CLK2.n442 4.65
R8341 CLK2.n439 CLK2.n438 4.65
R8342 CLK2.n435 CLK2.n434 4.65
R8343 CLK2.n431 CLK2.n430 4.65
R8344 CLK2.n426 CLK2.n425 4.65
R8345 CLK2.n422 CLK2.n421 4.65
R8346 CLK2.n418 CLK2.n417 4.65
R8347 CLK2.n414 CLK2.n413 4.65
R8348 CLK2.n410 CLK2.n407 4.65
R8349 CLK2.n406 CLK2.n405 4.65
R8350 CLK2.n402 CLK2.n401 4.65
R8351 CLK2.n397 CLK2.n396 4.65
R8352 CLK2.n393 CLK2.n392 4.65
R8353 CLK2.n380 CLK2.n379 4.65
R8354 CLK2.n455 CLK2.n103 4.65
R8355 CLK2.n454 CLK2.n453 4.65
R8356 CLK2.n461 CLK2.n460 4.65
R8357 CLK2.n547 CLK2.n546 4.65
R8358 CLK2.n470 CLK2.n469 4.65
R8359 CLK2.n474 CLK2.n473 4.65
R8360 CLK2.n478 CLK2.n477 4.65
R8361 CLK2.n482 CLK2.n481 4.65
R8362 CLK2.n486 CLK2.n485 4.65
R8363 CLK2.n490 CLK2.n489 4.65
R8364 CLK2.n495 CLK2.n494 4.65
R8365 CLK2.n499 CLK2.n498 4.65
R8366 CLK2.n503 CLK2.n502 4.65
R8367 CLK2.n507 CLK2.n504 4.65
R8368 CLK2.n511 CLK2.n510 4.65
R8369 CLK2.n515 CLK2.n514 4.65
R8370 CLK2.n519 CLK2.n518 4.65
R8371 CLK2.n524 CLK2.n523 4.65
R8372 CLK2.n528 CLK2.n527 4.65
R8373 CLK2.n532 CLK2.n531 4.65
R8374 CLK2.n536 CLK2.n535 4.65
R8375 CLK2.n541 CLK2.n540 4.65
R8376 CLK2.n545 CLK2.n544 4.65
R8377 CLK2.n613 CLK2.n612 4.65
R8378 CLK2.n608 CLK2.n607 4.65
R8379 CLK2.n604 CLK2.n603 4.65
R8380 CLK2.n600 CLK2.n599 4.65
R8381 CLK2.n595 CLK2.n594 4.65
R8382 CLK2.n591 CLK2.n590 4.65
R8383 CLK2.n587 CLK2.n586 4.65
R8384 CLK2.n583 CLK2.n582 4.65
R8385 CLK2.n579 CLK2.n576 4.65
R8386 CLK2.n575 CLK2.n574 4.65
R8387 CLK2.n571 CLK2.n570 4.65
R8388 CLK2.n566 CLK2.n565 4.65
R8389 CLK2.n562 CLK2.n561 4.65
R8390 CLK2.n558 CLK2.n557 4.65
R8391 CLK2.n554 CLK2.n553 4.65
R8392 CLK2.n617 CLK2.n98 4.65
R8393 CLK2.n616 CLK2.n615 4.65
R8394 CLK2.n621 CLK2.n620 4.65
R8395 CLK2.n687 CLK2.n686 4.65
R8396 CLK2.n683 CLK2.n682 4.65
R8397 CLK2.n679 CLK2.n678 4.65
R8398 CLK2.n675 CLK2.n674 4.65
R8399 CLK2.n670 CLK2.n669 4.65
R8400 CLK2.n666 CLK2.n665 4.65
R8401 CLK2.n662 CLK2.n661 4.65
R8402 CLK2.n658 CLK2.n657 4.65
R8403 CLK2.n654 CLK2.n651 4.65
R8404 CLK2.n650 CLK2.n649 4.65
R8405 CLK2.n646 CLK2.n645 4.65
R8406 CLK2.n641 CLK2.n640 4.65
R8407 CLK2.n637 CLK2.n636 4.65
R8408 CLK2.n633 CLK2.n632 4.65
R8409 CLK2.n629 CLK2.n628 4.65
R8410 CLK2.n689 CLK2.n92 4.65
R8411 CLK2.n690 CLK2.n91 4.65
R8412 CLK2.n769 CLK2.n768 4.65
R8413 CLK2.n765 CLK2.n764 4.65
R8414 CLK2.n761 CLK2.n760 4.65
R8415 CLK2.n757 CLK2.n756 4.65
R8416 CLK2.n753 CLK2.n752 4.65
R8417 CLK2.n749 CLK2.n748 4.65
R8418 CLK2.n744 CLK2.n743 4.65
R8419 CLK2.n740 CLK2.n739 4.65
R8420 CLK2.n736 CLK2.n735 4.65
R8421 CLK2.n732 CLK2.n731 4.65
R8422 CLK2.n728 CLK2.n725 4.65
R8423 CLK2.n724 CLK2.n723 4.65
R8424 CLK2.n720 CLK2.n719 4.65
R8425 CLK2.n715 CLK2.n714 4.65
R8426 CLK2.n711 CLK2.n710 4.65
R8427 CLK2.n707 CLK2.n706 4.65
R8428 CLK2.n703 CLK2.n702 4.65
R8429 CLK2.n698 CLK2.n697 4.65
R8430 CLK2.n694 CLK2.n693 4.65
R8431 CLK2.n773 CLK2.n87 4.65
R8432 CLK2.n772 CLK2.n771 4.65
R8433 CLK2.n779 CLK2.n778 4.65
R8434 CLK2.n788 CLK2.n787 4.65
R8435 CLK2.n792 CLK2.n791 4.65
R8436 CLK2.n796 CLK2.n795 4.65
R8437 CLK2.n800 CLK2.n799 4.65
R8438 CLK2.n804 CLK2.n803 4.65
R8439 CLK2.n808 CLK2.n807 4.65
R8440 CLK2.n813 CLK2.n812 4.65
R8441 CLK2.n817 CLK2.n816 4.65
R8442 CLK2.n821 CLK2.n820 4.65
R8443 CLK2.n823 CLK2.n822 4.65
R8444 CLK2.n827 CLK2.n826 4.65
R8445 CLK2.n831 CLK2.n830 4.65
R8446 CLK2.n835 CLK2.n834 4.65
R8447 CLK2.n840 CLK2.n839 4.65
R8448 CLK2.n844 CLK2.n843 4.65
R8449 CLK2.n848 CLK2.n847 4.65
R8450 CLK2.n852 CLK2.n851 4.65
R8451 CLK2.n939 CLK2.n938 4.65
R8452 CLK2.n935 CLK2.n934 4.65
R8453 CLK2.n931 CLK2.n930 4.65
R8454 CLK2.n927 CLK2.n926 4.65
R8455 CLK2.n923 CLK2.n922 4.65
R8456 CLK2.n919 CLK2.n918 4.65
R8457 CLK2.n914 CLK2.n913 4.65
R8458 CLK2.n910 CLK2.n909 4.65
R8459 CLK2.n906 CLK2.n905 4.65
R8460 CLK2.n902 CLK2.n901 4.65
R8461 CLK2.n898 CLK2.n895 4.65
R8462 CLK2.n894 CLK2.n893 4.65
R8463 CLK2.n890 CLK2.n889 4.65
R8464 CLK2.n885 CLK2.n884 4.65
R8465 CLK2.n881 CLK2.n880 4.65
R8466 CLK2.n877 CLK2.n876 4.65
R8467 CLK2.n873 CLK2.n872 4.65
R8468 CLK2.n868 CLK2.n867 4.65
R8469 CLK2.n944 CLK2.n943 4.65
R8470 CLK2.n942 CLK2.n941 4.65
R8471 CLK2.n953 CLK2.n74 4.65
R8472 CLK2.n952 CLK2.n951 4.65
R8473 CLK2.n6 CLK2.n5 4.65
R8474 CLK2.n10 CLK2.n9 4.65
R8475 CLK2.n14 CLK2.n13 4.65
R8476 CLK2.n18 CLK2.n17 4.65
R8477 CLK2.n22 CLK2.n21 4.65
R8478 CLK2.n26 CLK2.n25 4.65
R8479 CLK2.n31 CLK2.n30 4.65
R8480 CLK2.n35 CLK2.n34 4.65
R8481 CLK2.n39 CLK2.n38 4.65
R8482 CLK2.n43 CLK2.n40 4.65
R8483 CLK2.n47 CLK2.n46 4.65
R8484 CLK2.n51 CLK2.n50 4.65
R8485 CLK2.n55 CLK2.n54 4.65
R8486 CLK2.n60 CLK2.n59 4.65
R8487 CLK2.n64 CLK2.n63 4.65
R8488 CLK2.n68 CLK2.n67 4.65
R8489 CLK2.n72 CLK2.n71 4.65
R8490 EESPFAL_Sbox_0/CLK2 CLK2.n964 4.529
R8491 CLK2.n784 EESPFAL_Sbox_0/EESPFAL_s1_0/CLK2 4.509
R8492 EESPFAL_Sbox_0/EESPFAL_s3_0/CLK2 CLK2.n140 4.509
R8493 CLK2.n367 CLK2.n366 4.5
R8494 CLK2.n369 CLK2.n111 4.5
R8495 CLK2.n300 CLK2.n143 3.715
R8496 CLK2.n305 CLK2.n141 3.715
R8497 CLK2.n951 CLK2.n950 3.715
R8498 CLK2.n304 CLK2.n302 3.039
R8499 CLK2.n619 CLK2.n95 3.039
R8500 CLK2.n777 CLK2.n86 3.039
R8501 CLK2.n459 CLK2.n102 3.039
R8502 CLK2.n310 CLK2.n309 3.033
R8503 CLK2.n386 CLK2.n385 3.033
R8504 CLK2.n783 CLK2.n782 3.033
R8505 CLK2.n963 CLK2.n962 3.033
R8506 CLK2.n962 CLK2.n961 2.72
R8507 CLK2.n361 CLK2.n360 2.682
R8508 CLK2.n376 CLK2.n375 2.682
R8509 CLK2.n856 CLK2.n855 2.682
R8510 CLK2.n864 CLK2.n863 2.682
R8511 CLK2.n957 CLK2.n956 2.682
R8512 CLK2.n619 CLK2.n618 2.6
R8513 CLK2.n775 CLK2.n774 2.57
R8514 CLK2.n97 CLK2.n96 2.57
R8515 CLK2.n463 CLK2.n462 2.57
R8516 CLK2.n457 CLK2.n456 2.57
R8517 CLK2.n300 CLK2.n299 2.57
R8518 CLK2.n303 CLK2.n141 2.57
R8519 CLK2.n94 CLK2.n93 2.57
R8520 CLK2.n85 CLK2.n84 2.57
R8521 CLK2.n946 CLK2.n945 2.57
R8522 CLK2.n950 CLK2.n949 2.57
R8523 CLK2.n370 CLK2.n110 2.251
R8524 CLK2.n369 CLK2.n368 2.246
R8525 CLK2.n965 CLK2.n73 2.246
R8526 CLK2.n459 CLK2.n458 2.224
R8527 CLK2.n302 CLK2.n301 2.224
R8528 CLK2.n777 CLK2.n776 2.224
R8529 CLK2.n297 CLK2.n296 2.203
R8530 CLK2.n308 CLK2.n307 2.203
R8531 CLK2.n454 CLK2.n452 2.203
R8532 CLK2.n466 CLK2.n464 2.203
R8533 CLK2.n772 CLK2.n770 2.203
R8534 CLK2.n781 CLK2.n780 2.203
R8535 CLK2.n942 CLK2.n940 2.203
R8536 CLK2.n964 CLK2.n953 2.203
R8537 CLK2.n121 CLK2.n113 1.76
R8538 CLK2.n79 CLK2.n78 1.656
R8539 CLK2.n449 CLK2.n448 1.655
R8540 CLK2.n4 CLK2.n3 1.655
R8541 CLK2.n767 CLK2.n766 1.655
R8542 CLK2.n685 CLK2.n684 1.655
R8543 CLK2.n611 CLK2.n610 1.655
R8544 CLK2.n468 CLK2.n467 1.655
R8545 CLK2.n312 CLK2.n311 1.655
R8546 CLK2.n293 CLK2.n292 1.655
R8547 CLK2.n241 CLK2.n240 1.655
R8548 CLK2.n206 CLK2.n205 1.655
R8549 CLK2.n250 CLK2.n249 1.655
R8550 CLK2.n359 CLK2.n117 1.655
R8551 CLK2.n374 CLK2.n373 1.655
R8552 CLK2.n543 CLK2.n542 1.655
R8553 CLK2.n552 CLK2.n551 1.655
R8554 CLK2.n627 CLK2.n626 1.655
R8555 CLK2.n692 CLK2.n691 1.655
R8556 CLK2.n786 CLK2.n785 1.655
R8557 CLK2.n937 CLK2.n936 1.655
R8558 CLK2.n862 CLK2.n861 1.655
R8559 CLK2.n955 CLK2.n954 1.655
R8560 CLK2.n387 CLK2.n371 1.497
R8561 CLK2.n616 CLK2.n614 1.14
R8562 CLK2.n688 CLK2.n622 1.14
R8563 CLK2.n362 CLK2.n361 1.095
R8564 CLK2.n380 CLK2.n376 1.095
R8565 CLK2.n855 CLK2.n854 1.095
R8566 CLK2.n868 CLK2.n864 1.095
R8567 CLK2.n958 CLK2.n957 1.073
R8568 CLK2.n246 CLK2.n245 1.047
R8569 CLK2.n690 CLK2.n689 1.047
R8570 CLK2.n609 CLK2.n547 1.046
R8571 CLK2.n366 CLK2.n113 0.96
R8572 EESPFAL_Sbox_0/EESPFAL_s1_0/CLK2 CLK2.n783 0.928
R8573 CLK2.n309 EESPFAL_Sbox_0/EESPFAL_s3_0/CLK2 0.927
R8574 EESPFAL_Sbox_0/EESPFAL_s2_0/CLK2 CLK2.n370 0.648
R8575 CLK2.n297 CLK2.n142 0.125
R8576 CLK2.n307 CLK2.n306 0.125
R8577 CLK2.n455 CLK2.n454 0.125
R8578 CLK2.n464 CLK2.n461 0.125
R8579 CLK2.n617 CLK2.n616 0.125
R8580 CLK2.n622 CLK2.n621 0.125
R8581 CLK2.n773 CLK2.n772 0.125
R8582 CLK2.n780 CLK2.n779 0.125
R8583 CLK2.n944 CLK2.n942 0.125
R8584 CLK2.n953 CLK2.n952 0.125
R8585 CLK2.n952 CLK2.n948 0.125
R8586 CLK2.n306 CLK2.n302 0.12
R8587 CLK2.n621 CLK2.n619 0.12
R8588 CLK2.n779 CLK2.n777 0.12
R8589 CLK2.n461 CLK2.n459 0.119
R8590 CLK2.n618 CLK2.n617 0.119
R8591 CLK2.n301 CLK2.n142 0.119
R8592 CLK2.n776 CLK2.n773 0.119
R8593 CLK2.n458 CLK2.n455 0.117
R8594 CLK2.n243 CLK2.n179 0.1
R8595 CLK2.n235 CLK2.n179 0.1
R8596 CLK2.n235 CLK2.n234 0.1
R8597 CLK2.n232 CLK2.n185 0.1
R8598 CLK2.n224 CLK2.n185 0.1
R8599 CLK2.n224 CLK2.n223 0.1
R8600 CLK2.n222 CLK2.n191 0.1
R8601 CLK2.n214 CLK2.n191 0.1
R8602 CLK2.n212 CLK2.n211 0.1
R8603 CLK2.n211 CLK2.n198 0.1
R8604 CLK2.n203 CLK2.n198 0.1
R8605 CLK2.n295 CLK2.n145 0.1
R8606 CLK2.n287 CLK2.n145 0.1
R8607 CLK2.n287 CLK2.n286 0.1
R8608 CLK2.n286 CLK2.n285 0.1
R8609 CLK2.n285 CLK2.n151 0.1
R8610 CLK2.n277 CLK2.n276 0.1
R8611 CLK2.n276 CLK2.n275 0.1
R8612 CLK2.n275 CLK2.n158 0.1
R8613 CLK2.n267 CLK2.n266 0.1
R8614 CLK2.n266 CLK2.n265 0.1
R8615 CLK2.n257 CLK2.n171 0.1
R8616 CLK2.n257 CLK2.n256 0.1
R8617 CLK2.n256 CLK2.n255 0.1
R8618 CLK2.n247 CLK2.n177 0.1
R8619 CLK2.n247 CLK2.n246 0.1
R8620 CLK2.n315 CLK2.n314 0.1
R8621 CLK2.n316 CLK2.n315 0.1
R8622 CLK2.n316 CLK2.n134 0.1
R8623 CLK2.n324 CLK2.n134 0.1
R8624 CLK2.n325 CLK2.n324 0.1
R8625 CLK2.n327 CLK2.n128 0.1
R8626 CLK2.n336 CLK2.n128 0.1
R8627 CLK2.n337 CLK2.n336 0.1
R8628 CLK2.n338 CLK2.n122 0.1
R8629 CLK2.n347 CLK2.n122 0.1
R8630 CLK2.n351 CLK2.n349 0.1
R8631 CLK2.n451 CLK2.n447 0.1
R8632 CLK2.n447 CLK2.n443 0.1
R8633 CLK2.n443 CLK2.n439 0.1
R8634 CLK2.n439 CLK2.n435 0.1
R8635 CLK2.n435 CLK2.n431 0.1
R8636 CLK2.n426 CLK2.n422 0.1
R8637 CLK2.n422 CLK2.n418 0.1
R8638 CLK2.n418 CLK2.n414 0.1
R8639 CLK2.n407 CLK2.n406 0.1
R8640 CLK2.n406 CLK2.n402 0.1
R8641 CLK2.n397 CLK2.n393 0.1
R8642 CLK2.n393 CLK2.n389 0.1
R8643 CLK2.n474 CLK2.n470 0.1
R8644 CLK2.n478 CLK2.n474 0.1
R8645 CLK2.n482 CLK2.n478 0.1
R8646 CLK2.n486 CLK2.n482 0.1
R8647 CLK2.n490 CLK2.n486 0.1
R8648 CLK2.n499 CLK2.n495 0.1
R8649 CLK2.n503 CLK2.n499 0.1
R8650 CLK2.n504 CLK2.n503 0.1
R8651 CLK2.n515 CLK2.n511 0.1
R8652 CLK2.n519 CLK2.n515 0.1
R8653 CLK2.n528 CLK2.n524 0.1
R8654 CLK2.n532 CLK2.n528 0.1
R8655 CLK2.n536 CLK2.n532 0.1
R8656 CLK2.n545 CLK2.n541 0.1
R8657 CLK2.n547 CLK2.n545 0.1
R8658 CLK2.n608 CLK2.n604 0.1
R8659 CLK2.n604 CLK2.n600 0.1
R8660 CLK2.n595 CLK2.n591 0.1
R8661 CLK2.n591 CLK2.n587 0.1
R8662 CLK2.n587 CLK2.n583 0.1
R8663 CLK2.n576 CLK2.n575 0.1
R8664 CLK2.n575 CLK2.n571 0.1
R8665 CLK2.n566 CLK2.n562 0.1
R8666 CLK2.n562 CLK2.n558 0.1
R8667 CLK2.n558 CLK2.n554 0.1
R8668 CLK2.n687 CLK2.n683 0.1
R8669 CLK2.n683 CLK2.n679 0.1
R8670 CLK2.n679 CLK2.n675 0.1
R8671 CLK2.n670 CLK2.n666 0.1
R8672 CLK2.n666 CLK2.n662 0.1
R8673 CLK2.n662 CLK2.n658 0.1
R8674 CLK2.n651 CLK2.n650 0.1
R8675 CLK2.n650 CLK2.n646 0.1
R8676 CLK2.n641 CLK2.n637 0.1
R8677 CLK2.n637 CLK2.n633 0.1
R8678 CLK2.n633 CLK2.n629 0.1
R8679 CLK2.n769 CLK2.n765 0.1
R8680 CLK2.n765 CLK2.n761 0.1
R8681 CLK2.n761 CLK2.n757 0.1
R8682 CLK2.n757 CLK2.n753 0.1
R8683 CLK2.n753 CLK2.n749 0.1
R8684 CLK2.n744 CLK2.n740 0.1
R8685 CLK2.n740 CLK2.n736 0.1
R8686 CLK2.n736 CLK2.n732 0.1
R8687 CLK2.n725 CLK2.n724 0.1
R8688 CLK2.n724 CLK2.n720 0.1
R8689 CLK2.n715 CLK2.n711 0.1
R8690 CLK2.n711 CLK2.n707 0.1
R8691 CLK2.n707 CLK2.n703 0.1
R8692 CLK2.n698 CLK2.n694 0.1
R8693 CLK2.n694 CLK2.n690 0.1
R8694 CLK2.n792 CLK2.n788 0.1
R8695 CLK2.n796 CLK2.n792 0.1
R8696 CLK2.n800 CLK2.n796 0.1
R8697 CLK2.n804 CLK2.n800 0.1
R8698 CLK2.n808 CLK2.n804 0.1
R8699 CLK2.n817 CLK2.n813 0.1
R8700 CLK2.n821 CLK2.n817 0.1
R8701 CLK2.n822 CLK2.n821 0.1
R8702 CLK2.n831 CLK2.n827 0.1
R8703 CLK2.n835 CLK2.n831 0.1
R8704 CLK2.n844 CLK2.n840 0.1
R8705 CLK2.n848 CLK2.n844 0.1
R8706 CLK2.n852 CLK2.n848 0.1
R8707 CLK2.n939 CLK2.n935 0.1
R8708 CLK2.n935 CLK2.n931 0.1
R8709 CLK2.n931 CLK2.n927 0.1
R8710 CLK2.n927 CLK2.n923 0.1
R8711 CLK2.n923 CLK2.n919 0.1
R8712 CLK2.n914 CLK2.n910 0.1
R8713 CLK2.n910 CLK2.n906 0.1
R8714 CLK2.n906 CLK2.n902 0.1
R8715 CLK2.n895 CLK2.n894 0.1
R8716 CLK2.n894 CLK2.n890 0.1
R8717 CLK2.n885 CLK2.n881 0.1
R8718 CLK2.n881 CLK2.n877 0.1
R8719 CLK2.n877 CLK2.n873 0.1
R8720 CLK2.n10 CLK2.n6 0.1
R8721 CLK2.n14 CLK2.n10 0.1
R8722 CLK2.n18 CLK2.n14 0.1
R8723 CLK2.n22 CLK2.n18 0.1
R8724 CLK2.n26 CLK2.n22 0.1
R8725 CLK2.n35 CLK2.n31 0.1
R8726 CLK2.n39 CLK2.n35 0.1
R8727 CLK2.n40 CLK2.n39 0.1
R8728 CLK2.n51 CLK2.n47 0.1
R8729 CLK2.n55 CLK2.n51 0.1
R8730 CLK2.n64 CLK2.n60 0.1
R8731 CLK2.n68 CLK2.n64 0.1
R8732 CLK2.n72 CLK2.n68 0.1
R8733 CLK2.n244 CLK2.n243 0.087
R8734 CLK2.n203 CLK2.n202 0.087
R8735 CLK2.n255 CLK2.n173 0.087
R8736 CLK2.n364 CLK2.n363 0.087
R8737 CLK2.n537 CLK2.n536 0.087
R8738 CLK2.n614 CLK2.n613 0.087
R8739 CLK2.n554 CLK2.n550 0.087
R8740 CLK2.n688 CLK2.n687 0.087
R8741 CLK2.n629 CLK2.n625 0.087
R8742 CLK2.n703 CLK2.n699 0.087
R8743 CLK2.n853 CLK2.n852 0.087
R8744 CLK2.n873 CLK2.n869 0.087
R8745 CLK2.n351 CLK2.n350 0.086
R8746 CLK2.n73 CLK2.n72 0.077
R8747 CLK2.n233 CLK2.n232 0.075
R8748 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/CLK CLK2.n222 0.075
R8749 CLK2.n214 CLK2.n213 0.075
R8750 CLK2.n296 CLK2.n295 0.075
R8751 CLK2.n277 CLK2.n156 0.075
R8752 CLK2.n267 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/CLK 0.075
R8753 CLK2.n265 CLK2.n165 0.075
R8754 CLK2.n327 CLK2.n326 0.075
R8755 CLK2.n338 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/CLK 0.075
R8756 CLK2.n348 CLK2.n347 0.075
R8757 CLK2.n452 CLK2.n451 0.075
R8758 CLK2.n427 CLK2.n426 0.075
R8759 CLK2.n407 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/CLK 0.075
R8760 CLK2.n402 CLK2.n398 0.075
R8761 CLK2.n470 CLK2.n466 0.075
R8762 CLK2.n495 CLK2.n491 0.075
R8763 CLK2.n511 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/CLK 0.075
R8764 CLK2.n520 CLK2.n519 0.075
R8765 CLK2.n613 CLK2.n609 0.075
R8766 CLK2.n596 CLK2.n595 0.075
R8767 CLK2.n576 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/CLK 0.075
R8768 CLK2.n571 CLK2.n567 0.075
R8769 CLK2.n671 CLK2.n670 0.075
R8770 CLK2.n651 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/CLK 0.075
R8771 CLK2.n646 CLK2.n642 0.075
R8772 CLK2.n770 CLK2.n769 0.075
R8773 CLK2.n745 CLK2.n744 0.075
R8774 CLK2.n725 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/CLK 0.075
R8775 CLK2.n720 CLK2.n716 0.075
R8776 CLK2.n813 CLK2.n809 0.075
R8777 CLK2.n827 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/CLK 0.075
R8778 CLK2.n836 CLK2.n835 0.075
R8779 CLK2.n940 CLK2.n939 0.075
R8780 CLK2.n915 CLK2.n914 0.075
R8781 CLK2.n895 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/CLK 0.075
R8782 CLK2.n890 CLK2.n886 0.075
R8783 CLK2.n6 CLK2.n2 0.075
R8784 CLK2.n31 CLK2.n27 0.075
R8785 CLK2.n47 CLK2 0.075
R8786 CLK2.n56 CLK2.n55 0.075
R8787 CLK2.n382 CLK2.n381 0.074
R8788 CLK2.n314 CLK2.n140 0.072
R8789 CLK2.n389 CLK2.n388 0.072
R8790 CLK2.n788 CLK2.n784 0.072
R8791 CLK2.n947 CLK2.n944 0.062
R8792 CLK2.n364 CLK2.n111 0.06
R8793 CLK2.n371 EESPFAL_Sbox_0/EESPFAL_s2_0/CLK2 0.042
R8794 CLK2.n388 CLK2.n387 0.026
R8795 CLK2.n234 CLK2.n233 0.025
R8796 CLK2.n223 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/CLK 0.025
R8797 CLK2.n213 CLK2.n212 0.025
R8798 CLK2.n156 CLK2.n151 0.025
R8799 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/CLK CLK2.n158 0.025
R8800 CLK2.n171 CLK2.n165 0.025
R8801 CLK2.n309 CLK2.n308 0.025
R8802 CLK2.n326 CLK2.n325 0.025
R8803 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/CLK CLK2.n337 0.025
R8804 CLK2.n349 CLK2.n348 0.025
R8805 CLK2.n431 CLK2.n427 0.025
R8806 CLK2.n414 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/CLK 0.025
R8807 CLK2.n398 CLK2.n397 0.025
R8808 CLK2.n491 CLK2.n490 0.025
R8809 CLK2.n504 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/CLK 0.025
R8810 CLK2.n524 CLK2.n520 0.025
R8811 CLK2.n609 CLK2.n608 0.025
R8812 CLK2.n600 CLK2.n596 0.025
R8813 CLK2.n583 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/CLK 0.025
R8814 CLK2.n567 CLK2.n566 0.025
R8815 CLK2.n675 CLK2.n671 0.025
R8816 CLK2.n658 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/CLK 0.025
R8817 CLK2.n642 CLK2.n641 0.025
R8818 CLK2.n749 CLK2.n745 0.025
R8819 CLK2.n732 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/CLK 0.025
R8820 CLK2.n716 CLK2.n715 0.025
R8821 CLK2.n783 CLK2.n781 0.025
R8822 CLK2.n809 CLK2.n808 0.025
R8823 CLK2.n822 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/CLK 0.025
R8824 CLK2.n840 CLK2.n836 0.025
R8825 CLK2.n919 CLK2.n915 0.025
R8826 CLK2.n902 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/CLK 0.025
R8827 CLK2.n886 CLK2.n885 0.025
R8828 CLK2.n27 CLK2.n26 0.025
R8829 CLK2.n40 CLK2 0.025
R8830 CLK2.n60 CLK2.n56 0.025
R8831 EESPFAL_Sbox_0/EESPFAL_s0_0/CLK2 CLK2.n965 0.023
R8832 CLK2.n963 CLK2.n958 0.021
R8833 CLK2.n370 CLK2.n369 0.017
R8834 CLK2.n111 CLK2.n110 0.015
R8835 CLK2.n386 CLK2.n382 0.013
R8836 CLK2.n350 CLK2.n112 0.013
R8837 CLK2.n371 CLK2.n109 0.012
R8838 CLK2.n245 CLK2.n244 0.012
R8839 CLK2.n177 CLK2.n173 0.012
R8840 CLK2.n363 CLK2.n362 0.012
R8841 CLK2.n381 CLK2.n380 0.012
R8842 CLK2.n541 CLK2.n537 0.012
R8843 CLK2.n689 CLK2.n688 0.012
R8844 CLK2.n699 CLK2.n698 0.012
R8845 CLK2.n854 CLK2.n853 0.012
R8846 CLK2.n869 CLK2.n868 0.012
R8847 CLK2.n964 CLK2.n963 0.012
R8848 CLK2.n964 CLK2.n73 0.01
R8849 CLK2.n368 CLK2.n367 0.009
R8850 CLK2.n368 CLK2.n110 0.009
R8851 CLK2.n367 CLK2.n112 0.007
R8852 CLK2.n965 EESPFAL_Sbox_0/CLK2 0.004
R8853 CLK2.n308 CLK2.n140 0.002
R8854 CLK2.n784 CLK2.n781 0.002
R8855 CLK2.n387 CLK2.n386 0.001
R8856 x1.n0 x1.t1 1176.57
R8857 x1.n0 x1.t0 1149.49
R8858 x1 x1.n0 128
R8859 x1 EESPFAL_4in_XOR_0/x1 36.16
R8860 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t7 819.4
R8861 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t6 775.706
R8862 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t8 514.133
R8863 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t5 305.266
R8864 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n0 166.734
R8865 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 163.511
R8866 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n2 102.4
R8867 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n1 88.255
R8868 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t3 81.937
R8869 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n6 76
R8870 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n5 57.6
R8871 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n3 51.539
R8872 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t1 39.4
R8873 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t4 39.4
R8874 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t0 24
R8875 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t2 24
R8876 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n4 6.4
R8877 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n7 3.2
R8878 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 819.4
R8879 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 506.1
R8880 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 313.3
R8881 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 305.997
R8882 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 206.179
R8883 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 187.536
R8884 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 128.334
R8885 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 115.2
R8886 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 57.939
R8887 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 57.6
R8888 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 41.6
R8889 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 39.4
R8890 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 39.4
R8891 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 24
R8892 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 24
R8893 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 8.764
R8894 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 4.65
R8895 s3.t7 s3.t9 819.4
R8896 s3.n3 s3.t7 514.133
R8897 s3.n3 s3.t8 305.266
R8898 s3.n4 s3.n1 166.734
R8899 s3.n5 s3.n4 105.6
R8900 s3.n5 s3.t1 97.937
R8901 s3.n6 s3.n5 96
R8902 EESPFAL_Sbox_0/s3 s3.n6 83.597
R8903 s3 s3.n3 79.2
R8904 s3.n4 s3.n2 73.937
R8905 s3.n6 s3.n0 73.937
R8906 s3.n4 s3 54.4
R8907 s3.n1 s3.t3 39.4
R8908 s3.n1 s3.t6 39.4
R8909 s3.n2 s3.t2 24
R8910 s3.n2 s3.t0 24
R8911 s3.n0 s3.t4 24
R8912 s3.n0 s3.t5 24
R8913 EESPFAL_Sbox_0/s3 EESPFAL_Sbox_0/EESPFAL_s3_0/s3 0.087
R8914 Dis1.n1 Dis1 598.4
R8915 Dis1.n18 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/Dis 563.2
R8916 Dis1.n14 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/Dis 563.2
R8917 Dis1.n29 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/Dis 556.8
R8918 Dis1.n25 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/Dis 556.8
R8919 Dis1.n10 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/Dis 556.8
R8920 Dis1.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_1/Dis 556.8
R8921 Dis1.n0 Dis1.t18 504.5
R8922 Dis1.n32 Dis1.t7 504.5
R8923 Dis1.n28 Dis1.t14 504.5
R8924 Dis1.n24 Dis1.t34 504.5
R8925 Dis1.n21 Dis1.t21 504.5
R8926 Dis1.n17 Dis1.t9 504.5
R8927 Dis1.n13 Dis1.t4 504.5
R8928 Dis1.n9 Dis1.t17 504.5
R8929 Dis1.n5 Dis1.t8 504.5
R8930 Dis1.n4 Dis1.t2 504.5
R8931 Dis1.n3 Dis1.t22 504.5
R8932 Dis1.n2 Dis1.t5 389.3
R8933 Dis1.n1 Dis1.t26 389.3
R8934 Dis1.n0 Dis1.t23 389.3
R8935 Dis1.n32 Dis1.t24 389.3
R8936 Dis1.n30 Dis1.t10 389.3
R8937 Dis1.n29 Dis1.t31 389.3
R8938 Dis1.n28 Dis1.t33 389.3
R8939 Dis1.n26 Dis1.t28 389.3
R8940 Dis1.n25 Dis1.t11 389.3
R8941 Dis1.n24 Dis1.t13 389.3
R8942 Dis1.n21 Dis1.t12 389.3
R8943 Dis1.n19 Dis1.t19 389.3
R8944 Dis1.n18 Dis1.t32 389.3
R8945 Dis1.n17 Dis1.t20 389.3
R8946 Dis1.n15 Dis1.t35 389.3
R8947 Dis1.n14 Dis1.t27 389.3
R8948 Dis1.n13 Dis1.t15 389.3
R8949 Dis1.n11 Dis1.t0 389.3
R8950 Dis1.n10 Dis1.t16 389.3
R8951 Dis1.n9 Dis1.t1 389.3
R8952 Dis1.n7 Dis1.t29 389.3
R8953 Dis1.n6 Dis1.t6 389.3
R8954 Dis1.n5 Dis1.t30 389.3
R8955 Dis1.n4 Dis1.t25 389.3
R8956 Dis1.n3 Dis1.t3 389.3
R8957 Dis1.n22 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/Dis 281.856
R8958 Dis1.n33 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/Dis 241.216
R8959 Dis1.n34 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/Dis 240.897
R8960 Dis1.n8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/Dis 235.714
R8961 Dis1.n23 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/Dis 227.781
R8962 Dis1.n31 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/Dis 227.456
R8963 Dis1.n27 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/Dis 227.456
R8964 Dis1.n12 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/Dis 227.456
R8965 Dis1.n8 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/Dis 227.456
R8966 Dis1.n20 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/Dis 137.536
R8967 Dis1.n16 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/Dis 137.536
R8968 Dis1.n2 Dis1.n1 115.2
R8969 Dis1.n30 Dis1.n29 115.2
R8970 Dis1.n26 Dis1.n25 115.2
R8971 Dis1.n19 Dis1.n18 115.2
R8972 Dis1.n15 Dis1.n14 115.2
R8973 Dis1.n11 Dis1.n10 115.2
R8974 Dis1.n7 Dis1.n6 115.2
R8975 Dis1.n22 Dis1.n20 9.213
R8976 Dis1.n27 Dis1.n23 7.933
R8977 Dis1.n33 EESPFAL_Sbox_0/EESPFAL_s1_0/Dis1 4.681
R8978 Dis1.n16 EESPFAL_Sbox_0/EESPFAL_s2_0/Dis1 3.351
R8979 EESPFAL_Sbox_0/EESPFAL_s1_0/Dis1 Dis1.n31 3.266
R8980 EESPFAL_Sbox_0/EESPFAL_s3_0/Dis1 Dis1.n12 3.266
R8981 Dis1 Dis1.n0 3.2
R8982 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/Dis Dis1.n2 3.2
R8983 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/Dis Dis1.n32 3.2
R8984 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/Dis Dis1.n28 3.2
R8985 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/Dis Dis1.n30 3.2
R8986 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/Dis Dis1.n24 3.2
R8987 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/Dis Dis1.n26 3.2
R8988 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/Dis Dis1.n21 3.2
R8989 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/Dis Dis1.n17 3.2
R8990 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/Dis Dis1.n19 3.2
R8991 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/Dis Dis1.n13 3.2
R8992 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/Dis Dis1.n15 3.2
R8993 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/Dis Dis1.n9 3.2
R8994 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/Dis Dis1.n11 3.2
R8995 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_1/Dis Dis1.n5 3.2
R8996 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/Dis Dis1.n7 3.2
R8997 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/Dis Dis1.n4 3.2
R8998 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/Dis Dis1.n3 3.2
R8999 EESPFAL_Sbox_0/Dis1 Dis1.n34 3.049
R9000 EESPFAL_Sbox_0/EESPFAL_s2_0/Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/Dis1 2.199
R9001 Dis1.n23 Dis1.n22 1.174
R9002 Dis1.n12 Dis1.n8 0.627
R9003 Dis1.n20 Dis1.n16 0.627
R9004 Dis1.n31 Dis1.n27 0.627
R9005 Dis1.n34 Dis1.n33 0.625
R9006 EESPFAL_Sbox_0/Dis1 Dis1 0.165
R9007 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/Dis1 0.034
R9008 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t6 1074.82
R9009 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t7 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t9 819.4
R9010 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t8 506.1
R9011 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 442.013
R9012 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t7 313.3
R9013 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t1 273.936
R9014 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n0 128.334
R9015 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n1 105.6
R9016 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t3 81.937
R9017 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n2 57.939
R9018 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n4 57.6
R9019 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n3 41.6
R9020 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t4 39.4
R9021 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t2 39.4
R9022 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t5 24
R9023 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t0 24
R9024 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n5 8.764
R9025 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n6 4.65
R9026 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 819.4
R9027 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 506.1
R9028 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 313.3
R9029 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 305.997
R9030 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 210.945
R9031 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 187.536
R9032 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 128.334
R9033 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 115.2
R9034 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 57.937
R9035 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 57.6
R9036 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 41.6
R9037 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 39.4
R9038 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 39.4
R9039 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 24
R9040 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 24
R9041 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 8.764
R9042 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 4.65
R9043 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t5 819.4
R9044 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t7 775.706
R9045 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t6 514.133
R9046 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t8 305.266
R9047 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n4 166.736
R9048 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 163.511
R9049 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n2 102.4
R9050 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n1 88.292
R9051 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t4 81.937
R9052 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n6 76
R9053 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n5 57.6
R9054 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n0 51.537
R9055 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t1 39.4
R9056 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t2 39.4
R9057 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t0 24
R9058 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t3 24
R9059 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n3 6.4
R9060 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n7 3.2
R9061 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/A_bar 922.56
R9062 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t7 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t8 819.4
R9063 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t9 684.833
R9064 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t6 506.1
R9065 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t7 313.3
R9066 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t0 177.936
R9067 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n3 128.335
R9068 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n1 105.6
R9069 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t2 81.937
R9070 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n0 58.265
R9071 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n4 57.6
R9072 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n2 41.6
R9073 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t3 39.4
R9074 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t4 39.4
R9075 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t5 24
R9076 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t1 24
R9077 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n5 8.764
R9078 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n6 4.65
R9079 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t12 1077.04
R9080 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t14 1015.9
R9081 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t7 904.039
R9082 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t6 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t10 819.4
R9083 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t17 810.772
R9084 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t15 810.772
R9085 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t8 810.772
R9086 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/C_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t11 703.9
R9087 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t13 694.566
R9088 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t16 694.566
R9089 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t9 694.566
R9090 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t18 604.112
R9091 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t19 506.1
R9092 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B_bar 323.912
R9093 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n7 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C 314.248
R9094 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t6 313.3
R9095 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/B_bar 287.113
R9096 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/C_bar 285.185
R9097 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n8 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/B_bar 278.57
R9098 EESPFAL_Sbox_0/x0_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 274.313
R9099 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n11 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t3 273.936
R9100 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/B_bar 271.113
R9101 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_4in_XOR_0/XOR0_bar 220.08
R9102 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n14 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n13 128.335
R9103 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n11 105.6
R9104 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n11 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t4 81.937
R9105 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n0 81.6
R9106 EESPFAL_4in_XOR_0/XOR0_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n9 80.393
R9107 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n12 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n10 57.937
R9108 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n14 57.6
R9109 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n14 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n12 41.6
R9110 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t1 39.4
R9111 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n13 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t0 39.4
R9112 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n2 25.6
R9113 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n4 25.6
R9114 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n1 25.6
R9115 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n10 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t2 24
R9116 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n10 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t5 24
R9117 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n16 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n15 8.764
R9118 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n16 4.65
R9119 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n8 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n7 4.179
R9120 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n9 EESPFAL_Sbox_0/EESPFAL_s1_0/x0_bar 3.986
R9121 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/x0_bar 2.669
R9122 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n6 2.588
R9123 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n5 2.194
R9124 EESPFAL_Sbox_0/EESPFAL_s2_0/x0_bar EESPFAL_Sbox_0/EESPFAL_s3_0/x0_bar 1.39
R9125 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n9 EESPFAL_Sbox_0/x0_bar 0.387
R9126 EESPFAL_Sbox_0/EESPFAL_s1_0/x0_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n8 0.321
R9127 EESPFAL_Sbox_0/EESPFAL_s3_0/x0_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n3 0.314
R9128 s2_bar.t7 s2_bar.t6 819.4
R9129 s2_bar.n4 s2_bar.t5 506.1
R9130 s2_bar.n4 s2_bar.t7 313.3
R9131 s2_bar EESPFAL_Sbox_0/s2_bar 188.755
R9132 s2_bar.n1 s2_bar.t1 181.136
R9133 s2_bar.n3 s2_bar.n2 128.334
R9134 s2_bar.n1 s2_bar.n0 57.937
R9135 s2_bar.n5 s2_bar.n3 57.6
R9136 s2_bar.n3 s2_bar.n1 41.6
R9137 s2_bar.n2 s2_bar.t3 39.4
R9138 s2_bar.n2 s2_bar.t2 39.4
R9139 s2_bar.n0 s2_bar.t0 24
R9140 s2_bar.n0 s2_bar.t4 24
R9141 s2_bar.n5 s2_bar.n4 8.764
R9142 s2_bar s2_bar.n5 4.681
R9143 s2.t8 s2.t9 819.4
R9144 s2.n3 s2.t8 514.133
R9145 s2.n3 s2.t7 305.266
R9146 s2.n4 s2.n2 166.734
R9147 s2.n5 s2.n4 105.6
R9148 s2.n5 s2.t1 97.937
R9149 s2.n6 s2.n5 96
R9150 EESPFAL_Sbox_0/s2 s2.n6 83.731
R9151 s2 s2.n3 79.2
R9152 s2.n4 s2.n1 73.937
R9153 s2.n6 s2.n0 73.937
R9154 s2.n4 s2 54.4
R9155 s2.n2 s2.t4 39.4
R9156 s2.n2 s2.t5 39.4
R9157 s2.n1 s2.t6 24
R9158 s2.n1 s2.t0 24
R9159 s2.n0 s2.t2 24
R9160 s2.n0 s2.t3 24
R9161 EESPFAL_Sbox_0/s2 EESPFAL_Sbox_0/EESPFAL_s2_0/s2 0.081
R9162 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t7 1071.3
R9163 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t8 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t9 819.4
R9164 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 526.35
R9165 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t6 506.1
R9166 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t8 313.3
R9167 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t5 273.936
R9168 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n4 128.336
R9169 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n2 105.6
R9170 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t4 81.937
R9171 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n1 57.937
R9172 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n5 57.6
R9173 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n3 41.6
R9174 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t0 39.4
R9175 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t1 39.4
R9176 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t2 24
R9177 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t3 24
R9178 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n7 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n6 8.764
R9179 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n7 4.65
R9180 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 3.52
R9181 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n0 2.607
R9182 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t8 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t7 819.4
R9183 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t5 775.706
R9184 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t8 514.133
R9185 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t6 305.266
R9186 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n4 166.735
R9187 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C 163.511
R9188 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n2 102.4
R9189 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n1 88.255
R9190 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t1 81.937
R9191 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n6 76
R9192 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n5 57.6
R9193 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n0 51.537
R9194 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t2 39.4
R9195 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t3 39.4
R9196 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t0 24
R9197 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t4 24
R9198 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n3 6.4
R9199 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n7 3.2
R9200 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 819.4
R9201 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 506.1
R9202 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 313.3
R9203 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 305.997
R9204 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 206.179
R9205 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 187.536
R9206 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 128.335
R9207 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 115.2
R9208 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 57.937
R9209 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 57.6
R9210 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 41.6
R9211 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 39.4
R9212 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 39.4
R9213 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 24
R9214 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 24
R9215 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 8.764
R9216 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 4.65
R9217 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t8 819.4
R9218 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t7 736.033
R9219 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t6 514.133
R9220 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t9 305.266
R9221 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n5 192
R9222 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n3 166.735
R9223 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n4 105.6
R9224 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t0 97.937
R9225 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t2 97.937
R9226 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n1 76
R9227 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n0 73.937
R9228 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n2 57.6
R9229 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n6 53.658
R9230 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t3 39.4
R9231 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t4 39.4
R9232 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t1 24
R9233 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t5 24
R9234 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT 3.2
R9235 k1_bar.n0 k1_bar.t1 810.772
R9236 k1_bar.n0 k1_bar.t0 694.566
R9237 k1_bar EESPFAL_4in_XOR_0/k1_bar 36.16
R9238 k1_bar k1_bar.n0 25.6
R9239 s3_bar.t5 s3_bar.t6 819.4
R9240 s3_bar.n4 s3_bar.t7 506.1
R9241 s3_bar.n4 s3_bar.t5 313.3
R9242 EESPFAL_Sbox_0/s3_bar s3_bar 188.536
R9243 s3_bar.n2 s3_bar.t4 181.136
R9244 s3_bar.n3 s3_bar.n0 128.334
R9245 s3_bar.n2 s3_bar.n1 57.937
R9246 s3_bar.n5 s3_bar.n3 57.6
R9247 s3_bar.n3 s3_bar.n2 41.6
R9248 s3_bar.n0 s3_bar.t1 39.4
R9249 s3_bar.n0 s3_bar.t2 39.4
R9250 s3_bar.n1 s3_bar.t0 24
R9251 s3_bar.n1 s3_bar.t3 24
R9252 s3_bar.n5 s3_bar.n4 8.764
R9253 s3_bar s3_bar.n5 4.681
R9254 EESPFAL_Sbox_0/s3_bar EESPFAL_Sbox_0/EESPFAL_s3_0/s3_bar 0.09
R9255 s1.t7 s1.t8 819.4
R9256 s1.n3 s1.t7 514.133
R9257 s1.n3 s1.t9 305.266
R9258 s1.n4 s1.n1 166.734
R9259 s1.n5 s1.n4 105.6
R9260 s1.n5 s1.t5 97.937
R9261 s1.n6 s1.n5 96
R9262 EESPFAL_Sbox_0/s1 s1.n6 83.588
R9263 s1 s1.n3 79.2
R9264 s1.n4 s1.n2 73.937
R9265 s1.n6 s1.n0 73.937
R9266 s1.n4 s1 54.4
R9267 s1.n1 s1.t3 39.4
R9268 s1.n1 s1.t2 39.4
R9269 s1.n2 s1.t4 24
R9270 s1.n2 s1.t0 24
R9271 s1.n0 s1.t6 24
R9272 s1.n0 s1.t1 24
R9273 EESPFAL_Sbox_0/s1 EESPFAL_Sbox_0/EESPFAL_s1_0/s1 0.109
R9274 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t10 1074.82
R9275 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t8 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t6 819.4
R9276 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t9 736.033
R9277 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t8 514.133
R9278 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t7 305.266
R9279 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n5 192
R9280 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n0 166.734
R9281 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n4 105.6
R9282 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t0 97.939
R9283 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t3 97.937
R9284 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n7 76.565
R9285 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n2 76
R9286 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n1 73.937
R9287 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n3 57.6
R9288 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t5 39.4
R9289 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t4 39.4
R9290 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n6 25.6
R9291 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t1 24
R9292 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t2 24
R9293 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/A_bar 21.729
R9294 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT 3.2
R9295 x1_bar.n0 x1_bar.t1 1077.04
R9296 x1_bar.n0 x1_bar.t0 1015.9
R9297 x1_bar x1_bar.n0 81.6
R9298 x1_bar EESPFAL_4in_XOR_0/x1_bar 36.16
R9299 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t6 1074.82
R9300 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t9 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t10 819.4
R9301 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t8 736.033
R9302 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t7 506.1
R9303 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t9 313.3
R9304 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t0 273.936
R9305 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/A 180.175
R9306 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n0 161.141
R9307 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n4 128.335
R9308 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n2 105.6
R9309 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t2 81.937
R9310 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n5 64
R9311 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n1 57.937
R9312 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n3 41.6
R9313 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t3 39.4
R9314 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t4 39.4
R9315 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 24.135
R9316 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t5 24
R9317 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t1 24
R9318 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n7 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n6 8.764
R9319 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n7 4.65
R9320 k0.n0 k0.t0 800.452
R9321 k0.n0 k0.t1 787.997
R9322 k0 k0.n0 169.6
R9323 k0 EESPFAL_4in_XOR_0/k0 36.16
R9324 Dis0.n3 Dis0.t0 504.5
R9325 Dis0.n2 Dis0.t6 504.5
R9326 Dis0.n1 Dis0.t1 504.5
R9327 Dis0.n0 Dis0.t4 504.5
R9328 Dis0.n3 Dis0.t2 389.3
R9329 Dis0.n2 Dis0.t7 389.3
R9330 Dis0.n1 Dis0.t3 389.3
R9331 Dis0.n0 Dis0.t5 389.3
R9332 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/Dis Dis0.n6 220.138
R9333 Dis0.n4 Dis0 219.457
R9334 Dis0.n5 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_1/Dis 219.456
R9335 Dis0.n6 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_2/Dis 219.456
R9336 Dis0.n6 Dis0.n5 6.477
R9337 Dis0 Dis0.n3 3.2
R9338 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_1/Dis Dis0.n2 3.2
R9339 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_2/Dis Dis0.n1 3.2
R9340 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/Dis Dis0.n0 3.2
R9341 Dis0.n4 EESPFAL_4in_XOR_0/Dis 3.193
R9342 Dis0.n5 Dis0.n4 0.631
R9343 s0_bar.t7 s0_bar.t6 819.4
R9344 s0_bar.n4 s0_bar.t5 506.1
R9345 s0_bar.n4 s0_bar.t7 313.3
R9346 s0_bar.n1 s0_bar.t1 187.536
R9347 s0_bar.n3 s0_bar.n2 128.334
R9348 EESPFAL_Sbox_0/s0_bar s0_bar 114.151
R9349 s0_bar.n1 s0_bar.n0 57.937
R9350 s0_bar.n5 s0_bar.n3 57.6
R9351 s0_bar.n3 s0_bar.n1 41.6
R9352 s0_bar.n2 s0_bar.t2 39.4
R9353 s0_bar.n2 s0_bar.t3 39.4
R9354 s0_bar.n0 s0_bar.t0 24
R9355 s0_bar.n0 s0_bar.t4 24
R9356 s0_bar.n5 s0_bar.n4 8.764
R9357 s0_bar s0_bar.n5 4.681
R9358 EESPFAL_Sbox_0/s0_bar s0_bar 0.078
R9359 s0_bar EESPFAL_Sbox_0/EESPFAL_s0_0/s0_bar 0.003
R9360 k2.n0 k2.t0 800.452
R9361 k2.n0 k2.t1 787.997
R9362 k2 k2.n0 169.6
R9363 k2 EESPFAL_4in_XOR_0/k2 36.16
R9364 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t8 1074.82
R9365 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t9 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t6 819.4
R9366 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t7 506.1
R9367 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 442.013
R9368 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t9 313.3
R9369 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t0 273.939
R9370 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n0 128.334
R9371 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n2 105.6
R9372 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t4 81.937
R9373 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n1 57.937
R9374 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n4 57.6
R9375 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n3 41.6
R9376 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t5 39.4
R9377 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t2 39.4
R9378 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t3 24
R9379 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t1 24
R9380 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n5 8.764
R9381 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n6 4.65
R9382 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t9 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t8 819.4
R9383 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t6 736.033
R9384 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t9 514.133
R9385 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t7 305.266
R9386 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n5 192
R9387 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n3 166.735
R9388 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n4 105.6
R9389 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t0 97.937
R9390 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t2 97.937
R9391 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n1 76
R9392 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n0 73.937
R9393 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n2 57.6
R9394 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n6 56.157
R9395 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t4 39.4
R9396 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t3 39.4
R9397 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t1 24
R9398 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t5 24
R9399 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT 3.2
R9400 x3.n0 x3.t0 1176.57
R9401 x3.n0 x3.t1 1149.49
R9402 x3 x3.n0 128
R9403 x3 EESPFAL_4in_XOR_0/x3 35.84
R9404 k3.n0 k3.t1 800.452
R9405 k3.n0 k3.t0 787.997
R9406 k3 k3.n0 169.6
R9407 k3 EESPFAL_4in_XOR_0/k3 35.84
R9408 k0_bar.n0 k0_bar.t0 810.772
R9409 k0_bar.n0 k0_bar.t1 694.566
R9410 k0_bar EESPFAL_4in_XOR_0/k0_bar 36.16
R9411 k0_bar k0_bar.n0 25.6
R9412 k2_bar.n0 k2_bar.t0 810.772
R9413 k2_bar.n0 k2_bar.t1 694.566
R9414 k2_bar EESPFAL_4in_XOR_0/k2_bar 36.16
R9415 k2_bar k2_bar.n0 25.6
R9416 k1.n0 k1.t1 800.452
R9417 k1.n0 k1.t0 787.997
R9418 k1 k1.n0 169.6
R9419 k1 EESPFAL_4in_XOR_0/k1 36.16
R9420 x0.n0 x0.t1 1176.57
R9421 x0.n0 x0.t0 1149.49
R9422 x0 x0.n0 128
R9423 x0 EESPFAL_4in_XOR_0/x0 36.16
R9424 x2.n0 x2.t1 1176.57
R9425 x2.n0 x2.t0 1149.49
R9426 x2 x2.n0 128
R9427 x2 EESPFAL_4in_XOR_0/x2 36.16
R9428 k3_bar.n0 k3_bar.t0 810.772
R9429 k3_bar.n0 k3_bar.t1 694.566
R9430 k3_bar EESPFAL_4in_XOR_0/k3_bar 35.84
R9431 k3_bar k3_bar.n0 25.6
R9432 x0_bar.n0 x0_bar.t1 1077.04
R9433 x0_bar.n0 x0_bar.t0 1015.9
R9434 x0_bar x0_bar.n0 81.6
R9435 x0_bar EESPFAL_4in_XOR_0/x0_bar 36.16
R9436 x2_bar.n0 x2_bar.t1 1077.04
R9437 x2_bar.n0 x2_bar.t0 1015.9
R9438 x2_bar x2_bar.n0 81.6
R9439 x2_bar EESPFAL_4in_XOR_0/x2_bar 36.16
C0 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.04fF
C1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.03fF
C2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C3 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C4 a_6136_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C5 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C6 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar CLK1 7.33fF
C7 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C8 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C9 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.01fF
C10 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.10fF
C11 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C a_10377_n6134# 0.00fF
C12 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar a_4876_4548# 0.01fF
C13 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.32fF
C14 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.08fF
C15 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.03fF
C16 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar a_10206_5228# 0.00fF
C17 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.94fF
C18 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6136_n3313# 0.00fF
C19 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C20 a_10206_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C21 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_3040_7368# 0.00fF
C22 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.03fF
C23 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C24 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.23fF
C25 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar a_10596_1647# 0.00fF
C26 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C27 a_7196_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.00fF
C28 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4576_8048# 0.00fF
C29 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_10446_1647# 0.00fF
C30 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.03fF
C31 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.08fF
C32 a_4576_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C33 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_4616_n1173# 0.00fF
C34 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar CLK1 0.04fF
C35 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar a_6287_n6133# 0.00fF
C36 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A CLK1 1.43fF
C37 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.17fF
C38 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.07fF
C39 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.06fF
C40 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C41 a_6136_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C42 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4576_n3313# 0.00fF
C43 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.10fF
C44 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.04fF
C45 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_4616_n493# 0.00fF
C46 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.07fF
C47 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.01fF
C48 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6476_n493# 0.00fF
C49 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar a_10265_n493# 0.00fF
C50 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6136_7368# 0.01fF
C51 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.07fF
C52 a_6136_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C53 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.02fF
C54 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.01fF
C55 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C56 Dis2 a_10476_8048# 0.00fF
C57 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.01fF
C58 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C59 s0_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.01fF
C60 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_2740_8048# 0.00fF
C61 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C62 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.01fF
C63 a_10446_1647# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C64 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.36fF
C65 Dis1 a_6436_4548# 0.00fF
C66 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0.08fF
C67 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.91fF
C68 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 1.68fF
C69 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 3.63fF
C70 a_4576_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C71 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.06fF
C72 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4576_n3993# 0.00fF
C73 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.04fF
C74 a_4876_8048# CLK1 0.02fF
C75 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C76 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.02fF
C77 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.08fF
C78 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.01fF
C79 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.07fF
C80 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.09fF
C81 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C82 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6476_n1173# 0.00fF
C83 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.01fF
C84 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C85 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_4616_n1173# 0.00fF
C86 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.01fF
C87 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.02fF
C88 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4916_n493# 0.01fF
C89 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C90 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.03fF
C91 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C92 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B a_8456_7368# 0.01fF
C93 Dis1 a_3040_7368# 0.00fF
C94 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar a_6137_n6133# 0.00fF
C95 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.03fF
C96 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C97 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.04fF
C98 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 0.00fF
C99 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.04fF
C100 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C101 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.07fF
C102 a_10377_2407# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C103 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar a_6476_1648# 0.00fF
C104 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.29fF
C105 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4916_n1173# 0.01fF
C106 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_2740_5688# 0.00fF
C107 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_2740_5688# 0.00fF
C108 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar a_8456_7368# 0.01fF
C109 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_10227_2407# 0.00fF
C110 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.02fF
C111 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.00fF
C112 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4876_5228# 0.00fF
C113 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_2740_5008# 0.00fF
C114 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_6176_n493# 0.01fF
C115 a_4876_n3993# CLK1 0.02fF
C116 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.02fF
C117 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C118 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.07fF
C119 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_6136_5228# 0.00fF
C120 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.16fF
C121 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C122 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C123 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.03fF
C124 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 0.02fF
C125 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.01fF
C126 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6137_2408# 0.00fF
C127 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C128 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A 0.04fF
C129 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_1180_5688# 0.01fF
C130 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.09fF
C131 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C132 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C133 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C134 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.08fF
C135 a_4876_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C136 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.07fF
C137 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C 0.07fF
C138 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_6176_n1173# 0.00fF
C139 a_6176_n493# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C140 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4876_4548# 0.00fF
C141 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_1180_5008# 0.00fF
C142 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.48fF
C143 a_10227_2407# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C144 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_3040_5008# 0.00fF
C145 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.52fF
C146 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_4616_n493# 0.01fF
C147 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar s0_bar 0.15fF
C148 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar 0.29fF
C149 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar a_10377_n6134# 0.00fF
C150 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.16fF
C151 CLK1 a_3040_5688# 0.00fF
C152 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar a_6436_4548# 0.00fF
C153 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar 0.10fF
C154 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.22fF
C155 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar a_6436_n3993# 0.00fF
C156 a_4876_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C157 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.01fF
C158 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.31fF
C159 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.12fF
C160 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.73fF
C161 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.00fF
C162 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_6176_n1173# 0.01fF
C163 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C164 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C165 a_6136_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C166 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6136_8048# 0.00fF
C167 a_8456_7368# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.00fF
C168 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_4616_n1173# 0.00fF
C169 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.02fF
C170 a_4616_n493# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C171 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C172 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar CLK1 5.72fF
C173 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.01fF
C174 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C175 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar a_10377_n6134# 0.00fF
C176 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.17fF
C177 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.09fF
C178 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.07fF
C179 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.18fF
C180 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.10fF
C181 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6136_n3313# 0.00fF
C182 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_6176_n493# 0.00fF
C183 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.13fF
C184 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.08fF
C185 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.03fF
C186 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT a_10596_1647# 0.00fF
C187 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A a_6176_n493# 0.00fF
C188 a_7196_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C189 Dis2 a_10206_4548# 0.00fF
C190 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_4616_n1173# 0.01fF
C191 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.50fF
C192 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.15fF
C193 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4576_8048# 0.00fF
C194 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar CLK1 0.05fF
C195 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar CLK1 1.67fF
C196 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C197 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A s0 0.01fF
C198 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.14fF
C199 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.10fF
C200 CLK1 a_4576_4548# 0.01fF
C201 a_6436_8048# CLK1 0.01fF
C202 a_6136_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C203 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6136_n3993# 0.00fF
C204 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.33fF
C205 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4576_n3313# 0.00fF
C206 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C207 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C208 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.31fF
C209 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_6176_n1173# 0.00fF
C210 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.07fF
C211 a_6136_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.00fF
C212 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4616_n493# 0.00fF
C213 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT a_10265_n493# 0.01fF
C214 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.02fF
C215 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6476_n493# 0.01fF
C216 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B s0_bar 0.02fF
C217 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.99fF
C218 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.01fF
C219 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C220 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C221 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C222 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_2740_8048# 0.00fF
C223 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.01fF
C224 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.05fF
C225 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.02fF
C226 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.32fF
C227 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.03fF
C228 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C229 a_10446_1647# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C230 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_10227_n6134# 0.00fF
C231 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.10fF
C232 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0.04fF
C233 a_6137_n6133# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C234 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.00fF
C235 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.95fF
C236 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 2.67fF
C237 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.72fF
C238 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.07fF
C239 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.07fF
C240 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4576_n3993# 0.00fF
C241 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.01fF
C242 a_6176_1648# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.01fF
C243 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.07fF
C244 a_6287_2408# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.01fF
C245 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.03fF
C246 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4616_n1173# 0.00fF
C247 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C248 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.02fF
C249 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar a_6176_1648# 0.00fF
C250 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.01fF
C251 a_6287_2408# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.00fF
C252 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6476_n1173# 0.01fF
C253 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT a_10265_n1173# 0.01fF
C254 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.00fF
C255 a_4576_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C256 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.56fF
C257 a_6436_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.00fF
C258 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4916_n493# 0.00fF
C259 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.04fF
C260 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_4576_5228# 0.01fF
C261 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_1180_8048# 0.00fF
C262 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6436_5228# 0.01fF
C263 a_6436_n3993# CLK1 0.02fF
C264 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_10265_n493# 0.01fF
C265 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar a_8456_7368# 0.00fF
C266 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_10206_5228# 0.01fF
C267 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.98fF
C268 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.21fF
C269 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 0.01fF
C270 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C271 a_10377_2407# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C272 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.51fF
C273 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.07fF
C274 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4916_n1173# 0.00fF
C275 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_2740_5688# 0.00fF
C276 a_6436_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C277 a_4876_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C278 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.03fF
C279 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6436_4548# 0.00fF
C280 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_2740_5008# 0.01fF
C281 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_10265_n1173# 0.00fF
C282 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4876_5228# 0.00fF
C283 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_6176_n493# 0.00fF
C284 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C285 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.03fF
C286 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.02fF
C287 Dis1 a_4616_n493# 0.01fF
C288 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.74fF
C289 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C290 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.39fF
C291 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.03fF
C292 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6137_2408# 0.00fF
C293 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.01fF
C294 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.01fF
C295 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C296 a_6436_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C297 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A 0.00fF
C298 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C299 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C300 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_1180_5688# 0.00fF
C301 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.01fF
C302 a_4876_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.01fF
C303 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C304 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 0.34fF
C305 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_3040_7368# 0.01fF
C306 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A a_6287_2408# 0.01fF
C307 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_6176_n1173# 0.00fF
C308 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_4876_4548# 0.00fF
C309 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_7196_8048# 0.00fF
C310 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4876_4548# 0.00fF
C311 a_6176_n493# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C312 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_3040_5008# 0.00fF
C313 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.43fF
C314 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A 0.84fF
C315 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_6136_4548# 0.00fF
C316 Dis1 a_4616_n1173# 0.01fF
C317 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C318 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar a_6436_4548# 0.00fF
C319 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 0.73fF
C320 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar 0.02fF
C321 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.08fF
C322 a_4876_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.01fF
C323 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B a_8456_7368# 0.00fF
C324 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.00fF
C325 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.01fF
C326 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.23fF
C327 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.24fF
C328 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_1480_7368# 0.00fF
C329 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.00fF
C330 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_1480_7368# 0.00fF
C331 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.01fF
C332 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.00fF
C333 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_6176_n1173# 0.00fF
C334 a_3040_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C335 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C336 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C337 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C338 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6136_8048# 0.00fF
C339 Dis2 CLK1 0.32fF
C340 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C341 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_4576_4548# 0.00fF
C342 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6287_n6133# 0.00fF
C343 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C344 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.16fF
C345 CLK1 a_6136_4548# 0.02fF
C346 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.23fF
C347 Dis1 a_2740_5008# 0.00fF
C348 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.61fF
C349 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6136_n3313# 0.00fF
C350 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B s0 0.09fF
C351 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.01fF
C352 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6176_n493# 0.00fF
C353 a_10206_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.00fF
C354 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.14fF
C355 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.32fF
C356 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.01fF
C357 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT a_10596_1647# 0.00fF
C358 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar a_6176_n493# 0.00fF
C359 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.07fF
C360 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4576_8048# 0.01fF
C361 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B CLK1 0.83fF
C362 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar s0 0.01fF
C363 CLK1 a_2740_7368# 0.00fF
C364 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.21fF
C365 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.04fF
C366 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar a_10206_4548# 0.00fF
C367 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6136_n3993# 0.00fF
C368 a_6476_1648# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C369 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.01fF
C370 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6176_n1173# 0.00fF
C371 a_6136_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C372 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C373 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C374 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C375 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.02fF
C376 a_10206_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C377 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6476_n493# 0.00fF
C378 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C379 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar a_6476_1648# 0.00fF
C380 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.01fF
C381 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.08fF
C382 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar s0_bar 0.00fF
C383 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT a_10265_n493# 0.01fF
C384 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C385 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C386 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_6136_5228# 0.01fF
C387 s0_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.02fF
C388 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.21fF
C389 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.03fF
C390 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.06fF
C391 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_2740_8048# 0.00fF
C392 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A CLK1 1.05fF
C393 Dis1 a_4876_n3313# 0.01fF
C394 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.03fF
C395 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C396 a_6137_n6133# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C397 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.06fF
C398 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.05fF
C399 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 14.56fF
C400 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C401 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 2.26fF
C402 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.00fF
C403 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.13fF
C404 a_6287_2408# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C405 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4576_n3993# 0.00fF
C406 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.19fF
C407 a_6176_1648# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C408 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.14fF
C409 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6176_1648# 0.00fF
C410 a_6326_1648# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C411 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_1480_5688# 0.00fF
C412 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C413 a_6287_2408# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.00fF
C414 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT a_10265_n1173# 0.00fF
C415 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.00fF
C416 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6476_n1173# 0.00fF
C417 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C418 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C419 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.00fF
C420 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.07fF
C421 a_6436_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C422 a_4876_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.00fF
C423 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6436_5228# 0.00fF
C424 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4576_5228# 0.00fF
C425 s0_bar a_8456_7368# 0.00fF
C426 Dis1 a_6176_n493# 0.01fF
C427 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.07fF
C428 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.36fF
C429 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.41fF
C430 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.08fF
C431 s0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.00fF
C432 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_4576_n3993# 0.00fF
C433 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C434 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.09fF
C435 a_10377_2407# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C436 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_2740_5688# 0.01fF
C437 a_6436_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C438 a_3040_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C439 a_10265_n493# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C440 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4876_5228# 0.00fF
C441 a_6326_1648# CLK1 0.02fF
C442 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C443 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.01fF
C444 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.02fF
C445 Dis1 a_6176_n1173# 0.01fF
C446 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0.07fF
C447 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.00fF
C448 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.24fF
C449 a_6436_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.01fF
C450 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C451 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C452 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C453 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C454 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_1180_5688# 0.00fF
C455 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A 0.06fF
C456 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_3040_7368# 0.00fF
C457 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_3040_7368# 0.01fF
C458 a_4876_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C459 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_10265_n1173# 0.01fF
C460 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4876_4548# 0.01fF
C461 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_7196_8048# 0.00fF
C462 Dis1 a_6137_n6133# 0.00fF
C463 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B 0.71fF
C464 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C465 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_6136_4548# 0.00fF
C466 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C467 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B a_6436_4548# 0.00fF
C468 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.05fF
C469 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.07fF
C470 Dis1 a_4576_5228# 0.02fF
C471 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar 0.80fF
C472 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.69fF
C473 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar a_8456_7368# 0.00fF
C474 a_10265_n1173# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C475 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.08fF
C476 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.16fF
C477 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_1480_7368# 0.00fF
C478 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.06fF
C479 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4616_n493# 0.00fF
C480 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C481 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C482 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.00fF
C483 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.01fF
C484 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6136_8048# 0.01fF
C485 a_3040_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C486 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C487 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar CLK1 0.05fF
C488 CLK1 a_6136_7368# 0.02fF
C489 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.14fF
C490 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.22fF
C491 a_4876_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C492 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C493 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 19.73fF
C494 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 2.61fF
C495 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.05fF
C496 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar s0 0.69fF
C497 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 1.10fF
C498 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.04fF
C499 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.19fF
C500 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.01fF
C501 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4616_n1173# 0.00fF
C502 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.16fF
C503 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar 0.09fF
C504 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.01fF
C505 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.07fF
C506 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C507 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.00fF
C508 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4576_8048# 0.01fF
C509 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar CLK1 0.87fF
C510 Dis1 a_6436_n3313# 0.00fF
C511 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C512 a_6136_5228# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C513 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6136_n3993# 0.00fF
C514 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C515 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.03fF
C516 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C517 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_3040_5688# 0.00fF
C518 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.10fF
C519 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B a_6136_7368# 0.01fF
C520 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.05fF
C521 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.26fF
C522 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A s0_bar 0.12fF
C523 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C524 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.12fF
C525 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.26fF
C526 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6136_5228# 0.00fF
C527 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C528 a_6436_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.01fF
C529 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_2740_5008# 0.00fF
C530 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C531 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.01fF
C532 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar CLK1 1.42fF
C533 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C534 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 2.09fF
C535 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.05fF
C536 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.06fF
C537 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.99fF
C538 a_4576_5228# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C539 Dis1 a_3040_8048# 0.00fF
C540 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.31fF
C541 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4576_n3993# 0.01fF
C542 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.13fF
C543 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.02fF
C544 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6176_1648# 0.00fF
C545 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_6136_n3993# 0.01fF
C546 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.09fF
C547 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C548 a_6326_1648# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C549 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C550 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.02fF
C551 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C552 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.02fF
C553 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C554 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.10fF
C555 a_4876_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C556 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6436_5228# 0.00fF
C557 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C CLK1 0.10fF
C558 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 1.28fF
C559 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B s0 0.02fF
C560 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C561 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.07fF
C562 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.49fF
C563 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.23fF
C564 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.32fF
C565 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.10fF
C566 a_4876_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C567 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.10fF
C568 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.16fF
C569 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C570 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar a_4576_n3993# 0.01fF
C571 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_2740_5688# 0.00fF
C572 a_6436_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C573 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_8456_7368# 0.00fF
C574 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6436_4548# 0.01fF
C575 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_4576_4548# 0.01fF
C576 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar a_6176_n493# 0.00fF
C577 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_10206_4548# 0.00fF
C578 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.02fF
C579 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.03fF
C580 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B a_10206_5228# 0.00fF
C581 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.17fF
C582 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0.01fF
C583 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0.11fF
C584 Dis1 a_6136_5228# 0.00fF
C585 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C586 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C587 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C588 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C589 a_6436_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C590 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A 0.01fF
C591 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_3040_7368# 0.00fF
C592 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6176_n493# 0.00fF
C593 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_7196_8048# 0.01fF
C594 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4876_4548# 0.00fF
C595 a_4876_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.01fF
C596 a_1480_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C597 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar 0.93fF
C598 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C599 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.06fF
C600 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C601 a_6436_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C602 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.34fF
C603 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar 0.06fF
C604 Dis2 a_10206_n3313# 0.00fF
C605 a_4876_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C606 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6176_n1173# 0.00fF
C607 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_4616_n493# 0.00fF
C608 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.30fF
C609 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.12fF
C610 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4616_n493# 0.00fF
C611 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.03fF
C612 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.01fF
C613 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.00fF
C614 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.01fF
C615 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar a_6176_n1173# 0.00fF
C616 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6136_8048# 0.01fF
C617 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B CLK1 0.97fF
C618 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C619 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.28fF
C620 a_4576_n3313# CLK1 0.02fF
C621 a_10206_5228# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C622 a_4876_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.01fF
C623 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.05fF
C624 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.14fF
C625 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C626 a_6137_n6133# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.01fF
C627 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 3.28fF
C628 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 15.83fF
C629 s0_bar s0 1.62fF
C630 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar 0.00fF
C631 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C632 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C633 a_6287_2408# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C634 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C635 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_4616_n1173# 0.00fF
C636 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar a_6287_2408# 0.01fF
C637 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4616_n1173# 0.01fF
C638 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.29fF
C639 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C640 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.00fF
C641 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.16fF
C642 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C643 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C644 a_10476_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.01fF
C645 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4576_5228# 0.00fF
C646 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT CLK1 0.01fF
C647 a_10446_1647# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C648 CLK1 a_4916_n493# 0.01fF
C649 a_6136_5228# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C650 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6136_n3993# 0.01fF
C651 Dis1 a_4876_8048# 0.01fF
C652 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 2.14fF
C653 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6476_1648# 0.00fF
C654 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_10206_n3993# 0.01fF
C655 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar a_6136_7368# 0.01fF
C656 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_3040_5688# 0.00fF
C657 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.18fF
C658 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C659 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.02fF
C660 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.06fF
C661 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar s0_bar 0.05fF
C662 a_6436_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C663 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 3.15fF
C664 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 1.05fF
C665 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.00fF
C666 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.06fF
C667 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.01fF
C668 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C CLK1 0.11fF
C669 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_2740_5008# 0.00fF
C670 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_2740_5008# 0.00fF
C671 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.01fF
C672 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.01fF
C673 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar a_6136_5228# 0.00fF
C674 CLK1 a_4916_n1173# 0.02fF
C675 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0.00fF
C676 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 3.70fF
C677 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.02fF
C678 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.11fF
C679 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C680 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.07fF
C681 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar a_6136_n3993# 0.00fF
C682 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.04fF
C683 a_6436_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C684 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.02fF
C685 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C686 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 1.02fF
C687 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.02fF
C688 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C689 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C690 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C691 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_6136_4548# 0.01fF
C692 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_1180_5008# 0.00fF
C693 Dis1 a_4876_n3993# 0.01fF
C694 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar CLK1 0.15fF
C695 a_6137_2408# CLK1 0.02fF
C696 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar s0 0.01fF
C697 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 1.69fF
C698 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A a_4576_4548# 0.00fF
C699 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C700 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C701 s0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C702 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.14fF
C703 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.02fF
C704 CLK1 a_3040_5008# 0.00fF
C705 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C706 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.09fF
C707 a_4876_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C708 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4876_n3313# 0.00fF
C709 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_2740_7368# 0.00fF
C710 a_6436_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C711 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4576_4548# 0.00fF
C712 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C a_10446_1647# 0.00fF
C713 a_6436_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C714 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6436_4548# 0.00fF
C715 a_3040_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.01fF
C716 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 1.64fF
C717 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C718 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6287_n6133# 0.00fF
C719 Dis1 a_3040_5688# 0.00fF
C720 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.09fF
C721 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C722 s0 a_8456_7368# 0.00fF
C723 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C724 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 1.45fF
C725 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.10fF
C726 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C727 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C728 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C729 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A 0.05fF
C730 a_6436_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C731 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_6176_n493# 0.00fF
C732 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6176_n493# 0.01fF
C733 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_3040_7368# 0.00fF
C734 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4876_4548# 0.00fF
C735 a_10596_1647# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C736 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_7196_8048# 0.00fF
C737 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar 0.76fF
C738 a_1480_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.01fF
C739 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C740 a_6136_n3313# CLK1 0.02fF
C741 a_6436_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C742 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C743 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_6176_n1173# 0.00fF
C744 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6176_n1173# 0.01fF
C745 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar a_10206_n3313# 0.00fF
C746 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.04fF
C747 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.24fF
C748 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.01fF
C749 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C750 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_1480_7368# 0.01fF
C751 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4616_n493# 0.00fF
C752 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.02fF
C753 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar CLK1 1.26fF
C754 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C755 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6136_5228# 0.00fF
C756 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.32fF
C757 a_10476_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.00fF
C758 CLK1 a_6476_n493# 0.02fF
C759 Dis1 a_6436_8048# 0.00fF
C760 Dis1 a_4576_4548# 0.02fF
C761 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6137_n6133# 0.00fF
C762 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.11fF
C763 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.98fF
C764 a_2740_8048# CLK1 0.00fF
C765 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B 4.44fF
C766 a_6326_1648# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C767 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 2.27fF
C768 a_10227_2407# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C769 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A a_6326_1648# 0.01fF
C770 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6287_2408# 0.00fF
C771 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C772 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar 0.05fF
C773 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C774 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4616_n1173# 0.00fF
C775 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.01fF
C776 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.07fF
C777 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C778 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 2.13fF
C779 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_6287_2408# 0.00fF
C780 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A a_6136_7368# 0.00fF
C781 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.09fF
C782 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.02fF
C783 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C784 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4576_5228# 0.00fF
C785 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_4576_5228# 0.00fF
C786 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar CLK1 0.05fF
C787 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_4876_5228# 0.00fF
C788 CLK1 a_6476_n1173# 0.02fF
C789 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.76fF
C790 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0.10fF
C791 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.01fF
C792 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C793 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.02fF
C794 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.15fF
C795 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C796 a_10377_2407# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C797 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.05fF
C798 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.07fF
C799 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.07fF
C800 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.04fF
C801 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.04fF
C802 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar CLK1 0.16fF
C803 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_2740_5008# 0.00fF
C804 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 1.45fF
C805 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.01fF
C806 Dis1 a_6436_n3993# 0.00fF
C807 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_3040_5008# 0.00fF
C808 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT a_10227_n6134# 0.00fF
C809 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A a_6136_4548# 0.01fF
C810 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.01fF
C811 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0.00fF
C812 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.01fF
C813 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C814 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.03fF
C815 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C816 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.01fF
C817 CLK1 a_4876_5228# 0.02fF
C818 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6176_1648# 0.00fF
C819 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C820 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6436_n3313# 0.00fF
C821 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.05fF
C822 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C823 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C824 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_6136_7368# 0.00fF
C825 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C826 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A a_6326_1648# 0.00fF
C827 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C828 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6136_4548# 0.00fF
C829 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.03fF
C830 a_4876_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C831 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_10596_1647# 0.00fF
C832 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT CLK1 0.01fF
C833 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C a_10227_n6134# 0.00fF
C834 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A s0 0.06fF
C835 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar a_4576_4548# 0.01fF
C836 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.08fF
C837 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.12fF
C838 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.01fF
C839 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.02fF
C840 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4876_n3313# 0.00fF
C841 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.66fF
C842 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C843 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C844 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_2740_7368# 0.00fF
C845 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6436_4548# 0.00fF
C846 a_6436_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.00fF
C847 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar a_10446_1647# 0.00fF
C848 a_3040_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C849 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_3040_8048# 0.00fF
C850 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.09fF
C851 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6287_n6133# 0.01fF
C852 a_10377_n6134# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C853 CLK1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 1.47fF
C854 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.72fF
C855 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.01fF
C856 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.09fF
C857 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.08fF
C858 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.04fF
C859 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C860 a_4876_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C861 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6176_n493# 0.01fF
C862 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_3040_7368# 0.00fF
C863 Dis2 a_7196_8048# 0.00fF
C864 Dis1 Dis2 0.13fF
C865 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 1.24fF
C866 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C867 CLK1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 1.49fF
C868 Dis1 a_6136_4548# 0.00fF
C869 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 2.13fF
C870 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C871 a_4576_8048# CLK1 0.01fF
C872 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.05fF
C873 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_3040_5688# 0.00fF
C874 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.22fF
C875 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6176_n1173# 0.01fF
C876 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A a_10476_7368# 0.00fF
C877 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.03fF
C878 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4616_n493# 0.01fF
C879 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_10377_2407# 0.00fF
C880 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.05fF
C881 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.30fF
C882 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_6136_5228# 0.00fF
C883 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6136_5228# 0.00fF
C884 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.09fF
C885 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_6436_5228# 0.01fF
C886 a_10476_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.01fF
C887 CLK1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 1.38fF
C888 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C889 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.32fF
C890 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6137_n6133# 0.00fF
C891 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 1.23fF
C892 Dis2 a_10206_n3993# 0.00fF
C893 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar 1.23fF
C894 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 4.59fF
C895 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C896 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar 0.09fF
C897 a_10206_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C898 a_10227_2407# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C899 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar a_6326_1648# 0.00fF
C900 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_6287_2408# 0.00fF
C901 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.05fF
C902 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C903 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar a_6136_7368# 0.01fF
C904 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.33fF
C905 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4616_n1173# 0.00fF
C906 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.02fF
C907 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 6.89fF
C908 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.11fF
C909 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4576_5228# 0.00fF
C910 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_1480_5008# 0.01fF
C911 a_4576_n3993# CLK1 0.01fF
C912 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_4916_n493# 0.00fF
C913 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A CLK1 0.92fF
C914 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT a_10206_5228# 0.01fF
C915 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_4876_5228# 0.01fF
C916 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A a_10206_4548# 0.01fF
C917 CLK1 a_6436_5228# 0.02fF
C918 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6476_1648# 0.00fF
C919 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 1.45fF
C920 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C921 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.26fF
C922 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C923 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.05fF
C924 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C925 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.01fF
C926 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.02fF
C927 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.09fF
C928 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C929 a_4576_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C930 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.06fF
C931 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C932 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C933 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.33fF
C934 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4576_4548# 0.00fF
C935 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_2740_5008# 0.00fF
C936 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.04fF
C937 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.08fF
C938 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.02fF
C939 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar a_6136_4548# 0.00fF
C940 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.00fF
C941 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.07fF
C942 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C943 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.01fF
C944 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar a_6136_n3993# 0.00fF
C945 a_4576_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C946 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6436_n3313# 0.00fF
C947 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C948 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.07fF
C949 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.03fF
C950 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C951 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6136_7368# 0.00fF
C952 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C953 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.02fF
C954 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C955 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B a_6436_5228# 0.00fF
C956 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4876_8048# 0.00fF
C957 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_4916_n1173# 0.00fF
C958 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_10596_1647# 0.00fF
C959 a_4876_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C960 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C961 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C962 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT CLK1 0.01fF
C963 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar a_10227_n6134# 0.00fF
C964 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.15fF
C965 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar s0 0.10fF
C966 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A CLK1 1.07fF
C967 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.14fF
C968 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.01fF
C969 a_6436_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C970 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4876_n3313# 0.00fF
C971 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_4916_n493# 0.00fF
C972 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C973 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.01fF
C974 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT a_10446_1647# 0.00fF
C975 a_6436_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C976 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_3040_8048# 0.00fF
C977 a_10596_1647# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C978 CLK1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 1.98fF
C979 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.11fF
C980 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.16fF
C981 a_4876_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C982 a_6136_8048# CLK1 0.02fF
C983 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4876_n3993# 0.00fF
C984 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.22fF
C985 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_4916_n1173# 0.00fF
C986 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6176_n493# 0.01fF
C987 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 1.57fF
C988 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B a_10476_7368# 0.00fF
C989 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.02fF
C990 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C991 Dis1 a_6136_7368# 0.00fF
C992 CLK1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 1.87fF
C993 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C994 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C995 a_6137_2408# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C996 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.98fF
C997 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C998 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.31fF
C999 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.13fF
C1000 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_3040_5688# 0.00fF
C1001 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_3040_5688# 0.00fF
C1002 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.08fF
C1003 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_10377_2407# 0.00fF
C1004 a_6137_2408# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.00fF
C1005 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6176_n1173# 0.01fF
C1006 Dis2 s0_bar 0.01fF
C1007 a_6136_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.00fF
C1008 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.02fF
C1009 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4616_n493# 0.00fF
C1010 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.31fF
C1011 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_3040_5008# 0.00fF
C1012 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6136_5228# 0.00fF
C1013 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_6476_n493# 0.01fF
C1014 a_6136_n3993# CLK1 0.02fF
C1015 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.16fF
C1016 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar a_6136_7368# 0.00fF
C1017 CLK1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 1.93fF
C1018 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_6436_5228# 0.00fF
C1019 a_10476_8048# s0_bar 0.00fF
C1020 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.26fF
C1021 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 1.26fF
C1022 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C1023 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6137_n6133# 0.00fF
C1024 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1025 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 1.23fF
C1026 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar 21.74fF
C1027 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 1.44fF
C1028 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar 23.09fF
C1029 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6287_2408# 0.00fF
C1030 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar a_10206_n3993# 0.00fF
C1031 a_10206_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1032 a_10227_2407# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1033 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar 0.01fF
C1034 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C1035 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_1480_5688# 0.01fF
C1036 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C1037 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4616_n1173# 0.00fF
C1038 a_6136_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C1039 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.00fF
C1040 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A a_10206_5228# 0.00fF
C1041 a_6476_n493# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1042 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6136_4548# 0.00fF
C1043 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_6476_n1173# 0.00fF
C1044 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_1480_5008# 0.00fF
C1045 a_10377_2407# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1046 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4576_5228# 0.00fF
C1047 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 0.27fF
C1048 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 5.58fF
C1049 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_4916_n493# 0.01fF
C1050 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar CLK1 1.84fF
C1051 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.75fF
C1052 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.01fF
C1053 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C1054 a_6136_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.01fF
C1055 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.08fF
C1056 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.03fF
C1057 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.10fF
C1058 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 1.06fF
C1059 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1060 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C1061 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C1062 a_4576_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.01fF
C1063 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.15fF
C1064 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_2740_7368# 0.00fF
C1065 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A a_6137_2408# 0.01fF
C1066 a_6436_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C1067 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.03fF
C1068 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_4576_4548# 0.00fF
C1069 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6436_8048# 0.00fF
C1070 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_6476_n1173# 0.01fF
C1071 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1072 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4576_4548# 0.00fF
C1073 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.00fF
C1074 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_2740_5008# 0.00fF
C1075 a_4916_n493# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C1076 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_4916_n1173# 0.00fF
C1077 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.22fF
C1078 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1079 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.29fF
C1080 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.03fF
C1081 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.04fF
C1082 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.06fF
C1083 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.00fF
C1084 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1085 a_4576_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.01fF
C1086 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.03fF
C1087 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6436_n3313# 0.00fF
C1088 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.16fF
C1089 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1090 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.02fF
C1091 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_6476_n493# 0.00fF
C1092 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C1093 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C1094 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1095 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1096 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_1180_7368# 0.00fF
C1097 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1098 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A a_6476_n493# 0.00fF
C1099 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.08fF
C1100 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_1180_7368# 0.00fF
C1101 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.01fF
C1102 a_2740_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C1103 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1104 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_4916_n1173# 0.01fF
C1105 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4876_8048# 0.00fF
C1106 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1107 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C1108 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.09fF
C1109 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.66fF
C1110 CLK1 a_4876_4548# 0.02fF
C1111 a_7196_8048# CLK1 0.02fF
C1112 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6436_n3993# 0.00fF
C1113 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4876_n3313# 0.01fF
C1114 Dis1 CLK1 11.98fF
C1115 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4916_n493# 0.00fF
C1116 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.07fF
C1117 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_6476_n1173# 0.00fF
C1118 a_6436_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.00fF
C1119 Dis2 a_8456_7368# 0.02fF
C1120 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C1121 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT a_10446_1647# 0.01fF
C1122 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar a_10596_1647# 0.00fF
C1123 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_3040_8048# 0.01fF
C1124 a_10596_1647# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1125 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.19fF
C1126 CLK1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 1.04fF
C1127 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C1128 a_6326_1648# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1129 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4876_n3993# 0.00fF
C1130 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4916_n1173# 0.00fF
C1131 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar a_6326_1648# 0.00fF
C1132 a_4876_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1133 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar a_10265_n493# 0.00fF
C1134 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6176_n493# 0.00fF
C1135 a_7196_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.00fF
C1136 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_4876_5228# 0.01fF
C1137 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.13fF
C1138 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_1480_8048# 0.00fF
C1139 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C1140 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar a_10476_7368# 0.02fF
C1141 Dis1 a_4576_n3313# 0.03fF
C1142 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C1143 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.02fF
C1144 CLK1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.90fF
C1145 a_6137_2408# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C1146 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C1147 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1148 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar a_10265_n1173# 0.00fF
C1149 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.27fF
C1150 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_1180_5688# 0.00fF
C1151 a_6137_2408# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.00fF
C1152 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.00fF
C1153 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_3040_5688# 0.00fF
C1154 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.14fF
C1155 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6176_n1173# 0.00fF
C1156 a_6136_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C1157 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 1.00fF
C1158 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.38fF
C1159 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_3040_5008# 0.01fF
C1160 a_4576_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.00fF
C1161 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6136_5228# 0.00fF
C1162 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_6476_n493# 0.00fF
C1163 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1164 CLK1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.87fF
C1165 Dis1 a_4916_n493# 0.02fF
C1166 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.06fF
C1167 s0_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.03fF
C1168 a_10206_5228# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1169 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 1.68fF
C1170 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A Dis2 0.02fF
C1171 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar 1.14fF
C1172 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6287_2408# 0.00fF
C1173 a_10227_2407# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1174 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C 0.43fF
C1175 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_1480_5688# 0.00fF
C1176 a_6136_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C1177 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.03fF
C1178 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6136_7368# 0.00fF
C1179 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.07fF
C1180 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C1181 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_6136_4548# 0.00fF
C1182 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6136_4548# 0.00fF
C1183 a_2740_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1184 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_6476_n1173# 0.00fF
C1185 a_6476_n493# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C1186 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4576_5228# 0.00fF
C1187 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1188 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.83fF
C1189 a_10377_2407# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1190 a_6176_1648# CLK1 0.02fF
C1191 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_6436_4548# 0.00fF
C1192 Dis1 a_4916_n1173# 0.02fF
C1193 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 1.03fF
C1194 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.09fF
C1195 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1196 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT a_10206_n3993# 0.01fF
C1197 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 1.76fF
C1198 a_6136_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.01fF
C1199 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.07fF
C1200 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.04fF
C1201 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.16fF
C1202 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.09fF
C1203 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.06fF
C1204 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.09fF
C1205 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_2740_7368# 0.00fF
C1206 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_2740_7368# 0.01fF
C1207 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_6476_n1173# 0.00fF
C1208 a_4576_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C1209 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.06fF
C1210 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1211 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6436_8048# 0.00fF
C1212 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4576_4548# 0.01fF
C1213 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT a_10206_4548# 0.01fF
C1214 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C1215 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_4876_4548# 0.00fF
C1216 Dis1 a_6137_2408# 0.00fF
C1217 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.32fF
C1218 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B a_6136_4548# 0.00fF
C1219 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.05fF
C1220 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.02fF
C1221 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0.11fF
C1222 CLK1 a_6436_4548# 0.02fF
C1223 a_10206_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1224 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.06fF
C1225 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C1226 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.05fF
C1227 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C1228 Dis1 a_3040_5008# 0.00fF
C1229 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C1230 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6436_n3313# 0.01fF
C1231 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 1.02fF
C1232 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.02fF
C1233 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C1234 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C1235 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.03fF
C1236 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1237 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_1180_7368# 0.00fF
C1238 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar a_6476_n493# 0.00fF
C1239 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.01fF
C1240 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.06fF
C1241 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.01fF
C1242 a_10476_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0.01fF
C1243 a_2740_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C1244 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4876_8048# 0.01fF
C1245 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1246 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C1247 s0_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1248 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.87fF
C1249 CLK1 a_3040_7368# 0.00fF
C1250 a_4576_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C1251 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6436_n3993# 0.00fF
C1252 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1253 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.07fF
C1254 a_6436_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1255 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1256 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.04fF
C1257 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar a_10596_1647# 0.00fF
C1258 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.08fF
C1259 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_6436_5228# 0.01fF
C1260 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_3040_8048# 0.00fF
C1261 a_10227_2407# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C1262 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 1.18fF
C1263 Dis1 a_6136_n3313# 0.00fF
C1264 CLK1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.87fF
C1265 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C1266 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4876_n3993# 0.00fF
C1267 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6326_1648# 0.01fF
C1268 a_6476_1648# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1269 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.01fF
C1270 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_2740_5688# 0.00fF
C1271 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar a_10265_n493# 0.00fF
C1272 a_10206_n3313# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C1273 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.03fF
C1274 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.30fF
C1275 a_6136_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.01fF
C1276 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4876_5228# 0.01fF
C1277 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.04fF
C1278 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.02fF
C1279 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 4.22fF
C1280 s0_bar a_10476_7368# 0.00fF
C1281 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C1282 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C1283 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar CLK1 1.44fF
C1284 CLK1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 1.01fF
C1285 Dis1 a_6476_n493# 0.00fF
C1286 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 1.57fF
C1287 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_4876_n3993# 0.00fF
C1288 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.04fF
C1289 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar a_10265_n1173# 0.00fF
C1290 a_6176_1648# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C1291 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1292 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B s0_bar 0.00fF
C1293 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1294 a_10206_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.01fF
C1295 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_3040_5688# 0.01fF
C1296 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.09fF
C1297 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.01fF
C1298 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.03fF
C1299 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1300 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 2.86fF
C1301 a_4576_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C1302 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B a_6476_n493# 0.00fF
C1303 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6136_5228# 0.00fF
C1304 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1305 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_10206_4548# 0.00fF
C1306 a_6476_1648# CLK1 0.02fF
C1307 CLK1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 1.17fF
C1308 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A a_6287_n6133# 0.01fF
C1309 Dis1 a_6476_n1173# 0.00fF
C1310 a_10206_5228# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1311 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.02fF
C1312 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B Dis2 0.01fF
C1313 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar 15.98fF
C1314 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.70fF
C1315 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 0.25fF
C1316 a_4576_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1317 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_1480_5688# 0.00fF
C1318 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C1319 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.04fF
C1320 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6136_7368# 0.00fF
C1321 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_6136_7368# 0.00fF
C1322 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C1323 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.03fF
C1324 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.02fF
C1325 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6136_4548# 0.01fF
C1326 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C1327 a_6136_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C1328 a_8456_7368# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1329 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.79fF
C1330 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C1331 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_6436_4548# 0.00fF
C1332 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.10fF
C1333 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1334 Dis2 s0 0.02fF
C1335 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.32fF
C1336 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.08fF
C1337 Dis1 a_4876_5228# 0.01fF
C1338 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar a_10206_n3993# 0.00fF
C1339 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.06fF
C1340 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.33fF
C1341 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.20fF
C1342 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.00fF
C1343 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.14fF
C1344 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.04fF
C1345 a_6136_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1346 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.87fF
C1347 a_10476_8048# s0 0.00fF
C1348 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1349 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4916_n493# 0.01fF
C1350 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 3.16fF
C1351 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_2740_7368# 0.00fF
C1352 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C1353 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B a_6476_n1173# 0.00fF
C1354 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_4576_4548# 0.00fF
C1355 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar a_6436_5228# 0.00fF
C1356 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.13fF
C1357 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6436_8048# 0.01fF
C1358 a_4576_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C1359 a_1180_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1360 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1361 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C1362 CLK1 a_8456_7368# 0.00fF
C1363 Dis2 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.24fF
C1364 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A a_6137_n6133# 0.01fF
C1365 a_6136_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.01fF
C1366 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 0.04fF
C1367 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1368 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar 0.68fF
C1369 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.02fF
C1370 a_10206_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C1371 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.06fF
C1372 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.05fF
C1373 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 3.09fF
C1374 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.31fF
C1375 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.27fF
C1376 a_4576_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C1377 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4916_n1173# 0.00fF
C1378 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1379 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.02fF
C1380 a_10476_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.01fF
C1381 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.01fF
C1382 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.03fF
C1383 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C1384 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.13fF
C1385 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1386 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4876_8048# 0.01fF
C1387 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.02fF
C1388 s0_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C1389 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.29fF
C1390 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 20.59fF
C1391 a_4576_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C1392 a_6436_5228# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C1393 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.02fF
C1394 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.05fF
C1395 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1396 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1397 a_6137_2408# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1398 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.01fF
C1399 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.97fF
C1400 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C1401 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.07fF
C1402 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C1403 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.10fF
C1404 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1405 Dis2 a_10265_n493# 0.00fF
C1406 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.07fF
C1407 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar a_6137_2408# 0.01fF
C1408 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6436_5228# 0.00fF
C1409 a_7196_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.01fF
C1410 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.32fF
C1411 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_3040_5008# 0.00fF
C1412 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 1.02fF
C1413 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B a_6436_5228# 0.00fF
C1414 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.31fF
C1415 CLK1 a_4616_n493# 0.01fF
C1416 a_4876_5228# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1417 Dis1 a_4576_8048# 0.02fF
C1418 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4876_n3993# 0.01fF
C1419 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_6436_n3993# 0.01fF
C1420 a_6476_1648# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C1421 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6326_1648# 0.00fF
C1422 Dis2 a_10265_n1173# 0.00fF
C1423 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar a_3040_7368# 0.00fF
C1424 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_2740_5688# 0.00fF
C1425 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C1426 a_10206_n3313# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.00fF
C1427 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.11fF
C1428 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.10fF
C1429 a_6136_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C1430 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C1431 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.02fF
C1432 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.00fF
C1433 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.06fF
C1434 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 2.05fF
C1435 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A CLK1 8.62fF
C1436 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C CLK1 0.12fF
C1437 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.29fF
C1438 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C1439 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.00fF
C1440 CLK1 a_4616_n1173# 0.01fF
C1441 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar a_4876_n3993# 0.01fF
C1442 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.02fF
C1443 a_6136_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1444 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1445 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_3040_5688# 0.00fF
C1446 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.01fF
C1447 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_4876_4548# 0.01fF
C1448 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.04fF
C1449 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.34fF
C1450 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_10206_4548# 0.00fF
C1451 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar a_6476_n493# 0.00fF
C1452 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 1.08fF
C1453 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.12fF
C1454 Dis1 a_4576_n3993# 0.02fF
C1455 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar a_6287_n6133# 0.00fF
C1456 CLK1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1457 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.02fF
C1458 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.01fF
C1459 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.00fF
C1460 Dis1 a_6436_5228# 0.00fF
C1461 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.88fF
C1462 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar Dis2 0.00fF
C1463 a_4576_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C1464 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4576_n3313# 0.00fF
C1465 a_6136_n3313# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C1466 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.01fF
C1467 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6476_n493# 0.00fF
C1468 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_6136_7368# 0.00fF
C1469 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.00fF
C1470 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.01fF
C1471 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C1472 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.03fF
C1473 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1474 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.16fF
C1475 a_6136_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C1476 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6136_4548# 0.00fF
C1477 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0.00fF
C1478 a_8456_7368# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.00fF
C1479 a_2740_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.01fF
C1480 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.01fF
C1481 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.02fF
C1482 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT a_10206_4548# 0.01fF
C1483 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 1.05fF
C1484 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.19fF
C1485 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C1486 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.27fF
C1487 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.12fF
C1488 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C1489 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1490 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.04fF
C1491 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.00fF
C1492 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C1493 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.02fF
C1494 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6476_n1173# 0.00fF
C1495 a_6136_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C1496 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.00fF
C1497 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A a_10476_7368# 0.01fF
C1498 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.07fF
C1499 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4916_n493# 0.00fF
C1500 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_4916_n493# 0.00fF
C1501 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_2740_7368# 0.00fF
C1502 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.31fF
C1503 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_4576_4548# 0.00fF
C1504 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar a_6476_n1173# 0.00fF
C1505 Dis2 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.31fF
C1506 s0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C1507 a_10446_1647# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1508 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6436_8048# 0.01fF
C1509 a_1180_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.01fF
C1510 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1511 a_4876_n3313# CLK1 0.02fF
C1512 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A 0.11fF
C1513 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0.00fF
C1514 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar a_6137_n6133# 0.00fF
C1515 a_6136_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.00fF
C1516 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.03fF
C1517 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1518 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1519 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 0.08fF
C1520 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.09fF
C1521 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.08fF
C1522 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.13fF
C1523 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 1.06fF
C1524 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 1.64fF
C1525 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C1526 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_4916_n1173# 0.00fF
C1527 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4916_n1173# 0.01fF
C1528 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.08fF
C1529 CLK1 a_6287_n6133# 0.02fF
C1530 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_1180_7368# 0.01fF
C1531 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.07fF
C1532 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.39fF
C1533 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_4876_5228# 0.00fF
C1534 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C1535 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C1536 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar a_10377_n6134# 0.00fF
C1537 CLK1 a_6176_n493# 0.02fF
C1538 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.01fF
C1539 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.38fF
C1540 a_10596_1647# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C1541 a_6436_5228# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1542 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.00fF
C1543 Dis1 a_6136_8048# 0.00fF
C1544 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6436_n3993# 0.01fF
C1545 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1546 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.06fF
C1547 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.06fF
C1548 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C1549 a_6176_1648# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.00fF
C1550 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.08fF
C1551 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.04fF
C1552 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A a_6176_1648# 0.01fF
C1553 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.10fF
C1554 a_6137_2408# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C1555 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6137_2408# 0.01fF
C1556 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.31fF
C1557 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C1558 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C1559 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.01fF
C1560 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_6137_2408# 0.00fF
C1561 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.02fF
C1562 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C1563 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.07fF
C1564 a_7196_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C1565 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_3040_5008# 0.00fF
C1566 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_3040_5008# 0.00fF
C1567 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.08fF
C1568 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.38fF
C1569 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.78fF
C1570 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar a_6436_5228# 0.00fF
C1571 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_4576_5228# 0.00fF
C1572 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.90fF
C1573 CLK1 a_6176_n1173# 0.02fF
C1574 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.34fF
C1575 s0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1576 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar a_6436_n3993# 0.00fF
C1577 a_10227_2407# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1578 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.14fF
C1579 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.10fF
C1580 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A s0_bar 0.01fF
C1581 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_6436_4548# 0.00fF
C1582 Dis2 a_10206_5228# 0.00fF
C1583 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_1480_5008# 0.00fF
C1584 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.04fF
C1585 a_6137_n6133# CLK1 0.02fF
C1586 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.00fF
C1587 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C1588 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1589 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C1590 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B CLK1 6.23fF
C1591 Dis1 a_6136_n3993# 0.00fF
C1592 a_6287_2408# CLK1 0.02fF
C1593 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.00fF
C1594 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.01fF
C1595 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar CLK1 0.17fF
C1596 Dis1 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.33fF
C1597 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_2740_5008# 0.00fF
C1598 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A a_4876_4548# 0.00fF
C1599 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.28fF
C1600 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.04fF
C1601 CLK1 a_4576_5228# 0.01fF
C1602 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.06fF
C1603 a_6136_n3313# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.00fF
C1604 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6136_n3313# 0.00fF
C1605 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_3040_7368# 0.00fF
C1606 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A a_6176_1648# 0.00fF
C1607 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1608 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.03fF
C1609 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_4876_4548# 0.01fF
C1610 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C a_10596_1647# 0.00fF
C1611 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.96fF
C1612 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.42fF
C1613 a_4576_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1614 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0.81fF
C1615 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_10446_1647# 0.00fF
C1616 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0.39fF
C1617 a_10377_2407# EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C1618 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C a_6287_n6133# 0.00fF
C1619 Dis1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.10fF
C1620 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.10fF
C1621 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.03fF
C1622 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.01fF
C1623 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar Dis2 0.00fF
C1624 CLK1 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C1625 s0 a_10476_7368# 0.00fF
C1626 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4576_n3313# 0.00fF
C1627 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.09fF
C1628 a_10206_n3993# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C1629 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar a_6136_7368# 0.01fF
C1630 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.02fF
C1631 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.01fF
C1632 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6476_n493# 0.00fF
C1633 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C a_10265_n493# 0.00fF
C1634 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.03fF
C1635 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1636 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6136_4548# 0.00fF
C1637 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C1638 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.01fF
C1639 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.02fF
C1640 CLK1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0.02fF
C1641 a_2740_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0.01fF
C1642 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.01fF
C1643 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C1644 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_2740_8048# 0.00fF
C1645 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B s0 0.00fF
C1646 a_6436_n3313# CLK1 0.02fF
C1647 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar a_10206_4548# 0.00fF
C1648 a_10227_n6134# EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1649 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.41fF
C1650 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.08fF
C1651 Dis2 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar 0.28fF
C1652 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.37fF
C1653 Dis2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.04fF
C1654 a_4576_n3993# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1655 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C1656 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1657 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.01fF
C1658 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar a_10476_7368# 0.00fF
C1659 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.07fF
C1660 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.09fF
C1661 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.00fF
C1662 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C1663 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C1664 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_6476_n1173# 0.01fF
C1665 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0.01fF
C1666 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.01fF
C1667 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_2740_7368# 0.00fF
C1668 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.38fF
C1669 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4916_n493# 0.00fF
C1670 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 1.00fF
C1671 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_6436_5228# 0.00fF
C1672 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C1673 Dis1 a_4876_4548# 0.01fF
C1674 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C a_6137_n6133# 0.00fF
C1675 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 3.23fF
C1676 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C1677 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.00fF
C1678 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 1.02fF
C1679 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 0.09fF
C1680 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C1681 Dis1 a_7196_8048# 0.00fF
C1682 a_6476_1648# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0.01fF
C1683 a_3040_8048# CLK1 0.00fF
C1684 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.04fF
C1685 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.33fF
C1686 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.01fF
C1687 a_10377_2407# EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1688 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A a_6476_1648# 0.01fF
C1689 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.36fF
C1690 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_4916_n1173# 0.00fF
C1691 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A a_2740_5688# 0.00fF
C1692 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.09fF
C1693 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_10227_2407# 0.00fF
C1694 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A a_8456_7368# 0.00fF
C1695 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C1696 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.10fF
C1697 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C1698 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar a_4876_5228# 0.00fF
C1699 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A a_4876_5228# 0.00fF
C1700 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1701 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C1702 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_6136_5228# 0.01fF
C1703 a_7196_8048# EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.00fF
C1704 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.09fF
C1705 Dis1 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.02fF
C1706 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C1707 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0.00fF
C1708 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 0.01fF
C1709 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1710 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0.01fF
C1711 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1712 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.33fF
C1713 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C1714 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar a_6176_1648# 0.00fF
C1715 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0.00fF
C1716 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1717 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C1718 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_6137_2408# 0.00fF
C1719 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.13fF
C1720 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.05fF
C1721 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar 0.74fF
C1722 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.56fF
C1723 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar a_1180_5008# 0.01fF
C1724 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B a_3040_5008# 0.00fF
C1725 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.34fF
C1726 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_4616_n493# 0.00fF
C1727 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B s0_bar 0.90fF
C1728 Dis1 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.09fF
C1729 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_4576_5228# 0.01fF
C1730 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT a_10377_n6134# 0.00fF
C1731 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A a_6436_4548# 0.01fF
C1732 s0 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.01fF
C1733 CLK1 a_6136_5228# 0.02fF
C1734 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B a_6436_n3993# 0.00fF
C1735 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C1736 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar a_6326_1648# 0.00fF
C1737 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1738 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A a_6476_1648# 0.00fF
C1739 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar s0_bar 0.00fF
C1740 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.11fF
C1741 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.08fF
C1742 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.08fF
C1743 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B a_6436_4548# 0.00fF
C1744 a_10377_n6134# 0 0.02fF
C1745 a_10227_n6134# 0 0.02fF
C1746 a_6287_n6133# 0 0.02fF
C1747 a_6137_n6133# 0 0.02fF
C1748 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0 1.26fF $ **FLOATING
C1749 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0 1.22fF $ **FLOATING
C1750 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 0 1.22fF
C1751 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/A 0 1.36fF
C1752 a_10206_n3993# 0 0.02fF
C1753 a_6436_n3993# 0 0.01fF
C1754 a_6136_n3993# 0 0.01fF
C1755 a_4876_n3993# 0 0.01fF
C1756 a_4576_n3993# 0 0.01fF
C1757 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0 1.49fF
C1758 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0 1.14fF
C1759 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0 1.09fF
C1760 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0 1.28fF
C1761 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0 2.14fF $ **FLOATING
C1762 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0 2.42fF $ **FLOATING
C1763 a_10206_n3313# 0 0.02fF
C1764 a_6436_n3313# 0 0.01fF
C1765 a_6136_n3313# 0 0.01fF
C1766 a_4876_n3313# 0 0.01fF
C1767 a_4576_n3313# 0 0.01fF
C1768 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0 2.53fF $ **FLOATING
C1769 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0 1.73fF
C1770 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0 1.10fF
C1771 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0 1.34fF
C1772 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0 2.68fF $ **FLOATING
C1773 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0 1.93fF $ **FLOATING
C1774 a_10265_n1173# 0 0.02fF
C1775 a_6476_n1173# 0 0.01fF
C1776 a_6176_n1173# 0 0.01fF
C1777 a_4916_n1173# 0 0.02fF
C1778 a_4616_n1173# 0 0.01fF
C1779 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0 1.14fF
C1780 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0 1.34fF
C1781 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0 2.10fF $ **FLOATING
C1782 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0 1.65fF $ **FLOATING
C1783 a_10265_n493# 0 0.02fF
C1784 a_6476_n493# 0 0.01fF
C1785 a_6176_n493# 0 0.01fF
C1786 a_4916_n493# 0 0.02fF
C1787 a_4616_n493# 0 0.01fF
C1788 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0 1.09fF
C1789 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0 1.24fF
C1790 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0 1.57fF
C1791 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0 1.41fF
C1792 a_10596_1647# 0 0.02fF
C1793 a_10446_1647# 0 0.02fF
C1794 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar 0 2.57fF $ **FLOATING
C1795 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0 1.54fF
C1796 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0 1.14fF
C1797 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT 0 1.69fF
C1798 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0 1.28fF $ **FLOATING
C1799 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0 1.25fF $ **FLOATING
C1800 a_6476_1648# 0 0.02fF
C1801 a_6326_1648# 0 0.02fF
C1802 a_6176_1648# 0 0.02fF
C1803 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 0 1.70fF
C1804 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/A 0 1.69fF
C1805 a_10377_2407# 0 0.02fF
C1806 a_10227_2407# 0 0.02fF
C1807 a_6287_2408# 0 0.02fF
C1808 a_6137_2408# 0 0.02fF
C1809 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 0 1.28fF $ **FLOATING
C1810 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C 0 1.25fF $ **FLOATING
C1811 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A_bar 0 1.33fF
C1812 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/A 0 1.35fF
C1813 a_10206_4548# 0 0.02fF
C1814 a_6436_4548# 0 0.01fF
C1815 a_6136_4548# 0 0.01fF
C1816 a_4876_4548# 0 0.01fF
C1817 a_4576_4548# 0 0.01fF
C1818 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0 1.50fF
C1819 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0 1.14fF
C1820 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0 1.21fF
C1821 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0 1.11fF
C1822 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0 2.39fF $ **FLOATING
C1823 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0 2.46fF $ **FLOATING
C1824 a_10206_5228# 0 0.02fF
C1825 a_6436_5228# 0 0.01fF
C1826 a_6136_5228# 0 0.01fF
C1827 a_4876_5228# 0 0.02fF
C1828 a_4576_5228# 0 0.02fF
C1829 a_3040_5008# 0 0.02fF
C1830 a_2740_5008# 0 0.02fF
C1831 a_1480_5008# 0 0.02fF
C1832 a_1180_5008# 0 0.01fF
C1833 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0 2.53fF $ **FLOATING
C1834 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0 1.74fF
C1835 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0 1.10fF
C1836 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0 1.33fF
C1837 a_3040_5688# 0 0.01fF
C1838 a_2740_5688# 0 0.01fF
C1839 a_1480_5688# 0 0.02fF
C1840 a_1180_5688# 0 0.02fF
C1841 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0 2.64fF $ **FLOATING
C1842 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0 1.90fF $ **FLOATING
C1843 a_10476_7368# 0 0.01fF
C1844 a_8456_7368# 0 0.01fF
C1845 a_6136_7368# 0 0.02fF
C1846 a_3040_7368# 0 0.02fF
C1847 a_2740_7368# 0 0.02fF
C1848 a_1480_7368# 0 0.02fF
C1849 a_1180_7368# 0 0.02fF
C1850 s0 0 0.86fF
C1851 s0_bar 0 0.79fF
C1852 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0 1.44fF
C1853 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0 1.10fF
C1854 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0 1.32fF
C1855 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0 1.29fF
C1856 a_10476_8048# 0 0.02fF
C1857 a_7196_8048# 0 0.02fF
C1858 a_6436_8048# 0 0.01fF
C1859 a_6136_8048# 0 0.01fF
C1860 a_4876_8048# 0 0.01fF
C1861 a_4576_8048# 0 0.01fF
C1862 a_3040_8048# 0 0.01fF
C1863 a_2740_8048# 0 0.01fF
C1864 a_1480_8048# 0 0.01fF
C1865 a_1180_8048# 0 0.01fF
C1866 Dis2 0 17.25fF
C1867 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar 0 7.46fF $ **FLOATING
C1868 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar 0 7.31fF $ **FLOATING
C1869 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B 0 8.30fF $ **FLOATING
C1870 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A 0 7.24fF
C1871 Dis1 0 29.93fF
C1872 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar 0 1.73fF
C1873 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_0/A 0 1.61fF
C1874 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0 1.17fF
C1875 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/B 0 1.33fF
C1876 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B 0 6.58fF
C1877 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar 0 17.93fF $ **FLOATING
C1878 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0 2.49fF $ **FLOATING
C1879 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0 3.06fF $ **FLOATING
C1880 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar 0 7.54fF $ **FLOATING
C1881 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A 0 8.23fF
C1882 CLK1 0 61.04fF
C1883 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t6 0 0.08fF
C1884 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t2 0 0.24fF
C1885 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t0 0 0.24fF
C1886 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t1 0 0.05fF
C1887 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t5 0 0.05fF
C1888 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n0 0 0.18fF $ **FLOATING
C1889 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t8 0 0.07fF
C1890 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t9 0 0.08fF
C1891 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t7 0 0.04fF
C1892 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n1 0 0.08fF $ **FLOATING
C1893 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT 0 0.01fF $ **FLOATING
C1894 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n2 0 0.04fF $ **FLOATING
C1895 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t4 0 0.05fF
C1896 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t3 0 0.05fF
C1897 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n3 0 0.17fF $ **FLOATING
C1898 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n4 0 0.24fF $ **FLOATING
C1899 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n5 0 0.24fF $ **FLOATING
C1900 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n6 0 0.52fF $ **FLOATING
C1901 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT_bar 0 0.30fF $ **FLOATING
C1902 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t8 0 0.12fF
C1903 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t5 0 0.04fF
C1904 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t2 0 0.04fF
C1905 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n0 0 0.11fF $ **FLOATING
C1906 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t3 0 0.04fF
C1907 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t1 0 0.04fF
C1908 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n1 0 0.13fF $ **FLOATING
C1909 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t4 0 0.17fF
C1910 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t0 0 0.29fF
C1911 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n2 0 0.26fF $ **FLOATING
C1912 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n3 0 0.11fF $ **FLOATING
C1913 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n4 0 0.12fF $ **FLOATING
C1914 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t6 0 0.06fF
C1915 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t9 0 0.05fF
C1916 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t7 0 0.04fF
C1917 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n5 0 0.06fF $ **FLOATING
C1918 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n6 0 0.04fF $ **FLOATING
C1919 Dis0.t4 0 0.17fF
C1920 Dis0.t5 0 0.11fF
C1921 Dis0.n0 0 0.42fF $ **FLOATING
C1922 Dis0.t1 0 0.17fF
C1923 Dis0.t3 0 0.11fF
C1924 Dis0.n1 0 0.42fF $ **FLOATING
C1925 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_2/Dis 0 0.20fF $ **FLOATING
C1926 Dis0.t6 0 0.17fF
C1927 Dis0.t7 0 0.11fF
C1928 Dis0.n2 0 0.42fF $ **FLOATING
C1929 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_1/Dis 0 0.20fF $ **FLOATING
C1930 Dis0.t0 0 0.17fF
C1931 Dis0.t2 0 0.11fF
C1932 Dis0.n3 0 0.42fF $ **FLOATING
C1933 EESPFAL_4in_XOR_0/Dis 0 0.29fF $ **FLOATING
C1934 Dis0.n4 0 0.61fF $ **FLOATING
C1935 Dis0.n5 0 0.88fF $ **FLOATING
C1936 Dis0.n6 0 1.25fF $ **FLOATING
C1937 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/Dis 0 0.20fF $ **FLOATING
C1938 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT_bar 0 0.12fF $ **FLOATING
C1939 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t8 0 0.04fF
C1940 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t6 0 0.07fF
C1941 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/A 0 0.34fF $ **FLOATING
C1942 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n0 0 0.62fF $ **FLOATING
C1943 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t5 0 0.03fF
C1944 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t1 0 0.03fF
C1945 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n1 0 0.08fF $ **FLOATING
C1946 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t2 0 0.11fF
C1947 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t0 0 0.18fF
C1948 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n2 0 0.16fF $ **FLOATING
C1949 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n3 0 0.07fF $ **FLOATING
C1950 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t3 0 0.03fF
C1951 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t4 0 0.03fF
C1952 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n4 0 0.07fF $ **FLOATING
C1953 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n5 0 0.08fF $ **FLOATING
C1954 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t10 0 0.04fF
C1955 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t9 0 0.03fF
C1956 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t7 0 0.03fF
C1957 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n6 0 0.04fF $ **FLOATING
C1958 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n7 0 0.01fF $ **FLOATING
C1959 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t10 0 0.08fF
C1960 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t9 0 0.04fF
C1961 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/A_bar 0 0.16fF $ **FLOATING
C1962 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t3 0 0.12fF
C1963 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t5 0 0.03fF
C1964 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t4 0 0.03fF
C1965 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n0 0 0.09fF $ **FLOATING
C1966 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t1 0 0.03fF
C1967 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t2 0 0.03fF
C1968 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n1 0 0.10fF $ **FLOATING
C1969 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t6 0 0.04fF
C1970 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t8 0 0.04fF
C1971 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t7 0 0.02fF
C1972 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n2 0 0.04fF $ **FLOATING
C1973 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT 0 0.01fF $ **FLOATING
C1974 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n3 0 0.02fF $ **FLOATING
C1975 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n4 0 0.13fF $ **FLOATING
C1976 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t0 0 0.12fF
C1977 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n5 0 0.13fF $ **FLOATING
C1978 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n6 0 0.11fF $ **FLOATING
C1979 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n7 0 0.36fF $ **FLOATING
C1980 EESPFAL_Sbox_0/EESPFAL_s1_0/s1 0 0.01fF $ **FLOATING
C1981 s1.t6 0 0.04fF
C1982 s1.t1 0 0.04fF
C1983 s1.n0 0 0.15fF $ **FLOATING
C1984 s1.t5 0 0.19fF
C1985 s1.t3 0 0.04fF
C1986 s1.t2 0 0.04fF
C1987 s1.n1 0 0.14fF $ **FLOATING
C1988 s1.t4 0 0.04fF
C1989 s1.t0 0 0.04fF
C1990 s1.n2 0 0.15fF $ **FLOATING
C1991 s1.t8 0 0.06fF
C1992 s1.t7 0 0.06fF
C1993 s1.t9 0 0.03fF
C1994 s1.n3 0 0.06fF $ **FLOATING
C1995 s1.n4 0 0.19fF $ **FLOATING
C1996 s1.n5 0 0.16fF $ **FLOATING
C1997 s1.n6 0 0.13fF $ **FLOATING
C1998 EESPFAL_Sbox_0/s1 0 0.48fF $ **FLOATING
C1999 EESPFAL_Sbox_0/EESPFAL_s3_0/s3_bar 0 0.01fF $ **FLOATING
C2000 s3_bar.t1 0 0.05fF
C2001 s3_bar.t2 0 0.05fF
C2002 s3_bar.n0 0 0.12fF $ **FLOATING
C2003 s3_bar.t0 0 0.05fF
C2004 s3_bar.t3 0 0.05fF
C2005 s3_bar.n1 0 0.14fF $ **FLOATING
C2006 s3_bar.t4 0 0.27fF
C2007 s3_bar.n2 0 0.19fF $ **FLOATING
C2008 s3_bar.n3 0 0.13fF $ **FLOATING
C2009 s3_bar.t6 0 0.06fF
C2010 s3_bar.t5 0 0.06fF
C2011 s3_bar.t7 0 0.04fF
C2012 s3_bar.n4 0 0.07fF $ **FLOATING
C2013 s3_bar.n5 0 0.05fF $ **FLOATING
C2014 EESPFAL_Sbox_0/s3_bar 0 0.57fF $ **FLOATING
C2015 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t7 0 0.07fF
C2016 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t2 0 0.23fF
C2017 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t0 0 0.23fF
C2018 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t1 0 0.05fF
C2019 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t5 0 0.05fF
C2020 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n0 0 0.18fF $ **FLOATING
C2021 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t8 0 0.07fF
C2022 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t6 0 0.08fF
C2023 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t9 0 0.04fF
C2024 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n1 0 0.08fF $ **FLOATING
C2025 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT 0 0.01fF $ **FLOATING
C2026 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n2 0 0.04fF $ **FLOATING
C2027 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t3 0 0.05fF
C2028 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t4 0 0.05fF
C2029 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n3 0 0.16fF $ **FLOATING
C2030 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n4 0 0.24fF $ **FLOATING
C2031 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n5 0 0.24fF $ **FLOATING
C2032 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n6 0 0.56fF $ **FLOATING
C2033 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/OUT 0 0.23fF $ **FLOATING
C2034 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 0 0.03fF
C2035 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 0 0.63fF $ **FLOATING
C2036 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 0 0.04fF
C2037 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 0 0.04fF
C2038 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 0 0.13fF $ **FLOATING
C2039 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 0 0.25fF
C2040 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 0 0.17fF $ **FLOATING
C2041 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 0 0.04fF
C2042 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 0 0.04fF
C2043 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 0 0.11fF $ **FLOATING
C2044 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 0 0.12fF $ **FLOATING
C2045 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 0 0.06fF
C2046 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 0 0.05fF
C2047 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 0 0.04fF
C2048 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 0 0.06fF $ **FLOATING
C2049 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 0 0.04fF $ **FLOATING
C2050 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t0 0 0.04fF
C2051 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t4 0 0.04fF
C2052 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n0 0 0.12fF $ **FLOATING
C2053 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t1 0 0.16fF
C2054 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t5 0 0.05fF
C2055 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n1 0 0.77fF $ **FLOATING
C2056 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n2 0 0.18fF $ **FLOATING
C2057 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n3 0 0.11fF $ **FLOATING
C2058 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t2 0 0.04fF
C2059 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t3 0 0.04fF
C2060 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n4 0 0.13fF $ **FLOATING
C2061 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n5 0 0.11fF $ **FLOATING
C2062 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t7 0 0.06fF
C2063 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t8 0 0.06fF
C2064 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t6 0 0.03fF
C2065 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n6 0 0.06fF $ **FLOATING
C2066 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n7 0 0.03fF $ **FLOATING
C2067 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/OUT_bar 0 0.01fF $ **FLOATING
C2068 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT_bar 0 0.35fF $ **FLOATING
C2069 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t7 0 0.11fF
C2070 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n0 0 0.43fF $ **FLOATING
C2071 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t2 0 0.04fF
C2072 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t3 0 0.04fF
C2073 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n1 0 0.12fF $ **FLOATING
C2074 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t4 0 0.15fF
C2075 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t5 0 0.27fF
C2076 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n2 0 0.23fF $ **FLOATING
C2077 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n3 0 0.10fF $ **FLOATING
C2078 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t0 0 0.04fF
C2079 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t1 0 0.04fF
C2080 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n4 0 0.10fF $ **FLOATING
C2081 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n5 0 0.11fF $ **FLOATING
C2082 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t6 0 0.04fF
C2083 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t9 0 0.05fF
C2084 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.t8 0 0.05fF
C2085 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n6 0 0.06fF $ **FLOATING
C2086 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A.n7 0 0.04fF $ **FLOATING
C2087 EESPFAL_Sbox_0/x0_bar 0 0.87fF $ **FLOATING
C2088 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_0/OUT_bar 0 0.73fF $ **FLOATING
C2089 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t12 0 0.42fF
C2090 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t14 0 0.23fF
C2091 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n0 0 2.19fF $ **FLOATING
C2092 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t8 0 0.53fF
C2093 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t9 0 0.18fF
C2094 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n1 0 1.78fF $ **FLOATING
C2095 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/B_bar 0 0.33fF $ **FLOATING
C2096 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t18 0 0.20fF
C2097 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B_bar 0 0.77fF $ **FLOATING
C2098 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t17 0 0.53fF
C2099 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t13 0 0.18fF
C2100 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n2 0 1.78fF $ **FLOATING
C2101 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/B_bar 0 0.32fF $ **FLOATING
C2102 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n3 0 6.07fF $ **FLOATING
C2103 EESPFAL_Sbox_0/EESPFAL_s3_0/x0_bar 0 0.75fF $ **FLOATING
C2104 EESPFAL_Sbox_0/EESPFAL_s2_0/x0_bar 0 1.79fF $ **FLOATING
C2105 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t15 0 0.53fF
C2106 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t16 0 0.18fF
C2107 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n4 0 1.78fF $ **FLOATING
C2108 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/B_bar 0 0.34fF $ **FLOATING
C2109 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n5 0 2.63fF $ **FLOATING
C2110 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t11 0 0.21fF
C2111 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/C_bar 0 0.69fF $ **FLOATING
C2112 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n6 0 2.60fF $ **FLOATING
C2113 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t7 0 0.48fF
C2114 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C 0 1.90fF $ **FLOATING
C2115 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n7 0 3.52fF $ **FLOATING
C2116 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n8 0 2.36fF $ **FLOATING
C2117 EESPFAL_Sbox_0/EESPFAL_s1_0/x0_bar 0 1.89fF $ **FLOATING
C2118 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n9 0 2.20fF $ **FLOATING
C2119 EESPFAL_4in_XOR_0/XOR0_bar 0 0.33fF $ **FLOATING
C2120 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t2 0 0.15fF
C2121 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t5 0 0.15fF
C2122 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n10 0 0.47fF $ **FLOATING
C2123 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t4 0 0.59fF
C2124 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t3 0 1.02fF
C2125 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n11 0 0.90fF $ **FLOATING
C2126 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n12 0 0.38fF $ **FLOATING
C2127 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t1 0 0.15fF
C2128 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t0 0 0.15fF
C2129 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n13 0 0.39fF $ **FLOATING
C2130 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n14 0 0.43fF $ **FLOATING
C2131 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t10 0 0.20fF
C2132 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t6 0 0.19fF
C2133 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.t19 0 0.14fF
C2134 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n15 0 0.22fF $ **FLOATING
C2135 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar.n16 0 0.16fF $ **FLOATING
C2136 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t9 0 0.04fF
C2137 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/A_bar 0 0.53fF $ **FLOATING
C2138 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t5 0 0.04fF
C2139 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t1 0 0.04fF
C2140 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n0 0 0.11fF $ **FLOATING
C2141 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t2 0 0.13fF
C2142 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t0 0 0.20fF
C2143 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n1 0 0.19fF $ **FLOATING
C2144 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n2 0 0.09fF $ **FLOATING
C2145 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t3 0 0.04fF
C2146 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t4 0 0.04fF
C2147 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n3 0 0.09fF $ **FLOATING
C2148 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n4 0 0.10fF $ **FLOATING
C2149 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t8 0 0.05fF
C2150 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t7 0 0.04fF
C2151 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t6 0 0.03fF
C2152 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n5 0 0.05fF $ **FLOATING
C2153 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n6 0 0.04fF $ **FLOATING
C2154 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t0 0 0.04fF
C2155 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t3 0 0.04fF
C2156 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n0 0 0.12fF $ **FLOATING
C2157 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t4 0 0.17fF
C2158 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t7 0 0.05fF
C2159 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n1 0 0.78fF $ **FLOATING
C2160 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n2 0 0.18fF $ **FLOATING
C2161 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n3 0 0.11fF $ **FLOATING
C2162 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t1 0 0.04fF
C2163 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t2 0 0.04fF
C2164 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n4 0 0.13fF $ **FLOATING
C2165 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n5 0 0.11fF $ **FLOATING
C2166 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t8 0 0.03fF
C2167 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t5 0 0.06fF
C2168 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t6 0 0.06fF
C2169 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n6 0 0.06fF $ **FLOATING
C2170 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n7 0 0.03fF $ **FLOATING
C2171 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/OUT_bar 0 0.01fF $ **FLOATING
C2172 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/OUT 0 0.23fF $ **FLOATING
C2173 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 0 0.03fF
C2174 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 0 0.63fF $ **FLOATING
C2175 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 0 0.04fF
C2176 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 0 0.04fF
C2177 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 0 0.11fF $ **FLOATING
C2178 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 0 0.25fF
C2179 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 0 0.04fF
C2180 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 0 0.04fF
C2181 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 0 0.13fF $ **FLOATING
C2182 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 0 0.17fF $ **FLOATING
C2183 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 0 0.12fF $ **FLOATING
C2184 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 0 0.04fF
C2185 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 0 0.06fF
C2186 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 0 0.05fF
C2187 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 0 0.06fF $ **FLOATING
C2188 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 0 0.04fF $ **FLOATING
C2189 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT_bar 0 0.30fF $ **FLOATING
C2190 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t6 0 0.12fF
C2191 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t4 0 0.04fF
C2192 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t2 0 0.04fF
C2193 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n0 0 0.11fF $ **FLOATING
C2194 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t3 0 0.17fF
C2195 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t1 0 0.29fF
C2196 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n1 0 0.26fF $ **FLOATING
C2197 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t5 0 0.04fF
C2198 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t0 0 0.04fF
C2199 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n2 0 0.13fF $ **FLOATING
C2200 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n3 0 0.11fF $ **FLOATING
C2201 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n4 0 0.12fF $ **FLOATING
C2202 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t9 0 0.06fF
C2203 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t7 0 0.05fF
C2204 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t8 0 0.04fF
C2205 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n5 0 0.06fF $ **FLOATING
C2206 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n6 0 0.04fF $ **FLOATING
C2207 EESPFAL_Sbox_0/EESPFAL_s0_0/Dis1 0 0.03fF $ **FLOATING
C2208 Dis1.t18 0 0.21fF
C2209 Dis1.t23 0 0.14fF
C2210 Dis1.n0 0 0.53fF $ **FLOATING
C2211 Dis1.t26 0 0.14fF
C2212 Dis1.n1 0 0.91fF $ **FLOATING
C2213 Dis1.t5 0 0.14fF
C2214 Dis1.n2 0 0.28fF $ **FLOATING
C2215 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/Dis 0 0.28fF $ **FLOATING
C2216 Dis1.t22 0 0.21fF
C2217 Dis1.t3 0 0.14fF
C2218 Dis1.n3 0 0.53fF $ **FLOATING
C2219 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/Dis 0 0.27fF $ **FLOATING
C2220 Dis1.t2 0 0.21fF
C2221 Dis1.t25 0 0.14fF
C2222 Dis1.n4 0 0.53fF $ **FLOATING
C2223 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/Dis 0 0.31fF $ **FLOATING
C2224 Dis1.t8 0 0.21fF
C2225 Dis1.t30 0 0.14fF
C2226 Dis1.n5 0 0.53fF $ **FLOATING
C2227 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_1/Dis 0 0.60fF $ **FLOATING
C2228 Dis1.t6 0 0.14fF
C2229 Dis1.n6 0 0.87fF $ **FLOATING
C2230 Dis1.t29 0 0.14fF
C2231 Dis1.n7 0 0.28fF $ **FLOATING
C2232 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/Dis 0 0.26fF $ **FLOATING
C2233 Dis1.n8 0 2.57fF $ **FLOATING
C2234 Dis1.t17 0 0.21fF
C2235 Dis1.t1 0 0.14fF
C2236 Dis1.n9 0 0.53fF $ **FLOATING
C2237 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/Dis 0 0.60fF $ **FLOATING
C2238 Dis1.t16 0 0.14fF
C2239 Dis1.n10 0 0.87fF $ **FLOATING
C2240 Dis1.t0 0 0.14fF
C2241 Dis1.n11 0 0.28fF $ **FLOATING
C2242 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/Dis 0 0.26fF $ **FLOATING
C2243 Dis1.n12 0 0.80fF $ **FLOATING
C2244 EESPFAL_Sbox_0/EESPFAL_s3_0/Dis1 0 0.58fF $ **FLOATING
C2245 EESPFAL_Sbox_0/EESPFAL_s2_0/Dis1 0 0.59fF $ **FLOATING
C2246 Dis1.t4 0 0.21fF
C2247 Dis1.t15 0 0.14fF
C2248 Dis1.n13 0 0.53fF $ **FLOATING
C2249 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/Dis 0 0.60fF $ **FLOATING
C2250 Dis1.t27 0 0.14fF
C2251 Dis1.n14 0 0.88fF $ **FLOATING
C2252 Dis1.t35 0 0.14fF
C2253 Dis1.n15 0 0.28fF $ **FLOATING
C2254 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/Dis 0 0.17fF $ **FLOATING
C2255 Dis1.n16 0 0.54fF $ **FLOATING
C2256 Dis1.t9 0 0.21fF
C2257 Dis1.t20 0 0.14fF
C2258 Dis1.n17 0 0.53fF $ **FLOATING
C2259 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/Dis 0 0.60fF $ **FLOATING
C2260 Dis1.t32 0 0.14fF
C2261 Dis1.n18 0 0.88fF $ **FLOATING
C2262 Dis1.t19 0 0.14fF
C2263 Dis1.n19 0 0.28fF $ **FLOATING
C2264 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/Dis 0 0.17fF $ **FLOATING
C2265 Dis1.n20 0 1.16fF $ **FLOATING
C2266 Dis1.t21 0 0.21fF
C2267 Dis1.t12 0 0.14fF
C2268 Dis1.n21 0 0.53fF $ **FLOATING
C2269 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/Dis 0 0.32fF $ **FLOATING
C2270 Dis1.n22 0 1.64fF $ **FLOATING
C2271 Dis1.n23 0 1.46fF $ **FLOATING
C2272 Dis1.t34 0 0.21fF
C2273 Dis1.t13 0 0.14fF
C2274 Dis1.n24 0 0.53fF $ **FLOATING
C2275 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/Dis 0 0.60fF $ **FLOATING
C2276 Dis1.t11 0 0.14fF
C2277 Dis1.n25 0 0.87fF $ **FLOATING
C2278 Dis1.t28 0 0.14fF
C2279 Dis1.n26 0 0.28fF $ **FLOATING
C2280 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/Dis 0 0.26fF $ **FLOATING
C2281 Dis1.n27 0 1.28fF $ **FLOATING
C2282 Dis1.t14 0 0.21fF
C2283 Dis1.t33 0 0.14fF
C2284 Dis1.n28 0 0.53fF $ **FLOATING
C2285 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/Dis 0 0.60fF $ **FLOATING
C2286 Dis1.t31 0 0.14fF
C2287 Dis1.n29 0 0.87fF $ **FLOATING
C2288 Dis1.t10 0 0.14fF
C2289 Dis1.n30 0 0.28fF $ **FLOATING
C2290 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/Dis 0 0.26fF $ **FLOATING
C2291 Dis1.n31 0 0.80fF $ **FLOATING
C2292 EESPFAL_Sbox_0/EESPFAL_s1_0/Dis1 0 0.84fF $ **FLOATING
C2293 Dis1.t7 0 0.21fF
C2294 Dis1.t24 0 0.14fF
C2295 Dis1.n32 0 0.53fF $ **FLOATING
C2296 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/Dis 0 0.28fF $ **FLOATING
C2297 Dis1.n33 0 1.07fF $ **FLOATING
C2298 Dis1.n34 0 0.82fF $ **FLOATING
C2299 EESPFAL_Sbox_0/Dis1 0 0.33fF $ **FLOATING
C2300 EESPFAL_Sbox_0/EESPFAL_s3_0/s3 0 0.01fF $ **FLOATING
C2301 s3.t4 0 0.04fF
C2302 s3.t5 0 0.04fF
C2303 s3.n0 0 0.15fF $ **FLOATING
C2304 s3.t1 0 0.19fF
C2305 s3.t3 0 0.04fF
C2306 s3.t6 0 0.04fF
C2307 s3.n1 0 0.14fF $ **FLOATING
C2308 s3.t2 0 0.04fF
C2309 s3.t0 0 0.04fF
C2310 s3.n2 0 0.15fF $ **FLOATING
C2311 s3.t9 0 0.06fF
C2312 s3.t7 0 0.06fF
C2313 s3.t8 0 0.03fF
C2314 s3.n3 0 0.06fF $ **FLOATING
C2315 s3.n4 0 0.20fF $ **FLOATING
C2316 s3.n5 0 0.17fF $ **FLOATING
C2317 s3.n6 0 0.14fF $ **FLOATING
C2318 EESPFAL_Sbox_0/s3 0 0.48fF $ **FLOATING
C2319 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/OUT 0 0.23fF $ **FLOATING
C2320 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 0 0.03fF
C2321 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 0 0.63fF $ **FLOATING
C2322 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 0 0.04fF
C2323 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 0 0.04fF
C2324 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 0 0.11fF $ **FLOATING
C2325 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 0 0.25fF
C2326 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 0 0.04fF
C2327 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 0 0.04fF
C2328 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 0 0.13fF $ **FLOATING
C2329 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 0 0.17fF $ **FLOATING
C2330 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 0 0.12fF $ **FLOATING
C2331 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 0 0.06fF
C2332 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 0 0.05fF
C2333 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 0 0.04fF
C2334 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 0 0.06fF $ **FLOATING
C2335 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 0 0.04fF $ **FLOATING
C2336 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t1 0 0.04fF
C2337 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t4 0 0.04fF
C2338 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n0 0 0.13fF $ **FLOATING
C2339 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t3 0 0.16fF
C2340 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t6 0 0.05fF
C2341 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n1 0 0.77fF $ **FLOATING
C2342 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n2 0 0.18fF $ **FLOATING
C2343 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t0 0 0.04fF
C2344 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t2 0 0.04fF
C2345 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n3 0 0.12fF $ **FLOATING
C2346 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n4 0 0.11fF $ **FLOATING
C2347 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n5 0 0.11fF $ **FLOATING
C2348 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t7 0 0.06fF
C2349 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t8 0 0.06fF
C2350 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t5 0 0.03fF
C2351 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n6 0 0.06fF $ **FLOATING
C2352 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n7 0 0.03fF $ **FLOATING
C2353 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/OUT_bar 0 0.01fF $ **FLOATING
C2354 CLK2.t61 0 0.04fF
C2355 CLK2.t86 0 0.03fF
C2356 CLK2.t59 0 0.03fF
C2357 CLK2.n0 0 0.08fF $ **FLOATING
C2358 CLK2.t84 0 0.04fF
C2359 CLK2.t98 0 0.06fF
C2360 CLK2.n1 0 0.09fF $ **FLOATING
C2361 CLK2.n2 0 0.26fF $ **FLOATING
C2362 CLK2.n3 0 0.05fF $ **FLOATING
C2363 CLK2.n4 0 0.02fF $ **FLOATING
C2364 CLK2.n5 0 0.02fF $ **FLOATING
C2365 CLK2.n6 0 0.02fF $ **FLOATING
C2366 CLK2.n7 0 0.04fF $ **FLOATING
C2367 CLK2.n8 0 0.02fF $ **FLOATING
C2368 CLK2.n9 0 0.02fF $ **FLOATING
C2369 CLK2.n10 0 0.02fF $ **FLOATING
C2370 CLK2.n11 0 0.04fF $ **FLOATING
C2371 CLK2.n12 0 0.02fF $ **FLOATING
C2372 CLK2.n13 0 0.02fF $ **FLOATING
C2373 CLK2.n14 0 0.02fF $ **FLOATING
C2374 CLK2.n15 0 0.04fF $ **FLOATING
C2375 CLK2.n16 0 0.02fF $ **FLOATING
C2376 CLK2.n17 0 0.02fF $ **FLOATING
C2377 CLK2.n18 0 0.02fF $ **FLOATING
C2378 CLK2.n19 0 0.10fF $ **FLOATING
C2379 CLK2.n20 0 0.02fF $ **FLOATING
C2380 CLK2.n21 0 0.02fF $ **FLOATING
C2381 CLK2.n22 0 0.02fF $ **FLOATING
C2382 CLK2.n23 0 0.13fF $ **FLOATING
C2383 CLK2.n24 0 0.02fF $ **FLOATING
C2384 CLK2.n25 0 0.02fF $ **FLOATING
C2385 CLK2.n26 0 0.01fF $ **FLOATING
C2386 CLK2.n27 0 0.21fF $ **FLOATING
C2387 CLK2.t83 0 0.06fF
C2388 CLK2.n28 0 0.08fF $ **FLOATING
C2389 CLK2.n29 0 0.02fF $ **FLOATING
C2390 CLK2.n30 0 0.02fF $ **FLOATING
C2391 CLK2.n31 0 0.02fF $ **FLOATING
C2392 CLK2.n32 0 0.12fF $ **FLOATING
C2393 CLK2.n33 0 0.02fF $ **FLOATING
C2394 CLK2.n34 0 0.02fF $ **FLOATING
C2395 CLK2.n35 0 0.02fF $ **FLOATING
C2396 CLK2.t85 0 0.06fF
C2397 CLK2.n36 0 0.07fF $ **FLOATING
C2398 CLK2.n37 0 0.02fF $ **FLOATING
C2399 CLK2.n38 0 0.02fF $ **FLOATING
C2400 CLK2.n39 0 0.02fF $ **FLOATING
C2401 CLK2.n40 0 0.13fF $ **FLOATING
C2402 CLK2.n41 0 0.12fF $ **FLOATING
C2403 CLK2.n42 0 0.02fF $ **FLOATING
C2404 CLK2.n43 0 0.02fF $ **FLOATING
C2405 CLK2.t58 0 0.06fF
C2406 CLK2.n44 0 0.07fF $ **FLOATING
C2407 CLK2.n45 0 0.02fF $ **FLOATING
C2408 CLK2.n46 0 0.02fF $ **FLOATING
C2409 CLK2.n47 0 0.02fF $ **FLOATING
C2410 CLK2.n48 0 0.12fF $ **FLOATING
C2411 CLK2.n49 0 0.02fF $ **FLOATING
C2412 CLK2.n50 0 0.02fF $ **FLOATING
C2413 CLK2.n51 0 0.02fF $ **FLOATING
C2414 CLK2.t60 0 0.06fF
C2415 CLK2.n52 0 0.08fF $ **FLOATING
C2416 CLK2.n53 0 0.02fF $ **FLOATING
C2417 CLK2.n54 0 0.02fF $ **FLOATING
C2418 CLK2.n55 0 0.02fF $ **FLOATING
C2419 CLK2.n56 0 0.21fF $ **FLOATING
C2420 CLK2.n57 0 0.13fF $ **FLOATING
C2421 CLK2.n58 0 0.02fF $ **FLOATING
C2422 CLK2.n59 0 0.02fF $ **FLOATING
C2423 CLK2.n60 0 0.01fF $ **FLOATING
C2424 CLK2.n61 0 0.10fF $ **FLOATING
C2425 CLK2.n62 0 0.02fF $ **FLOATING
C2426 CLK2.n63 0 0.02fF $ **FLOATING
C2427 CLK2.n64 0 0.02fF $ **FLOATING
C2428 CLK2.n65 0 0.04fF $ **FLOATING
C2429 CLK2.n66 0 0.02fF $ **FLOATING
C2430 CLK2.n67 0 0.02fF $ **FLOATING
C2431 CLK2.n68 0 0.02fF $ **FLOATING
C2432 CLK2.n69 0 0.04fF $ **FLOATING
C2433 CLK2.n70 0 0.02fF $ **FLOATING
C2434 CLK2.n71 0 0.02fF $ **FLOATING
C2435 CLK2.n72 0 0.02fF $ **FLOATING
C2436 CLK2.n73 0 0.01fF $ **FLOATING
C2437 CLK2.n74 0 0.02fF $ **FLOATING
C2438 CLK2.n75 0 0.04fF $ **FLOATING
C2439 CLK2.n76 0 0.02fF $ **FLOATING
C2440 CLK2.n77 0 0.01fF $ **FLOATING
C2441 CLK2.n78 0 0.05fF $ **FLOATING
C2442 CLK2.n79 0 0.02fF $ **FLOATING
C2443 CLK2.t19 0 0.03fF
C2444 CLK2.t0 0 0.03fF
C2445 CLK2.n80 0 0.11fF $ **FLOATING
C2446 CLK2.t31 0 0.04fF
C2447 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/CLK 0 0.01fF $ **FLOATING
C2448 CLK2.n81 0 0.12fF $ **FLOATING
C2449 CLK2.n82 0 0.02fF $ **FLOATING
C2450 CLK2.t93 0 0.03fF
C2451 CLK2.t29 0 0.03fF
C2452 CLK2.n83 0 0.08fF $ **FLOATING
C2453 CLK2.t91 0 0.04fF
C2454 CLK2.t56 0 0.03fF
C2455 CLK2.n84 0 0.08fF $ **FLOATING
C2456 CLK2.n85 0 0.01fF $ **FLOATING
C2457 CLK2.n86 0 0.02fF $ **FLOATING
C2458 CLK2.n87 0 0.02fF $ **FLOATING
C2459 CLK2.n88 0 0.09fF $ **FLOATING
C2460 CLK2.t42 0 0.04fF
C2461 CLK2.t44 0 0.03fF
C2462 CLK2.t108 0 0.03fF
C2463 CLK2.n89 0 0.08fF $ **FLOATING
C2464 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/CLK 0 0.01fF $ **FLOATING
C2465 CLK2.t110 0 0.04fF
C2466 CLK2.t62 0 0.03fF
C2467 CLK2.t4 0 0.03fF
C2468 CLK2.n90 0 0.11fF $ **FLOATING
C2469 CLK2.n91 0 0.09fF $ **FLOATING
C2470 CLK2.n92 0 0.11fF $ **FLOATING
C2471 CLK2.t3 0 0.03fF
C2472 CLK2.n93 0 0.08fF $ **FLOATING
C2473 CLK2.n94 0 0.01fF $ **FLOATING
C2474 CLK2.n95 0 0.02fF $ **FLOATING
C2475 CLK2.t51 0 0.03fF
C2476 CLK2.n96 0 0.08fF $ **FLOATING
C2477 CLK2.n97 0 0.01fF $ **FLOATING
C2478 CLK2.n98 0 0.02fF $ **FLOATING
C2479 CLK2.n99 0 0.11fF $ **FLOATING
C2480 CLK2.t2 0 0.03fF
C2481 CLK2.t55 0 0.03fF
C2482 CLK2.n100 0 0.11fF $ **FLOATING
C2483 CLK2.t21 0 0.04fF
C2484 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/CLK 0 0.01fF $ **FLOATING
C2485 CLK2.t25 0 0.03fF
C2486 CLK2.t23 0 0.03fF
C2487 CLK2.n101 0 0.08fF $ **FLOATING
C2488 CLK2.t27 0 0.04fF
C2489 CLK2.n102 0 0.02fF $ **FLOATING
C2490 CLK2.n103 0 0.02fF $ **FLOATING
C2491 CLK2.n104 0 0.09fF $ **FLOATING
C2492 CLK2.t112 0 0.04fF
C2493 CLK2.t114 0 0.03fF
C2494 CLK2.t34 0 0.03fF
C2495 CLK2.n105 0 0.08fF $ **FLOATING
C2496 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/CLK 0 0.01fF $ **FLOATING
C2497 CLK2.t36 0 0.04fF
C2498 CLK2.n106 0 0.04fF $ **FLOATING
C2499 CLK2.n107 0 0.02fF $ **FLOATING
C2500 CLK2.n108 0 0.02fF $ **FLOATING
C2501 CLK2.n109 0 0.01fF $ **FLOATING
C2502 CLK2.n110 0 0.00fF $ **FLOATING
C2503 CLK2.n111 0 0.01fF $ **FLOATING
C2504 CLK2.n112 0 0.00fF $ **FLOATING
C2505 CLK2.n113 0 0.00fF $ **FLOATING
C2506 CLK2.n114 0 0.02fF $ **FLOATING
C2507 CLK2.n115 0 0.02fF $ **FLOATING
C2508 CLK2.t52 0 0.03fF
C2509 CLK2.t82 0 0.03fF
C2510 CLK2.n116 0 0.11fF $ **FLOATING
C2511 CLK2.n117 0 0.05fF $ **FLOATING
C2512 CLK2.n118 0 0.10fF $ **FLOATING
C2513 CLK2.n119 0 0.02fF $ **FLOATING
C2514 CLK2.n120 0 0.02fF $ **FLOATING
C2515 CLK2.n121 0 0.01fF $ **FLOATING
C2516 CLK2.t75 0 0.04fF
C2517 CLK2.n122 0 0.02fF $ **FLOATING
C2518 CLK2.n123 0 0.02fF $ **FLOATING
C2519 CLK2.n124 0 0.02fF $ **FLOATING
C2520 CLK2.t72 0 0.06fF
C2521 CLK2.n125 0 0.02fF $ **FLOATING
C2522 CLK2.n126 0 0.02fF $ **FLOATING
C2523 CLK2.t14 0 0.03fF
C2524 CLK2.t73 0 0.03fF
C2525 CLK2.n127 0 0.08fF $ **FLOATING
C2526 CLK2.n128 0 0.02fF $ **FLOATING
C2527 CLK2.n129 0 0.02fF $ **FLOATING
C2528 CLK2.n130 0 0.02fF $ **FLOATING
C2529 CLK2.n131 0 0.13fF $ **FLOATING
C2530 CLK2.n132 0 0.02fF $ **FLOATING
C2531 CLK2.n133 0 0.02fF $ **FLOATING
C2532 CLK2.t12 0 0.04fF
C2533 CLK2.n134 0 0.02fF $ **FLOATING
C2534 CLK2.n135 0 0.02fF $ **FLOATING
C2535 CLK2.n136 0 0.02fF $ **FLOATING
C2536 CLK2.n137 0 0.04fF $ **FLOATING
C2537 CLK2.n138 0 0.02fF $ **FLOATING
C2538 CLK2.n139 0 0.02fF $ **FLOATING
C2539 CLK2.n140 0 0.01fF $ **FLOATING
C2540 CLK2.n141 0 0.01fF $ **FLOATING
C2541 CLK2.n142 0 0.02fF $ **FLOATING
C2542 CLK2.n143 0 0.02fF $ **FLOATING
C2543 CLK2.t106 0 0.03fF
C2544 CLK2.n144 0 0.09fF $ **FLOATING
C2545 CLK2.n145 0 0.02fF $ **FLOATING
C2546 CLK2.n146 0 0.02fF $ **FLOATING
C2547 CLK2.n147 0 0.02fF $ **FLOATING
C2548 CLK2.n148 0 0.04fF $ **FLOATING
C2549 CLK2.n149 0 0.02fF $ **FLOATING
C2550 CLK2.n150 0 0.02fF $ **FLOATING
C2551 CLK2.n151 0 0.01fF $ **FLOATING
C2552 CLK2.n152 0 0.02fF $ **FLOATING
C2553 CLK2.n153 0 0.02fF $ **FLOATING
C2554 CLK2.t45 0 0.06fF
C2555 CLK2.n154 0 0.02fF $ **FLOATING
C2556 CLK2.n155 0 0.02fF $ **FLOATING
C2557 CLK2.t46 0 0.04fF
C2558 CLK2.n156 0 0.21fF $ **FLOATING
C2559 CLK2.t48 0 0.03fF
C2560 CLK2.t68 0 0.03fF
C2561 CLK2.n157 0 0.08fF $ **FLOATING
C2562 CLK2.n158 0 0.13fF $ **FLOATING
C2563 CLK2.n159 0 0.02fF $ **FLOATING
C2564 CLK2.n160 0 0.02fF $ **FLOATING
C2565 CLK2.n161 0 0.12fF $ **FLOATING
C2566 CLK2.n162 0 0.12fF $ **FLOATING
C2567 CLK2.n163 0 0.02fF $ **FLOATING
C2568 CLK2.n164 0 0.02fF $ **FLOATING
C2569 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/CLK 0 0.01fF $ **FLOATING
C2570 CLK2.t70 0 0.04fF
C2571 CLK2.n165 0 0.21fF $ **FLOATING
C2572 CLK2.n166 0 0.02fF $ **FLOATING
C2573 CLK2.n167 0 0.02fF $ **FLOATING
C2574 CLK2.t69 0 0.06fF
C2575 CLK2.n168 0 0.04fF $ **FLOATING
C2576 CLK2.n169 0 0.02fF $ **FLOATING
C2577 CLK2.n170 0 0.02fF $ **FLOATING
C2578 CLK2.n171 0 0.01fF $ **FLOATING
C2579 CLK2.t7 0 0.03fF
C2580 CLK2.t15 0 0.03fF
C2581 CLK2.n172 0 0.11fF $ **FLOATING
C2582 CLK2.n173 0 0.14fF $ **FLOATING
C2583 CLK2.n174 0 0.02fF $ **FLOATING
C2584 CLK2.n175 0 0.02fF $ **FLOATING
C2585 CLK2.n176 0 0.09fF $ **FLOATING
C2586 CLK2.n177 0 0.01fF $ **FLOATING
C2587 CLK2.n178 0 0.11fF $ **FLOATING
C2588 CLK2.t87 0 0.05fF
C2589 CLK2.n179 0 0.02fF $ **FLOATING
C2590 CLK2.n180 0 0.02fF $ **FLOATING
C2591 CLK2.n181 0 0.02fF $ **FLOATING
C2592 CLK2.n182 0 0.13fF $ **FLOATING
C2593 CLK2.n183 0 0.02fF $ **FLOATING
C2594 CLK2.n184 0 0.02fF $ **FLOATING
C2595 CLK2.t6 0 0.04fF
C2596 CLK2.n185 0 0.02fF $ **FLOATING
C2597 CLK2.n186 0 0.02fF $ **FLOATING
C2598 CLK2.n187 0 0.02fF $ **FLOATING
C2599 CLK2.t116 0 0.06fF
C2600 CLK2.n188 0 0.02fF $ **FLOATING
C2601 CLK2.n189 0 0.02fF $ **FLOATING
C2602 CLK2.t117 0 0.03fF
C2603 CLK2.t97 0 0.03fF
C2604 CLK2.n190 0 0.08fF $ **FLOATING
C2605 CLK2.n191 0 0.02fF $ **FLOATING
C2606 CLK2.n192 0 0.02fF $ **FLOATING
C2607 CLK2.n193 0 0.02fF $ **FLOATING
C2608 CLK2.n194 0 0.12fF $ **FLOATING
C2609 CLK2.t96 0 0.06fF
C2610 CLK2.n195 0 0.13fF $ **FLOATING
C2611 CLK2.n196 0 0.02fF $ **FLOATING
C2612 CLK2.n197 0 0.02fF $ **FLOATING
C2613 CLK2.t18 0 0.04fF
C2614 CLK2.n198 0 0.02fF $ **FLOATING
C2615 CLK2.n199 0 0.02fF $ **FLOATING
C2616 CLK2.n200 0 0.02fF $ **FLOATING
C2617 CLK2.n201 0 0.11fF $ **FLOATING
C2618 CLK2.t65 0 0.05fF
C2619 CLK2.n202 0 0.34fF $ **FLOATING
C2620 CLK2.n203 0 0.02fF $ **FLOATING
C2621 CLK2.n204 0 0.02fF $ **FLOATING
C2622 CLK2.n205 0 0.02fF $ **FLOATING
C2623 CLK2.n206 0 0.05fF $ **FLOATING
C2624 CLK2.n207 0 0.04fF $ **FLOATING
C2625 CLK2.n208 0 0.10fF $ **FLOATING
C2626 CLK2.n209 0 0.02fF $ **FLOATING
C2627 CLK2.n210 0 0.02fF $ **FLOATING
C2628 CLK2.n211 0 0.02fF $ **FLOATING
C2629 CLK2.n212 0 0.01fF $ **FLOATING
C2630 CLK2.n213 0 0.21fF $ **FLOATING
C2631 CLK2.n214 0 0.02fF $ **FLOATING
C2632 CLK2.n215 0 0.02fF $ **FLOATING
C2633 CLK2.n216 0 0.02fF $ **FLOATING
C2634 CLK2.n217 0 0.08fF $ **FLOATING
C2635 CLK2.t17 0 0.06fF
C2636 CLK2.n218 0 0.12fF $ **FLOATING
C2637 CLK2.n219 0 0.07fF $ **FLOATING
C2638 CLK2.n220 0 0.02fF $ **FLOATING
C2639 CLK2.n221 0 0.02fF $ **FLOATING
C2640 CLK2.n222 0 0.02fF $ **FLOATING
C2641 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/CLK 0 0.01fF $ **FLOATING
C2642 CLK2.n223 0 0.13fF $ **FLOATING
C2643 CLK2.n224 0 0.02fF $ **FLOATING
C2644 CLK2.n225 0 0.02fF $ **FLOATING
C2645 CLK2.n226 0 0.02fF $ **FLOATING
C2646 CLK2.n227 0 0.07fF $ **FLOATING
C2647 CLK2.n228 0 0.12fF $ **FLOATING
C2648 CLK2.t5 0 0.06fF
C2649 CLK2.n229 0 0.08fF $ **FLOATING
C2650 CLK2.n230 0 0.02fF $ **FLOATING
C2651 CLK2.n231 0 0.02fF $ **FLOATING
C2652 CLK2.n232 0 0.02fF $ **FLOATING
C2653 CLK2.n233 0 0.21fF $ **FLOATING
C2654 CLK2.n234 0 0.01fF $ **FLOATING
C2655 CLK2.n235 0 0.02fF $ **FLOATING
C2656 CLK2.n236 0 0.02fF $ **FLOATING
C2657 CLK2.n237 0 0.02fF $ **FLOATING
C2658 CLK2.n238 0 0.10fF $ **FLOATING
C2659 CLK2.n239 0 0.04fF $ **FLOATING
C2660 CLK2.n240 0 0.05fF $ **FLOATING
C2661 CLK2.n241 0 0.02fF $ **FLOATING
C2662 CLK2.n242 0 0.02fF $ **FLOATING
C2663 CLK2.n243 0 0.02fF $ **FLOATING
C2664 CLK2.n244 0 0.32fF $ **FLOATING
C2665 CLK2.n245 0 0.15fF $ **FLOATING
C2666 CLK2.n246 0 0.15fF $ **FLOATING
C2667 CLK2.n247 0 0.02fF $ **FLOATING
C2668 CLK2.n248 0 0.02fF $ **FLOATING
C2669 CLK2.n249 0 0.02fF $ **FLOATING
C2670 CLK2.n250 0 0.05fF $ **FLOATING
C2671 CLK2.n251 0 0.04fF $ **FLOATING
C2672 CLK2.n252 0 0.04fF $ **FLOATING
C2673 CLK2.n253 0 0.02fF $ **FLOATING
C2674 CLK2.n254 0 0.02fF $ **FLOATING
C2675 CLK2.n255 0 0.02fF $ **FLOATING
C2676 CLK2.n256 0 0.02fF $ **FLOATING
C2677 CLK2.n257 0 0.02fF $ **FLOATING
C2678 CLK2.n258 0 0.02fF $ **FLOATING
C2679 CLK2.n259 0 0.02fF $ **FLOATING
C2680 CLK2.n260 0 0.10fF $ **FLOATING
C2681 CLK2.n261 0 0.13fF $ **FLOATING
C2682 CLK2.n262 0 0.08fF $ **FLOATING
C2683 CLK2.n263 0 0.02fF $ **FLOATING
C2684 CLK2.n264 0 0.02fF $ **FLOATING
C2685 CLK2.n265 0 0.02fF $ **FLOATING
C2686 CLK2.n266 0 0.02fF $ **FLOATING
C2687 CLK2.n267 0 0.02fF $ **FLOATING
C2688 CLK2.n268 0 0.02fF $ **FLOATING
C2689 CLK2.n269 0 0.02fF $ **FLOATING
C2690 CLK2.n270 0 0.07fF $ **FLOATING
C2691 CLK2.t67 0 0.06fF
C2692 CLK2.n271 0 0.12fF $ **FLOATING
C2693 CLK2.t47 0 0.06fF
C2694 CLK2.n272 0 0.07fF $ **FLOATING
C2695 CLK2.n273 0 0.02fF $ **FLOATING
C2696 CLK2.n274 0 0.02fF $ **FLOATING
C2697 CLK2.n275 0 0.02fF $ **FLOATING
C2698 CLK2.n276 0 0.02fF $ **FLOATING
C2699 CLK2.n277 0 0.02fF $ **FLOATING
C2700 CLK2.n278 0 0.02fF $ **FLOATING
C2701 CLK2.n279 0 0.02fF $ **FLOATING
C2702 CLK2.n280 0 0.08fF $ **FLOATING
C2703 CLK2.n281 0 0.13fF $ **FLOATING
C2704 CLK2.n282 0 0.10fF $ **FLOATING
C2705 CLK2.n283 0 0.02fF $ **FLOATING
C2706 CLK2.n284 0 0.02fF $ **FLOATING
C2707 CLK2.n285 0 0.02fF $ **FLOATING
C2708 CLK2.n286 0 0.02fF $ **FLOATING
C2709 CLK2.n287 0 0.02fF $ **FLOATING
C2710 CLK2.n288 0 0.02fF $ **FLOATING
C2711 CLK2.n289 0 0.02fF $ **FLOATING
C2712 CLK2.n290 0 0.04fF $ **FLOATING
C2713 CLK2.n291 0 0.04fF $ **FLOATING
C2714 CLK2.n292 0 0.05fF $ **FLOATING
C2715 CLK2.n293 0 0.02fF $ **FLOATING
C2716 CLK2.n294 0 0.02fF $ **FLOATING
C2717 CLK2.n295 0 0.02fF $ **FLOATING
C2718 CLK2.n296 0 0.06fF $ **FLOATING
C2719 CLK2.n297 0 0.06fF $ **FLOATING
C2720 CLK2.n298 0 0.02fF $ **FLOATING
C2721 CLK2.n299 0 0.08fF $ **FLOATING
C2722 CLK2.n300 0 0.01fF $ **FLOATING
C2723 CLK2.n301 0 0.09fF $ **FLOATING
C2724 CLK2.n302 0 0.08fF $ **FLOATING
C2725 CLK2.t8 0 0.03fF
C2726 CLK2.n303 0 0.08fF $ **FLOATING
C2727 CLK2.n304 0 0.02fF $ **FLOATING
C2728 CLK2.n305 0 0.02fF $ **FLOATING
C2729 CLK2.n306 0 0.02fF $ **FLOATING
C2730 CLK2.n307 0 0.07fF $ **FLOATING
C2731 CLK2.n308 0 0.04fF $ **FLOATING
C2732 EESPFAL_Sbox_0/EESPFAL_s3_0/CLK2 0 0.02fF $ **FLOATING
C2733 CLK2.n309 0 0.01fF $ **FLOATING
C2734 CLK2.n310 0 0.09fF $ **FLOATING
C2735 CLK2.n311 0 0.05fF $ **FLOATING
C2736 CLK2.n312 0 0.02fF $ **FLOATING
C2737 CLK2.n313 0 0.02fF $ **FLOATING
C2738 CLK2.n314 0 0.02fF $ **FLOATING
C2739 CLK2.n315 0 0.02fF $ **FLOATING
C2740 CLK2.n316 0 0.02fF $ **FLOATING
C2741 CLK2.n317 0 0.02fF $ **FLOATING
C2742 CLK2.n318 0 0.02fF $ **FLOATING
C2743 CLK2.n319 0 0.04fF $ **FLOATING
C2744 CLK2.n320 0 0.04fF $ **FLOATING
C2745 CLK2.n321 0 0.10fF $ **FLOATING
C2746 CLK2.n322 0 0.02fF $ **FLOATING
C2747 CLK2.n323 0 0.02fF $ **FLOATING
C2748 CLK2.n324 0 0.02fF $ **FLOATING
C2749 CLK2.n325 0 0.01fF $ **FLOATING
C2750 CLK2.n326 0 0.21fF $ **FLOATING
C2751 CLK2.n327 0 0.02fF $ **FLOATING
C2752 CLK2.n328 0 0.02fF $ **FLOATING
C2753 CLK2.n329 0 0.02fF $ **FLOATING
C2754 CLK2.n330 0 0.08fF $ **FLOATING
C2755 CLK2.t11 0 0.06fF
C2756 CLK2.n331 0 0.12fF $ **FLOATING
C2757 CLK2.n332 0 0.12fF $ **FLOATING
C2758 CLK2.t13 0 0.06fF
C2759 CLK2.n333 0 0.07fF $ **FLOATING
C2760 CLK2.n334 0 0.02fF $ **FLOATING
C2761 CLK2.n335 0 0.02fF $ **FLOATING
C2762 CLK2.n336 0 0.02fF $ **FLOATING
C2763 CLK2.n337 0 0.13fF $ **FLOATING
C2764 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/CLK 0 0.01fF $ **FLOATING
C2765 CLK2.n338 0 0.02fF $ **FLOATING
C2766 CLK2.n339 0 0.02fF $ **FLOATING
C2767 CLK2.n340 0 0.02fF $ **FLOATING
C2768 CLK2.n341 0 0.07fF $ **FLOATING
C2769 CLK2.n342 0 0.12fF $ **FLOATING
C2770 CLK2.t74 0 0.06fF
C2771 CLK2.n343 0 0.13fF $ **FLOATING
C2772 CLK2.n344 0 0.08fF $ **FLOATING
C2773 CLK2.n345 0 0.02fF $ **FLOATING
C2774 CLK2.n346 0 0.02fF $ **FLOATING
C2775 CLK2.n347 0 0.02fF $ **FLOATING
C2776 CLK2.n348 0 0.21fF $ **FLOATING
C2777 CLK2.n349 0 0.01fF $ **FLOATING
C2778 CLK2.n350 0 0.01fF $ **FLOATING
C2779 CLK2.n351 0 0.02fF $ **FLOATING
C2780 CLK2.n352 0 0.02fF $ **FLOATING
C2781 CLK2.n353 0 0.02fF $ **FLOATING
C2782 CLK2.n354 0 0.02fF $ **FLOATING
C2783 CLK2.n355 0 0.04fF $ **FLOATING
C2784 CLK2.n356 0 0.04fF $ **FLOATING
C2785 CLK2.n357 0 0.04fF $ **FLOATING
C2786 CLK2.n358 0 0.02fF $ **FLOATING
C2787 CLK2.n359 0 0.02fF $ **FLOATING
C2788 CLK2.n360 0 0.02fF $ **FLOATING
C2789 CLK2.n361 0 0.09fF $ **FLOATING
C2790 CLK2.n362 0 0.05fF $ **FLOATING
C2791 CLK2.n363 0 0.14fF $ **FLOATING
C2792 CLK2.n364 0 0.02fF $ **FLOATING
C2793 CLK2.n365 0 0.02fF $ **FLOATING
C2794 CLK2.n366 0 0.01fF $ **FLOATING
C2795 CLK2.n367 0 0.00fF $ **FLOATING
C2796 CLK2.n369 0 0.01fF $ **FLOATING
C2797 CLK2.n370 0 0.05fF $ **FLOATING
C2798 EESPFAL_Sbox_0/EESPFAL_s2_0/CLK2 0 0.05fF $ **FLOATING
C2799 CLK2.n371 0 0.00fF $ **FLOATING
C2800 CLK2.t1 0 0.03fF
C2801 CLK2.t50 0 0.03fF
C2802 CLK2.n372 0 0.11fF $ **FLOATING
C2803 CLK2.n373 0 0.05fF $ **FLOATING
C2804 CLK2.n374 0 0.02fF $ **FLOATING
C2805 CLK2.n375 0 0.02fF $ **FLOATING
C2806 CLK2.n376 0 0.09fF $ **FLOATING
C2807 CLK2.n377 0 0.04fF $ **FLOATING
C2808 CLK2.n378 0 0.02fF $ **FLOATING
C2809 CLK2.n379 0 0.02fF $ **FLOATING
C2810 CLK2.n380 0 0.05fF $ **FLOATING
C2811 CLK2.n381 0 0.14fF $ **FLOATING
C2812 CLK2.n382 0 0.01fF $ **FLOATING
C2813 CLK2.n383 0 0.04fF $ **FLOATING
C2814 CLK2.n384 0 0.02fF $ **FLOATING
C2815 CLK2.n385 0 0.02fF $ **FLOATING
C2816 CLK2.n386 0 0.00fF $ **FLOATING
C2817 CLK2.n387 0 0.00fF $ **FLOATING
C2818 CLK2.n388 0 0.01fF $ **FLOATING
C2819 CLK2.n389 0 0.02fF $ **FLOATING
C2820 CLK2.n390 0 0.10fF $ **FLOATING
C2821 CLK2.n391 0 0.02fF $ **FLOATING
C2822 CLK2.n392 0 0.02fF $ **FLOATING
C2823 CLK2.n393 0 0.02fF $ **FLOATING
C2824 CLK2.n394 0 0.13fF $ **FLOATING
C2825 CLK2.n395 0 0.02fF $ **FLOATING
C2826 CLK2.n396 0 0.02fF $ **FLOATING
C2827 CLK2.n397 0 0.01fF $ **FLOATING
C2828 CLK2.n398 0 0.21fF $ **FLOATING
C2829 CLK2.t35 0 0.06fF
C2830 CLK2.n399 0 0.08fF $ **FLOATING
C2831 CLK2.n400 0 0.02fF $ **FLOATING
C2832 CLK2.n401 0 0.02fF $ **FLOATING
C2833 CLK2.n402 0 0.02fF $ **FLOATING
C2834 CLK2.n403 0 0.12fF $ **FLOATING
C2835 CLK2.n404 0 0.02fF $ **FLOATING
C2836 CLK2.n405 0 0.02fF $ **FLOATING
C2837 CLK2.n406 0 0.02fF $ **FLOATING
C2838 CLK2.n407 0 0.02fF $ **FLOATING
C2839 CLK2.t33 0 0.06fF
C2840 CLK2.n408 0 0.07fF $ **FLOATING
C2841 CLK2.n409 0 0.02fF $ **FLOATING
C2842 CLK2.n410 0 0.02fF $ **FLOATING
C2843 CLK2.n411 0 0.12fF $ **FLOATING
C2844 CLK2.n412 0 0.02fF $ **FLOATING
C2845 CLK2.n413 0 0.02fF $ **FLOATING
C2846 CLK2.n414 0 0.13fF $ **FLOATING
C2847 CLK2.t113 0 0.06fF
C2848 CLK2.n415 0 0.07fF $ **FLOATING
C2849 CLK2.n416 0 0.02fF $ **FLOATING
C2850 CLK2.n417 0 0.02fF $ **FLOATING
C2851 CLK2.n418 0 0.02fF $ **FLOATING
C2852 CLK2.n419 0 0.12fF $ **FLOATING
C2853 CLK2.n420 0 0.02fF $ **FLOATING
C2854 CLK2.n421 0 0.02fF $ **FLOATING
C2855 CLK2.n422 0 0.02fF $ **FLOATING
C2856 CLK2.t111 0 0.06fF
C2857 CLK2.n423 0 0.08fF $ **FLOATING
C2858 CLK2.n424 0 0.02fF $ **FLOATING
C2859 CLK2.n425 0 0.02fF $ **FLOATING
C2860 CLK2.n426 0 0.02fF $ **FLOATING
C2861 CLK2.n427 0 0.21fF $ **FLOATING
C2862 CLK2.n428 0 0.13fF $ **FLOATING
C2863 CLK2.n429 0 0.02fF $ **FLOATING
C2864 CLK2.n430 0 0.02fF $ **FLOATING
C2865 CLK2.n431 0 0.01fF $ **FLOATING
C2866 CLK2.n432 0 0.10fF $ **FLOATING
C2867 CLK2.n433 0 0.02fF $ **FLOATING
C2868 CLK2.n434 0 0.02fF $ **FLOATING
C2869 CLK2.n435 0 0.02fF $ **FLOATING
C2870 CLK2.n436 0 0.04fF $ **FLOATING
C2871 CLK2.n437 0 0.02fF $ **FLOATING
C2872 CLK2.n438 0 0.02fF $ **FLOATING
C2873 CLK2.n439 0 0.02fF $ **FLOATING
C2874 CLK2.n440 0 0.04fF $ **FLOATING
C2875 CLK2.n441 0 0.02fF $ **FLOATING
C2876 CLK2.n442 0 0.02fF $ **FLOATING
C2877 CLK2.n443 0 0.02fF $ **FLOATING
C2878 CLK2.n444 0 0.04fF $ **FLOATING
C2879 CLK2.n445 0 0.02fF $ **FLOATING
C2880 CLK2.n446 0 0.02fF $ **FLOATING
C2881 CLK2.n447 0 0.02fF $ **FLOATING
C2882 CLK2.n448 0 0.05fF $ **FLOATING
C2883 CLK2.n449 0 0.02fF $ **FLOATING
C2884 CLK2.n450 0 0.02fF $ **FLOATING
C2885 CLK2.n451 0 0.02fF $ **FLOATING
C2886 CLK2.n452 0 0.06fF $ **FLOATING
C2887 CLK2.n453 0 0.02fF $ **FLOATING
C2888 CLK2.n454 0 0.06fF $ **FLOATING
C2889 CLK2.n455 0 0.02fF $ **FLOATING
C2890 CLK2.t115 0 0.03fF
C2891 CLK2.n456 0 0.08fF $ **FLOATING
C2892 CLK2.n457 0 0.01fF $ **FLOATING
C2893 CLK2.n458 0 0.09fF $ **FLOATING
C2894 CLK2.n459 0 0.08fF $ **FLOATING
C2895 CLK2.n460 0 0.02fF $ **FLOATING
C2896 CLK2.n461 0 0.02fF $ **FLOATING
C2897 CLK2.t16 0 0.03fF
C2898 CLK2.n462 0 0.08fF $ **FLOATING
C2899 CLK2.n463 0 0.01fF $ **FLOATING
C2900 CLK2.n464 0 0.07fF $ **FLOATING
C2901 CLK2.n465 0 0.09fF $ **FLOATING
C2902 CLK2.n466 0 0.06fF $ **FLOATING
C2903 CLK2.n467 0 0.05fF $ **FLOATING
C2904 CLK2.n468 0 0.02fF $ **FLOATING
C2905 CLK2.n469 0 0.02fF $ **FLOATING
C2906 CLK2.n470 0 0.02fF $ **FLOATING
C2907 CLK2.n471 0 0.04fF $ **FLOATING
C2908 CLK2.n472 0 0.02fF $ **FLOATING
C2909 CLK2.n473 0 0.02fF $ **FLOATING
C2910 CLK2.n474 0 0.02fF $ **FLOATING
C2911 CLK2.n475 0 0.04fF $ **FLOATING
C2912 CLK2.n476 0 0.02fF $ **FLOATING
C2913 CLK2.n477 0 0.02fF $ **FLOATING
C2914 CLK2.n478 0 0.02fF $ **FLOATING
C2915 CLK2.n479 0 0.04fF $ **FLOATING
C2916 CLK2.n480 0 0.02fF $ **FLOATING
C2917 CLK2.n481 0 0.02fF $ **FLOATING
C2918 CLK2.n482 0 0.02fF $ **FLOATING
C2919 CLK2.n483 0 0.10fF $ **FLOATING
C2920 CLK2.n484 0 0.02fF $ **FLOATING
C2921 CLK2.n485 0 0.02fF $ **FLOATING
C2922 CLK2.n486 0 0.02fF $ **FLOATING
C2923 CLK2.n487 0 0.13fF $ **FLOATING
C2924 CLK2.n488 0 0.02fF $ **FLOATING
C2925 CLK2.n489 0 0.02fF $ **FLOATING
C2926 CLK2.n490 0 0.01fF $ **FLOATING
C2927 CLK2.n491 0 0.21fF $ **FLOATING
C2928 CLK2.t26 0 0.06fF
C2929 CLK2.n492 0 0.08fF $ **FLOATING
C2930 CLK2.n493 0 0.02fF $ **FLOATING
C2931 CLK2.n494 0 0.02fF $ **FLOATING
C2932 CLK2.n495 0 0.02fF $ **FLOATING
C2933 CLK2.n496 0 0.12fF $ **FLOATING
C2934 CLK2.n497 0 0.02fF $ **FLOATING
C2935 CLK2.n498 0 0.02fF $ **FLOATING
C2936 CLK2.n499 0 0.02fF $ **FLOATING
C2937 CLK2.t24 0 0.06fF
C2938 CLK2.n500 0 0.07fF $ **FLOATING
C2939 CLK2.n501 0 0.02fF $ **FLOATING
C2940 CLK2.n502 0 0.02fF $ **FLOATING
C2941 CLK2.n503 0 0.02fF $ **FLOATING
C2942 CLK2.n504 0 0.13fF $ **FLOATING
C2943 CLK2.n505 0 0.12fF $ **FLOATING
C2944 CLK2.n506 0 0.02fF $ **FLOATING
C2945 CLK2.n507 0 0.02fF $ **FLOATING
C2946 CLK2.t22 0 0.06fF
C2947 CLK2.n508 0 0.07fF $ **FLOATING
C2948 CLK2.n509 0 0.02fF $ **FLOATING
C2949 CLK2.n510 0 0.02fF $ **FLOATING
C2950 CLK2.n511 0 0.02fF $ **FLOATING
C2951 CLK2.n512 0 0.12fF $ **FLOATING
C2952 CLK2.n513 0 0.02fF $ **FLOATING
C2953 CLK2.n514 0 0.02fF $ **FLOATING
C2954 CLK2.n515 0 0.02fF $ **FLOATING
C2955 CLK2.t20 0 0.06fF
C2956 CLK2.n516 0 0.08fF $ **FLOATING
C2957 CLK2.n517 0 0.02fF $ **FLOATING
C2958 CLK2.n518 0 0.02fF $ **FLOATING
C2959 CLK2.n519 0 0.02fF $ **FLOATING
C2960 CLK2.n520 0 0.21fF $ **FLOATING
C2961 CLK2.n521 0 0.13fF $ **FLOATING
C2962 CLK2.n522 0 0.02fF $ **FLOATING
C2963 CLK2.n523 0 0.02fF $ **FLOATING
C2964 CLK2.n524 0 0.01fF $ **FLOATING
C2965 CLK2.n525 0 0.10fF $ **FLOATING
C2966 CLK2.n526 0 0.02fF $ **FLOATING
C2967 CLK2.n527 0 0.02fF $ **FLOATING
C2968 CLK2.n528 0 0.02fF $ **FLOATING
C2969 CLK2.n529 0 0.04fF $ **FLOATING
C2970 CLK2.n530 0 0.02fF $ **FLOATING
C2971 CLK2.n531 0 0.02fF $ **FLOATING
C2972 CLK2.n532 0 0.02fF $ **FLOATING
C2973 CLK2.n533 0 0.04fF $ **FLOATING
C2974 CLK2.n534 0 0.02fF $ **FLOATING
C2975 CLK2.n535 0 0.02fF $ **FLOATING
C2976 CLK2.n536 0 0.02fF $ **FLOATING
C2977 CLK2.n537 0 0.14fF $ **FLOATING
C2978 CLK2.n538 0 0.04fF $ **FLOATING
C2979 CLK2.n539 0 0.02fF $ **FLOATING
C2980 CLK2.n540 0 0.02fF $ **FLOATING
C2981 CLK2.n541 0 0.01fF $ **FLOATING
C2982 CLK2.n542 0 0.05fF $ **FLOATING
C2983 CLK2.n543 0 0.02fF $ **FLOATING
C2984 CLK2.n544 0 0.02fF $ **FLOATING
C2985 CLK2.n545 0 0.02fF $ **FLOATING
C2986 CLK2.n546 0 0.09fF $ **FLOATING
C2987 CLK2.n547 0 0.15fF $ **FLOATING
C2988 CLK2.t105 0 0.04fF
C2989 CLK2.t101 0 0.03fF
C2990 CLK2.t81 0 0.03fF
C2991 CLK2.n548 0 0.08fF $ **FLOATING
C2992 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/CLK 0 0.01fF $ **FLOATING
C2993 CLK2.t89 0 0.04fF
C2994 CLK2.t9 0 0.05fF
C2995 CLK2.n549 0 0.11fF $ **FLOATING
C2996 CLK2.n550 0 0.34fF $ **FLOATING
C2997 CLK2.n551 0 0.05fF $ **FLOATING
C2998 CLK2.n552 0 0.02fF $ **FLOATING
C2999 CLK2.n553 0 0.02fF $ **FLOATING
C3000 CLK2.n554 0 0.02fF $ **FLOATING
C3001 CLK2.n555 0 0.04fF $ **FLOATING
C3002 CLK2.n556 0 0.02fF $ **FLOATING
C3003 CLK2.n557 0 0.02fF $ **FLOATING
C3004 CLK2.n558 0 0.02fF $ **FLOATING
C3005 CLK2.n559 0 0.10fF $ **FLOATING
C3006 CLK2.n560 0 0.02fF $ **FLOATING
C3007 CLK2.n561 0 0.02fF $ **FLOATING
C3008 CLK2.n562 0 0.02fF $ **FLOATING
C3009 CLK2.n563 0 0.13fF $ **FLOATING
C3010 CLK2.n564 0 0.02fF $ **FLOATING
C3011 CLK2.n565 0 0.02fF $ **FLOATING
C3012 CLK2.n566 0 0.01fF $ **FLOATING
C3013 CLK2.n567 0 0.21fF $ **FLOATING
C3014 CLK2.t88 0 0.06fF
C3015 CLK2.n568 0 0.08fF $ **FLOATING
C3016 CLK2.n569 0 0.02fF $ **FLOATING
C3017 CLK2.n570 0 0.02fF $ **FLOATING
C3018 CLK2.n571 0 0.02fF $ **FLOATING
C3019 CLK2.n572 0 0.12fF $ **FLOATING
C3020 CLK2.n573 0 0.02fF $ **FLOATING
C3021 CLK2.n574 0 0.02fF $ **FLOATING
C3022 CLK2.n575 0 0.02fF $ **FLOATING
C3023 CLK2.n576 0 0.02fF $ **FLOATING
C3024 CLK2.t80 0 0.06fF
C3025 CLK2.n577 0 0.07fF $ **FLOATING
C3026 CLK2.n578 0 0.02fF $ **FLOATING
C3027 CLK2.n579 0 0.02fF $ **FLOATING
C3028 CLK2.n580 0 0.12fF $ **FLOATING
C3029 CLK2.n581 0 0.02fF $ **FLOATING
C3030 CLK2.n582 0 0.02fF $ **FLOATING
C3031 CLK2.n583 0 0.13fF $ **FLOATING
C3032 CLK2.t100 0 0.06fF
C3033 CLK2.n584 0 0.07fF $ **FLOATING
C3034 CLK2.n585 0 0.02fF $ **FLOATING
C3035 CLK2.n586 0 0.02fF $ **FLOATING
C3036 CLK2.n587 0 0.02fF $ **FLOATING
C3037 CLK2.n588 0 0.12fF $ **FLOATING
C3038 CLK2.n589 0 0.02fF $ **FLOATING
C3039 CLK2.n590 0 0.02fF $ **FLOATING
C3040 CLK2.n591 0 0.02fF $ **FLOATING
C3041 CLK2.t104 0 0.06fF
C3042 CLK2.n592 0 0.08fF $ **FLOATING
C3043 CLK2.n593 0 0.02fF $ **FLOATING
C3044 CLK2.n594 0 0.02fF $ **FLOATING
C3045 CLK2.n595 0 0.02fF $ **FLOATING
C3046 CLK2.n596 0 0.21fF $ **FLOATING
C3047 CLK2.n597 0 0.13fF $ **FLOATING
C3048 CLK2.n598 0 0.02fF $ **FLOATING
C3049 CLK2.n599 0 0.02fF $ **FLOATING
C3050 CLK2.n600 0 0.01fF $ **FLOATING
C3051 CLK2.n601 0 0.10fF $ **FLOATING
C3052 CLK2.n602 0 0.02fF $ **FLOATING
C3053 CLK2.n603 0 0.02fF $ **FLOATING
C3054 CLK2.n604 0 0.02fF $ **FLOATING
C3055 CLK2.n605 0 0.04fF $ **FLOATING
C3056 CLK2.n606 0 0.02fF $ **FLOATING
C3057 CLK2.n607 0 0.02fF $ **FLOATING
C3058 CLK2.n608 0 0.01fF $ **FLOATING
C3059 CLK2.n609 0 0.15fF $ **FLOATING
C3060 CLK2.n610 0 0.05fF $ **FLOATING
C3061 CLK2.n611 0 0.02fF $ **FLOATING
C3062 CLK2.n612 0 0.02fF $ **FLOATING
C3063 CLK2.n613 0 0.02fF $ **FLOATING
C3064 CLK2.n614 0 0.11fF $ **FLOATING
C3065 CLK2.n615 0 0.02fF $ **FLOATING
C3066 CLK2.n616 0 0.09fF $ **FLOATING
C3067 CLK2.n617 0 0.02fF $ **FLOATING
C3068 CLK2.n618 0 0.12fF $ **FLOATING
C3069 CLK2.n619 0 0.11fF $ **FLOATING
C3070 CLK2.n620 0 0.02fF $ **FLOATING
C3071 CLK2.n621 0 0.02fF $ **FLOATING
C3072 CLK2.n622 0 0.10fF $ **FLOATING
C3073 CLK2.t103 0 0.04fF
C3074 CLK2.t54 0 0.03fF
C3075 CLK2.t95 0 0.03fF
C3076 CLK2.n623 0 0.08fF $ **FLOATING
C3077 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/CLK 0 0.01fF $ **FLOATING
C3078 CLK2.t64 0 0.04fF
C3079 CLK2.t57 0 0.05fF
C3080 CLK2.n624 0 0.11fF $ **FLOATING
C3081 CLK2.n625 0 0.34fF $ **FLOATING
C3082 CLK2.n626 0 0.05fF $ **FLOATING
C3083 CLK2.n627 0 0.02fF $ **FLOATING
C3084 CLK2.n628 0 0.02fF $ **FLOATING
C3085 CLK2.n629 0 0.02fF $ **FLOATING
C3086 CLK2.n630 0 0.04fF $ **FLOATING
C3087 CLK2.n631 0 0.02fF $ **FLOATING
C3088 CLK2.n632 0 0.02fF $ **FLOATING
C3089 CLK2.n633 0 0.02fF $ **FLOATING
C3090 CLK2.n634 0 0.10fF $ **FLOATING
C3091 CLK2.n635 0 0.02fF $ **FLOATING
C3092 CLK2.n636 0 0.02fF $ **FLOATING
C3093 CLK2.n637 0 0.02fF $ **FLOATING
C3094 CLK2.n638 0 0.13fF $ **FLOATING
C3095 CLK2.n639 0 0.02fF $ **FLOATING
C3096 CLK2.n640 0 0.02fF $ **FLOATING
C3097 CLK2.n641 0 0.01fF $ **FLOATING
C3098 CLK2.n642 0 0.21fF $ **FLOATING
C3099 CLK2.t63 0 0.06fF
C3100 CLK2.n643 0 0.08fF $ **FLOATING
C3101 CLK2.n644 0 0.02fF $ **FLOATING
C3102 CLK2.n645 0 0.02fF $ **FLOATING
C3103 CLK2.n646 0 0.02fF $ **FLOATING
C3104 CLK2.n647 0 0.12fF $ **FLOATING
C3105 CLK2.n648 0 0.02fF $ **FLOATING
C3106 CLK2.n649 0 0.02fF $ **FLOATING
C3107 CLK2.n650 0 0.02fF $ **FLOATING
C3108 CLK2.n651 0 0.02fF $ **FLOATING
C3109 CLK2.t94 0 0.06fF
C3110 CLK2.n652 0 0.07fF $ **FLOATING
C3111 CLK2.n653 0 0.02fF $ **FLOATING
C3112 CLK2.n654 0 0.02fF $ **FLOATING
C3113 CLK2.n655 0 0.12fF $ **FLOATING
C3114 CLK2.n656 0 0.02fF $ **FLOATING
C3115 CLK2.n657 0 0.02fF $ **FLOATING
C3116 CLK2.n658 0 0.13fF $ **FLOATING
C3117 CLK2.t53 0 0.06fF
C3118 CLK2.n659 0 0.07fF $ **FLOATING
C3119 CLK2.n660 0 0.02fF $ **FLOATING
C3120 CLK2.n661 0 0.02fF $ **FLOATING
C3121 CLK2.n662 0 0.02fF $ **FLOATING
C3122 CLK2.n663 0 0.12fF $ **FLOATING
C3123 CLK2.n664 0 0.02fF $ **FLOATING
C3124 CLK2.n665 0 0.02fF $ **FLOATING
C3125 CLK2.n666 0 0.02fF $ **FLOATING
C3126 CLK2.t102 0 0.06fF
C3127 CLK2.n667 0 0.08fF $ **FLOATING
C3128 CLK2.n668 0 0.02fF $ **FLOATING
C3129 CLK2.n669 0 0.02fF $ **FLOATING
C3130 CLK2.n670 0 0.02fF $ **FLOATING
C3131 CLK2.n671 0 0.21fF $ **FLOATING
C3132 CLK2.n672 0 0.13fF $ **FLOATING
C3133 CLK2.n673 0 0.02fF $ **FLOATING
C3134 CLK2.n674 0 0.02fF $ **FLOATING
C3135 CLK2.n675 0 0.01fF $ **FLOATING
C3136 CLK2.n676 0 0.10fF $ **FLOATING
C3137 CLK2.n677 0 0.02fF $ **FLOATING
C3138 CLK2.n678 0 0.02fF $ **FLOATING
C3139 CLK2.n679 0 0.02fF $ **FLOATING
C3140 CLK2.n680 0 0.04fF $ **FLOATING
C3141 CLK2.n681 0 0.02fF $ **FLOATING
C3142 CLK2.n682 0 0.02fF $ **FLOATING
C3143 CLK2.n683 0 0.02fF $ **FLOATING
C3144 CLK2.n684 0 0.05fF $ **FLOATING
C3145 CLK2.n685 0 0.02fF $ **FLOATING
C3146 CLK2.n686 0 0.02fF $ **FLOATING
C3147 CLK2.n687 0 0.02fF $ **FLOATING
C3148 CLK2.n688 0 0.09fF $ **FLOATING
C3149 CLK2.n689 0 0.15fF $ **FLOATING
C3150 CLK2.n690 0 0.15fF $ **FLOATING
C3151 CLK2.n691 0 0.05fF $ **FLOATING
C3152 CLK2.n692 0 0.02fF $ **FLOATING
C3153 CLK2.n693 0 0.02fF $ **FLOATING
C3154 CLK2.n694 0 0.02fF $ **FLOATING
C3155 CLK2.n695 0 0.04fF $ **FLOATING
C3156 CLK2.n696 0 0.02fF $ **FLOATING
C3157 CLK2.n697 0 0.02fF $ **FLOATING
C3158 CLK2.n698 0 0.01fF $ **FLOATING
C3159 CLK2.n699 0 0.14fF $ **FLOATING
C3160 CLK2.n700 0 0.04fF $ **FLOATING
C3161 CLK2.n701 0 0.02fF $ **FLOATING
C3162 CLK2.n702 0 0.02fF $ **FLOATING
C3163 CLK2.n703 0 0.02fF $ **FLOATING
C3164 CLK2.n704 0 0.04fF $ **FLOATING
C3165 CLK2.n705 0 0.02fF $ **FLOATING
C3166 CLK2.n706 0 0.02fF $ **FLOATING
C3167 CLK2.n707 0 0.02fF $ **FLOATING
C3168 CLK2.n708 0 0.10fF $ **FLOATING
C3169 CLK2.n709 0 0.02fF $ **FLOATING
C3170 CLK2.n710 0 0.02fF $ **FLOATING
C3171 CLK2.n711 0 0.02fF $ **FLOATING
C3172 CLK2.n712 0 0.13fF $ **FLOATING
C3173 CLK2.n713 0 0.02fF $ **FLOATING
C3174 CLK2.n714 0 0.02fF $ **FLOATING
C3175 CLK2.n715 0 0.01fF $ **FLOATING
C3176 CLK2.n716 0 0.21fF $ **FLOATING
C3177 CLK2.t109 0 0.06fF
C3178 CLK2.n717 0 0.08fF $ **FLOATING
C3179 CLK2.n718 0 0.02fF $ **FLOATING
C3180 CLK2.n719 0 0.02fF $ **FLOATING
C3181 CLK2.n720 0 0.02fF $ **FLOATING
C3182 CLK2.n721 0 0.12fF $ **FLOATING
C3183 CLK2.n722 0 0.02fF $ **FLOATING
C3184 CLK2.n723 0 0.02fF $ **FLOATING
C3185 CLK2.n724 0 0.02fF $ **FLOATING
C3186 CLK2.n725 0 0.02fF $ **FLOATING
C3187 CLK2.t107 0 0.06fF
C3188 CLK2.n726 0 0.07fF $ **FLOATING
C3189 CLK2.n727 0 0.02fF $ **FLOATING
C3190 CLK2.n728 0 0.02fF $ **FLOATING
C3191 CLK2.n729 0 0.12fF $ **FLOATING
C3192 CLK2.n730 0 0.02fF $ **FLOATING
C3193 CLK2.n731 0 0.02fF $ **FLOATING
C3194 CLK2.n732 0 0.13fF $ **FLOATING
C3195 CLK2.t43 0 0.06fF
C3196 CLK2.n733 0 0.07fF $ **FLOATING
C3197 CLK2.n734 0 0.02fF $ **FLOATING
C3198 CLK2.n735 0 0.02fF $ **FLOATING
C3199 CLK2.n736 0 0.02fF $ **FLOATING
C3200 CLK2.n737 0 0.12fF $ **FLOATING
C3201 CLK2.n738 0 0.02fF $ **FLOATING
C3202 CLK2.n739 0 0.02fF $ **FLOATING
C3203 CLK2.n740 0 0.02fF $ **FLOATING
C3204 CLK2.t41 0 0.06fF
C3205 CLK2.n741 0 0.08fF $ **FLOATING
C3206 CLK2.n742 0 0.02fF $ **FLOATING
C3207 CLK2.n743 0 0.02fF $ **FLOATING
C3208 CLK2.n744 0 0.02fF $ **FLOATING
C3209 CLK2.n745 0 0.21fF $ **FLOATING
C3210 CLK2.n746 0 0.13fF $ **FLOATING
C3211 CLK2.n747 0 0.02fF $ **FLOATING
C3212 CLK2.n748 0 0.02fF $ **FLOATING
C3213 CLK2.n749 0 0.01fF $ **FLOATING
C3214 CLK2.n750 0 0.10fF $ **FLOATING
C3215 CLK2.n751 0 0.02fF $ **FLOATING
C3216 CLK2.n752 0 0.02fF $ **FLOATING
C3217 CLK2.n753 0 0.02fF $ **FLOATING
C3218 CLK2.n754 0 0.04fF $ **FLOATING
C3219 CLK2.n755 0 0.02fF $ **FLOATING
C3220 CLK2.n756 0 0.02fF $ **FLOATING
C3221 CLK2.n757 0 0.02fF $ **FLOATING
C3222 CLK2.n758 0 0.04fF $ **FLOATING
C3223 CLK2.n759 0 0.02fF $ **FLOATING
C3224 CLK2.n760 0 0.02fF $ **FLOATING
C3225 CLK2.n761 0 0.02fF $ **FLOATING
C3226 CLK2.n762 0 0.04fF $ **FLOATING
C3227 CLK2.n763 0 0.02fF $ **FLOATING
C3228 CLK2.n764 0 0.02fF $ **FLOATING
C3229 CLK2.n765 0 0.02fF $ **FLOATING
C3230 CLK2.n766 0 0.05fF $ **FLOATING
C3231 CLK2.n767 0 0.02fF $ **FLOATING
C3232 CLK2.n768 0 0.02fF $ **FLOATING
C3233 CLK2.n769 0 0.02fF $ **FLOATING
C3234 CLK2.n770 0 0.06fF $ **FLOATING
C3235 CLK2.n771 0 0.02fF $ **FLOATING
C3236 CLK2.n772 0 0.06fF $ **FLOATING
C3237 CLK2.n773 0 0.02fF $ **FLOATING
C3238 CLK2.t66 0 0.03fF
C3239 CLK2.n774 0 0.08fF $ **FLOATING
C3240 CLK2.n775 0 0.01fF $ **FLOATING
C3241 CLK2.n776 0 0.09fF $ **FLOATING
C3242 CLK2.n777 0 0.08fF $ **FLOATING
C3243 CLK2.n778 0 0.02fF $ **FLOATING
C3244 CLK2.n779 0 0.02fF $ **FLOATING
C3245 CLK2.n780 0 0.07fF $ **FLOATING
C3246 CLK2.n781 0 0.04fF $ **FLOATING
C3247 CLK2.n782 0 0.09fF $ **FLOATING
C3248 CLK2.n783 0 0.01fF $ **FLOATING
C3249 EESPFAL_Sbox_0/EESPFAL_s1_0/CLK2 0 0.02fF $ **FLOATING
C3250 CLK2.n784 0 0.01fF $ **FLOATING
C3251 CLK2.n785 0 0.05fF $ **FLOATING
C3252 CLK2.n786 0 0.02fF $ **FLOATING
C3253 CLK2.n787 0 0.02fF $ **FLOATING
C3254 CLK2.n788 0 0.02fF $ **FLOATING
C3255 CLK2.n789 0 0.04fF $ **FLOATING
C3256 CLK2.n790 0 0.02fF $ **FLOATING
C3257 CLK2.n791 0 0.02fF $ **FLOATING
C3258 CLK2.n792 0 0.02fF $ **FLOATING
C3259 CLK2.n793 0 0.04fF $ **FLOATING
C3260 CLK2.n794 0 0.02fF $ **FLOATING
C3261 CLK2.n795 0 0.02fF $ **FLOATING
C3262 CLK2.n796 0 0.02fF $ **FLOATING
C3263 CLK2.n797 0 0.04fF $ **FLOATING
C3264 CLK2.n798 0 0.02fF $ **FLOATING
C3265 CLK2.n799 0 0.02fF $ **FLOATING
C3266 CLK2.n800 0 0.02fF $ **FLOATING
C3267 CLK2.n801 0 0.10fF $ **FLOATING
C3268 CLK2.n802 0 0.02fF $ **FLOATING
C3269 CLK2.n803 0 0.02fF $ **FLOATING
C3270 CLK2.n804 0 0.02fF $ **FLOATING
C3271 CLK2.n805 0 0.13fF $ **FLOATING
C3272 CLK2.n806 0 0.02fF $ **FLOATING
C3273 CLK2.n807 0 0.02fF $ **FLOATING
C3274 CLK2.n808 0 0.01fF $ **FLOATING
C3275 CLK2.n809 0 0.21fF $ **FLOATING
C3276 CLK2.t90 0 0.06fF
C3277 CLK2.n810 0 0.08fF $ **FLOATING
C3278 CLK2.n811 0 0.02fF $ **FLOATING
C3279 CLK2.n812 0 0.02fF $ **FLOATING
C3280 CLK2.n813 0 0.02fF $ **FLOATING
C3281 CLK2.n814 0 0.12fF $ **FLOATING
C3282 CLK2.n815 0 0.02fF $ **FLOATING
C3283 CLK2.n816 0 0.02fF $ **FLOATING
C3284 CLK2.n817 0 0.02fF $ **FLOATING
C3285 CLK2.t92 0 0.06fF
C3286 CLK2.n818 0 0.07fF $ **FLOATING
C3287 CLK2.n819 0 0.02fF $ **FLOATING
C3288 CLK2.n820 0 0.02fF $ **FLOATING
C3289 CLK2.n821 0 0.02fF $ **FLOATING
C3290 CLK2.n822 0 0.13fF $ **FLOATING
C3291 CLK2.n823 0 0.02fF $ **FLOATING
C3292 CLK2.t28 0 0.06fF
C3293 CLK2.n824 0 0.07fF $ **FLOATING
C3294 CLK2.n825 0 0.02fF $ **FLOATING
C3295 CLK2.n826 0 0.02fF $ **FLOATING
C3296 CLK2.n827 0 0.02fF $ **FLOATING
C3297 CLK2.n828 0 0.12fF $ **FLOATING
C3298 CLK2.n829 0 0.02fF $ **FLOATING
C3299 CLK2.n830 0 0.02fF $ **FLOATING
C3300 CLK2.n831 0 0.02fF $ **FLOATING
C3301 CLK2.t30 0 0.06fF
C3302 CLK2.n832 0 0.08fF $ **FLOATING
C3303 CLK2.n833 0 0.02fF $ **FLOATING
C3304 CLK2.n834 0 0.02fF $ **FLOATING
C3305 CLK2.n835 0 0.02fF $ **FLOATING
C3306 CLK2.n836 0 0.21fF $ **FLOATING
C3307 CLK2.n837 0 0.13fF $ **FLOATING
C3308 CLK2.n838 0 0.02fF $ **FLOATING
C3309 CLK2.n839 0 0.02fF $ **FLOATING
C3310 CLK2.n840 0 0.01fF $ **FLOATING
C3311 CLK2.n841 0 0.10fF $ **FLOATING
C3312 CLK2.n842 0 0.02fF $ **FLOATING
C3313 CLK2.n843 0 0.02fF $ **FLOATING
C3314 CLK2.n844 0 0.02fF $ **FLOATING
C3315 CLK2.n845 0 0.04fF $ **FLOATING
C3316 CLK2.n846 0 0.02fF $ **FLOATING
C3317 CLK2.n847 0 0.02fF $ **FLOATING
C3318 CLK2.n848 0 0.02fF $ **FLOATING
C3319 CLK2.n849 0 0.04fF $ **FLOATING
C3320 CLK2.n850 0 0.02fF $ **FLOATING
C3321 CLK2.n851 0 0.02fF $ **FLOATING
C3322 CLK2.n852 0 0.02fF $ **FLOATING
C3323 CLK2.n853 0 0.14fF $ **FLOATING
C3324 CLK2.n854 0 0.05fF $ **FLOATING
C3325 CLK2.n855 0 0.09fF $ **FLOATING
C3326 CLK2.n856 0 0.01fF $ **FLOATING
C3327 CLK2.n857 0 0.09fF $ **FLOATING
C3328 CLK2.n858 0 0.16fF $ **FLOATING
C3329 CLK2.t40 0 0.04fF
C3330 CLK2.t38 0 0.03fF
C3331 CLK2.t77 0 0.03fF
C3332 CLK2.n859 0 0.08fF $ **FLOATING
C3333 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/CLK 0 0.01fF $ **FLOATING
C3334 CLK2.t79 0 0.04fF
C3335 CLK2.t99 0 0.03fF
C3336 CLK2.t32 0 0.03fF
C3337 CLK2.n860 0 0.11fF $ **FLOATING
C3338 CLK2.n861 0 0.05fF $ **FLOATING
C3339 CLK2.n862 0 0.02fF $ **FLOATING
C3340 CLK2.n863 0 0.02fF $ **FLOATING
C3341 CLK2.n864 0 0.09fF $ **FLOATING
C3342 CLK2.n865 0 0.04fF $ **FLOATING
C3343 CLK2.n866 0 0.02fF $ **FLOATING
C3344 CLK2.n867 0 0.02fF $ **FLOATING
C3345 CLK2.n868 0 0.05fF $ **FLOATING
C3346 CLK2.n869 0 0.14fF $ **FLOATING
C3347 CLK2.n870 0 0.04fF $ **FLOATING
C3348 CLK2.n871 0 0.02fF $ **FLOATING
C3349 CLK2.n872 0 0.02fF $ **FLOATING
C3350 CLK2.n873 0 0.02fF $ **FLOATING
C3351 CLK2.n874 0 0.04fF $ **FLOATING
C3352 CLK2.n875 0 0.02fF $ **FLOATING
C3353 CLK2.n876 0 0.02fF $ **FLOATING
C3354 CLK2.n877 0 0.02fF $ **FLOATING
C3355 CLK2.n878 0 0.10fF $ **FLOATING
C3356 CLK2.n879 0 0.02fF $ **FLOATING
C3357 CLK2.n880 0 0.02fF $ **FLOATING
C3358 CLK2.n881 0 0.02fF $ **FLOATING
C3359 CLK2.n882 0 0.13fF $ **FLOATING
C3360 CLK2.n883 0 0.02fF $ **FLOATING
C3361 CLK2.n884 0 0.02fF $ **FLOATING
C3362 CLK2.n885 0 0.01fF $ **FLOATING
C3363 CLK2.n886 0 0.21fF $ **FLOATING
C3364 CLK2.t78 0 0.06fF
C3365 CLK2.n887 0 0.08fF $ **FLOATING
C3366 CLK2.n888 0 0.02fF $ **FLOATING
C3367 CLK2.n889 0 0.02fF $ **FLOATING
C3368 CLK2.n890 0 0.02fF $ **FLOATING
C3369 CLK2.n891 0 0.12fF $ **FLOATING
C3370 CLK2.n892 0 0.02fF $ **FLOATING
C3371 CLK2.n893 0 0.02fF $ **FLOATING
C3372 CLK2.n894 0 0.02fF $ **FLOATING
C3373 CLK2.n895 0 0.02fF $ **FLOATING
C3374 CLK2.t76 0 0.06fF
C3375 CLK2.n896 0 0.07fF $ **FLOATING
C3376 CLK2.n897 0 0.02fF $ **FLOATING
C3377 CLK2.n898 0 0.02fF $ **FLOATING
C3378 CLK2.n899 0 0.12fF $ **FLOATING
C3379 CLK2.n900 0 0.02fF $ **FLOATING
C3380 CLK2.n901 0 0.02fF $ **FLOATING
C3381 CLK2.n902 0 0.13fF $ **FLOATING
C3382 CLK2.t37 0 0.06fF
C3383 CLK2.n903 0 0.07fF $ **FLOATING
C3384 CLK2.n904 0 0.02fF $ **FLOATING
C3385 CLK2.n905 0 0.02fF $ **FLOATING
C3386 CLK2.n906 0 0.02fF $ **FLOATING
C3387 CLK2.n907 0 0.12fF $ **FLOATING
C3388 CLK2.n908 0 0.02fF $ **FLOATING
C3389 CLK2.n909 0 0.02fF $ **FLOATING
C3390 CLK2.n910 0 0.02fF $ **FLOATING
C3391 CLK2.t39 0 0.06fF
C3392 CLK2.n911 0 0.08fF $ **FLOATING
C3393 CLK2.n912 0 0.02fF $ **FLOATING
C3394 CLK2.n913 0 0.02fF $ **FLOATING
C3395 CLK2.n914 0 0.02fF $ **FLOATING
C3396 CLK2.n915 0 0.21fF $ **FLOATING
C3397 CLK2.n916 0 0.13fF $ **FLOATING
C3398 CLK2.n917 0 0.02fF $ **FLOATING
C3399 CLK2.n918 0 0.02fF $ **FLOATING
C3400 CLK2.n919 0 0.01fF $ **FLOATING
C3401 CLK2.n920 0 0.10fF $ **FLOATING
C3402 CLK2.n921 0 0.02fF $ **FLOATING
C3403 CLK2.n922 0 0.02fF $ **FLOATING
C3404 CLK2.n923 0 0.02fF $ **FLOATING
C3405 CLK2.n924 0 0.04fF $ **FLOATING
C3406 CLK2.n925 0 0.02fF $ **FLOATING
C3407 CLK2.n926 0 0.02fF $ **FLOATING
C3408 CLK2.n927 0 0.02fF $ **FLOATING
C3409 CLK2.n928 0 0.04fF $ **FLOATING
C3410 CLK2.n929 0 0.02fF $ **FLOATING
C3411 CLK2.n930 0 0.02fF $ **FLOATING
C3412 CLK2.n931 0 0.02fF $ **FLOATING
C3413 CLK2.n932 0 0.04fF $ **FLOATING
C3414 CLK2.n933 0 0.02fF $ **FLOATING
C3415 CLK2.n934 0 0.02fF $ **FLOATING
C3416 CLK2.n935 0 0.02fF $ **FLOATING
C3417 CLK2.n936 0 0.05fF $ **FLOATING
C3418 CLK2.n937 0 0.02fF $ **FLOATING
C3419 CLK2.n938 0 0.02fF $ **FLOATING
C3420 CLK2.n939 0 0.02fF $ **FLOATING
C3421 CLK2.n940 0 0.06fF $ **FLOATING
C3422 CLK2.n941 0 0.02fF $ **FLOATING
C3423 CLK2.n942 0 0.06fF $ **FLOATING
C3424 CLK2.n943 0 0.02fF $ **FLOATING
C3425 CLK2.n944 0 0.01fF $ **FLOATING
C3426 CLK2.t71 0 0.03fF
C3427 CLK2.n945 0 0.08fF $ **FLOATING
C3428 CLK2.n946 0 0.01fF $ **FLOATING
C3429 CLK2.n947 0 0.11fF $ **FLOATING
C3430 CLK2.n948 0 0.12fF $ **FLOATING
C3431 CLK2.t49 0 0.03fF
C3432 CLK2.t10 0 0.03fF
C3433 CLK2.n949 0 0.05fF $ **FLOATING
C3434 CLK2.n950 0 0.01fF $ **FLOATING
C3435 CLK2.n951 0 0.02fF $ **FLOATING
C3436 CLK2.n952 0 0.02fF $ **FLOATING
C3437 CLK2.n953 0 0.06fF $ **FLOATING
C3438 CLK2.n954 0 0.05fF $ **FLOATING
C3439 CLK2.n955 0 0.02fF $ **FLOATING
C3440 CLK2.n956 0 0.02fF $ **FLOATING
C3441 CLK2.n957 0 0.09fF $ **FLOATING
C3442 CLK2.n958 0 0.05fF $ **FLOATING
C3443 CLK2.n959 0 0.04fF $ **FLOATING
C3444 CLK2.n960 0 0.02fF $ **FLOATING
C3445 CLK2.n961 0 0.01fF $ **FLOATING
C3446 CLK2.n962 0 0.01fF $ **FLOATING
C3447 CLK2.n963 0 0.00fF $ **FLOATING
C3448 CLK2.n964 0 0.04fF $ **FLOATING
C3449 EESPFAL_Sbox_0/CLK2 0 0.01fF $ **FLOATING
C3450 CLK2.n965 0 0.00fF $ **FLOATING
C3451 EESPFAL_Sbox_0/EESPFAL_s0_0/CLK2 0 0.01fF $ **FLOATING
C3452 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_2/OUT_bar 0 0.72fF $ **FLOATING
C3453 EESPFAL_Sbox_0/EESPFAL_s1_0/x2_bar 0 1.25fF $ **FLOATING
C3454 EESPFAL_Sbox_0/x2_bar 0 0.24fF $ **FLOATING
C3455 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t18 0 0.40fF
C3456 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n0 0 4.46fF $ **FLOATING
C3457 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t9 0 0.21fF
C3458 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/A_bar 0 0.62fF $ **FLOATING
C3459 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n1 0 2.03fF $ **FLOATING
C3460 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t14 0 0.41fF
C3461 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t15 0 0.23fF
C3462 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n2 0 2.13fF $ **FLOATING
C3463 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/A_bar 0 0.23fF $ **FLOATING
C3464 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t12 0 0.16fF
C3465 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/D_bar 0 0.42fF $ **FLOATING
C3466 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t17 0 0.52fF
C3467 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t11 0 0.18fF
C3468 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n3 0 1.73fF $ **FLOATING
C3469 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/B_bar 0 0.18fF $ **FLOATING
C3470 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t7 0 0.41fF
C3471 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t19 0 0.23fF
C3472 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n4 0 2.13fF $ **FLOATING
C3473 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/A_bar 0 0.22fF $ **FLOATING
C3474 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t6 0 0.45fF
C3475 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A 0 2.03fF $ **FLOATING
C3476 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n5 0 4.52fF $ **FLOATING
C3477 EESPFAL_Sbox_0/EESPFAL_s3_0/x2_bar 0 1.84fF $ **FLOATING
C3478 EESPFAL_Sbox_0/EESPFAL_s2_0/x2_bar 0 0.78fF $ **FLOATING
C3479 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n6 0 1.72fF $ **FLOATING
C3480 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t16 0 0.19fF
C3481 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/A 0 0.86fF $ **FLOATING
C3482 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n7 0 6.77fF $ **FLOATING
C3483 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n8 0 3.16fF $ **FLOATING
C3484 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t10 0 0.14fF
C3485 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/A_bar 0 0.47fF $ **FLOATING
C3486 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n9 0 6.72fF $ **FLOATING
C3487 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n10 0 1.09fF $ **FLOATING
C3488 EESPFAL_4in_XOR_0/XOR2_bar 0 0.50fF $ **FLOATING
C3489 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t2 0 0.15fF
C3490 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t3 0 0.15fF
C3491 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n11 0 0.45fF $ **FLOATING
C3492 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t5 0 0.58fF
C3493 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t4 0 1.00fF
C3494 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n12 0 0.87fF $ **FLOATING
C3495 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n13 0 0.37fF $ **FLOATING
C3496 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t1 0 0.15fF
C3497 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t0 0 0.15fF
C3498 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n14 0 0.38fF $ **FLOATING
C3499 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n15 0 0.42fF $ **FLOATING
C3500 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t13 0 0.20fF
C3501 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t8 0 0.19fF
C3502 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.t20 0 0.14fF
C3503 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n16 0 0.22fF $ **FLOATING
C3504 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B.n17 0 0.15fF $ **FLOATING
C3505 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t9 0 0.04fF
C3506 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/A_bar 0 0.53fF $ **FLOATING
C3507 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t3 0 0.04fF
C3508 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t2 0 0.04fF
C3509 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n0 0 0.09fF $ **FLOATING
C3510 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t1 0 0.14fF
C3511 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t5 0 0.20fF
C3512 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n1 0 0.19fF $ **FLOATING
C3513 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t4 0 0.04fF
C3514 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t0 0 0.04fF
C3515 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n2 0 0.11fF $ **FLOATING
C3516 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n3 0 0.09fF $ **FLOATING
C3517 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n4 0 0.10fF $ **FLOATING
C3518 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t6 0 0.03fF
C3519 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t8 0 0.05fF
C3520 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.t7 0 0.04fF
C3521 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n5 0 0.05fF $ **FLOATING
C3522 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar.n6 0 0.04fF $ **FLOATING
C3523 EESPFAL_Sbox_0/EESPFAL_s2_0/x1_bar 0 1.36fF $ **FLOATING
C3524 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_1/OUT_bar 0 0.71fF $ **FLOATING
C3525 EESPFAL_Sbox_0/EESPFAL_s3_0/x1_bar 0 9.85fF $ **FLOATING
C3526 EESPFAL_Sbox_0/x1_bar 0 0.68fF $ **FLOATING
C3527 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t18 0 0.39fF
C3528 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/B 0 1.77fF $ **FLOATING
C3529 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t10 0 0.16fF
C3530 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n0 0 4.86fF $ **FLOATING
C3531 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t6 0 0.41fF
C3532 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t7 0 0.23fF
C3533 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n1 0 2.13fF $ **FLOATING
C3534 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/A_bar 0 0.30fF $ **FLOATING
C3535 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t11 0 0.20fF
C3536 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B_bar 0 0.63fF $ **FLOATING
C3537 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t20 0 0.41fF
C3538 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t16 0 0.23fF
C3539 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n2 0 2.13fF $ **FLOATING
C3540 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/A_bar 0 0.32fF $ **FLOATING
C3541 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t9 0 0.19fF
C3542 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/A 0 0.76fF $ **FLOATING
C3543 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n3 0 5.10fF $ **FLOATING
C3544 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t13 0 0.41fF
C3545 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t8 0 0.23fF
C3546 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n4 0 2.13fF $ **FLOATING
C3547 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/A_bar 0 0.30fF $ **FLOATING
C3548 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t14 0 0.14fF
C3549 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_1/A_bar 0 0.56fF $ **FLOATING
C3550 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n5 0 0.59fF $ **FLOATING
C3551 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n6 0 2.28fF $ **FLOATING
C3552 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t17 0 0.25fF
C3553 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/B_bar 0 0.71fF $ **FLOATING
C3554 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n7 0 2.17fF $ **FLOATING
C3555 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n8 0 2.32fF $ **FLOATING
C3556 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n9 0 2.43fF $ **FLOATING
C3557 EESPFAL_Sbox_0/EESPFAL_s1_0/x1_bar 0 1.98fF $ **FLOATING
C3558 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n10 0 1.38fF $ **FLOATING
C3559 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n11 0 0.71fF $ **FLOATING
C3560 EESPFAL_4in_XOR_0/XOR1_bar 0 0.44fF $ **FLOATING
C3561 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t2 0 0.15fF
C3562 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t4 0 0.15fF
C3563 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n12 0 0.45fF $ **FLOATING
C3564 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t3 0 0.58fF
C3565 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t5 0 1.00fF
C3566 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n13 0 0.87fF $ **FLOATING
C3567 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n14 0 0.37fF $ **FLOATING
C3568 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t1 0 0.15fF
C3569 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t0 0 0.15fF
C3570 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n15 0 0.38fF $ **FLOATING
C3571 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n16 0 0.42fF $ **FLOATING
C3572 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t12 0 0.14fF
C3573 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t19 0 0.20fF
C3574 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.t15 0 0.19fF
C3575 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n17 0 0.22fF $ **FLOATING
C3576 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar.n18 0 0.15fF $ **FLOATING
C3577 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT_bar 0 0.32fF $ **FLOATING
C3578 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t9 0 0.07fF
C3579 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t3 0 0.05fF
C3580 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t5 0 0.05fF
C3581 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n0 0 0.16fF $ **FLOATING
C3582 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t4 0 0.20fF
C3583 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t0 0 0.34fF
C3584 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n1 0 0.30fF $ **FLOATING
C3585 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n2 0 0.13fF $ **FLOATING
C3586 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t1 0 0.05fF
C3587 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t2 0 0.05fF
C3588 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n3 0 0.13fF $ **FLOATING
C3589 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n4 0 0.14fF $ **FLOATING
C3590 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t6 0 0.05fF
C3591 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t8 0 0.07fF
C3592 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t7 0 0.06fF
C3593 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n5 0 0.07fF $ **FLOATING
C3594 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n6 0 0.05fF $ **FLOATING
C3595 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t7 0 0.13fF
C3596 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t4 0 0.21fF
C3597 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t1 0 0.05fF
C3598 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t2 0 0.05fF
C3599 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n0 0 0.16fF $ **FLOATING
C3600 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t3 0 0.05fF
C3601 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t5 0 0.05fF
C3602 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n1 0 0.15fF $ **FLOATING
C3603 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t6 0 0.04fF
C3604 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t8 0 0.06fF
C3605 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t9 0 0.07fF
C3606 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n2 0 0.07fF $ **FLOATING
C3607 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT 0 0.01fF $ **FLOATING
C3608 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n3 0 0.04fF $ **FLOATING
C3609 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n4 0 0.22fF $ **FLOATING
C3610 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t0 0 0.21fF
C3611 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n5 0 0.22fF $ **FLOATING
C3612 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n6 0 0.31fF $ **FLOATING
C3613 EESPFAL_Sbox_0/EESPFAL_s0_0/Dis2 0 0.03fF $ **FLOATING
C3614 Dis2.t7 0 0.24fF
C3615 Dis2.t20 0 0.15fF
C3616 Dis2.n0 0 0.61fF $ **FLOATING
C3617 Dis2.t11 0 0.15fF
C3618 Dis2.t18 0 0.15fF
C3619 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_1/Dis 0 -0.29fF $ **FLOATING
C3620 Dis2.n1 0 0.32fF $ **FLOATING
C3621 Dis2.n2 0 0.55fF $ **FLOATING
C3622 Dis2.t5 0 0.15fF
C3623 Dis2.t10 0 0.15fF
C3624 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_2/Dis 0 -0.29fF $ **FLOATING
C3625 Dis2.n3 0 0.32fF $ **FLOATING
C3626 Dis2.n4 0 1.49fF $ **FLOATING
C3627 Dis2.t16 0 0.24fF
C3628 Dis2.t21 0 0.15fF
C3629 Dis2.n5 0 0.61fF $ **FLOATING
C3630 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/Dis 0 0.25fF $ **FLOATING
C3631 Dis2.n6 0 2.97fF $ **FLOATING
C3632 Dis2.t1 0 0.24fF
C3633 Dis2.t6 0 0.15fF
C3634 Dis2.n7 0 0.61fF $ **FLOATING
C3635 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/Dis 0 0.25fF $ **FLOATING
C3636 Dis2.n8 0 0.96fF $ **FLOATING
C3637 EESPFAL_Sbox_0/EESPFAL_s3_0/Dis2 0 0.75fF $ **FLOATING
C3638 EESPFAL_Sbox_0/EESPFAL_s2_0/Dis2 0 0.76fF $ **FLOATING
C3639 Dis2.t2 0 0.24fF
C3640 Dis2.t9 0 0.15fF
C3641 Dis2.n9 0 0.61fF $ **FLOATING
C3642 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/Dis 0 0.24fF $ **FLOATING
C3643 Dis2.n10 0 0.97fF $ **FLOATING
C3644 Dis2.t17 0 0.24fF
C3645 Dis2.t13 0 0.15fF
C3646 Dis2.n11 0 0.61fF $ **FLOATING
C3647 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_1/Dis 0 0.25fF $ **FLOATING
C3648 Dis2.n12 0 2.09fF $ **FLOATING
C3649 Dis2.n13 0 1.96fF $ **FLOATING
C3650 Dis2.t15 0 0.15fF
C3651 Dis2.t12 0 0.15fF
C3652 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_2/Dis 0 -0.29fF $ **FLOATING
C3653 Dis2.n14 0 0.32fF $ **FLOATING
C3654 Dis2.n15 0 0.68fF $ **FLOATING
C3655 Dis2.n16 0 1.90fF $ **FLOATING
C3656 Dis2.t14 0 0.24fF
C3657 Dis2.t8 0 0.15fF
C3658 Dis2.n17 0 0.61fF $ **FLOATING
C3659 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_1/Dis 0 0.25fF $ **FLOATING
C3660 Dis2.n18 0 2.11fF $ **FLOATING
C3661 Dis2.t3 0 0.24fF
C3662 Dis2.t19 0 0.15fF
C3663 Dis2.n19 0 0.61fF $ **FLOATING
C3664 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_NAND_v3_0/Dis 0 0.25fF $ **FLOATING
C3665 Dis2.n20 0 0.96fF $ **FLOATING
C3666 EESPFAL_Sbox_0/EESPFAL_s1_0/Dis2 0 1.40fF $ **FLOATING
C3667 Dis2.t0 0 0.15fF
C3668 Dis2.t4 0 0.15fF
C3669 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_1/Dis 0 -0.40fF $ **FLOATING
C3670 Dis2.n21 0 0.32fF $ **FLOATING
C3671 Dis2.n22 0 0.50fF $ **FLOATING
C3672 Dis2.n23 0 1.09fF $ **FLOATING
C3673 Dis2.n24 0 0.87fF $ **FLOATING
C3674 EESPFAL_Sbox_0/Dis2 0 0.70fF $ **FLOATING
C3675 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/OUT_bar 0 0.66fF $ **FLOATING
C3676 EESPFAL_Sbox_0/x3_bar 0 0.30fF $ **FLOATING
C3677 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t7 0 0.48fF
C3678 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t8 0 0.16fF
C3679 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n0 0 1.60fF $ **FLOATING
C3680 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n1 0 1.95fF $ **FLOATING
C3681 EESPFAL_Sbox_0/EESPFAL_s1_0/x3_bar 0 1.94fF $ **FLOATING
C3682 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t19 0 0.13fF
C3683 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0 0.43fF $ **FLOATING
C3684 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n2 0 3.97fF $ **FLOATING
C3685 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t17 0 0.48fF
C3686 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t18 0 0.16fF
C3687 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n3 0 1.60fF $ **FLOATING
C3688 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/B_bar 0 0.09fF $ **FLOATING
C3689 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t12 0 0.41fF
C3690 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A 0 1.79fF $ **FLOATING
C3691 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t10 0 0.38fF
C3692 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t11 0 0.21fF
C3693 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n4 0 1.97fF $ **FLOATING
C3694 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/A_bar 0 0.16fF $ **FLOATING
C3695 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t14 0 0.48fF
C3696 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t6 0 0.16fF
C3697 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n5 0 1.60fF $ **FLOATING
C3698 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/B_bar 0 0.09fF $ **FLOATING
C3699 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t16 0 0.14fF
C3700 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C_bar 0 0.38fF $ **FLOATING
C3701 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n6 0 4.12fF $ **FLOATING
C3702 EESPFAL_Sbox_0/EESPFAL_s3_0/x3_bar 0 1.13fF $ **FLOATING
C3703 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t13 0 0.18fF
C3704 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/A 0 0.76fF $ **FLOATING
C3705 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n7 0 4.72fF $ **FLOATING
C3706 EESPFAL_Sbox_0/EESPFAL_s2_0/x3_bar 0 0.48fF $ **FLOATING
C3707 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n8 0 1.63fF $ **FLOATING
C3708 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t20 0 0.31fF
C3709 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/A 0 2.36fF $ **FLOATING
C3710 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n9 0 3.28fF $ **FLOATING
C3711 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n10 0 2.48fF $ **FLOATING
C3712 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n11 0 1.16fF $ **FLOATING
C3713 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n12 0 1.15fF $ **FLOATING
C3714 EESPFAL_4in_XOR_0/XOR3_bar 0 0.50fF $ **FLOATING
C3715 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t4 0 0.14fF
C3716 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t0 0 0.14fF
C3717 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n13 0 0.42fF $ **FLOATING
C3718 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t1 0 0.53fF
C3719 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t5 0 0.92fF
C3720 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n14 0 0.81fF $ **FLOATING
C3721 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n15 0 0.35fF $ **FLOATING
C3722 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t2 0 0.14fF
C3723 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t3 0 0.14fF
C3724 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n16 0 0.35fF $ **FLOATING
C3725 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n17 0 0.38fF $ **FLOATING
C3726 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t9 0 0.13fF
C3727 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t21 0 0.18fF
C3728 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.t15 0 0.17fF
C3729 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n18 0 0.20fF $ **FLOATING
C3730 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar.n19 0 0.14fF $ **FLOATING
C3731 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t8 0 0.07fF
C3732 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t2 0 0.21fF
C3733 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t4 0 0.05fF
C3734 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t5 0 0.05fF
C3735 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n0 0 0.17fF $ **FLOATING
C3736 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t3 0 0.05fF
C3737 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t1 0 0.05fF
C3738 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n1 0 0.15fF $ **FLOATING
C3739 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t9 0 0.04fF
C3740 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t6 0 0.07fF
C3741 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t7 0 0.07fF
C3742 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n2 0 0.07fF $ **FLOATING
C3743 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT 0 0.01fF $ **FLOATING
C3744 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n3 0 0.04fF $ **FLOATING
C3745 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n4 0 0.22fF $ **FLOATING
C3746 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n5 0 0.22fF $ **FLOATING
C3747 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.t0 0 0.21fF
C3748 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar.n6 0 0.76fF $ **FLOATING
C3749 EESPFAL_Sbox_0/EESPFAL_s1_0/x2 0 2.02fF $ **FLOATING
C3750 EESPFAL_Sbox_0/x2 0 0.48fF $ **FLOATING
C3751 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t13 0 0.29fF
C3752 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t14 0 0.25fF
C3753 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n0 0 2.18fF $ **FLOATING
C3754 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/A 0 0.31fF $ **FLOATING
C3755 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t10 0 0.21fF
C3756 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n1 0 4.97fF $ **FLOATING
C3757 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t18 0 0.40fF
C3758 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/A 0 1.92fF $ **FLOATING
C3759 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n2 0 1.96fF $ **FLOATING
C3760 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t11 0 0.29fF
C3761 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_4in_NAND_0/D 0 2.20fF $ **FLOATING
C3762 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t7 0 0.29fF
C3763 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t17 0 0.25fF
C3764 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n3 0 2.18fF $ **FLOATING
C3765 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/A 0 0.31fF $ **FLOATING
C3766 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t12 0 0.24fF
C3767 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A_bar 0 0.73fF $ **FLOATING
C3768 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n4 0 4.63fF $ **FLOATING
C3769 EESPFAL_Sbox_0/EESPFAL_s3_0/x2 0 1.89fF $ **FLOATING
C3770 EESPFAL_Sbox_0/EESPFAL_s2_0/x2 0 0.67fF $ **FLOATING
C3771 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t6 0 0.20fF
C3772 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t20 0 0.19fF
C3773 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n5 0 2.27fF $ **FLOATING
C3774 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/B 0 0.37fF $ **FLOATING
C3775 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n6 0 1.32fF $ **FLOATING
C3776 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t9 0 0.14fF
C3777 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/A_bar 0 0.49fF $ **FLOATING
C3778 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n7 0 5.82fF $ **FLOATING
C3779 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n8 0 3.26fF $ **FLOATING
C3780 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t16 0 0.19fF
C3781 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/A 0 0.88fF $ **FLOATING
C3782 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n9 0 8.19fF $ **FLOATING
C3783 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n10 0 0.46fF $ **FLOATING
C3784 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t5 0 0.65fF
C3785 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t4 0 0.15fF
C3786 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t2 0 0.15fF
C3787 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n11 0 0.47fF $ **FLOATING
C3788 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t3 0 0.15fF
C3789 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t1 0 0.15fF
C3790 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n12 0 0.51fF $ **FLOATING
C3791 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t15 0 0.20fF
C3792 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t8 0 0.22fF
C3793 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t19 0 0.11fF
C3794 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n13 0 0.22fF $ **FLOATING
C3795 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_2/OUT 0 0.04fF $ **FLOATING
C3796 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n14 0 0.11fF $ **FLOATING
C3797 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n15 0 0.67fF $ **FLOATING
C3798 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n16 0 0.67fF $ **FLOATING
C3799 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.t0 0 0.65fF
C3800 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar.n17 0 0.57fF $ **FLOATING
C3801 EESPFAL_4in_XOR_0/XOR2 0 0.21fF $ **FLOATING
C3802 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t7 0 0.04fF
C3803 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/A_bar 0 0.53fF $ **FLOATING
C3804 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t4 0 0.04fF
C3805 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t2 0 0.04fF
C3806 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n0 0 0.09fF $ **FLOATING
C3807 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t3 0 0.04fF
C3808 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t1 0 0.04fF
C3809 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n1 0 0.11fF $ **FLOATING
C3810 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t5 0 0.20fF
C3811 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t0 0 0.13fF
C3812 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n2 0 0.19fF $ **FLOATING
C3813 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n3 0 0.09fF $ **FLOATING
C3814 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n4 0 0.10fF $ **FLOATING
C3815 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t9 0 0.05fF
C3816 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t8 0 0.04fF
C3817 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t6 0 0.03fF
C3818 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n5 0 0.05fF $ **FLOATING
C3819 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n6 0 0.04fF $ **FLOATING
C3820 EESPFAL_Sbox_0/EESPFAL_s1_0/s1_bar 0 0.01fF $ **FLOATING
C3821 s1_bar.t2 0 0.05fF
C3822 s1_bar.t3 0 0.05fF
C3823 s1_bar.n0 0 0.12fF $ **FLOATING
C3824 s1_bar.t0 0 0.05fF
C3825 s1_bar.t1 0 0.05fF
C3826 s1_bar.n1 0 0.14fF $ **FLOATING
C3827 s1_bar.t4 0 0.27fF
C3828 s1_bar.n2 0 0.19fF $ **FLOATING
C3829 s1_bar.n3 0 0.13fF $ **FLOATING
C3830 s1_bar.t7 0 0.06fF
C3831 s1_bar.t5 0 0.06fF
C3832 s1_bar.t6 0 0.04fF
C3833 s1_bar.n4 0 0.07fF $ **FLOATING
C3834 s1_bar.n5 0 0.05fF $ **FLOATING
C3835 EESPFAL_Sbox_0/s1_bar 0 0.56fF $ **FLOATING
C3836 Dis3.t6 0 0.14fF
C3837 Dis3.t2 0 0.15fF
C3838 Dis3.n0 0 0.44fF $ **FLOATING
C3839 Dis3.t4 0 0.14fF
C3840 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/Dis 0 -0.17fF $ **FLOATING
C3841 Dis3.t1 0 0.15fF
C3842 Dis3.n1 0 0.72fF $ **FLOATING
C3843 EESPFAL_Sbox_0/EESPFAL_s3_0/Dis3 0 3.46fF $ **FLOATING
C3844 EESPFAL_Sbox_0/EESPFAL_s2_0/Dis3 0 0.20fF $ **FLOATING
C3845 Dis3.n2 0 1.38fF $ **FLOATING
C3846 Dis3.t5 0 0.14fF
C3847 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/Dis 0 -0.17fF $ **FLOATING
C3848 Dis3.t7 0 0.15fF
C3849 Dis3.n3 0 0.64fF $ **FLOATING
C3850 Dis3.n4 0 2.12fF $ **FLOATING
C3851 Dis3.t0 0 0.14fF
C3852 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/Dis 0 -0.17fF $ **FLOATING
C3853 Dis3.t3 0 0.15fF
C3854 Dis3.n5 0 0.64fF $ **FLOATING
C3855 Dis3.n6 0 2.14fF $ **FLOATING
C3856 EESPFAL_Sbox_0/EESPFAL_s1_0/Dis3 0 2.12fF $ **FLOATING
C3857 Dis3.n7 0 1.74fF $ **FLOATING
C3858 EESPFAL_Sbox_0/Dis3 0 0.54fF $ **FLOATING
C3859 EESPFAL_Sbox_0/EESPFAL_s0_0/Dis3 0 0.02fF $ **FLOATING
C3860 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT_bar 0 0.50fF $ **FLOATING
C3861 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t9 0 0.07fF
C3862 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t5 0 0.05fF
C3863 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t1 0 0.05fF
C3864 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n0 0 0.15fF $ **FLOATING
C3865 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t0 0 0.19fF
C3866 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t2 0 0.33fF
C3867 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n1 0 0.29fF $ **FLOATING
C3868 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n2 0 0.12fF $ **FLOATING
C3869 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t3 0 0.05fF
C3870 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t4 0 0.05fF
C3871 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n3 0 0.13fF $ **FLOATING
C3872 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n4 0 0.14fF $ **FLOATING
C3873 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t7 0 0.05fF
C3874 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t6 0 0.06fF
C3875 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t8 0 0.06fF
C3876 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n5 0 0.07fF $ **FLOATING
C3877 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n6 0 0.05fF $ **FLOATING
C3878 CLK1.t80 0 0.03fF
C3879 CLK1.t154 0 0.03fF
C3880 CLK1.n0 0 0.15fF $ **FLOATING
C3881 CLK1.t176 0 0.05fF
C3882 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_XOR_v3_0/CLK 0 0.02fF $ **FLOATING
C3883 CLK1.n1 0 0.17fF $ **FLOATING
C3884 CLK1.n2 0 0.03fF $ **FLOATING
C3885 CLK1.t188 0 0.03fF
C3886 CLK1.t174 0 0.03fF
C3887 CLK1.n3 0 0.10fF $ **FLOATING
C3888 CLK1.t194 0 0.05fF
C3889 CLK1.t137 0 0.03fF
C3890 CLK1.t79 0 0.03fF
C3891 CLK1.n4 0 0.15fF $ **FLOATING
C3892 CLK1.t177 0 0.08fF
C3893 CLK1.t93 0 0.05fF
C3894 CLK1.n5 0 0.17fF $ **FLOATING
C3895 CLK1.n6 0 0.03fF $ **FLOATING
C3896 CLK1.t56 0 0.03fF
C3897 CLK1.t95 0 0.03fF
C3898 CLK1.n7 0 0.10fF $ **FLOATING
C3899 CLK1.t54 0 0.05fF
C3900 CLK1.t33 0 0.03fF
C3901 CLK1.t102 0 0.03fF
C3902 CLK1.n8 0 0.15fF $ **FLOATING
C3903 CLK1.n9 0 0.08fF $ **FLOATING
C3904 CLK1.n10 0 0.03fF $ **FLOATING
C3905 CLK1.n11 0 0.02fF $ **FLOATING
C3906 CLK1.n12 0 0.13fF $ **FLOATING
C3907 CLK1.n13 0 0.06fF $ **FLOATING
C3908 CLK1.n14 0 0.03fF $ **FLOATING
C3909 CLK1.n15 0 0.02fF $ **FLOATING
C3910 CLK1.n16 0 0.07fF $ **FLOATING
C3911 CLK1.n17 0 0.19fF $ **FLOATING
C3912 CLK1.n18 0 0.06fF $ **FLOATING
C3913 CLK1.n19 0 0.03fF $ **FLOATING
C3914 CLK1.n20 0 0.02fF $ **FLOATING
C3915 CLK1.n21 0 0.03fF $ **FLOATING
C3916 CLK1.n22 0 0.06fF $ **FLOATING
C3917 CLK1.n23 0 0.03fF $ **FLOATING
C3918 CLK1.n24 0 0.02fF $ **FLOATING
C3919 CLK1.n25 0 0.03fF $ **FLOATING
C3920 CLK1.n26 0 0.14fF $ **FLOATING
C3921 CLK1.n27 0 0.03fF $ **FLOATING
C3922 CLK1.n28 0 0.02fF $ **FLOATING
C3923 CLK1.n29 0 0.03fF $ **FLOATING
C3924 CLK1.n30 0 0.18fF $ **FLOATING
C3925 CLK1.n31 0 0.03fF $ **FLOATING
C3926 CLK1.n32 0 0.02fF $ **FLOATING
C3927 CLK1.n33 0 0.02fF $ **FLOATING
C3928 CLK1.n34 0 0.29fF $ **FLOATING
C3929 CLK1.t53 0 0.09fF
C3930 CLK1.n35 0 0.11fF $ **FLOATING
C3931 CLK1.n36 0 0.03fF $ **FLOATING
C3932 CLK1.n37 0 0.02fF $ **FLOATING
C3933 CLK1.n38 0 0.03fF $ **FLOATING
C3934 CLK1.n39 0 0.16fF $ **FLOATING
C3935 CLK1.n40 0 0.03fF $ **FLOATING
C3936 CLK1.n41 0 0.02fF $ **FLOATING
C3937 CLK1.n42 0 0.03fF $ **FLOATING
C3938 CLK1.t55 0 0.09fF
C3939 CLK1.n43 0 0.09fF $ **FLOATING
C3940 CLK1.n44 0 0.03fF $ **FLOATING
C3941 CLK1.n45 0 0.02fF $ **FLOATING
C3942 CLK1.n46 0 0.03fF $ **FLOATING
C3943 CLK1.n47 0 0.17fF $ **FLOATING
C3944 CLK1.n48 0 0.02fF $ **FLOATING
C3945 CLK1.t94 0 0.09fF
C3946 CLK1.n49 0 0.09fF $ **FLOATING
C3947 CLK1.n50 0 0.03fF $ **FLOATING
C3948 CLK1.n51 0 0.02fF $ **FLOATING
C3949 CLK1.n52 0 0.03fF $ **FLOATING
C3950 CLK1.n53 0 0.16fF $ **FLOATING
C3951 CLK1.n54 0 0.03fF $ **FLOATING
C3952 CLK1.n55 0 0.02fF $ **FLOATING
C3953 CLK1.n56 0 0.03fF $ **FLOATING
C3954 CLK1.t92 0 0.09fF
C3955 CLK1.n57 0 0.11fF $ **FLOATING
C3956 CLK1.n58 0 0.03fF $ **FLOATING
C3957 CLK1.n59 0 0.02fF $ **FLOATING
C3958 CLK1.n60 0 0.03fF $ **FLOATING
C3959 CLK1.n61 0 0.29fF $ **FLOATING
C3960 CLK1.n62 0 0.18fF $ **FLOATING
C3961 CLK1.n63 0 0.03fF $ **FLOATING
C3962 CLK1.n64 0 0.02fF $ **FLOATING
C3963 CLK1.n65 0 0.02fF $ **FLOATING
C3964 CLK1.n66 0 0.14fF $ **FLOATING
C3965 CLK1.n67 0 0.03fF $ **FLOATING
C3966 CLK1.n68 0 0.02fF $ **FLOATING
C3967 CLK1.n69 0 0.03fF $ **FLOATING
C3968 CLK1.n70 0 0.06fF $ **FLOATING
C3969 CLK1.n71 0 0.03fF $ **FLOATING
C3970 CLK1.n72 0 0.02fF $ **FLOATING
C3971 CLK1.n73 0 0.03fF $ **FLOATING
C3972 CLK1.n74 0 0.06fF $ **FLOATING
C3973 CLK1.n75 0 0.03fF $ **FLOATING
C3974 CLK1.n76 0 0.02fF $ **FLOATING
C3975 CLK1.n77 0 0.03fF $ **FLOATING
C3976 CLK1.n78 0 0.06fF $ **FLOATING
C3977 CLK1.n79 0 0.03fF $ **FLOATING
C3978 CLK1.n80 0 0.02fF $ **FLOATING
C3979 CLK1.n81 0 0.03fF $ **FLOATING
C3980 CLK1.n82 0 0.07fF $ **FLOATING
C3981 CLK1.n83 0 0.03fF $ **FLOATING
C3982 CLK1.n84 0 0.02fF $ **FLOATING
C3983 CLK1.n85 0 0.03fF $ **FLOATING
C3984 CLK1.n86 0 0.34fF $ **FLOATING
C3985 CLK1.n87 0 0.13fF $ **FLOATING
C3986 CLK1.n88 0 0.10fF $ **FLOATING
C3987 CLK1.n89 0 0.21fF $ **FLOATING
C3988 CLK1.n90 0 0.11fF $ **FLOATING
C3989 CLK1.n91 0 0.08fF $ **FLOATING
C3990 CLK1.n92 0 0.03fF $ **FLOATING
C3991 CLK1.n93 0 0.02fF $ **FLOATING
C3992 CLK1.n94 0 0.03fF $ **FLOATING
C3993 CLK1.n95 0 0.06fF $ **FLOATING
C3994 CLK1.n96 0 0.03fF $ **FLOATING
C3995 CLK1.n97 0 0.02fF $ **FLOATING
C3996 CLK1.n98 0 0.03fF $ **FLOATING
C3997 CLK1.n99 0 0.06fF $ **FLOATING
C3998 CLK1.n100 0 0.03fF $ **FLOATING
C3999 CLK1.n101 0 0.02fF $ **FLOATING
C4000 CLK1.n102 0 0.02fF $ **FLOATING
C4001 CLK1.n103 0 0.19fF $ **FLOATING
C4002 CLK1.n104 0 0.06fF $ **FLOATING
C4003 CLK1.n105 0 0.03fF $ **FLOATING
C4004 CLK1.n106 0 0.02fF $ **FLOATING
C4005 CLK1.n107 0 0.03fF $ **FLOATING
C4006 CLK1.n108 0 0.06fF $ **FLOATING
C4007 CLK1.n109 0 0.03fF $ **FLOATING
C4008 CLK1.n110 0 0.02fF $ **FLOATING
C4009 CLK1.n111 0 0.03fF $ **FLOATING
C4010 CLK1.n112 0 0.06fF $ **FLOATING
C4011 CLK1.n113 0 0.03fF $ **FLOATING
C4012 CLK1.n114 0 0.02fF $ **FLOATING
C4013 CLK1.n115 0 0.03fF $ **FLOATING
C4014 CLK1.n116 0 0.06fF $ **FLOATING
C4015 CLK1.n117 0 0.03fF $ **FLOATING
C4016 CLK1.n118 0 0.02fF $ **FLOATING
C4017 CLK1.n119 0 0.03fF $ **FLOATING
C4018 CLK1.n120 0 0.14fF $ **FLOATING
C4019 CLK1.n121 0 0.03fF $ **FLOATING
C4020 CLK1.n122 0 0.02fF $ **FLOATING
C4021 CLK1.n123 0 0.03fF $ **FLOATING
C4022 CLK1.n124 0 0.18fF $ **FLOATING
C4023 CLK1.n125 0 0.03fF $ **FLOATING
C4024 CLK1.n126 0 0.02fF $ **FLOATING
C4025 CLK1.n127 0 0.02fF $ **FLOATING
C4026 CLK1.n128 0 0.29fF $ **FLOATING
C4027 CLK1.t193 0 0.09fF
C4028 CLK1.n129 0 0.11fF $ **FLOATING
C4029 CLK1.n130 0 0.03fF $ **FLOATING
C4030 CLK1.n131 0 0.02fF $ **FLOATING
C4031 CLK1.n132 0 0.03fF $ **FLOATING
C4032 CLK1.n133 0 0.16fF $ **FLOATING
C4033 CLK1.n134 0 0.03fF $ **FLOATING
C4034 CLK1.n135 0 0.02fF $ **FLOATING
C4035 CLK1.n136 0 0.03fF $ **FLOATING
C4036 CLK1.t187 0 0.09fF
C4037 CLK1.n137 0 0.09fF $ **FLOATING
C4038 CLK1.n138 0 0.03fF $ **FLOATING
C4039 CLK1.n139 0 0.02fF $ **FLOATING
C4040 CLK1.n140 0 0.03fF $ **FLOATING
C4041 CLK1.n141 0 0.17fF $ **FLOATING
C4042 CLK1.n142 0 0.02fF $ **FLOATING
C4043 CLK1.t173 0 0.09fF
C4044 CLK1.n143 0 0.09fF $ **FLOATING
C4045 CLK1.n144 0 0.03fF $ **FLOATING
C4046 CLK1.n145 0 0.02fF $ **FLOATING
C4047 CLK1.n146 0 0.03fF $ **FLOATING
C4048 CLK1.n147 0 0.16fF $ **FLOATING
C4049 CLK1.n148 0 0.03fF $ **FLOATING
C4050 CLK1.n149 0 0.02fF $ **FLOATING
C4051 CLK1.n150 0 0.03fF $ **FLOATING
C4052 CLK1.t175 0 0.09fF
C4053 CLK1.n151 0 0.11fF $ **FLOATING
C4054 CLK1.n152 0 0.03fF $ **FLOATING
C4055 CLK1.n153 0 0.02fF $ **FLOATING
C4056 CLK1.n154 0 0.03fF $ **FLOATING
C4057 CLK1.n155 0 0.29fF $ **FLOATING
C4058 CLK1.n156 0 0.18fF $ **FLOATING
C4059 CLK1.n157 0 0.03fF $ **FLOATING
C4060 CLK1.n158 0 0.02fF $ **FLOATING
C4061 CLK1.n159 0 0.02fF $ **FLOATING
C4062 CLK1.n160 0 0.14fF $ **FLOATING
C4063 CLK1.n161 0 0.03fF $ **FLOATING
C4064 CLK1.n162 0 0.02fF $ **FLOATING
C4065 CLK1.n163 0 0.03fF $ **FLOATING
C4066 CLK1.n164 0 0.06fF $ **FLOATING
C4067 CLK1.n165 0 0.03fF $ **FLOATING
C4068 CLK1.n166 0 0.02fF $ **FLOATING
C4069 CLK1.n167 0 0.03fF $ **FLOATING
C4070 CLK1.n168 0 0.06fF $ **FLOATING
C4071 CLK1.n169 0 0.03fF $ **FLOATING
C4072 CLK1.n170 0 0.02fF $ **FLOATING
C4073 CLK1.n171 0 0.03fF $ **FLOATING
C4074 CLK1.n172 0 0.06fF $ **FLOATING
C4075 CLK1.n173 0 0.03fF $ **FLOATING
C4076 CLK1.n174 0 0.02fF $ **FLOATING
C4077 CLK1.n175 0 0.03fF $ **FLOATING
C4078 CLK1.n176 0 0.06fF $ **FLOATING
C4079 CLK1.n177 0 0.03fF $ **FLOATING
C4080 CLK1.n178 0 0.02fF $ **FLOATING
C4081 CLK1.n179 0 0.03fF $ **FLOATING
C4082 CLK1.n180 0 0.19fF $ **FLOATING
C4083 CLK1.n181 0 0.06fF $ **FLOATING
C4084 CLK1.n182 0 0.03fF $ **FLOATING
C4085 CLK1.n183 0 0.02fF $ **FLOATING
C4086 CLK1.n184 0 0.02fF $ **FLOATING
C4087 CLK1.n185 0 0.06fF $ **FLOATING
C4088 CLK1.n186 0 0.03fF $ **FLOATING
C4089 CLK1.n187 0 0.02fF $ **FLOATING
C4090 CLK1.n188 0 0.03fF $ **FLOATING
C4091 CLK1.n189 0 0.08fF $ **FLOATING
C4092 CLK1.n190 0 0.03fF $ **FLOATING
C4093 CLK1.n191 0 0.02fF $ **FLOATING
C4094 CLK1.n192 0 0.03fF $ **FLOATING
C4095 CLK1.n193 0 0.21fF $ **FLOATING
C4096 CLK1.n194 0 0.05fF $ **FLOATING
C4097 CLK1.n195 0 0.03fF $ **FLOATING
C4098 CLK1.n196 0 0.02fF $ **FLOATING
C4099 CLK1.n197 0 0.03fF $ **FLOATING
C4100 CLK1.n198 0 0.06fF $ **FLOATING
C4101 CLK1.n199 0 0.03fF $ **FLOATING
C4102 CLK1.n200 0 0.02fF $ **FLOATING
C4103 CLK1.t150 0 0.03fF
C4104 CLK1.t32 0 0.03fF
C4105 CLK1.n201 0 0.15fF $ **FLOATING
C4106 CLK1.n202 0 0.03fF $ **FLOATING
C4107 CLK1.n203 0 0.02fF $ **FLOATING
C4108 CLK1.n204 0 0.03fF $ **FLOATING
C4109 CLK1.n205 0 0.11fF $ **FLOATING
C4110 CLK1.n206 0 0.03fF $ **FLOATING
C4111 CLK1.n207 0 0.02fF $ **FLOATING
C4112 CLK1.t139 0 0.05fF
C4113 CLK1.n208 0 0.03fF $ **FLOATING
C4114 CLK1.n209 0 0.02fF $ **FLOATING
C4115 CLK1.n210 0 0.03fF $ **FLOATING
C4116 CLK1.t89 0 0.09fF
C4117 CLK1.n211 0 0.03fF $ **FLOATING
C4118 CLK1.n212 0 0.02fF $ **FLOATING
C4119 CLK1.t90 0 0.03fF
C4120 CLK1.t141 0 0.03fF
C4121 CLK1.n213 0 0.10fF $ **FLOATING
C4122 CLK1.n214 0 0.03fF $ **FLOATING
C4123 CLK1.n215 0 0.02fF $ **FLOATING
C4124 CLK1.n216 0 0.03fF $ **FLOATING
C4125 CLK1.n217 0 0.14fF $ **FLOATING
C4126 CLK1.n218 0 0.03fF $ **FLOATING
C4127 CLK1.n219 0 0.02fF $ **FLOATING
C4128 CLK1.n220 0 0.03fF $ **FLOATING
C4129 CLK1.n221 0 0.02fF $ **FLOATING
C4130 CLK1.n222 0 0.03fF $ **FLOATING
C4131 CLK1.n223 0 0.07fF $ **FLOATING
C4132 CLK1.n224 0 0.03fF $ **FLOATING
C4133 CLK1.n225 0 0.02fF $ **FLOATING
C4134 CLK1.t113 0 0.08fF
C4135 CLK1.n226 0 0.13fF $ **FLOATING
C4136 CLK1.n227 0 0.36fF $ **FLOATING
C4137 CLK1.n228 0 0.03fF $ **FLOATING
C4138 CLK1.n229 0 0.03fF $ **FLOATING
C4139 CLK1.n230 0 0.02fF $ **FLOATING
C4140 CLK1.n231 0 0.03fF $ **FLOATING
C4141 CLK1.n232 0 0.06fF $ **FLOATING
C4142 CLK1.n233 0 0.06fF $ **FLOATING
C4143 CLK1.n234 0 0.06fF $ **FLOATING
C4144 CLK1.n235 0 0.03fF $ **FLOATING
C4145 CLK1.n236 0 0.02fF $ **FLOATING
C4146 CLK1.n237 0 0.03fF $ **FLOATING
C4147 CLK1.n238 0 0.03fF $ **FLOATING
C4148 CLK1.t88 0 0.05fF
C4149 CLK1.n239 0 0.29fF $ **FLOATING
C4150 CLK1.n240 0 0.02fF $ **FLOATING
C4151 CLK1.n241 0 0.02fF $ **FLOATING
C4152 CLK1.n242 0 0.03fF $ **FLOATING
C4153 CLK1.n243 0 0.18fF $ **FLOATING
C4154 CLK1.n244 0 0.11fF $ **FLOATING
C4155 CLK1.t87 0 0.09fF
C4156 CLK1.n245 0 0.09fF $ **FLOATING
C4157 CLK1.n246 0 0.16fF $ **FLOATING
C4158 CLK1.n247 0 0.03fF $ **FLOATING
C4159 CLK1.n248 0 0.02fF $ **FLOATING
C4160 CLK1.n249 0 0.03fF $ **FLOATING
C4161 CLK1.n250 0 0.03fF $ **FLOATING
C4162 EESPFAL_Sbox_0/EESPFAL_s0_0/EESPFAL_NAND_v3_2/CLK 0 0.02fF $ **FLOATING
C4163 CLK1.n251 0 0.17fF $ **FLOATING
C4164 CLK1.n252 0 0.02fF $ **FLOATING
C4165 CLK1.n253 0 0.03fF $ **FLOATING
C4166 CLK1.n254 0 0.17fF $ **FLOATING
C4167 CLK1.t140 0 0.09fF
C4168 CLK1.n255 0 0.09fF $ **FLOATING
C4169 CLK1.t138 0 0.09fF
C4170 CLK1.n256 0 0.16fF $ **FLOATING
C4171 CLK1.n257 0 0.03fF $ **FLOATING
C4172 CLK1.n258 0 0.02fF $ **FLOATING
C4173 CLK1.n259 0 0.03fF $ **FLOATING
C4174 CLK1.n260 0 0.03fF $ **FLOATING
C4175 CLK1.n261 0 0.29fF $ **FLOATING
C4176 CLK1.n262 0 0.02fF $ **FLOATING
C4177 CLK1.n263 0 0.02fF $ **FLOATING
C4178 CLK1.n264 0 0.03fF $ **FLOATING
C4179 CLK1.n265 0 0.18fF $ **FLOATING
C4180 CLK1.n266 0 0.14fF $ **FLOATING
C4181 CLK1.n267 0 0.06fF $ **FLOATING
C4182 CLK1.n268 0 0.03fF $ **FLOATING
C4183 CLK1.n269 0 0.02fF $ **FLOATING
C4184 CLK1.n270 0 0.03fF $ **FLOATING
C4185 CLK1.n271 0 0.03fF $ **FLOATING
C4186 CLK1.n272 0 0.19fF $ **FLOATING
C4187 CLK1.n273 0 0.02fF $ **FLOATING
C4188 CLK1.n274 0 0.02fF $ **FLOATING
C4189 CLK1.n275 0 0.03fF $ **FLOATING
C4190 CLK1.n276 0 0.06fF $ **FLOATING
C4191 CLK1.n277 0 0.07fF $ **FLOATING
C4192 CLK1.n278 0 0.13fF $ **FLOATING
C4193 CLK1.n279 0 0.14fF $ **FLOATING
C4194 CLK1.n280 0 0.00fF $ **FLOATING
C4195 EESPFAL_Sbox_0/EESPFAL_s1_0/CLK1 0 0.00fF $ **FLOATING
C4196 CLK1.n281 0 0.01fF $ **FLOATING
C4197 CLK1.t81 0 0.08fF
C4198 CLK1.n282 0 0.34fF $ **FLOATING
C4199 CLK1.n283 0 0.02fF $ **FLOATING
C4200 CLK1.n284 0 0.03fF $ **FLOATING
C4201 CLK1.n285 0 0.06fF $ **FLOATING
C4202 CLK1.n286 0 0.03fF $ **FLOATING
C4203 CLK1.n287 0 0.02fF $ **FLOATING
C4204 CLK1.t167 0 0.03fF
C4205 CLK1.t178 0 0.03fF
C4206 CLK1.n288 0 0.15fF $ **FLOATING
C4207 CLK1.n289 0 0.19fF $ **FLOATING
C4208 CLK1.n290 0 0.02fF $ **FLOATING
C4209 CLK1.n291 0 0.03fF $ **FLOATING
C4210 CLK1.n292 0 0.14fF $ **FLOATING
C4211 CLK1.n293 0 0.03fF $ **FLOATING
C4212 CLK1.n294 0 0.02fF $ **FLOATING
C4213 CLK1.t17 0 0.05fF
C4214 CLK1.n295 0 0.29fF $ **FLOATING
C4215 CLK1.n296 0 0.02fF $ **FLOATING
C4216 CLK1.n297 0 0.03fF $ **FLOATING
C4217 CLK1.n298 0 0.09fF $ **FLOATING
C4218 CLK1.n299 0 0.03fF $ **FLOATING
C4219 CLK1.n300 0 0.02fF $ **FLOATING
C4220 CLK1.t130 0 0.03fF
C4221 CLK1.t15 0 0.03fF
C4222 CLK1.n301 0 0.10fF $ **FLOATING
C4223 CLK1.n302 0 0.03fF $ **FLOATING
C4224 CLK1.n303 0 0.02fF $ **FLOATING
C4225 CLK1.n304 0 0.03fF $ **FLOATING
C4226 CLK1.t131 0 0.09fF
C4227 CLK1.n305 0 0.03fF $ **FLOATING
C4228 CLK1.n306 0 0.02fF $ **FLOATING
C4229 CLK1.t132 0 0.05fF
C4230 CLK1.n307 0 0.03fF $ **FLOATING
C4231 CLK1.n308 0 0.02fF $ **FLOATING
C4232 CLK1.n309 0 0.03fF $ **FLOATING
C4233 CLK1.n310 0 0.06fF $ **FLOATING
C4234 CLK1.n311 0 0.03fF $ **FLOATING
C4235 CLK1.n312 0 0.02fF $ **FLOATING
C4236 CLK1.n313 0 0.03fF $ **FLOATING
C4237 CLK1.n314 0 0.02fF $ **FLOATING
C4238 CLK1.n315 0 0.03fF $ **FLOATING
C4239 CLK1.n316 0 0.07fF $ **FLOATING
C4240 CLK1.n317 0 0.03fF $ **FLOATING
C4241 CLK1.n318 0 0.02fF $ **FLOATING
C4242 CLK1.n319 0 0.02fF $ **FLOATING
C4243 CLK1.n320 0 0.02fF $ **FLOATING
C4244 CLK1.n321 0 0.02fF $ **FLOATING
C4245 CLK1.t198 0 0.03fF
C4246 CLK1.t122 0 0.07fF
C4247 CLK1.n322 0 0.45fF $ **FLOATING
C4248 CLK1.n323 0 0.02fF $ **FLOATING
C4249 CLK1.n324 0 0.03fF $ **FLOATING
C4250 CLK1.n325 0 0.14fF $ **FLOATING
C4251 CLK1.n326 0 0.03fF $ **FLOATING
C4252 CLK1.n327 0 0.02fF $ **FLOATING
C4253 CLK1.t182 0 0.05fF
C4254 CLK1.n328 0 0.29fF $ **FLOATING
C4255 CLK1.n329 0 0.02fF $ **FLOATING
C4256 CLK1.n330 0 0.03fF $ **FLOATING
C4257 CLK1.n331 0 0.09fF $ **FLOATING
C4258 CLK1.n332 0 0.03fF $ **FLOATING
C4259 CLK1.n333 0 0.02fF $ **FLOATING
C4260 CLK1.t126 0 0.03fF
C4261 CLK1.t180 0 0.03fF
C4262 CLK1.n334 0 0.10fF $ **FLOATING
C4263 CLK1.n335 0 0.03fF $ **FLOATING
C4264 CLK1.n336 0 0.02fF $ **FLOATING
C4265 CLK1.n337 0 0.03fF $ **FLOATING
C4266 CLK1.t127 0 0.09fF
C4267 CLK1.n338 0 0.03fF $ **FLOATING
C4268 CLK1.n339 0 0.02fF $ **FLOATING
C4269 CLK1.t128 0 0.05fF
C4270 CLK1.n340 0 0.03fF $ **FLOATING
C4271 CLK1.n341 0 0.02fF $ **FLOATING
C4272 CLK1.n342 0 0.03fF $ **FLOATING
C4273 CLK1.n343 0 0.07fF $ **FLOATING
C4274 CLK1.n344 0 0.03fF $ **FLOATING
C4275 CLK1.n345 0 0.02fF $ **FLOATING
C4276 CLK1.t22 0 0.07fF
C4277 CLK1.n346 0 0.15fF $ **FLOATING
C4278 CLK1.n347 0 0.47fF $ **FLOATING
C4279 CLK1.n348 0 0.03fF $ **FLOATING
C4280 CLK1.n349 0 0.03fF $ **FLOATING
C4281 CLK1.n350 0 0.02fF $ **FLOATING
C4282 CLK1.n351 0 0.03fF $ **FLOATING
C4283 CLK1.n352 0 0.06fF $ **FLOATING
C4284 CLK1.n353 0 0.14fF $ **FLOATING
C4285 CLK1.n354 0 0.11fF $ **FLOATING
C4286 CLK1.n355 0 0.18fF $ **FLOATING
C4287 CLK1.n356 0 0.03fF $ **FLOATING
C4288 CLK1.n357 0 0.02fF $ **FLOATING
C4289 CLK1.n358 0 0.02fF $ **FLOATING
C4290 CLK1.n359 0 0.29fF $ **FLOATING
C4291 CLK1.n360 0 0.03fF $ **FLOATING
C4292 CLK1.n361 0 0.03fF $ **FLOATING
C4293 CLK1.n362 0 0.02fF $ **FLOATING
C4294 CLK1.n363 0 0.03fF $ **FLOATING
C4295 CLK1.n364 0 0.16fF $ **FLOATING
C4296 CLK1.n365 0 0.09fF $ **FLOATING
C4297 CLK1.t125 0 0.09fF
C4298 CLK1.t179 0 0.09fF
C4299 CLK1.n366 0 0.17fF $ **FLOATING
C4300 CLK1.n367 0 0.03fF $ **FLOATING
C4301 CLK1.n368 0 0.02fF $ **FLOATING
C4302 CLK1.n369 0 0.17fF $ **FLOATING
C4303 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_2/CLK 0 0.02fF $ **FLOATING
C4304 CLK1.n370 0 0.03fF $ **FLOATING
C4305 CLK1.n371 0 0.03fF $ **FLOATING
C4306 CLK1.n372 0 0.03fF $ **FLOATING
C4307 CLK1.n373 0 0.02fF $ **FLOATING
C4308 CLK1.n374 0 0.03fF $ **FLOATING
C4309 CLK1.n375 0 0.16fF $ **FLOATING
C4310 CLK1.t181 0 0.09fF
C4311 CLK1.n376 0 0.11fF $ **FLOATING
C4312 CLK1.n377 0 0.18fF $ **FLOATING
C4313 CLK1.n378 0 0.03fF $ **FLOATING
C4314 CLK1.n379 0 0.02fF $ **FLOATING
C4315 CLK1.n380 0 0.02fF $ **FLOATING
C4316 CLK1.n381 0 0.03fF $ **FLOATING
C4317 CLK1.n382 0 0.03fF $ **FLOATING
C4318 CLK1.n383 0 0.03fF $ **FLOATING
C4319 CLK1.n384 0 0.02fF $ **FLOATING
C4320 CLK1.n385 0 0.03fF $ **FLOATING
C4321 CLK1.n386 0 0.06fF $ **FLOATING
C4322 CLK1.n387 0 0.07fF $ **FLOATING
C4323 CLK1.n388 0 0.15fF $ **FLOATING
C4324 CLK1.n389 0 0.08fF $ **FLOATING
C4325 CLK1.n390 0 0.13fF $ **FLOATING
C4326 CLK1.n391 0 0.07fF $ **FLOATING
C4327 CLK1.n392 0 0.26fF $ **FLOATING
C4328 CLK1.n393 0 0.07fF $ **FLOATING
C4329 CLK1.n394 0 0.07fF $ **FLOATING
C4330 CLK1.n395 0 0.10fF $ **FLOATING
C4331 CLK1.n396 0 0.07fF $ **FLOATING
C4332 CLK1.n397 0 0.07fF $ **FLOATING
C4333 CLK1.n398 0 0.03fF $ **FLOATING
C4334 CLK1.n399 0 0.02fF $ **FLOATING
C4335 CLK1.n400 0 0.02fF $ **FLOATING
C4336 CLK1.t96 0 0.03fF
C4337 CLK1.n401 0 0.02fF $ **FLOATING
C4338 CLK1.n402 0 0.03fF $ **FLOATING
C4339 CLK1.n403 0 0.02fF $ **FLOATING
C4340 CLK1.n404 0 0.02fF $ **FLOATING
C4341 CLK1.n405 0 0.03fF $ **FLOATING
C4342 CLK1.n406 0 0.03fF $ **FLOATING
C4343 CLK1.n407 0 0.08fF $ **FLOATING
C4344 CLK1.n408 0 0.03fF $ **FLOATING
C4345 CLK1.n409 0 0.02fF $ **FLOATING
C4346 CLK1.t36 0 0.07fF
C4347 CLK1.n410 0 0.45fF $ **FLOATING
C4348 CLK1.n411 0 0.02fF $ **FLOATING
C4349 CLK1.n412 0 0.03fF $ **FLOATING
C4350 CLK1.n413 0 0.14fF $ **FLOATING
C4351 CLK1.n414 0 0.03fF $ **FLOATING
C4352 CLK1.n415 0 0.02fF $ **FLOATING
C4353 CLK1.t63 0 0.05fF
C4354 CLK1.n416 0 0.29fF $ **FLOATING
C4355 CLK1.n417 0 0.02fF $ **FLOATING
C4356 CLK1.n418 0 0.03fF $ **FLOATING
C4357 CLK1.n419 0 0.09fF $ **FLOATING
C4358 CLK1.n420 0 0.03fF $ **FLOATING
C4359 CLK1.n421 0 0.02fF $ **FLOATING
C4360 CLK1.t115 0 0.03fF
C4361 CLK1.t61 0 0.03fF
C4362 CLK1.n422 0 0.10fF $ **FLOATING
C4363 CLK1.n423 0 0.03fF $ **FLOATING
C4364 CLK1.n424 0 0.02fF $ **FLOATING
C4365 CLK1.n425 0 0.03fF $ **FLOATING
C4366 CLK1.t116 0 0.09fF
C4367 CLK1.n426 0 0.03fF $ **FLOATING
C4368 CLK1.n427 0 0.02fF $ **FLOATING
C4369 CLK1.t117 0 0.05fF
C4370 CLK1.n428 0 0.03fF $ **FLOATING
C4371 CLK1.n429 0 0.02fF $ **FLOATING
C4372 CLK1.n430 0 0.03fF $ **FLOATING
C4373 CLK1.n431 0 0.07fF $ **FLOATING
C4374 CLK1.n432 0 0.03fF $ **FLOATING
C4375 CLK1.n433 0 0.02fF $ **FLOATING
C4376 CLK1.t40 0 0.07fF
C4377 CLK1.n434 0 0.15fF $ **FLOATING
C4378 CLK1.n435 0 0.47fF $ **FLOATING
C4379 CLK1.n436 0 0.03fF $ **FLOATING
C4380 CLK1.n437 0 0.03fF $ **FLOATING
C4381 CLK1.n438 0 0.02fF $ **FLOATING
C4382 CLK1.n439 0 0.03fF $ **FLOATING
C4383 CLK1.n440 0 0.06fF $ **FLOATING
C4384 CLK1.n441 0 0.14fF $ **FLOATING
C4385 CLK1.n442 0 0.11fF $ **FLOATING
C4386 CLK1.n443 0 0.18fF $ **FLOATING
C4387 CLK1.n444 0 0.03fF $ **FLOATING
C4388 CLK1.n445 0 0.02fF $ **FLOATING
C4389 CLK1.n446 0 0.02fF $ **FLOATING
C4390 CLK1.n447 0 0.29fF $ **FLOATING
C4391 CLK1.n448 0 0.03fF $ **FLOATING
C4392 CLK1.n449 0 0.03fF $ **FLOATING
C4393 CLK1.n450 0 0.02fF $ **FLOATING
C4394 CLK1.n451 0 0.03fF $ **FLOATING
C4395 CLK1.n452 0 0.16fF $ **FLOATING
C4396 CLK1.n453 0 0.09fF $ **FLOATING
C4397 CLK1.t114 0 0.09fF
C4398 CLK1.t60 0 0.09fF
C4399 CLK1.n454 0 0.17fF $ **FLOATING
C4400 CLK1.n455 0 0.03fF $ **FLOATING
C4401 CLK1.n456 0 0.02fF $ **FLOATING
C4402 CLK1.n457 0 0.17fF $ **FLOATING
C4403 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_INV4_0/CLK 0 0.02fF $ **FLOATING
C4404 CLK1.n458 0 0.03fF $ **FLOATING
C4405 CLK1.n459 0 0.03fF $ **FLOATING
C4406 CLK1.n460 0 0.03fF $ **FLOATING
C4407 CLK1.n461 0 0.02fF $ **FLOATING
C4408 CLK1.n462 0 0.03fF $ **FLOATING
C4409 CLK1.n463 0 0.16fF $ **FLOATING
C4410 CLK1.t62 0 0.09fF
C4411 CLK1.n464 0 0.11fF $ **FLOATING
C4412 CLK1.n465 0 0.18fF $ **FLOATING
C4413 CLK1.n466 0 0.03fF $ **FLOATING
C4414 CLK1.n467 0 0.02fF $ **FLOATING
C4415 CLK1.n468 0 0.02fF $ **FLOATING
C4416 CLK1.n469 0 0.03fF $ **FLOATING
C4417 CLK1.n470 0 0.03fF $ **FLOATING
C4418 CLK1.n471 0 0.03fF $ **FLOATING
C4419 CLK1.n472 0 0.02fF $ **FLOATING
C4420 CLK1.n473 0 0.03fF $ **FLOATING
C4421 CLK1.n474 0 0.06fF $ **FLOATING
C4422 CLK1.n475 0 0.07fF $ **FLOATING
C4423 CLK1.n476 0 0.15fF $ **FLOATING
C4424 CLK1.n477 0 0.10fF $ **FLOATING
C4425 CLK1.n478 0 0.21fF $ **FLOATING
C4426 CLK1.n479 0 0.12fF $ **FLOATING
C4427 CLK1.n480 0 0.03fF $ **FLOATING
C4428 CLK1.n481 0 0.03fF $ **FLOATING
C4429 CLK1.n482 0 0.02fF $ **FLOATING
C4430 CLK1.n483 0 0.03fF $ **FLOATING
C4431 CLK1.n484 0 0.06fF $ **FLOATING
C4432 CLK1.n485 0 0.06fF $ **FLOATING
C4433 CLK1.n486 0 0.06fF $ **FLOATING
C4434 CLK1.n487 0 0.03fF $ **FLOATING
C4435 CLK1.n488 0 0.02fF $ **FLOATING
C4436 CLK1.n489 0 0.02fF $ **FLOATING
C4437 CLK1.n490 0 0.02fF $ **FLOATING
C4438 CLK1.n491 0 0.03fF $ **FLOATING
C4439 CLK1.t123 0 0.09fF
C4440 CLK1.n492 0 0.03fF $ **FLOATING
C4441 CLK1.n493 0 0.02fF $ **FLOATING
C4442 CLK1.t124 0 0.05fF
C4443 CLK1.n494 0 0.29fF $ **FLOATING
C4444 CLK1.t65 0 0.03fF
C4445 CLK1.t44 0 0.03fF
C4446 CLK1.n495 0 0.10fF $ **FLOATING
C4447 CLK1.n496 0 0.17fF $ **FLOATING
C4448 CLK1.n497 0 0.02fF $ **FLOATING
C4449 CLK1.n498 0 0.03fF $ **FLOATING
C4450 CLK1.n499 0 0.16fF $ **FLOATING
C4451 CLK1.n500 0 0.16fF $ **FLOATING
C4452 CLK1.n501 0 0.03fF $ **FLOATING
C4453 CLK1.n502 0 0.02fF $ **FLOATING
C4454 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_0/CLK 0 0.02fF $ **FLOATING
C4455 CLK1.t170 0 0.05fF
C4456 CLK1.n503 0 0.29fF $ **FLOATING
C4457 CLK1.n504 0 0.02fF $ **FLOATING
C4458 CLK1.n505 0 0.03fF $ **FLOATING
C4459 CLK1.t169 0 0.09fF
C4460 CLK1.n506 0 0.06fF $ **FLOATING
C4461 CLK1.n507 0 0.03fF $ **FLOATING
C4462 CLK1.n508 0 0.02fF $ **FLOATING
C4463 CLK1.n509 0 0.02fF $ **FLOATING
C4464 CLK1.n510 0 0.03fF $ **FLOATING
C4465 CLK1.n511 0 0.02fF $ **FLOATING
C4466 CLK1.n512 0 0.03fF $ **FLOATING
C4467 CLK1.n513 0 0.06fF $ **FLOATING
C4468 CLK1.n514 0 0.03fF $ **FLOATING
C4469 CLK1.n515 0 0.02fF $ **FLOATING
C4470 CLK1.t166 0 0.03fF
C4471 CLK1.t97 0 0.03fF
C4472 CLK1.n516 0 0.15fF $ **FLOATING
C4473 CLK1.n517 0 0.03fF $ **FLOATING
C4474 CLK1.n518 0 0.02fF $ **FLOATING
C4475 CLK1.n519 0 0.03fF $ **FLOATING
C4476 CLK1.n520 0 0.00fF $ **FLOATING
C4477 EESPFAL_Sbox_0/EESPFAL_s3_0/CLK1 0 0.00fF $ **FLOATING
C4478 CLK1.n521 0 0.01fF $ **FLOATING
C4479 CLK1.t41 0 0.08fF
C4480 CLK1.n522 0 0.34fF $ **FLOATING
C4481 CLK1.n523 0 0.02fF $ **FLOATING
C4482 CLK1.n524 0 0.03fF $ **FLOATING
C4483 CLK1.n525 0 0.06fF $ **FLOATING
C4484 CLK1.n526 0 0.03fF $ **FLOATING
C4485 CLK1.n527 0 0.02fF $ **FLOATING
C4486 CLK1.t191 0 0.03fF
C4487 CLK1.t42 0 0.03fF
C4488 CLK1.n528 0 0.15fF $ **FLOATING
C4489 CLK1.n529 0 0.19fF $ **FLOATING
C4490 CLK1.n530 0 0.02fF $ **FLOATING
C4491 CLK1.n531 0 0.03fF $ **FLOATING
C4492 CLK1.n532 0 0.14fF $ **FLOATING
C4493 CLK1.n533 0 0.03fF $ **FLOATING
C4494 CLK1.n534 0 0.02fF $ **FLOATING
C4495 CLK1.t162 0 0.05fF
C4496 CLK1.n535 0 0.29fF $ **FLOATING
C4497 CLK1.n536 0 0.02fF $ **FLOATING
C4498 CLK1.n537 0 0.03fF $ **FLOATING
C4499 CLK1.n538 0 0.09fF $ **FLOATING
C4500 CLK1.n539 0 0.03fF $ **FLOATING
C4501 CLK1.n540 0 0.02fF $ **FLOATING
C4502 CLK1.t143 0 0.03fF
C4503 CLK1.t160 0 0.03fF
C4504 CLK1.n541 0 0.10fF $ **FLOATING
C4505 CLK1.n542 0 0.03fF $ **FLOATING
C4506 CLK1.n543 0 0.02fF $ **FLOATING
C4507 CLK1.n544 0 0.03fF $ **FLOATING
C4508 CLK1.t144 0 0.09fF
C4509 CLK1.n545 0 0.03fF $ **FLOATING
C4510 CLK1.n546 0 0.02fF $ **FLOATING
C4511 CLK1.t145 0 0.05fF
C4512 CLK1.n547 0 0.03fF $ **FLOATING
C4513 CLK1.n548 0 0.02fF $ **FLOATING
C4514 CLK1.n549 0 0.03fF $ **FLOATING
C4515 CLK1.n550 0 0.06fF $ **FLOATING
C4516 CLK1.n551 0 0.03fF $ **FLOATING
C4517 CLK1.n552 0 0.02fF $ **FLOATING
C4518 CLK1.n553 0 0.03fF $ **FLOATING
C4519 CLK1.n554 0 0.02fF $ **FLOATING
C4520 CLK1.n555 0 0.03fF $ **FLOATING
C4521 CLK1.n556 0 0.07fF $ **FLOATING
C4522 CLK1.n557 0 0.03fF $ **FLOATING
C4523 CLK1.n558 0 0.02fF $ **FLOATING
C4524 CLK1.t66 0 0.08fF
C4525 CLK1.n559 0 0.13fF $ **FLOATING
C4526 CLK1.n560 0 0.36fF $ **FLOATING
C4527 CLK1.n561 0 0.03fF $ **FLOATING
C4528 CLK1.n562 0 0.03fF $ **FLOATING
C4529 CLK1.n563 0 0.02fF $ **FLOATING
C4530 CLK1.n564 0 0.03fF $ **FLOATING
C4531 CLK1.n565 0 0.06fF $ **FLOATING
C4532 CLK1.n566 0 0.06fF $ **FLOATING
C4533 CLK1.n567 0 0.06fF $ **FLOATING
C4534 CLK1.n568 0 0.03fF $ **FLOATING
C4535 CLK1.n569 0 0.02fF $ **FLOATING
C4536 CLK1.n570 0 0.03fF $ **FLOATING
C4537 CLK1.n571 0 0.03fF $ **FLOATING
C4538 CLK1.n572 0 0.03fF $ **FLOATING
C4539 CLK1.n573 0 0.02fF $ **FLOATING
C4540 CLK1.n574 0 0.03fF $ **FLOATING
C4541 CLK1.n575 0 0.06fF $ **FLOATING
C4542 CLK1.n576 0 0.14fF $ **FLOATING
C4543 CLK1.n577 0 0.11fF $ **FLOATING
C4544 CLK1.n578 0 0.18fF $ **FLOATING
C4545 CLK1.n579 0 0.03fF $ **FLOATING
C4546 CLK1.n580 0 0.02fF $ **FLOATING
C4547 CLK1.n581 0 0.02fF $ **FLOATING
C4548 CLK1.n582 0 0.29fF $ **FLOATING
C4549 CLK1.n583 0 0.03fF $ **FLOATING
C4550 CLK1.n584 0 0.03fF $ **FLOATING
C4551 CLK1.n585 0 0.02fF $ **FLOATING
C4552 CLK1.n586 0 0.03fF $ **FLOATING
C4553 CLK1.n587 0 0.16fF $ **FLOATING
C4554 CLK1.n588 0 0.09fF $ **FLOATING
C4555 CLK1.t142 0 0.09fF
C4556 CLK1.t159 0 0.09fF
C4557 CLK1.n589 0 0.17fF $ **FLOATING
C4558 CLK1.n590 0 0.03fF $ **FLOATING
C4559 CLK1.n591 0 0.02fF $ **FLOATING
C4560 CLK1.n592 0 0.17fF $ **FLOATING
C4561 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/CLK 0 0.02fF $ **FLOATING
C4562 CLK1.n593 0 0.03fF $ **FLOATING
C4563 CLK1.n594 0 0.03fF $ **FLOATING
C4564 CLK1.n595 0 0.03fF $ **FLOATING
C4565 CLK1.n596 0 0.02fF $ **FLOATING
C4566 CLK1.n597 0 0.03fF $ **FLOATING
C4567 CLK1.n598 0 0.16fF $ **FLOATING
C4568 CLK1.t161 0 0.09fF
C4569 CLK1.n599 0 0.11fF $ **FLOATING
C4570 CLK1.n600 0 0.18fF $ **FLOATING
C4571 CLK1.n601 0 0.03fF $ **FLOATING
C4572 CLK1.n602 0 0.02fF $ **FLOATING
C4573 CLK1.n603 0 0.02fF $ **FLOATING
C4574 CLK1.n604 0 0.03fF $ **FLOATING
C4575 CLK1.n605 0 0.03fF $ **FLOATING
C4576 CLK1.n606 0 0.03fF $ **FLOATING
C4577 CLK1.n607 0 0.02fF $ **FLOATING
C4578 CLK1.n608 0 0.03fF $ **FLOATING
C4579 CLK1.n609 0 0.06fF $ **FLOATING
C4580 CLK1.n610 0 0.06fF $ **FLOATING
C4581 CLK1.n611 0 0.06fF $ **FLOATING
C4582 CLK1.n612 0 0.03fF $ **FLOATING
C4583 CLK1.n613 0 0.02fF $ **FLOATING
C4584 CLK1.n614 0 0.02fF $ **FLOATING
C4585 CLK1.n615 0 0.03fF $ **FLOATING
C4586 CLK1.n616 0 0.03fF $ **FLOATING
C4587 CLK1.n617 0 0.03fF $ **FLOATING
C4588 CLK1.n618 0 0.02fF $ **FLOATING
C4589 CLK1.n619 0 0.03fF $ **FLOATING
C4590 CLK1.n620 0 0.06fF $ **FLOATING
C4591 CLK1.n621 0 0.07fF $ **FLOATING
C4592 CLK1.n622 0 0.13fF $ **FLOATING
C4593 CLK1.n623 0 0.08fF $ **FLOATING
C4594 CLK1.n624 0 0.13fF $ **FLOATING
C4595 CLK1.n625 0 0.02fF $ **FLOATING
C4596 CLK1.n626 0 0.01fF $ **FLOATING
C4597 CLK1.n627 0 0.03fF $ **FLOATING
C4598 CLK1.n628 0 0.06fF $ **FLOATING
C4599 CLK1.n629 0 0.03fF $ **FLOATING
C4600 CLK1.n630 0 0.02fF $ **FLOATING
C4601 CLK1.n631 0 0.02fF $ **FLOATING
C4602 CLK1.t112 0 0.03fF
C4603 CLK1.t118 0 0.03fF
C4604 CLK1.n632 0 0.15fF $ **FLOATING
C4605 CLK1.n633 0 0.03fF $ **FLOATING
C4606 CLK1.n634 0 0.02fF $ **FLOATING
C4607 CLK1.n635 0 0.03fF $ **FLOATING
C4608 CLK1.n636 0 0.06fF $ **FLOATING
C4609 CLK1.n637 0 0.03fF $ **FLOATING
C4610 CLK1.n638 0 0.02fF $ **FLOATING
C4611 CLK1.n639 0 0.02fF $ **FLOATING
C4612 CLK1.n640 0 0.02fF $ **FLOATING
C4613 CLK1.n641 0 0.03fF $ **FLOATING
C4614 CLK1.t185 0 0.09fF
C4615 CLK1.n642 0 0.03fF $ **FLOATING
C4616 CLK1.n643 0 0.02fF $ **FLOATING
C4617 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/CLK 0 0.02fF $ **FLOATING
C4618 CLK1.n644 0 0.02fF $ **FLOATING
C4619 CLK1.n645 0 0.03fF $ **FLOATING
C4620 CLK1.n646 0 0.16fF $ **FLOATING
C4621 CLK1.n647 0 0.03fF $ **FLOATING
C4622 CLK1.n648 0 0.02fF $ **FLOATING
C4623 CLK1.t13 0 0.05fF
C4624 CLK1.n649 0 0.29fF $ **FLOATING
C4625 CLK1.n650 0 0.02fF $ **FLOATING
C4626 CLK1.n651 0 0.03fF $ **FLOATING
C4627 CLK1.n652 0 0.06fF $ **FLOATING
C4628 CLK1.n653 0 0.03fF $ **FLOATING
C4629 CLK1.n654 0 0.02fF $ **FLOATING
C4630 CLK1.n655 0 0.03fF $ **FLOATING
C4631 CLK1.n656 0 0.02fF $ **FLOATING
C4632 CLK1.n657 0 0.03fF $ **FLOATING
C4633 CLK1.n658 0 0.06fF $ **FLOATING
C4634 CLK1.n659 0 0.03fF $ **FLOATING
C4635 CLK1.n660 0 0.02fF $ **FLOATING
C4636 CLK1.t151 0 0.03fF
C4637 CLK1.t82 0 0.03fF
C4638 CLK1.n661 0 0.15fF $ **FLOATING
C4639 CLK1.n662 0 0.03fF $ **FLOATING
C4640 CLK1.n663 0 0.02fF $ **FLOATING
C4641 CLK1.n664 0 0.03fF $ **FLOATING
C4642 CLK1.t197 0 0.07fF
C4643 CLK1.n665 0 0.45fF $ **FLOATING
C4644 CLK1.n666 0 0.02fF $ **FLOATING
C4645 CLK1.n667 0 0.03fF $ **FLOATING
C4646 CLK1.n668 0 0.14fF $ **FLOATING
C4647 CLK1.n669 0 0.03fF $ **FLOATING
C4648 CLK1.n670 0 0.02fF $ **FLOATING
C4649 CLK1.t74 0 0.05fF
C4650 CLK1.n671 0 0.29fF $ **FLOATING
C4651 CLK1.n672 0 0.02fF $ **FLOATING
C4652 CLK1.n673 0 0.03fF $ **FLOATING
C4653 CLK1.n674 0 0.09fF $ **FLOATING
C4654 CLK1.n675 0 0.03fF $ **FLOATING
C4655 CLK1.n676 0 0.02fF $ **FLOATING
C4656 CLK1.t68 0 0.03fF
C4657 CLK1.t72 0 0.03fF
C4658 CLK1.n677 0 0.10fF $ **FLOATING
C4659 CLK1.n678 0 0.03fF $ **FLOATING
C4660 CLK1.n679 0 0.02fF $ **FLOATING
C4661 CLK1.n680 0 0.03fF $ **FLOATING
C4662 CLK1.t69 0 0.09fF
C4663 CLK1.n681 0 0.03fF $ **FLOATING
C4664 CLK1.n682 0 0.02fF $ **FLOATING
C4665 CLK1.t70 0 0.05fF
C4666 CLK1.n683 0 0.03fF $ **FLOATING
C4667 CLK1.n684 0 0.02fF $ **FLOATING
C4668 CLK1.n685 0 0.03fF $ **FLOATING
C4669 CLK1.n686 0 0.07fF $ **FLOATING
C4670 CLK1.n687 0 0.03fF $ **FLOATING
C4671 CLK1.n688 0 0.02fF $ **FLOATING
C4672 CLK1.t31 0 0.07fF
C4673 CLK1.n689 0 0.15fF $ **FLOATING
C4674 CLK1.n690 0 0.47fF $ **FLOATING
C4675 CLK1.n691 0 0.03fF $ **FLOATING
C4676 CLK1.n692 0 0.03fF $ **FLOATING
C4677 CLK1.n693 0 0.02fF $ **FLOATING
C4678 CLK1.n694 0 0.03fF $ **FLOATING
C4679 CLK1.n695 0 0.06fF $ **FLOATING
C4680 CLK1.n696 0 0.14fF $ **FLOATING
C4681 CLK1.n697 0 0.11fF $ **FLOATING
C4682 CLK1.n698 0 0.18fF $ **FLOATING
C4683 CLK1.n699 0 0.03fF $ **FLOATING
C4684 CLK1.n700 0 0.02fF $ **FLOATING
C4685 CLK1.n701 0 0.02fF $ **FLOATING
C4686 CLK1.n702 0 0.29fF $ **FLOATING
C4687 CLK1.n703 0 0.03fF $ **FLOATING
C4688 CLK1.n704 0 0.03fF $ **FLOATING
C4689 CLK1.n705 0 0.02fF $ **FLOATING
C4690 CLK1.n706 0 0.03fF $ **FLOATING
C4691 CLK1.n707 0 0.16fF $ **FLOATING
C4692 CLK1.n708 0 0.09fF $ **FLOATING
C4693 CLK1.t67 0 0.09fF
C4694 CLK1.t71 0 0.09fF
C4695 CLK1.n709 0 0.17fF $ **FLOATING
C4696 CLK1.n710 0 0.03fF $ **FLOATING
C4697 CLK1.n711 0 0.02fF $ **FLOATING
C4698 CLK1.n712 0 0.17fF $ **FLOATING
C4699 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_1/CLK 0 0.02fF $ **FLOATING
C4700 CLK1.n713 0 0.03fF $ **FLOATING
C4701 CLK1.n714 0 0.03fF $ **FLOATING
C4702 CLK1.n715 0 0.03fF $ **FLOATING
C4703 CLK1.n716 0 0.02fF $ **FLOATING
C4704 CLK1.n717 0 0.03fF $ **FLOATING
C4705 CLK1.n718 0 0.16fF $ **FLOATING
C4706 CLK1.t73 0 0.09fF
C4707 CLK1.n719 0 0.11fF $ **FLOATING
C4708 CLK1.n720 0 0.18fF $ **FLOATING
C4709 CLK1.n721 0 0.03fF $ **FLOATING
C4710 CLK1.n722 0 0.02fF $ **FLOATING
C4711 CLK1.n723 0 0.02fF $ **FLOATING
C4712 CLK1.n724 0 0.03fF $ **FLOATING
C4713 CLK1.n725 0 0.03fF $ **FLOATING
C4714 CLK1.n726 0 0.03fF $ **FLOATING
C4715 CLK1.n727 0 0.02fF $ **FLOATING
C4716 CLK1.n728 0 0.03fF $ **FLOATING
C4717 CLK1.n729 0 0.06fF $ **FLOATING
C4718 CLK1.n730 0 0.07fF $ **FLOATING
C4719 CLK1.n731 0 0.15fF $ **FLOATING
C4720 CLK1.n732 0 0.10fF $ **FLOATING
C4721 CLK1.n733 0 0.11fF $ **FLOATING
C4722 CLK1.n734 0 0.21fF $ **FLOATING
C4723 CLK1.n735 0 0.08fF $ **FLOATING
C4724 CLK1.n736 0 0.06fF $ **FLOATING
C4725 CLK1.n737 0 0.03fF $ **FLOATING
C4726 CLK1.n738 0 0.02fF $ **FLOATING
C4727 CLK1.n739 0 0.03fF $ **FLOATING
C4728 CLK1.n740 0 0.02fF $ **FLOATING
C4729 CLK1.n741 0 0.19fF $ **FLOATING
C4730 CLK1.n742 0 0.03fF $ **FLOATING
C4731 CLK1.n743 0 0.02fF $ **FLOATING
C4732 CLK1.n744 0 0.03fF $ **FLOATING
C4733 CLK1.n745 0 0.06fF $ **FLOATING
C4734 CLK1.n746 0 0.06fF $ **FLOATING
C4735 CLK1.n747 0 0.06fF $ **FLOATING
C4736 CLK1.n748 0 0.03fF $ **FLOATING
C4737 CLK1.n749 0 0.02fF $ **FLOATING
C4738 CLK1.n750 0 0.03fF $ **FLOATING
C4739 CLK1.n751 0 0.03fF $ **FLOATING
C4740 CLK1.n752 0 0.02fF $ **FLOATING
C4741 CLK1.n753 0 0.03fF $ **FLOATING
C4742 CLK1.n754 0 0.02fF $ **FLOATING
C4743 CLK1.n755 0 0.03fF $ **FLOATING
C4744 CLK1.n756 0 0.14fF $ **FLOATING
C4745 CLK1.n757 0 0.18fF $ **FLOATING
C4746 CLK1.t12 0 0.09fF
C4747 CLK1.n758 0 0.11fF $ **FLOATING
C4748 CLK1.n759 0 0.03fF $ **FLOATING
C4749 CLK1.n760 0 0.02fF $ **FLOATING
C4750 CLK1.n761 0 0.03fF $ **FLOATING
C4751 CLK1.n762 0 0.03fF $ **FLOATING
C4752 CLK1.t47 0 0.03fF
C4753 CLK1.t184 0 0.03fF
C4754 CLK1.n763 0 0.10fF $ **FLOATING
C4755 CLK1.n764 0 0.17fF $ **FLOATING
C4756 CLK1.n765 0 0.03fF $ **FLOATING
C4757 CLK1.n766 0 0.02fF $ **FLOATING
C4758 CLK1.n767 0 0.03fF $ **FLOATING
C4759 CLK1.n768 0 0.09fF $ **FLOATING
C4760 CLK1.t46 0 0.09fF
C4761 CLK1.n769 0 0.17fF $ **FLOATING
C4762 CLK1.t183 0 0.09fF
C4763 CLK1.n770 0 0.16fF $ **FLOATING
C4764 CLK1.n771 0 0.09fF $ **FLOATING
C4765 CLK1.n772 0 0.03fF $ **FLOATING
C4766 CLK1.n773 0 0.02fF $ **FLOATING
C4767 CLK1.n774 0 0.03fF $ **FLOATING
C4768 CLK1.n775 0 0.03fF $ **FLOATING
C4769 CLK1.t186 0 0.05fF
C4770 CLK1.n776 0 0.29fF $ **FLOATING
C4771 CLK1.n777 0 0.03fF $ **FLOATING
C4772 CLK1.n778 0 0.02fF $ **FLOATING
C4773 CLK1.n779 0 0.03fF $ **FLOATING
C4774 CLK1.n780 0 0.11fF $ **FLOATING
C4775 CLK1.n781 0 0.18fF $ **FLOATING
C4776 CLK1.n782 0 0.14fF $ **FLOATING
C4777 CLK1.n783 0 0.03fF $ **FLOATING
C4778 CLK1.n784 0 0.02fF $ **FLOATING
C4779 CLK1.n785 0 0.03fF $ **FLOATING
C4780 CLK1.n786 0 0.03fF $ **FLOATING
C4781 CLK1.n787 0 0.03fF $ **FLOATING
C4782 CLK1.n788 0 0.02fF $ **FLOATING
C4783 CLK1.n789 0 0.03fF $ **FLOATING
C4784 CLK1.n790 0 0.06fF $ **FLOATING
C4785 CLK1.n791 0 0.06fF $ **FLOATING
C4786 CLK1.n792 0 0.06fF $ **FLOATING
C4787 CLK1.n793 0 0.03fF $ **FLOATING
C4788 CLK1.n794 0 0.02fF $ **FLOATING
C4789 CLK1.n795 0 0.03fF $ **FLOATING
C4790 CLK1.n796 0 0.19fF $ **FLOATING
C4791 CLK1.n797 0 0.02fF $ **FLOATING
C4792 CLK1.n798 0 0.03fF $ **FLOATING
C4793 CLK1.n799 0 0.03fF $ **FLOATING
C4794 CLK1.n800 0 0.02fF $ **FLOATING
C4795 CLK1.n801 0 0.03fF $ **FLOATING
C4796 CLK1.n802 0 0.06fF $ **FLOATING
C4797 CLK1.n803 0 0.08fF $ **FLOATING
C4798 CLK1.n804 0 0.19fF $ **FLOATING
C4799 CLK1.n805 0 0.01fF $ **FLOATING
C4800 CLK1.n806 0 0.00fF $ **FLOATING
C4801 CLK1.n807 0 0.03fF $ **FLOATING
C4802 CLK1.n808 0 0.36fF $ **FLOATING
C4803 CLK1.n809 0 0.36fF $ **FLOATING
C4804 CLK1.n810 0 0.02fF $ **FLOATING
C4805 CLK1.n811 0 0.01fF $ **FLOATING
C4806 CLK1.n812 0 0.03fF $ **FLOATING
C4807 CLK1.n813 0 0.06fF $ **FLOATING
C4808 CLK1.n814 0 0.03fF $ **FLOATING
C4809 CLK1.n815 0 0.02fF $ **FLOATING
C4810 CLK1.n816 0 0.02fF $ **FLOATING
C4811 CLK1.t34 0 0.03fF
C4812 CLK1.t39 0 0.03fF
C4813 CLK1.n817 0 0.15fF $ **FLOATING
C4814 CLK1.n818 0 0.03fF $ **FLOATING
C4815 CLK1.n819 0 0.02fF $ **FLOATING
C4816 CLK1.n820 0 0.03fF $ **FLOATING
C4817 CLK1.n821 0 0.06fF $ **FLOATING
C4818 CLK1.n822 0 0.03fF $ **FLOATING
C4819 CLK1.n823 0 0.02fF $ **FLOATING
C4820 CLK1.n824 0 0.02fF $ **FLOATING
C4821 CLK1.n825 0 0.02fF $ **FLOATING
C4822 CLK1.n826 0 0.03fF $ **FLOATING
C4823 CLK1.t57 0 0.09fF
C4824 CLK1.n827 0 0.03fF $ **FLOATING
C4825 CLK1.n828 0 0.02fF $ **FLOATING
C4826 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/CLK 0 0.02fF $ **FLOATING
C4827 CLK1.n829 0 0.02fF $ **FLOATING
C4828 CLK1.n830 0 0.03fF $ **FLOATING
C4829 CLK1.n831 0 0.16fF $ **FLOATING
C4830 CLK1.n832 0 0.03fF $ **FLOATING
C4831 CLK1.n833 0 0.02fF $ **FLOATING
C4832 CLK1.t134 0 0.05fF
C4833 CLK1.n834 0 0.29fF $ **FLOATING
C4834 CLK1.n835 0 0.02fF $ **FLOATING
C4835 CLK1.n836 0 0.03fF $ **FLOATING
C4836 CLK1.n837 0 0.06fF $ **FLOATING
C4837 CLK1.n838 0 0.03fF $ **FLOATING
C4838 CLK1.n839 0 0.02fF $ **FLOATING
C4839 CLK1.n840 0 0.03fF $ **FLOATING
C4840 CLK1.n841 0 0.02fF $ **FLOATING
C4841 CLK1.n842 0 0.03fF $ **FLOATING
C4842 CLK1.n843 0 0.06fF $ **FLOATING
C4843 CLK1.n844 0 0.03fF $ **FLOATING
C4844 CLK1.n845 0 0.02fF $ **FLOATING
C4845 CLK1.t91 0 0.03fF
C4846 CLK1.t35 0 0.03fF
C4847 CLK1.n846 0 0.15fF $ **FLOATING
C4848 CLK1.n847 0 0.03fF $ **FLOATING
C4849 CLK1.n848 0 0.02fF $ **FLOATING
C4850 CLK1.n849 0 0.03fF $ **FLOATING
C4851 CLK1.t168 0 0.07fF
C4852 CLK1.n850 0 0.45fF $ **FLOATING
C4853 CLK1.n851 0 0.02fF $ **FLOATING
C4854 CLK1.n852 0 0.03fF $ **FLOATING
C4855 CLK1.n853 0 0.14fF $ **FLOATING
C4856 CLK1.n854 0 0.03fF $ **FLOATING
C4857 CLK1.n855 0 0.02fF $ **FLOATING
C4858 CLK1.t5 0 0.05fF
C4859 CLK1.n856 0 0.29fF $ **FLOATING
C4860 CLK1.n857 0 0.02fF $ **FLOATING
C4861 CLK1.n858 0 0.03fF $ **FLOATING
C4862 CLK1.n859 0 0.09fF $ **FLOATING
C4863 CLK1.n860 0 0.03fF $ **FLOATING
C4864 CLK1.n861 0 0.02fF $ **FLOATING
C4865 CLK1.t158 0 0.03fF
C4866 CLK1.t7 0 0.03fF
C4867 CLK1.n862 0 0.10fF $ **FLOATING
C4868 CLK1.n863 0 0.03fF $ **FLOATING
C4869 CLK1.n864 0 0.02fF $ **FLOATING
C4870 CLK1.n865 0 0.03fF $ **FLOATING
C4871 CLK1.t155 0 0.09fF
C4872 CLK1.n866 0 0.03fF $ **FLOATING
C4873 CLK1.n867 0 0.02fF $ **FLOATING
C4874 CLK1.t156 0 0.05fF
C4875 CLK1.n868 0 0.03fF $ **FLOATING
C4876 CLK1.n869 0 0.02fF $ **FLOATING
C4877 CLK1.n870 0 0.03fF $ **FLOATING
C4878 CLK1.n871 0 0.07fF $ **FLOATING
C4879 CLK1.n872 0 0.03fF $ **FLOATING
C4880 CLK1.n873 0 0.02fF $ **FLOATING
C4881 CLK1.t101 0 0.07fF
C4882 CLK1.n874 0 0.15fF $ **FLOATING
C4883 CLK1.n875 0 0.47fF $ **FLOATING
C4884 CLK1.n876 0 0.03fF $ **FLOATING
C4885 CLK1.n877 0 0.03fF $ **FLOATING
C4886 CLK1.n878 0 0.02fF $ **FLOATING
C4887 CLK1.n879 0 0.03fF $ **FLOATING
C4888 CLK1.n880 0 0.06fF $ **FLOATING
C4889 CLK1.n881 0 0.14fF $ **FLOATING
C4890 CLK1.n882 0 0.11fF $ **FLOATING
C4891 CLK1.n883 0 0.18fF $ **FLOATING
C4892 CLK1.n884 0 0.03fF $ **FLOATING
C4893 CLK1.n885 0 0.02fF $ **FLOATING
C4894 CLK1.n886 0 0.02fF $ **FLOATING
C4895 CLK1.n887 0 0.29fF $ **FLOATING
C4896 CLK1.n888 0 0.03fF $ **FLOATING
C4897 CLK1.n889 0 0.03fF $ **FLOATING
C4898 CLK1.n890 0 0.02fF $ **FLOATING
C4899 CLK1.n891 0 0.03fF $ **FLOATING
C4900 CLK1.n892 0 0.16fF $ **FLOATING
C4901 CLK1.n893 0 0.09fF $ **FLOATING
C4902 CLK1.t157 0 0.09fF
C4903 CLK1.t6 0 0.09fF
C4904 CLK1.n894 0 0.17fF $ **FLOATING
C4905 CLK1.n895 0 0.03fF $ **FLOATING
C4906 CLK1.n896 0 0.02fF $ **FLOATING
C4907 CLK1.n897 0 0.17fF $ **FLOATING
C4908 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_INV4_0/CLK 0 0.02fF $ **FLOATING
C4909 CLK1.n898 0 0.03fF $ **FLOATING
C4910 CLK1.n899 0 0.03fF $ **FLOATING
C4911 CLK1.n900 0 0.03fF $ **FLOATING
C4912 CLK1.n901 0 0.02fF $ **FLOATING
C4913 CLK1.n902 0 0.03fF $ **FLOATING
C4914 CLK1.n903 0 0.16fF $ **FLOATING
C4915 CLK1.t4 0 0.09fF
C4916 CLK1.n904 0 0.11fF $ **FLOATING
C4917 CLK1.n905 0 0.18fF $ **FLOATING
C4918 CLK1.n906 0 0.03fF $ **FLOATING
C4919 CLK1.n907 0 0.02fF $ **FLOATING
C4920 CLK1.n908 0 0.02fF $ **FLOATING
C4921 CLK1.n909 0 0.03fF $ **FLOATING
C4922 CLK1.n910 0 0.03fF $ **FLOATING
C4923 CLK1.n911 0 0.03fF $ **FLOATING
C4924 CLK1.n912 0 0.02fF $ **FLOATING
C4925 CLK1.n913 0 0.03fF $ **FLOATING
C4926 CLK1.n914 0 0.06fF $ **FLOATING
C4927 CLK1.n915 0 0.07fF $ **FLOATING
C4928 CLK1.n916 0 0.15fF $ **FLOATING
C4929 CLK1.n917 0 0.10fF $ **FLOATING
C4930 CLK1.n918 0 0.11fF $ **FLOATING
C4931 CLK1.n919 0 0.21fF $ **FLOATING
C4932 CLK1.n920 0 0.08fF $ **FLOATING
C4933 CLK1.n921 0 0.06fF $ **FLOATING
C4934 CLK1.n922 0 0.03fF $ **FLOATING
C4935 CLK1.n923 0 0.02fF $ **FLOATING
C4936 CLK1.n924 0 0.03fF $ **FLOATING
C4937 CLK1.n925 0 0.02fF $ **FLOATING
C4938 CLK1.n926 0 0.19fF $ **FLOATING
C4939 CLK1.n927 0 0.03fF $ **FLOATING
C4940 CLK1.n928 0 0.02fF $ **FLOATING
C4941 CLK1.n929 0 0.03fF $ **FLOATING
C4942 CLK1.n930 0 0.06fF $ **FLOATING
C4943 CLK1.n931 0 0.06fF $ **FLOATING
C4944 CLK1.n932 0 0.06fF $ **FLOATING
C4945 CLK1.n933 0 0.03fF $ **FLOATING
C4946 CLK1.n934 0 0.02fF $ **FLOATING
C4947 CLK1.n935 0 0.03fF $ **FLOATING
C4948 CLK1.n936 0 0.03fF $ **FLOATING
C4949 CLK1.n937 0 0.02fF $ **FLOATING
C4950 CLK1.n938 0 0.03fF $ **FLOATING
C4951 CLK1.n939 0 0.02fF $ **FLOATING
C4952 CLK1.n940 0 0.03fF $ **FLOATING
C4953 CLK1.n941 0 0.14fF $ **FLOATING
C4954 CLK1.n942 0 0.18fF $ **FLOATING
C4955 CLK1.t133 0 0.09fF
C4956 CLK1.n943 0 0.11fF $ **FLOATING
C4957 CLK1.n944 0 0.03fF $ **FLOATING
C4958 CLK1.n945 0 0.02fF $ **FLOATING
C4959 CLK1.n946 0 0.03fF $ **FLOATING
C4960 CLK1.n947 0 0.03fF $ **FLOATING
C4961 CLK1.t136 0 0.03fF
C4962 CLK1.t104 0 0.03fF
C4963 CLK1.n948 0 0.10fF $ **FLOATING
C4964 CLK1.n949 0 0.17fF $ **FLOATING
C4965 CLK1.n950 0 0.03fF $ **FLOATING
C4966 CLK1.n951 0 0.02fF $ **FLOATING
C4967 CLK1.n952 0 0.03fF $ **FLOATING
C4968 CLK1.n953 0 0.09fF $ **FLOATING
C4969 CLK1.t135 0 0.09fF
C4970 CLK1.n954 0 0.17fF $ **FLOATING
C4971 CLK1.t103 0 0.09fF
C4972 CLK1.n955 0 0.16fF $ **FLOATING
C4973 CLK1.n956 0 0.09fF $ **FLOATING
C4974 CLK1.n957 0 0.03fF $ **FLOATING
C4975 CLK1.n958 0 0.02fF $ **FLOATING
C4976 CLK1.n959 0 0.03fF $ **FLOATING
C4977 CLK1.n960 0 0.03fF $ **FLOATING
C4978 CLK1.t58 0 0.05fF
C4979 CLK1.n961 0 0.29fF $ **FLOATING
C4980 CLK1.n962 0 0.03fF $ **FLOATING
C4981 CLK1.n963 0 0.02fF $ **FLOATING
C4982 CLK1.n964 0 0.03fF $ **FLOATING
C4983 CLK1.n965 0 0.11fF $ **FLOATING
C4984 CLK1.n966 0 0.18fF $ **FLOATING
C4985 CLK1.n967 0 0.14fF $ **FLOATING
C4986 CLK1.n968 0 0.03fF $ **FLOATING
C4987 CLK1.n969 0 0.02fF $ **FLOATING
C4988 CLK1.n970 0 0.03fF $ **FLOATING
C4989 CLK1.n971 0 0.03fF $ **FLOATING
C4990 CLK1.n972 0 0.03fF $ **FLOATING
C4991 CLK1.n973 0 0.02fF $ **FLOATING
C4992 CLK1.n974 0 0.03fF $ **FLOATING
C4993 CLK1.n975 0 0.06fF $ **FLOATING
C4994 CLK1.n976 0 0.06fF $ **FLOATING
C4995 CLK1.n977 0 0.06fF $ **FLOATING
C4996 CLK1.n978 0 0.03fF $ **FLOATING
C4997 CLK1.n979 0 0.02fF $ **FLOATING
C4998 CLK1.n980 0 0.03fF $ **FLOATING
C4999 CLK1.n981 0 0.19fF $ **FLOATING
C5000 CLK1.n982 0 0.02fF $ **FLOATING
C5001 CLK1.n983 0 0.03fF $ **FLOATING
C5002 CLK1.n984 0 0.03fF $ **FLOATING
C5003 CLK1.n985 0 0.02fF $ **FLOATING
C5004 CLK1.n986 0 0.03fF $ **FLOATING
C5005 CLK1.n987 0 0.06fF $ **FLOATING
C5006 CLK1.n988 0 0.08fF $ **FLOATING
C5007 CLK1.n989 0 0.19fF $ **FLOATING
C5008 CLK1.n990 0 0.01fF $ **FLOATING
C5009 CLK1.n991 0 0.00fF $ **FLOATING
C5010 CLK1.n992 0 0.03fF $ **FLOATING
C5011 CLK1.n993 0 0.07fF $ **FLOATING
C5012 CLK1.n994 0 0.08fF $ **FLOATING
C5013 EESPFAL_Sbox_0/EESPFAL_s2_0/CLK1 0 0.02fF $ **FLOATING
C5014 CLK1.n995 0 0.01fF $ **FLOATING
C5015 CLK1.n996 0 0.04fF $ **FLOATING
C5016 CLK1.n997 0 0.21fF $ **FLOATING
C5017 CLK1.n998 0 0.08fF $ **FLOATING
C5018 CLK1.n999 0 0.06fF $ **FLOATING
C5019 CLK1.n1000 0 0.03fF $ **FLOATING
C5020 CLK1.n1001 0 0.02fF $ **FLOATING
C5021 CLK1.n1002 0 0.03fF $ **FLOATING
C5022 CLK1.n1003 0 0.02fF $ **FLOATING
C5023 CLK1.n1004 0 0.19fF $ **FLOATING
C5024 CLK1.n1005 0 0.03fF $ **FLOATING
C5025 CLK1.n1006 0 0.02fF $ **FLOATING
C5026 CLK1.n1007 0 0.03fF $ **FLOATING
C5027 CLK1.n1008 0 0.06fF $ **FLOATING
C5028 CLK1.n1009 0 0.06fF $ **FLOATING
C5029 CLK1.n1010 0 0.06fF $ **FLOATING
C5030 CLK1.n1011 0 0.03fF $ **FLOATING
C5031 CLK1.n1012 0 0.02fF $ **FLOATING
C5032 CLK1.n1013 0 0.03fF $ **FLOATING
C5033 CLK1.n1014 0 0.03fF $ **FLOATING
C5034 CLK1.n1015 0 0.03fF $ **FLOATING
C5035 CLK1.n1016 0 0.02fF $ **FLOATING
C5036 CLK1.n1017 0 0.03fF $ **FLOATING
C5037 CLK1.n1018 0 0.14fF $ **FLOATING
C5038 CLK1.n1019 0 0.18fF $ **FLOATING
C5039 CLK1.n1020 0 0.11fF $ **FLOATING
C5040 CLK1.n1021 0 0.03fF $ **FLOATING
C5041 CLK1.n1022 0 0.02fF $ **FLOATING
C5042 CLK1.n1023 0 0.03fF $ **FLOATING
C5043 CLK1.n1024 0 0.03fF $ **FLOATING
C5044 CLK1.n1025 0 0.03fF $ **FLOATING
C5045 CLK1.n1026 0 0.02fF $ **FLOATING
C5046 CLK1.n1027 0 0.03fF $ **FLOATING
C5047 CLK1.n1028 0 0.09fF $ **FLOATING
C5048 CLK1.t43 0 0.09fF
C5049 CLK1.n1029 0 0.17fF $ **FLOATING
C5050 CLK1.t64 0 0.09fF
C5051 CLK1.n1030 0 0.09fF $ **FLOATING
C5052 CLK1.n1031 0 0.03fF $ **FLOATING
C5053 CLK1.n1032 0 0.02fF $ **FLOATING
C5054 CLK1.n1033 0 0.03fF $ **FLOATING
C5055 CLK1.n1034 0 0.03fF $ **FLOATING
C5056 CLK1.n1035 0 0.03fF $ **FLOATING
C5057 CLK1.n1036 0 0.02fF $ **FLOATING
C5058 CLK1.n1037 0 0.03fF $ **FLOATING
C5059 CLK1.n1038 0 0.11fF $ **FLOATING
C5060 CLK1.n1039 0 0.18fF $ **FLOATING
C5061 CLK1.n1040 0 0.14fF $ **FLOATING
C5062 CLK1.n1041 0 0.03fF $ **FLOATING
C5063 CLK1.n1042 0 0.02fF $ **FLOATING
C5064 CLK1.n1043 0 0.03fF $ **FLOATING
C5065 CLK1.n1044 0 0.03fF $ **FLOATING
C5066 CLK1.n1045 0 0.03fF $ **FLOATING
C5067 CLK1.n1046 0 0.02fF $ **FLOATING
C5068 CLK1.n1047 0 0.03fF $ **FLOATING
C5069 CLK1.n1048 0 0.06fF $ **FLOATING
C5070 CLK1.n1049 0 0.06fF $ **FLOATING
C5071 CLK1.n1050 0 0.06fF $ **FLOATING
C5072 CLK1.n1051 0 0.03fF $ **FLOATING
C5073 CLK1.n1052 0 0.02fF $ **FLOATING
C5074 CLK1.n1053 0 0.03fF $ **FLOATING
C5075 CLK1.n1054 0 0.07fF $ **FLOATING
C5076 CLK1.n1055 0 0.09fF $ **FLOATING
C5077 CLK1.n1056 0 0.02fF $ **FLOATING
C5078 CLK1.t165 0 0.03fF
C5079 CLK1.n1057 0 0.07fF $ **FLOATING
C5080 CLK1.n1058 0 0.02fF $ **FLOATING
C5081 CLK1.n1059 0 0.08fF $ **FLOATING
C5082 CLK1.n1060 0 0.09fF $ **FLOATING
C5083 CLK1.t48 0 0.03fF
C5084 CLK1.t37 0 0.03fF
C5085 CLK1.n1061 0 0.07fF $ **FLOATING
C5086 CLK1.n1062 0 0.01fF $ **FLOATING
C5087 CLK1.n1063 0 0.02fF $ **FLOATING
C5088 CLK1.n1064 0 0.02fF $ **FLOATING
C5089 CLK1.n1065 0 0.08fF $ **FLOATING
C5090 CLK1.n1066 0 0.07fF $ **FLOATING
C5091 CLK1.n1067 0 0.07fF $ **FLOATING
C5092 CLK1.n1068 0 0.07fF $ **FLOATING
C5093 CLK1.n1069 0 0.10fF $ **FLOATING
C5094 CLK1.n1070 0 0.07fF $ **FLOATING
C5095 CLK1.n1071 0 0.07fF $ **FLOATING
C5096 CLK1.n1072 0 0.05fF $ **FLOATING
C5097 CLK1.n1073 0 0.07fF $ **FLOATING
C5098 CLK1.n1074 0 0.25fF $ **FLOATING
C5099 CLK1.n1075 0 0.34fF $ **FLOATING
C5100 CLK1.n1076 0 0.20fF $ **FLOATING
C5101 CLK1.n1077 0 0.07fF $ **FLOATING
C5102 CLK1.n1078 0 0.07fF $ **FLOATING
C5103 CLK1.t51 0 0.05fF
C5104 CLK1.t11 0 0.05fF
C5105 CLK1.n1079 0 0.60fF $ **FLOATING
C5106 CLK1.t52 0 0.03fF
C5107 CLK1.t120 0 0.03fF
C5108 CLK1.n1080 0 0.10fF $ **FLOATING
C5109 CLK1.t9 0 0.03fF
C5110 CLK1.t76 0 0.03fF
C5111 CLK1.n1081 0 0.10fF $ **FLOATING
C5112 CLK1.n1082 0 0.36fF $ **FLOATING
C5113 CLK1.n1083 0 0.07fF $ **FLOATING
C5114 CLK1.t10 0 0.17fF
C5115 CLK1.n1084 0 0.31fF $ **FLOATING
C5116 CLK1.n1085 0 0.18fF $ **FLOATING
C5117 CLK1.t8 0 0.17fF
C5118 CLK1.n1086 0 0.32fF $ **FLOATING
C5119 CLK1.t75 0 0.17fF
C5120 CLK1.n1087 0 0.18fF $ **FLOATING
C5121 CLK1.n1088 0 0.07fF $ **FLOATING
C5122 CLK1.n1089 0 0.07fF $ **FLOATING
C5123 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_XOR_v3_1/CLK 0 0.04fF $ **FLOATING
C5124 CLK1.t121 0 0.05fF
C5125 CLK1.t78 0 0.05fF
C5126 CLK1.n1090 0 0.60fF $ **FLOATING
C5127 CLK1.n1091 0 0.07fF $ **FLOATING
C5128 CLK1.n1092 0 0.31fF $ **FLOATING
C5129 CLK1.t77 0 0.17fF
C5130 CLK1.n1093 0 0.20fF $ **FLOATING
C5131 CLK1.n1094 0 0.34fF $ **FLOATING
C5132 CLK1.n1095 0 0.25fF $ **FLOATING
C5133 CLK1.n1096 0 0.07fF $ **FLOATING
C5134 CLK1.n1097 0 0.07fF $ **FLOATING
C5135 CLK1.n1098 0 0.05fF $ **FLOATING
C5136 CLK1.t163 0 0.03fF
C5137 CLK1.t190 0 0.03fF
C5138 CLK1.n1099 0 0.18fF $ **FLOATING
C5139 CLK1.n1100 0 0.23fF $ **FLOATING
C5140 CLK1.n1101 0 0.07fF $ **FLOATING
C5141 CLK1.n1102 0 0.07fF $ **FLOATING
C5142 CLK1.n1103 0 0.10fF $ **FLOATING
C5143 CLK1.n1104 0 0.10fF $ **FLOATING
C5144 CLK1.n1105 0 0.07fF $ **FLOATING
C5145 CLK1.n1106 0 0.07fF $ **FLOATING
C5146 CLK1.n1107 0 0.04fF $ **FLOATING
C5147 CLK1.t38 0 0.03fF
C5148 CLK1.t189 0 0.03fF
C5149 CLK1.n1108 0 0.15fF $ **FLOATING
C5150 CLK1.t24 0 0.03fF
C5151 CLK1.t45 0 0.03fF
C5152 CLK1.n1109 0 0.18fF $ **FLOATING
C5153 CLK1.n1110 0 0.23fF $ **FLOATING
C5154 CLK1.n1111 0 0.07fF $ **FLOATING
C5155 CLK1.n1112 0 0.07fF $ **FLOATING
C5156 CLK1.n1113 0 0.19fF $ **FLOATING
C5157 CLK1.n1114 0 0.29fF $ **FLOATING
C5158 CLK1.n1115 0 0.07fF $ **FLOATING
C5159 CLK1.n1116 0 0.07fF $ **FLOATING
C5160 CLK1.n1117 0 0.14fF $ **FLOATING
C5161 CLK1.n1118 0 0.10fF $ **FLOATING
C5162 CLK1.n1119 0 0.10fF $ **FLOATING
C5163 CLK1.n1120 0 0.07fF $ **FLOATING
C5164 CLK1.n1121 0 0.07fF $ **FLOATING
C5165 CLK1.n1122 0 0.06fF $ **FLOATING
C5166 CLK1.n1123 0 0.05fF $ **FLOATING
C5167 CLK1.n1124 0 0.21fF $ **FLOATING
C5168 CLK1.n1125 0 0.06fF $ **FLOATING
C5169 CLK1.n1126 0 0.07fF $ **FLOATING
C5170 CLK1.n1127 0 0.07fF $ **FLOATING
C5171 CLK1.n1128 0 0.10fF $ **FLOATING
C5172 CLK1.n1129 0 0.10fF $ **FLOATING
C5173 CLK1.n1130 0 0.10fF $ **FLOATING
C5174 CLK1.n1131 0 0.07fF $ **FLOATING
C5175 CLK1.n1132 0 0.07fF $ **FLOATING
C5176 CLK1.n1133 0 0.07fF $ **FLOATING
C5177 CLK1.n1134 0 0.07fF $ **FLOATING
C5178 CLK1.n1135 0 0.07fF $ **FLOATING
C5179 CLK1.n1136 0 0.07fF $ **FLOATING
C5180 CLK1.n1137 0 0.07fF $ **FLOATING
C5181 CLK1.n1138 0 0.07fF $ **FLOATING
C5182 CLK1.n1139 0 0.07fF $ **FLOATING
C5183 CLK1.n1140 0 0.07fF $ **FLOATING
C5184 CLK1.n1141 0 0.06fF $ **FLOATING
C5185 CLK1.n1142 0 0.07fF $ **FLOATING
C5186 CLK1.n1143 0 0.06fF $ **FLOATING
C5187 CLK1.n1144 0 0.07fF $ **FLOATING
C5188 CLK1.n1145 0 0.07fF $ **FLOATING
C5189 CLK1.n1146 0 0.07fF $ **FLOATING
C5190 CLK1.n1147 0 0.07fF $ **FLOATING
C5191 CLK1.n1148 0 0.07fF $ **FLOATING
C5192 CLK1.n1149 0 0.07fF $ **FLOATING
C5193 CLK1.n1150 0 0.07fF $ **FLOATING
C5194 CLK1.n1151 0 0.06fF $ **FLOATING
C5195 CLK1.n1152 0 0.07fF $ **FLOATING
C5196 CLK1.n1153 0 0.07fF $ **FLOATING
C5197 CLK1.n1154 0 0.07fF $ **FLOATING
C5198 CLK1.n1155 0 0.07fF $ **FLOATING
C5199 CLK1.n1156 0 0.07fF $ **FLOATING
C5200 CLK1.n1157 0 0.07fF $ **FLOATING
C5201 CLK1.n1158 0 0.07fF $ **FLOATING
C5202 CLK1.n1159 0 0.07fF $ **FLOATING
C5203 CLK1.n1160 0 0.07fF $ **FLOATING
C5204 CLK1.n1161 0 0.07fF $ **FLOATING
C5205 CLK1.n1162 0 0.10fF $ **FLOATING
C5206 CLK1.n1163 0 0.10fF $ **FLOATING
C5207 CLK1.n1164 0 0.10fF $ **FLOATING
C5208 CLK1.n1165 0 0.07fF $ **FLOATING
C5209 CLK1.n1166 0 0.07fF $ **FLOATING
C5210 CLK1.n1167 0 0.06fF $ **FLOATING
C5211 CLK1.n1168 0 0.09fF $ **FLOATING
C5212 CLK1.n1169 0 0.05fF $ **FLOATING
C5213 CLK1.n1170 0 0.07fF $ **FLOATING
C5214 CLK1.n1171 0 0.07fF $ **FLOATING
C5215 CLK1.n1172 0 0.07fF $ **FLOATING
C5216 CLK1.n1173 0 0.10fF $ **FLOATING
C5217 CLK1.n1174 0 0.10fF $ **FLOATING
C5218 CLK1.n1175 0 0.13fF $ **FLOATING
C5219 CLK1.n1176 0 0.07fF $ **FLOATING
C5220 CLK1.n1177 0 0.07fF $ **FLOATING
C5221 CLK1.n1178 0 0.06fF $ **FLOATING
C5222 CLK1.n1179 0 0.12fF $ **FLOATING
C5223 CLK1.n1180 0 0.10fF $ **FLOATING
C5224 CLK1.n1181 0 0.03fF $ **FLOATING
C5225 CLK1.n1182 0 0.10fF $ **FLOATING
C5226 CLK1.n1183 0 0.01fF $ **FLOATING
C5227 CLK1.n1184 0 0.11fF $ **FLOATING
C5228 CLK1.n1185 0 0.10fF $ **FLOATING
C5229 CLK1.t100 0 0.03fF
C5230 CLK1.n1186 0 0.10fF $ **FLOATING
C5231 CLK1.n1187 0 0.02fF $ **FLOATING
C5232 CLK1.n1188 0 0.02fF $ **FLOATING
C5233 CLK1.n1189 0 0.02fF $ **FLOATING
C5234 CLK1.n1190 0 0.09fF $ **FLOATING
C5235 CLK1.n1191 0 0.13fF $ **FLOATING
C5236 CLK1.n1192 0 0.09fF $ **FLOATING
C5237 CLK1.n1193 0 0.03fF $ **FLOATING
C5238 CLK1.n1194 0 0.03fF $ **FLOATING
C5239 CLK1.n1195 0 0.02fF $ **FLOATING
C5240 CLK1.n1196 0 0.03fF $ **FLOATING
C5241 CLK1.n1197 0 0.06fF $ **FLOATING
C5242 CLK1.n1198 0 0.06fF $ **FLOATING
C5243 CLK1.n1199 0 0.06fF $ **FLOATING
C5244 CLK1.n1200 0 0.03fF $ **FLOATING
C5245 CLK1.n1201 0 0.02fF $ **FLOATING
C5246 CLK1.n1202 0 0.03fF $ **FLOATING
C5247 CLK1.n1203 0 0.03fF $ **FLOATING
C5248 CLK1.n1204 0 0.03fF $ **FLOATING
C5249 CLK1.n1205 0 0.02fF $ **FLOATING
C5250 CLK1.n1206 0 0.03fF $ **FLOATING
C5251 CLK1.n1207 0 0.06fF $ **FLOATING
C5252 CLK1.n1208 0 0.14fF $ **FLOATING
C5253 CLK1.n1209 0 0.11fF $ **FLOATING
C5254 CLK1.n1210 0 0.18fF $ **FLOATING
C5255 CLK1.n1211 0 0.03fF $ **FLOATING
C5256 CLK1.n1212 0 0.02fF $ **FLOATING
C5257 CLK1.n1213 0 0.02fF $ **FLOATING
C5258 CLK1.n1214 0 0.29fF $ **FLOATING
C5259 CLK1.n1215 0 0.03fF $ **FLOATING
C5260 CLK1.n1216 0 0.03fF $ **FLOATING
C5261 CLK1.n1217 0 0.02fF $ **FLOATING
C5262 CLK1.n1218 0 0.03fF $ **FLOATING
C5263 CLK1.n1219 0 0.16fF $ **FLOATING
C5264 CLK1.n1220 0 0.09fF $ **FLOATING
C5265 CLK1.t129 0 0.09fF
C5266 CLK1.t14 0 0.09fF
C5267 CLK1.n1221 0 0.17fF $ **FLOATING
C5268 CLK1.n1222 0 0.03fF $ **FLOATING
C5269 CLK1.n1223 0 0.02fF $ **FLOATING
C5270 CLK1.n1224 0 0.17fF $ **FLOATING
C5271 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/CLK 0 0.02fF $ **FLOATING
C5272 CLK1.n1225 0 0.03fF $ **FLOATING
C5273 CLK1.n1226 0 0.03fF $ **FLOATING
C5274 CLK1.n1227 0 0.03fF $ **FLOATING
C5275 CLK1.n1228 0 0.02fF $ **FLOATING
C5276 CLK1.n1229 0 0.03fF $ **FLOATING
C5277 CLK1.n1230 0 0.16fF $ **FLOATING
C5278 CLK1.t16 0 0.09fF
C5279 CLK1.n1231 0 0.11fF $ **FLOATING
C5280 CLK1.n1232 0 0.18fF $ **FLOATING
C5281 CLK1.n1233 0 0.03fF $ **FLOATING
C5282 CLK1.n1234 0 0.02fF $ **FLOATING
C5283 CLK1.n1235 0 0.02fF $ **FLOATING
C5284 CLK1.n1236 0 0.03fF $ **FLOATING
C5285 CLK1.n1237 0 0.03fF $ **FLOATING
C5286 CLK1.n1238 0 0.03fF $ **FLOATING
C5287 CLK1.n1239 0 0.02fF $ **FLOATING
C5288 CLK1.n1240 0 0.03fF $ **FLOATING
C5289 CLK1.n1241 0 0.06fF $ **FLOATING
C5290 CLK1.n1242 0 0.06fF $ **FLOATING
C5291 CLK1.n1243 0 0.06fF $ **FLOATING
C5292 CLK1.n1244 0 0.03fF $ **FLOATING
C5293 CLK1.n1245 0 0.02fF $ **FLOATING
C5294 CLK1.n1246 0 0.02fF $ **FLOATING
C5295 CLK1.n1247 0 0.03fF $ **FLOATING
C5296 CLK1.n1248 0 0.03fF $ **FLOATING
C5297 CLK1.n1249 0 0.03fF $ **FLOATING
C5298 CLK1.n1250 0 0.02fF $ **FLOATING
C5299 CLK1.n1251 0 0.03fF $ **FLOATING
C5300 CLK1.n1252 0 0.06fF $ **FLOATING
C5301 CLK1.n1253 0 0.07fF $ **FLOATING
C5302 CLK1.n1254 0 0.13fF $ **FLOATING
C5303 CLK1.n1255 0 0.08fF $ **FLOATING
C5304 CLK1.n1256 0 0.13fF $ **FLOATING
C5305 CLK1.n1257 0 0.02fF $ **FLOATING
C5306 CLK1.n1258 0 0.01fF $ **FLOATING
C5307 CLK1.n1259 0 0.03fF $ **FLOATING
C5308 CLK1.n1260 0 0.06fF $ **FLOATING
C5309 CLK1.n1261 0 0.03fF $ **FLOATING
C5310 CLK1.n1262 0 0.02fF $ **FLOATING
C5311 CLK1.n1263 0 0.02fF $ **FLOATING
C5312 CLK1.t30 0 0.03fF
C5313 CLK1.t106 0 0.03fF
C5314 CLK1.n1264 0 0.15fF $ **FLOATING
C5315 CLK1.n1265 0 0.03fF $ **FLOATING
C5316 CLK1.n1266 0 0.02fF $ **FLOATING
C5317 CLK1.n1267 0 0.03fF $ **FLOATING
C5318 CLK1.n1268 0 0.06fF $ **FLOATING
C5319 CLK1.n1269 0 0.03fF $ **FLOATING
C5320 CLK1.n1270 0 0.02fF $ **FLOATING
C5321 CLK1.n1271 0 0.02fF $ **FLOATING
C5322 CLK1.n1272 0 0.02fF $ **FLOATING
C5323 CLK1.n1273 0 0.03fF $ **FLOATING
C5324 CLK1.t195 0 0.09fF
C5325 CLK1.n1274 0 0.03fF $ **FLOATING
C5326 CLK1.n1275 0 0.02fF $ **FLOATING
C5327 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_1/CLK 0 0.02fF $ **FLOATING
C5328 CLK1.n1276 0 0.02fF $ **FLOATING
C5329 CLK1.n1277 0 0.03fF $ **FLOATING
C5330 CLK1.n1278 0 0.16fF $ **FLOATING
C5331 CLK1.n1279 0 0.03fF $ **FLOATING
C5332 CLK1.n1280 0 0.02fF $ **FLOATING
C5333 CLK1.t147 0 0.05fF
C5334 CLK1.n1281 0 0.29fF $ **FLOATING
C5335 CLK1.n1282 0 0.02fF $ **FLOATING
C5336 CLK1.n1283 0 0.03fF $ **FLOATING
C5337 CLK1.n1284 0 0.06fF $ **FLOATING
C5338 CLK1.n1285 0 0.03fF $ **FLOATING
C5339 CLK1.n1286 0 0.02fF $ **FLOATING
C5340 CLK1.n1287 0 0.03fF $ **FLOATING
C5341 CLK1.n1288 0 0.02fF $ **FLOATING
C5342 CLK1.n1289 0 0.03fF $ **FLOATING
C5343 CLK1.n1290 0 0.06fF $ **FLOATING
C5344 CLK1.n1291 0 0.03fF $ **FLOATING
C5345 CLK1.n1292 0 0.02fF $ **FLOATING
C5346 CLK1.t105 0 0.03fF
C5347 CLK1.t29 0 0.03fF
C5348 CLK1.n1293 0 0.15fF $ **FLOATING
C5349 CLK1.n1294 0 0.03fF $ **FLOATING
C5350 CLK1.n1295 0 0.02fF $ **FLOATING
C5351 CLK1.n1296 0 0.03fF $ **FLOATING
C5352 CLK1.t99 0 0.07fF
C5353 CLK1.n1297 0 0.45fF $ **FLOATING
C5354 CLK1.n1298 0 0.02fF $ **FLOATING
C5355 CLK1.n1299 0 0.03fF $ **FLOATING
C5356 CLK1.n1300 0 0.14fF $ **FLOATING
C5357 CLK1.n1301 0 0.03fF $ **FLOATING
C5358 CLK1.n1302 0 0.02fF $ **FLOATING
C5359 CLK1.t19 0 0.05fF
C5360 CLK1.n1303 0 0.29fF $ **FLOATING
C5361 CLK1.n1304 0 0.02fF $ **FLOATING
C5362 CLK1.n1305 0 0.03fF $ **FLOATING
C5363 CLK1.n1306 0 0.09fF $ **FLOATING
C5364 CLK1.n1307 0 0.03fF $ **FLOATING
C5365 CLK1.n1308 0 0.02fF $ **FLOATING
C5366 CLK1.t28 0 0.03fF
C5367 CLK1.t21 0 0.03fF
C5368 CLK1.n1309 0 0.10fF $ **FLOATING
C5369 CLK1.n1310 0 0.03fF $ **FLOATING
C5370 CLK1.n1311 0 0.02fF $ **FLOATING
C5371 CLK1.n1312 0 0.03fF $ **FLOATING
C5372 CLK1.t25 0 0.09fF
C5373 CLK1.n1313 0 0.03fF $ **FLOATING
C5374 CLK1.n1314 0 0.02fF $ **FLOATING
C5375 CLK1.t26 0 0.05fF
C5376 CLK1.n1315 0 0.03fF $ **FLOATING
C5377 CLK1.n1316 0 0.02fF $ **FLOATING
C5378 CLK1.n1317 0 0.03fF $ **FLOATING
C5379 CLK1.n1318 0 0.07fF $ **FLOATING
C5380 CLK1.n1319 0 0.03fF $ **FLOATING
C5381 CLK1.n1320 0 0.02fF $ **FLOATING
C5382 CLK1.t111 0 0.07fF
C5383 CLK1.n1321 0 0.15fF $ **FLOATING
C5384 CLK1.n1322 0 0.47fF $ **FLOATING
C5385 CLK1.n1323 0 0.03fF $ **FLOATING
C5386 CLK1.n1324 0 0.03fF $ **FLOATING
C5387 CLK1.n1325 0 0.02fF $ **FLOATING
C5388 CLK1.n1326 0 0.03fF $ **FLOATING
C5389 CLK1.n1327 0 0.06fF $ **FLOATING
C5390 CLK1.n1328 0 0.14fF $ **FLOATING
C5391 CLK1.n1329 0 0.11fF $ **FLOATING
C5392 CLK1.n1330 0 0.18fF $ **FLOATING
C5393 CLK1.n1331 0 0.03fF $ **FLOATING
C5394 CLK1.n1332 0 0.02fF $ **FLOATING
C5395 CLK1.n1333 0 0.02fF $ **FLOATING
C5396 CLK1.n1334 0 0.29fF $ **FLOATING
C5397 CLK1.n1335 0 0.03fF $ **FLOATING
C5398 CLK1.n1336 0 0.03fF $ **FLOATING
C5399 CLK1.n1337 0 0.02fF $ **FLOATING
C5400 CLK1.n1338 0 0.03fF $ **FLOATING
C5401 CLK1.n1339 0 0.16fF $ **FLOATING
C5402 CLK1.n1340 0 0.09fF $ **FLOATING
C5403 CLK1.t27 0 0.09fF
C5404 CLK1.t20 0 0.09fF
C5405 CLK1.n1341 0 0.17fF $ **FLOATING
C5406 CLK1.n1342 0 0.03fF $ **FLOATING
C5407 CLK1.n1343 0 0.02fF $ **FLOATING
C5408 CLK1.n1344 0 0.17fF $ **FLOATING
C5409 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_1/CLK 0 0.02fF $ **FLOATING
C5410 CLK1.n1345 0 0.03fF $ **FLOATING
C5411 CLK1.n1346 0 0.03fF $ **FLOATING
C5412 CLK1.n1347 0 0.03fF $ **FLOATING
C5413 CLK1.n1348 0 0.02fF $ **FLOATING
C5414 CLK1.n1349 0 0.03fF $ **FLOATING
C5415 CLK1.n1350 0 0.16fF $ **FLOATING
C5416 CLK1.t18 0 0.09fF
C5417 CLK1.n1351 0 0.11fF $ **FLOATING
C5418 CLK1.n1352 0 0.18fF $ **FLOATING
C5419 CLK1.n1353 0 0.03fF $ **FLOATING
C5420 CLK1.n1354 0 0.02fF $ **FLOATING
C5421 CLK1.n1355 0 0.02fF $ **FLOATING
C5422 CLK1.n1356 0 0.03fF $ **FLOATING
C5423 CLK1.n1357 0 0.03fF $ **FLOATING
C5424 CLK1.n1358 0 0.03fF $ **FLOATING
C5425 CLK1.n1359 0 0.02fF $ **FLOATING
C5426 CLK1.n1360 0 0.03fF $ **FLOATING
C5427 CLK1.n1361 0 0.06fF $ **FLOATING
C5428 CLK1.n1362 0 0.07fF $ **FLOATING
C5429 CLK1.n1363 0 0.15fF $ **FLOATING
C5430 CLK1.n1364 0 0.10fF $ **FLOATING
C5431 CLK1.n1365 0 0.11fF $ **FLOATING
C5432 CLK1.n1366 0 0.21fF $ **FLOATING
C5433 CLK1.n1367 0 0.08fF $ **FLOATING
C5434 CLK1.n1368 0 0.06fF $ **FLOATING
C5435 CLK1.n1369 0 0.03fF $ **FLOATING
C5436 CLK1.n1370 0 0.02fF $ **FLOATING
C5437 CLK1.n1371 0 0.03fF $ **FLOATING
C5438 CLK1.n1372 0 0.02fF $ **FLOATING
C5439 CLK1.n1373 0 0.19fF $ **FLOATING
C5440 CLK1.n1374 0 0.03fF $ **FLOATING
C5441 CLK1.n1375 0 0.02fF $ **FLOATING
C5442 CLK1.n1376 0 0.03fF $ **FLOATING
C5443 CLK1.n1377 0 0.06fF $ **FLOATING
C5444 CLK1.n1378 0 0.06fF $ **FLOATING
C5445 CLK1.n1379 0 0.06fF $ **FLOATING
C5446 CLK1.n1380 0 0.03fF $ **FLOATING
C5447 CLK1.n1381 0 0.02fF $ **FLOATING
C5448 CLK1.n1382 0 0.03fF $ **FLOATING
C5449 CLK1.n1383 0 0.03fF $ **FLOATING
C5450 CLK1.n1384 0 0.02fF $ **FLOATING
C5451 CLK1.n1385 0 0.03fF $ **FLOATING
C5452 CLK1.n1386 0 0.02fF $ **FLOATING
C5453 CLK1.n1387 0 0.03fF $ **FLOATING
C5454 CLK1.n1388 0 0.14fF $ **FLOATING
C5455 CLK1.n1389 0 0.18fF $ **FLOATING
C5456 CLK1.t146 0 0.09fF
C5457 CLK1.n1390 0 0.11fF $ **FLOATING
C5458 CLK1.n1391 0 0.03fF $ **FLOATING
C5459 CLK1.n1392 0 0.02fF $ **FLOATING
C5460 CLK1.n1393 0 0.03fF $ **FLOATING
C5461 CLK1.n1394 0 0.03fF $ **FLOATING
C5462 CLK1.t172 0 0.03fF
C5463 CLK1.t149 0 0.03fF
C5464 CLK1.n1395 0 0.10fF $ **FLOATING
C5465 CLK1.n1396 0 0.17fF $ **FLOATING
C5466 CLK1.n1397 0 0.03fF $ **FLOATING
C5467 CLK1.n1398 0 0.02fF $ **FLOATING
C5468 CLK1.n1399 0 0.03fF $ **FLOATING
C5469 CLK1.n1400 0 0.09fF $ **FLOATING
C5470 CLK1.t171 0 0.09fF
C5471 CLK1.n1401 0 0.17fF $ **FLOATING
C5472 CLK1.t148 0 0.09fF
C5473 CLK1.n1402 0 0.16fF $ **FLOATING
C5474 CLK1.n1403 0 0.09fF $ **FLOATING
C5475 CLK1.n1404 0 0.03fF $ **FLOATING
C5476 CLK1.n1405 0 0.02fF $ **FLOATING
C5477 CLK1.n1406 0 0.03fF $ **FLOATING
C5478 CLK1.n1407 0 0.03fF $ **FLOATING
C5479 CLK1.t196 0 0.05fF
C5480 CLK1.n1408 0 0.29fF $ **FLOATING
C5481 CLK1.n1409 0 0.03fF $ **FLOATING
C5482 CLK1.n1410 0 0.02fF $ **FLOATING
C5483 CLK1.n1411 0 0.03fF $ **FLOATING
C5484 CLK1.n1412 0 0.11fF $ **FLOATING
C5485 CLK1.n1413 0 0.18fF $ **FLOATING
C5486 CLK1.n1414 0 0.14fF $ **FLOATING
C5487 CLK1.n1415 0 0.03fF $ **FLOATING
C5488 CLK1.n1416 0 0.02fF $ **FLOATING
C5489 CLK1.n1417 0 0.03fF $ **FLOATING
C5490 CLK1.n1418 0 0.03fF $ **FLOATING
C5491 CLK1.n1419 0 0.03fF $ **FLOATING
C5492 CLK1.n1420 0 0.02fF $ **FLOATING
C5493 CLK1.n1421 0 0.03fF $ **FLOATING
C5494 CLK1.n1422 0 0.06fF $ **FLOATING
C5495 CLK1.n1423 0 0.06fF $ **FLOATING
C5496 CLK1.n1424 0 0.06fF $ **FLOATING
C5497 CLK1.n1425 0 0.03fF $ **FLOATING
C5498 CLK1.n1426 0 0.02fF $ **FLOATING
C5499 CLK1.n1427 0 0.03fF $ **FLOATING
C5500 CLK1.n1428 0 0.19fF $ **FLOATING
C5501 CLK1.n1429 0 0.02fF $ **FLOATING
C5502 CLK1.n1430 0 0.03fF $ **FLOATING
C5503 CLK1.n1431 0 0.03fF $ **FLOATING
C5504 CLK1.n1432 0 0.02fF $ **FLOATING
C5505 CLK1.n1433 0 0.03fF $ **FLOATING
C5506 CLK1.n1434 0 0.06fF $ **FLOATING
C5507 CLK1.n1435 0 0.08fF $ **FLOATING
C5508 CLK1.n1436 0 0.19fF $ **FLOATING
C5509 CLK1.n1437 0 0.01fF $ **FLOATING
C5510 CLK1.n1438 0 0.00fF $ **FLOATING
C5511 CLK1.n1439 0 0.03fF $ **FLOATING
C5512 CLK1.n1440 0 0.36fF $ **FLOATING
C5513 CLK1.n1441 0 0.36fF $ **FLOATING
C5514 CLK1.n1442 0 0.02fF $ **FLOATING
C5515 CLK1.n1443 0 0.01fF $ **FLOATING
C5516 CLK1.n1444 0 0.03fF $ **FLOATING
C5517 CLK1.n1445 0 0.06fF $ **FLOATING
C5518 CLK1.n1446 0 0.03fF $ **FLOATING
C5519 CLK1.n1447 0 0.02fF $ **FLOATING
C5520 CLK1.n1448 0 0.02fF $ **FLOATING
C5521 CLK1.t119 0 0.03fF
C5522 CLK1.t23 0 0.03fF
C5523 CLK1.n1449 0 0.15fF $ **FLOATING
C5524 CLK1.n1450 0 0.03fF $ **FLOATING
C5525 CLK1.n1451 0 0.02fF $ **FLOATING
C5526 CLK1.n1452 0 0.03fF $ **FLOATING
C5527 CLK1.n1453 0 0.06fF $ **FLOATING
C5528 CLK1.n1454 0 0.03fF $ **FLOATING
C5529 CLK1.n1455 0 0.02fF $ **FLOATING
C5530 CLK1.n1456 0 0.02fF $ **FLOATING
C5531 CLK1.n1457 0 0.02fF $ **FLOATING
C5532 CLK1.n1458 0 0.03fF $ **FLOATING
C5533 CLK1.t49 0 0.09fF
C5534 CLK1.n1459 0 0.03fF $ **FLOATING
C5535 CLK1.n1460 0 0.02fF $ **FLOATING
C5536 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_XOR_v3_0/CLK 0 0.02fF $ **FLOATING
C5537 CLK1.n1461 0 0.02fF $ **FLOATING
C5538 CLK1.n1462 0 0.03fF $ **FLOATING
C5539 CLK1.n1463 0 0.16fF $ **FLOATING
C5540 CLK1.n1464 0 0.03fF $ **FLOATING
C5541 CLK1.n1465 0 0.02fF $ **FLOATING
C5542 CLK1.t108 0 0.05fF
C5543 CLK1.n1466 0 0.29fF $ **FLOATING
C5544 CLK1.n1467 0 0.02fF $ **FLOATING
C5545 CLK1.n1468 0 0.03fF $ **FLOATING
C5546 CLK1.n1469 0 0.06fF $ **FLOATING
C5547 CLK1.n1470 0 0.03fF $ **FLOATING
C5548 CLK1.n1471 0 0.02fF $ **FLOATING
C5549 CLK1.n1472 0 0.03fF $ **FLOATING
C5550 CLK1.n1473 0 0.02fF $ **FLOATING
C5551 CLK1.n1474 0 0.03fF $ **FLOATING
C5552 CLK1.n1475 0 0.06fF $ **FLOATING
C5553 CLK1.n1476 0 0.03fF $ **FLOATING
C5554 CLK1.n1477 0 0.02fF $ **FLOATING
C5555 CLK1.t59 0 0.03fF
C5556 CLK1.t192 0 0.03fF
C5557 CLK1.n1478 0 0.15fF $ **FLOATING
C5558 CLK1.n1479 0 0.03fF $ **FLOATING
C5559 CLK1.n1480 0 0.02fF $ **FLOATING
C5560 CLK1.n1481 0 0.03fF $ **FLOATING
C5561 CLK1.t98 0 0.07fF
C5562 CLK1.n1482 0 0.45fF $ **FLOATING
C5563 CLK1.n1483 0 0.02fF $ **FLOATING
C5564 CLK1.n1484 0 0.03fF $ **FLOATING
C5565 CLK1.n1485 0 0.14fF $ **FLOATING
C5566 CLK1.n1486 0 0.03fF $ **FLOATING
C5567 CLK1.n1487 0 0.02fF $ **FLOATING
C5568 CLK1.t86 0 0.05fF
C5569 CLK1.n1488 0 0.29fF $ **FLOATING
C5570 CLK1.n1489 0 0.02fF $ **FLOATING
C5571 CLK1.n1490 0 0.03fF $ **FLOATING
C5572 CLK1.n1491 0 0.09fF $ **FLOATING
C5573 CLK1.n1492 0 0.03fF $ **FLOATING
C5574 CLK1.n1493 0 0.02fF $ **FLOATING
C5575 CLK1.t3 0 0.03fF
C5576 CLK1.t84 0 0.03fF
C5577 CLK1.n1494 0 0.10fF $ **FLOATING
C5578 CLK1.n1495 0 0.03fF $ **FLOATING
C5579 CLK1.n1496 0 0.02fF $ **FLOATING
C5580 CLK1.n1497 0 0.03fF $ **FLOATING
C5581 CLK1.t0 0 0.09fF
C5582 CLK1.n1498 0 0.03fF $ **FLOATING
C5583 CLK1.n1499 0 0.02fF $ **FLOATING
C5584 CLK1.t1 0 0.05fF
C5585 CLK1.n1500 0 0.03fF $ **FLOATING
C5586 CLK1.n1501 0 0.02fF $ **FLOATING
C5587 CLK1.n1502 0 0.03fF $ **FLOATING
C5588 CLK1.n1503 0 0.07fF $ **FLOATING
C5589 CLK1.n1504 0 0.03fF $ **FLOATING
C5590 CLK1.n1505 0 0.02fF $ **FLOATING
C5591 CLK1.t164 0 0.07fF
C5592 CLK1.n1506 0 0.15fF $ **FLOATING
C5593 CLK1.n1507 0 0.47fF $ **FLOATING
C5594 CLK1.n1508 0 0.03fF $ **FLOATING
C5595 CLK1.n1509 0 0.03fF $ **FLOATING
C5596 CLK1.n1510 0 0.02fF $ **FLOATING
C5597 CLK1.n1511 0 0.03fF $ **FLOATING
C5598 CLK1.n1512 0 0.06fF $ **FLOATING
C5599 CLK1.n1513 0 0.14fF $ **FLOATING
C5600 CLK1.n1514 0 0.11fF $ **FLOATING
C5601 CLK1.n1515 0 0.18fF $ **FLOATING
C5602 CLK1.n1516 0 0.03fF $ **FLOATING
C5603 CLK1.n1517 0 0.02fF $ **FLOATING
C5604 CLK1.n1518 0 0.02fF $ **FLOATING
C5605 CLK1.n1519 0 0.29fF $ **FLOATING
C5606 CLK1.n1520 0 0.03fF $ **FLOATING
C5607 CLK1.n1521 0 0.03fF $ **FLOATING
C5608 CLK1.n1522 0 0.02fF $ **FLOATING
C5609 CLK1.n1523 0 0.03fF $ **FLOATING
C5610 CLK1.n1524 0 0.16fF $ **FLOATING
C5611 CLK1.n1525 0 0.09fF $ **FLOATING
C5612 CLK1.t2 0 0.09fF
C5613 CLK1.t83 0 0.09fF
C5614 CLK1.n1526 0 0.17fF $ **FLOATING
C5615 CLK1.n1527 0 0.03fF $ **FLOATING
C5616 CLK1.n1528 0 0.02fF $ **FLOATING
C5617 CLK1.n1529 0 0.17fF $ **FLOATING
C5618 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_INV4_0/CLK 0 0.02fF $ **FLOATING
C5619 CLK1.n1530 0 0.03fF $ **FLOATING
C5620 CLK1.n1531 0 0.03fF $ **FLOATING
C5621 CLK1.n1532 0 0.03fF $ **FLOATING
C5622 CLK1.n1533 0 0.02fF $ **FLOATING
C5623 CLK1.n1534 0 0.03fF $ **FLOATING
C5624 CLK1.n1535 0 0.16fF $ **FLOATING
C5625 CLK1.t85 0 0.09fF
C5626 CLK1.n1536 0 0.11fF $ **FLOATING
C5627 CLK1.n1537 0 0.18fF $ **FLOATING
C5628 CLK1.n1538 0 0.03fF $ **FLOATING
C5629 CLK1.n1539 0 0.02fF $ **FLOATING
C5630 CLK1.n1540 0 0.02fF $ **FLOATING
C5631 CLK1.n1541 0 0.03fF $ **FLOATING
C5632 CLK1.n1542 0 0.03fF $ **FLOATING
C5633 CLK1.n1543 0 0.03fF $ **FLOATING
C5634 CLK1.n1544 0 0.02fF $ **FLOATING
C5635 CLK1.n1545 0 0.03fF $ **FLOATING
C5636 CLK1.n1546 0 0.06fF $ **FLOATING
C5637 CLK1.n1547 0 0.07fF $ **FLOATING
C5638 CLK1.n1548 0 0.15fF $ **FLOATING
C5639 CLK1.n1549 0 0.10fF $ **FLOATING
C5640 CLK1.n1550 0 0.11fF $ **FLOATING
C5641 CLK1.n1551 0 0.21fF $ **FLOATING
C5642 CLK1.n1552 0 0.08fF $ **FLOATING
C5643 CLK1.n1553 0 0.06fF $ **FLOATING
C5644 CLK1.n1554 0 0.03fF $ **FLOATING
C5645 CLK1.n1555 0 0.02fF $ **FLOATING
C5646 CLK1.n1556 0 0.03fF $ **FLOATING
C5647 CLK1.n1557 0 0.02fF $ **FLOATING
C5648 CLK1.n1558 0 0.19fF $ **FLOATING
C5649 CLK1.n1559 0 0.03fF $ **FLOATING
C5650 CLK1.n1560 0 0.02fF $ **FLOATING
C5651 CLK1.n1561 0 0.03fF $ **FLOATING
C5652 CLK1.n1562 0 0.06fF $ **FLOATING
C5653 CLK1.n1563 0 0.06fF $ **FLOATING
C5654 CLK1.n1564 0 0.06fF $ **FLOATING
C5655 CLK1.n1565 0 0.03fF $ **FLOATING
C5656 CLK1.n1566 0 0.02fF $ **FLOATING
C5657 CLK1.n1567 0 0.03fF $ **FLOATING
C5658 CLK1.n1568 0 0.03fF $ **FLOATING
C5659 CLK1.n1569 0 0.02fF $ **FLOATING
C5660 CLK1.n1570 0 0.03fF $ **FLOATING
C5661 CLK1.n1571 0 0.02fF $ **FLOATING
C5662 CLK1.n1572 0 0.03fF $ **FLOATING
C5663 CLK1.n1573 0 0.14fF $ **FLOATING
C5664 CLK1.n1574 0 0.18fF $ **FLOATING
C5665 CLK1.t107 0 0.09fF
C5666 CLK1.n1575 0 0.11fF $ **FLOATING
C5667 CLK1.n1576 0 0.03fF $ **FLOATING
C5668 CLK1.n1577 0 0.02fF $ **FLOATING
C5669 CLK1.n1578 0 0.03fF $ **FLOATING
C5670 CLK1.n1579 0 0.03fF $ **FLOATING
C5671 CLK1.t110 0 0.03fF
C5672 CLK1.t153 0 0.03fF
C5673 CLK1.n1580 0 0.10fF $ **FLOATING
C5674 CLK1.n1581 0 0.17fF $ **FLOATING
C5675 CLK1.n1582 0 0.03fF $ **FLOATING
C5676 CLK1.n1583 0 0.02fF $ **FLOATING
C5677 CLK1.n1584 0 0.03fF $ **FLOATING
C5678 CLK1.n1585 0 0.09fF $ **FLOATING
C5679 CLK1.t109 0 0.09fF
C5680 CLK1.n1586 0 0.17fF $ **FLOATING
C5681 CLK1.t152 0 0.09fF
C5682 CLK1.n1587 0 0.16fF $ **FLOATING
C5683 CLK1.n1588 0 0.09fF $ **FLOATING
C5684 CLK1.n1589 0 0.03fF $ **FLOATING
C5685 CLK1.n1590 0 0.02fF $ **FLOATING
C5686 CLK1.n1591 0 0.03fF $ **FLOATING
C5687 CLK1.n1592 0 0.03fF $ **FLOATING
C5688 CLK1.t50 0 0.05fF
C5689 CLK1.n1593 0 0.29fF $ **FLOATING
C5690 CLK1.n1594 0 0.03fF $ **FLOATING
C5691 CLK1.n1595 0 0.02fF $ **FLOATING
C5692 CLK1.n1596 0 0.03fF $ **FLOATING
C5693 CLK1.n1597 0 0.11fF $ **FLOATING
C5694 CLK1.n1598 0 0.18fF $ **FLOATING
C5695 CLK1.n1599 0 0.14fF $ **FLOATING
C5696 CLK1.n1600 0 0.03fF $ **FLOATING
C5697 CLK1.n1601 0 0.02fF $ **FLOATING
C5698 CLK1.n1602 0 0.03fF $ **FLOATING
C5699 CLK1.n1603 0 0.03fF $ **FLOATING
C5700 CLK1.n1604 0 0.03fF $ **FLOATING
C5701 CLK1.n1605 0 0.02fF $ **FLOATING
C5702 CLK1.n1606 0 0.03fF $ **FLOATING
C5703 CLK1.n1607 0 0.06fF $ **FLOATING
C5704 CLK1.n1608 0 0.06fF $ **FLOATING
C5705 CLK1.n1609 0 0.06fF $ **FLOATING
C5706 CLK1.n1610 0 0.03fF $ **FLOATING
C5707 CLK1.n1611 0 0.02fF $ **FLOATING
C5708 CLK1.n1612 0 0.03fF $ **FLOATING
C5709 CLK1.n1613 0 0.19fF $ **FLOATING
C5710 CLK1.n1614 0 0.02fF $ **FLOATING
C5711 CLK1.n1615 0 0.03fF $ **FLOATING
C5712 CLK1.n1616 0 0.03fF $ **FLOATING
C5713 CLK1.n1617 0 0.02fF $ **FLOATING
C5714 CLK1.n1618 0 0.03fF $ **FLOATING
C5715 CLK1.n1619 0 0.06fF $ **FLOATING
C5716 CLK1.n1620 0 0.08fF $ **FLOATING
C5717 CLK1.n1621 0 0.19fF $ **FLOATING
C5718 CLK1.n1622 0 0.01fF $ **FLOATING
C5719 CLK1.n1623 0 0.00fF $ **FLOATING
C5720 CLK1.n1624 0 0.03fF $ **FLOATING
C5721 CLK1.n1625 0 0.07fF $ **FLOATING
C5722 CLK1.n1626 0 0.43fF $ **FLOATING
C5723 EESPFAL_Sbox_0/CLK1 0 0.36fF $ **FLOATING
C5724 EESPFAL_Sbox_0/EESPFAL_s0_0/CLK1 0 0.02fF $ **FLOATING
C5725 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t9 0 0.12fF
C5726 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t3 0 0.20fF
C5727 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t5 0 0.05fF
C5728 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t4 0 0.05fF
C5729 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n0 0 0.16fF $ **FLOATING
C5730 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t0 0 0.05fF
C5731 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t2 0 0.05fF
C5732 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n1 0 0.14fF $ **FLOATING
C5733 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t7 0 0.03fF
C5734 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t6 0 0.06fF
C5735 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t8 0 0.07fF
C5736 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n2 0 0.07fF $ **FLOATING
C5737 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT 0 0.01fF $ **FLOATING
C5738 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n3 0 0.03fF $ **FLOATING
C5739 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n4 0 0.21fF $ **FLOATING
C5740 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t1 0 0.20fF
C5741 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n5 0 0.21fF $ **FLOATING
C5742 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n6 0 0.30fF $ **FLOATING
C5743 CLK0.t18 0 0.02fF
C5744 CLK0.t16 0 0.02fF
C5745 CLK0.n0 0 0.06fF $ **FLOATING
C5746 CLK0.t12 0 0.03fF
C5747 CLK0.n1 0 0.02fF $ **FLOATING
C5748 CLK0.t19 0 0.02fF
C5749 CLK0.t26 0 0.02fF
C5750 CLK0.n2 0 0.04fF $ **FLOATING
C5751 CLK0.n3 0 0.01fF $ **FLOATING
C5752 CLK0.t10 0 0.02fF
C5753 CLK0.t21 0 0.02fF
C5754 CLK0.n4 0 0.04fF $ **FLOATING
C5755 CLK0.n5 0 0.01fF $ **FLOATING
C5756 CLK0.n6 0 0.01fF $ **FLOATING
C5757 CLK0.n7 0 0.02fF $ **FLOATING
C5758 CLK0.t30 0 0.02fF
C5759 CLK0.t32 0 0.02fF
C5760 CLK0.n8 0 0.04fF $ **FLOATING
C5761 CLK0.n9 0 0.01fF $ **FLOATING
C5762 CLK0.t34 0 0.02fF
C5763 CLK0.t1 0 0.02fF
C5764 CLK0.n10 0 0.04fF $ **FLOATING
C5765 CLK0.n11 0 0.01fF $ **FLOATING
C5766 CLK0.n12 0 0.01fF $ **FLOATING
C5767 CLK0.n13 0 0.05fF $ **FLOATING
C5768 CLK0.n14 0 0.02fF $ **FLOATING
C5769 CLK0.n15 0 0.01fF $ **FLOATING
C5770 CLK0.n16 0 0.12fF $ **FLOATING
C5771 CLK0.n17 0 0.03fF $ **FLOATING
C5772 CLK0.n18 0 0.02fF $ **FLOATING
C5773 CLK0.n19 0 0.01fF $ **FLOATING
C5774 CLK0.n20 0 0.06fF $ **FLOATING
C5775 CLK0.n21 0 0.03fF $ **FLOATING
C5776 CLK0.n22 0 0.02fF $ **FLOATING
C5777 CLK0.n23 0 0.01fF $ **FLOATING
C5778 CLK0.n24 0 0.01fF $ **FLOATING
C5779 CLK0.t43 0 0.03fF
C5780 CLK0.t8 0 0.02fF
C5781 CLK0.t36 0 0.02fF
C5782 CLK0.n25 0 0.06fF $ **FLOATING
C5783 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_3/CLK 0 0.01fF $ **FLOATING
C5784 CLK0.t38 0 0.03fF
C5785 CLK0.t9 0 0.02fF
C5786 CLK0.t33 0 0.02fF
C5787 CLK0.n26 0 0.09fF $ **FLOATING
C5788 CLK0.n27 0 0.05fF $ **FLOATING
C5789 CLK0.n28 0 0.02fF $ **FLOATING
C5790 CLK0.n29 0 0.01fF $ **FLOATING
C5791 CLK0.n30 0 0.12fF $ **FLOATING
C5792 CLK0.n31 0 0.03fF $ **FLOATING
C5793 CLK0.n32 0 0.02fF $ **FLOATING
C5794 CLK0.n33 0 0.01fF $ **FLOATING
C5795 CLK0.n34 0 0.06fF $ **FLOATING
C5796 CLK0.n35 0 0.03fF $ **FLOATING
C5797 CLK0.n36 0 0.02fF $ **FLOATING
C5798 CLK0.n37 0 0.01fF $ **FLOATING
C5799 CLK0.n38 0 0.01fF $ **FLOATING
C5800 CLK0.n39 0 0.11fF $ **FLOATING
C5801 CLK0.n40 0 0.03fF $ **FLOATING
C5802 CLK0.n41 0 0.02fF $ **FLOATING
C5803 CLK0.n42 0 0.01fF $ **FLOATING
C5804 CLK0.n43 0 0.02fF $ **FLOATING
C5805 CLK0.n44 0 0.03fF $ **FLOATING
C5806 CLK0.n45 0 0.02fF $ **FLOATING
C5807 CLK0.n46 0 0.01fF $ **FLOATING
C5808 CLK0.n47 0 0.02fF $ **FLOATING
C5809 CLK0.n48 0 0.03fF $ **FLOATING
C5810 CLK0.n49 0 0.02fF $ **FLOATING
C5811 CLK0.n50 0 0.01fF $ **FLOATING
C5812 CLK0.n51 0 0.02fF $ **FLOATING
C5813 CLK0.n52 0 0.03fF $ **FLOATING
C5814 CLK0.n53 0 0.02fF $ **FLOATING
C5815 CLK0.n54 0 0.01fF $ **FLOATING
C5816 CLK0.n55 0 0.02fF $ **FLOATING
C5817 CLK0.n56 0 0.08fF $ **FLOATING
C5818 CLK0.n57 0 0.02fF $ **FLOATING
C5819 CLK0.n58 0 0.01fF $ **FLOATING
C5820 CLK0.n59 0 0.02fF $ **FLOATING
C5821 CLK0.n60 0 0.10fF $ **FLOATING
C5822 CLK0.n61 0 0.02fF $ **FLOATING
C5823 CLK0.n62 0 0.01fF $ **FLOATING
C5824 CLK0.n63 0 0.01fF $ **FLOATING
C5825 CLK0.n64 0 0.17fF $ **FLOATING
C5826 CLK0.t37 0 0.05fF
C5827 CLK0.n65 0 0.06fF $ **FLOATING
C5828 CLK0.n66 0 0.02fF $ **FLOATING
C5829 CLK0.n67 0 0.01fF $ **FLOATING
C5830 CLK0.n68 0 0.02fF $ **FLOATING
C5831 CLK0.n69 0 0.09fF $ **FLOATING
C5832 CLK0.n70 0 0.02fF $ **FLOATING
C5833 CLK0.n71 0 0.01fF $ **FLOATING
C5834 CLK0.n72 0 0.02fF $ **FLOATING
C5835 CLK0.n73 0 0.02fF $ **FLOATING
C5836 CLK0.t35 0 0.05fF
C5837 CLK0.n74 0 0.05fF $ **FLOATING
C5838 CLK0.n75 0 0.02fF $ **FLOATING
C5839 CLK0.n76 0 0.01fF $ **FLOATING
C5840 CLK0.n77 0 0.10fF $ **FLOATING
C5841 CLK0.n78 0 0.02fF $ **FLOATING
C5842 CLK0.n79 0 0.01fF $ **FLOATING
C5843 CLK0.n80 0 0.10fF $ **FLOATING
C5844 CLK0.t7 0 0.05fF
C5845 CLK0.n81 0 0.05fF $ **FLOATING
C5846 CLK0.n82 0 0.02fF $ **FLOATING
C5847 CLK0.n83 0 0.01fF $ **FLOATING
C5848 CLK0.n84 0 0.02fF $ **FLOATING
C5849 CLK0.n85 0 0.09fF $ **FLOATING
C5850 CLK0.n86 0 0.02fF $ **FLOATING
C5851 CLK0.n87 0 0.01fF $ **FLOATING
C5852 CLK0.n88 0 0.02fF $ **FLOATING
C5853 CLK0.t42 0 0.05fF
C5854 CLK0.n89 0 0.06fF $ **FLOATING
C5855 CLK0.n90 0 0.02fF $ **FLOATING
C5856 CLK0.n91 0 0.01fF $ **FLOATING
C5857 CLK0.n92 0 0.02fF $ **FLOATING
C5858 CLK0.n93 0 0.17fF $ **FLOATING
C5859 CLK0.n94 0 0.10fF $ **FLOATING
C5860 CLK0.n95 0 0.02fF $ **FLOATING
C5861 CLK0.n96 0 0.01fF $ **FLOATING
C5862 CLK0.n97 0 0.01fF $ **FLOATING
C5863 CLK0.n98 0 0.08fF $ **FLOATING
C5864 CLK0.n99 0 0.02fF $ **FLOATING
C5865 CLK0.n100 0 0.01fF $ **FLOATING
C5866 CLK0.n101 0 0.02fF $ **FLOATING
C5867 CLK0.n102 0 0.03fF $ **FLOATING
C5868 CLK0.n103 0 0.02fF $ **FLOATING
C5869 CLK0.n104 0 0.01fF $ **FLOATING
C5870 CLK0.n105 0 0.02fF $ **FLOATING
C5871 CLK0.n106 0 0.03fF $ **FLOATING
C5872 CLK0.n107 0 0.02fF $ **FLOATING
C5873 CLK0.n108 0 0.01fF $ **FLOATING
C5874 CLK0.n109 0 0.02fF $ **FLOATING
C5875 CLK0.n110 0 0.03fF $ **FLOATING
C5876 CLK0.n111 0 0.02fF $ **FLOATING
C5877 CLK0.n112 0 0.01fF $ **FLOATING
C5878 CLK0.n113 0 0.02fF $ **FLOATING
C5879 CLK0.n114 0 0.03fF $ **FLOATING
C5880 CLK0.n115 0 0.02fF $ **FLOATING
C5881 CLK0.n116 0 0.01fF $ **FLOATING
C5882 CLK0.n117 0 0.02fF $ **FLOATING
C5883 CLK0.n118 0 0.04fF $ **FLOATING
C5884 CLK0.n119 0 0.05fF $ **FLOATING
C5885 CLK0.n120 0 0.01fF $ **FLOATING
C5886 CLK0.n121 0 0.01fF $ **FLOATING
C5887 CLK0.n122 0 0.06fF $ **FLOATING
C5888 CLK0.n123 0 0.07fF $ **FLOATING
C5889 CLK0.n124 0 0.01fF $ **FLOATING
C5890 CLK0.n125 0 0.01fF $ **FLOATING
C5891 CLK0.n126 0 0.04fF $ **FLOATING
C5892 CLK0.n127 0 0.05fF $ **FLOATING
C5893 CLK0.n128 0 0.02fF $ **FLOATING
C5894 CLK0.n129 0 0.01fF $ **FLOATING
C5895 CLK0.n130 0 0.12fF $ **FLOATING
C5896 CLK0.n131 0 0.04fF $ **FLOATING
C5897 CLK0.n132 0 0.02fF $ **FLOATING
C5898 CLK0.n133 0 0.01fF $ **FLOATING
C5899 CLK0.n134 0 0.06fF $ **FLOATING
C5900 CLK0.n135 0 0.04fF $ **FLOATING
C5901 CLK0.n136 0 0.02fF $ **FLOATING
C5902 CLK0.n137 0 0.01fF $ **FLOATING
C5903 CLK0.n138 0 0.01fF $ **FLOATING
C5904 CLK0.t23 0 0.03fF
C5905 CLK0.t31 0 0.03fF
C5906 CLK0.t39 0 0.02fF
C5907 CLK0.t5 0 0.02fF
C5908 CLK0.n139 0 0.06fF $ **FLOATING
C5909 CLK0.t25 0 0.02fF
C5910 CLK0.t29 0 0.02fF
C5911 CLK0.n140 0 0.06fF $ **FLOATING
C5912 EESPFAL_4in_XOR_0/EESPFAL_XOR_v3_1/CLK 0 0.01fF $ **FLOATING
C5913 CLK0.t3 0 0.03fF
C5914 CLK0.t28 0 0.03fF
C5915 CLK0.t41 0 0.02fF
C5916 CLK0.t40 0 0.02fF
C5917 CLK0.n141 0 0.09fF $ **FLOATING
C5918 CLK0.t6 0 0.02fF
C5919 CLK0.t27 0 0.02fF
C5920 CLK0.n142 0 0.09fF $ **FLOATING
C5921 CLK0.n143 0 0.05fF $ **FLOATING
C5922 CLK0.n144 0 0.02fF $ **FLOATING
C5923 CLK0.n145 0 0.01fF $ **FLOATING
C5924 CLK0.n146 0 0.12fF $ **FLOATING
C5925 CLK0.n147 0 0.04fF $ **FLOATING
C5926 CLK0.n148 0 0.02fF $ **FLOATING
C5927 CLK0.n149 0 0.01fF $ **FLOATING
C5928 CLK0.n150 0 0.06fF $ **FLOATING
C5929 CLK0.n151 0 0.04fF $ **FLOATING
C5930 CLK0.n152 0 0.02fF $ **FLOATING
C5931 CLK0.n153 0 0.01fF $ **FLOATING
C5932 CLK0.n154 0 0.01fF $ **FLOATING
C5933 CLK0.n155 0 0.21fF $ **FLOATING
C5934 CLK0.n156 0 0.04fF $ **FLOATING
C5935 CLK0.n157 0 0.02fF $ **FLOATING
C5936 CLK0.n158 0 0.01fF $ **FLOATING
C5937 CLK0.n159 0 0.02fF $ **FLOATING
C5938 CLK0.n160 0 0.04fF $ **FLOATING
C5939 CLK0.n161 0 0.02fF $ **FLOATING
C5940 CLK0.n162 0 0.01fF $ **FLOATING
C5941 CLK0.n163 0 0.02fF $ **FLOATING
C5942 CLK0.n164 0 0.04fF $ **FLOATING
C5943 CLK0.n165 0 0.02fF $ **FLOATING
C5944 CLK0.n166 0 0.01fF $ **FLOATING
C5945 CLK0.n167 0 0.02fF $ **FLOATING
C5946 CLK0.n168 0 0.03fF $ **FLOATING
C5947 CLK0.n169 0 0.02fF $ **FLOATING
C5948 CLK0.n170 0 0.01fF $ **FLOATING
C5949 CLK0.n171 0 0.02fF $ **FLOATING
C5950 CLK0.n172 0 0.12fF $ **FLOATING
C5951 CLK0.n173 0 0.02fF $ **FLOATING
C5952 CLK0.n174 0 0.01fF $ **FLOATING
C5953 CLK0.n175 0 0.02fF $ **FLOATING
C5954 CLK0.n176 0 0.17fF $ **FLOATING
C5955 CLK0.n177 0 0.02fF $ **FLOATING
C5956 CLK0.n178 0 0.01fF $ **FLOATING
C5957 CLK0.n179 0 0.01fF $ **FLOATING
C5958 CLK0.n180 0 0.33fF $ **FLOATING
C5959 CLK0.t2 0 0.08fF
C5960 CLK0.n181 0 0.10fF $ **FLOATING
C5961 CLK0.n182 0 0.02fF $ **FLOATING
C5962 CLK0.n183 0 0.01fF $ **FLOATING
C5963 CLK0.n184 0 0.02fF $ **FLOATING
C5964 CLK0.n185 0 0.15fF $ **FLOATING
C5965 CLK0.n186 0 0.02fF $ **FLOATING
C5966 CLK0.n187 0 0.01fF $ **FLOATING
C5967 CLK0.n188 0 0.02fF $ **FLOATING
C5968 CLK0.n189 0 0.02fF $ **FLOATING
C5969 CLK0.t4 0 0.08fF
C5970 CLK0.n190 0 0.09fF $ **FLOATING
C5971 CLK0.n191 0 0.02fF $ **FLOATING
C5972 CLK0.n192 0 0.01fF $ **FLOATING
C5973 CLK0.n193 0 0.16fF $ **FLOATING
C5974 CLK0.n194 0 0.02fF $ **FLOATING
C5975 CLK0.n195 0 0.01fF $ **FLOATING
C5976 CLK0.n196 0 0.19fF $ **FLOATING
C5977 CLK0.t24 0 0.08fF
C5978 CLK0.n197 0 0.09fF $ **FLOATING
C5979 CLK0.n198 0 0.02fF $ **FLOATING
C5980 CLK0.n199 0 0.01fF $ **FLOATING
C5981 CLK0.n200 0 0.02fF $ **FLOATING
C5982 CLK0.n201 0 0.15fF $ **FLOATING
C5983 CLK0.n202 0 0.02fF $ **FLOATING
C5984 CLK0.n203 0 0.01fF $ **FLOATING
C5985 CLK0.n204 0 0.02fF $ **FLOATING
C5986 CLK0.t22 0 0.08fF
C5987 CLK0.n205 0 0.10fF $ **FLOATING
C5988 CLK0.n206 0 0.02fF $ **FLOATING
C5989 CLK0.n207 0 0.01fF $ **FLOATING
C5990 CLK0.n208 0 0.02fF $ **FLOATING
C5991 CLK0.n209 0 0.33fF $ **FLOATING
C5992 CLK0.n210 0 0.17fF $ **FLOATING
C5993 CLK0.n211 0 0.02fF $ **FLOATING
C5994 CLK0.n212 0 0.01fF $ **FLOATING
C5995 CLK0.n213 0 0.01fF $ **FLOATING
C5996 CLK0.n214 0 0.12fF $ **FLOATING
C5997 CLK0.n215 0 0.02fF $ **FLOATING
C5998 CLK0.n216 0 0.01fF $ **FLOATING
C5999 CLK0.n217 0 0.02fF $ **FLOATING
C6000 CLK0.n218 0 0.03fF $ **FLOATING
C6001 CLK0.n219 0 0.02fF $ **FLOATING
C6002 CLK0.n220 0 0.01fF $ **FLOATING
C6003 CLK0.n221 0 0.02fF $ **FLOATING
C6004 CLK0.n222 0 0.04fF $ **FLOATING
C6005 CLK0.n223 0 0.02fF $ **FLOATING
C6006 CLK0.n224 0 0.01fF $ **FLOATING
C6007 CLK0.n225 0 0.02fF $ **FLOATING
C6008 CLK0.n226 0 0.04fF $ **FLOATING
C6009 CLK0.n227 0 0.02fF $ **FLOATING
C6010 CLK0.n228 0 0.01fF $ **FLOATING
C6011 CLK0.n229 0 0.02fF $ **FLOATING
C6012 CLK0.n230 0 0.04fF $ **FLOATING
C6013 CLK0.n231 0 0.02fF $ **FLOATING
C6014 CLK0.n232 0 0.01fF $ **FLOATING
C6015 CLK0.n233 0 0.02fF $ **FLOATING
C6016 CLK0.n234 0 0.07fF $ **FLOATING
C6017 CLK0.n235 0 0.05fF $ **FLOATING
C6018 CLK0.n236 0 0.01fF $ **FLOATING
C6019 CLK0.n237 0 0.01fF $ **FLOATING
C6020 CLK0.n238 0 0.06fF $ **FLOATING
C6021 CLK0.n239 0 0.07fF $ **FLOATING
C6022 CLK0.n240 0 0.01fF $ **FLOATING
C6023 CLK0.n241 0 0.01fF $ **FLOATING
C6024 CLK0.n242 0 0.04fF $ **FLOATING
C6025 CLK0.n243 0 0.05fF $ **FLOATING
C6026 CLK0.n244 0 0.02fF $ **FLOATING
C6027 CLK0.n245 0 0.01fF $ **FLOATING
C6028 CLK0.n246 0 0.12fF $ **FLOATING
C6029 CLK0.n247 0 0.03fF $ **FLOATING
C6030 CLK0.n248 0 0.02fF $ **FLOATING
C6031 CLK0.n249 0 0.01fF $ **FLOATING
C6032 CLK0.n250 0 0.06fF $ **FLOATING
C6033 CLK0.n251 0 0.03fF $ **FLOATING
C6034 CLK0.n252 0 0.02fF $ **FLOATING
C6035 CLK0.n253 0 0.01fF $ **FLOATING
C6036 CLK0.n254 0 0.01fF $ **FLOATING
C6037 CLK0.n255 0 0.04fF $ **FLOATING
C6038 CLK0.n256 0 0.03fF $ **FLOATING
C6039 CLK0.n257 0 0.02fF $ **FLOATING
C6040 CLK0.n258 0 0.01fF $ **FLOATING
C6041 CLK0.n259 0 0.02fF $ **FLOATING
C6042 CLK0.n260 0 0.03fF $ **FLOATING
C6043 CLK0.n261 0 0.02fF $ **FLOATING
C6044 CLK0.n262 0 0.01fF $ **FLOATING
C6045 CLK0.n263 0 0.02fF $ **FLOATING
C6046 CLK0.n264 0 0.03fF $ **FLOATING
C6047 CLK0.n265 0 0.02fF $ **FLOATING
C6048 CLK0.n266 0 0.01fF $ **FLOATING
C6049 CLK0.n267 0 0.02fF $ **FLOATING
C6050 CLK0.n268 0 0.03fF $ **FLOATING
C6051 CLK0.n269 0 0.02fF $ **FLOATING
C6052 CLK0.n270 0 0.01fF $ **FLOATING
C6053 CLK0.n271 0 0.02fF $ **FLOATING
C6054 CLK0.n272 0 0.08fF $ **FLOATING
C6055 CLK0.n273 0 0.02fF $ **FLOATING
C6056 CLK0.n274 0 0.01fF $ **FLOATING
C6057 CLK0.n275 0 0.02fF $ **FLOATING
C6058 CLK0.n276 0 0.10fF $ **FLOATING
C6059 CLK0.n277 0 0.02fF $ **FLOATING
C6060 CLK0.n278 0 0.01fF $ **FLOATING
C6061 CLK0.n279 0 0.01fF $ **FLOATING
C6062 CLK0.n280 0 0.17fF $ **FLOATING
C6063 CLK0.t11 0 0.05fF
C6064 CLK0.n281 0 0.06fF $ **FLOATING
C6065 CLK0.n282 0 0.02fF $ **FLOATING
C6066 CLK0.n283 0 0.01fF $ **FLOATING
C6067 CLK0.n284 0 0.02fF $ **FLOATING
C6068 CLK0.n285 0 0.09fF $ **FLOATING
C6069 CLK0.n286 0 0.02fF $ **FLOATING
C6070 CLK0.n287 0 0.01fF $ **FLOATING
C6071 CLK0.n288 0 0.02fF $ **FLOATING
C6072 CLK0.t17 0 0.05fF
C6073 CLK0.n289 0 0.05fF $ **FLOATING
C6074 CLK0.n290 0 0.02fF $ **FLOATING
C6075 CLK0.n291 0 0.01fF $ **FLOATING
C6076 CLK0.n292 0 0.02fF $ **FLOATING
C6077 CLK0.n293 0 0.10fF $ **FLOATING
C6078 CLK0.n294 0 0.02fF $ **FLOATING
C6079 CLK0.n295 0 0.01fF $ **FLOATING
C6080 CLK0.n296 0 0.10fF $ **FLOATING
C6081 CLK0.t14 0 0.03fF
C6082 CLK0.t0 0 0.02fF
C6083 CLK0.t20 0 0.02fF
C6084 CLK0.n297 0 0.09fF $ **FLOATING
C6085 CLK0.n298 0 0.12fF $ **FLOATING
C6086 EESPFAL_4in_XOR_0/CLK 0 0.01fF $ **FLOATING
C6087 CLK0.n299 0 0.03fF $ **FLOATING
C6088 CLK0.n300 0 0.05fF $ **FLOATING
C6089 CLK0.n301 0 0.02fF $ **FLOATING
C6090 CLK0.n302 0 0.01fF $ **FLOATING
C6091 CLK0.n303 0 0.02fF $ **FLOATING
C6092 CLK0.n304 0 0.03fF $ **FLOATING
C6093 CLK0.n305 0 0.02fF $ **FLOATING
C6094 CLK0.n306 0 0.01fF $ **FLOATING
C6095 CLK0.n307 0 0.02fF $ **FLOATING
C6096 CLK0.n308 0 0.03fF $ **FLOATING
C6097 CLK0.n309 0 0.02fF $ **FLOATING
C6098 CLK0.n310 0 0.01fF $ **FLOATING
C6099 CLK0.n311 0 0.01fF $ **FLOATING
C6100 CLK0.n312 0 0.11fF $ **FLOATING
C6101 CLK0.n313 0 0.03fF $ **FLOATING
C6102 CLK0.n314 0 0.02fF $ **FLOATING
C6103 CLK0.n315 0 0.01fF $ **FLOATING
C6104 CLK0.n316 0 0.02fF $ **FLOATING
C6105 CLK0.n317 0 0.03fF $ **FLOATING
C6106 CLK0.n318 0 0.02fF $ **FLOATING
C6107 CLK0.n319 0 0.01fF $ **FLOATING
C6108 CLK0.n320 0 0.02fF $ **FLOATING
C6109 CLK0.n321 0 0.03fF $ **FLOATING
C6110 CLK0.n322 0 0.02fF $ **FLOATING
C6111 CLK0.n323 0 0.01fF $ **FLOATING
C6112 CLK0.n324 0 0.02fF $ **FLOATING
C6113 CLK0.n325 0 0.03fF $ **FLOATING
C6114 CLK0.n326 0 0.02fF $ **FLOATING
C6115 CLK0.n327 0 0.01fF $ **FLOATING
C6116 CLK0.n328 0 0.02fF $ **FLOATING
C6117 CLK0.n329 0 0.08fF $ **FLOATING
C6118 CLK0.n330 0 0.02fF $ **FLOATING
C6119 CLK0.n331 0 0.01fF $ **FLOATING
C6120 CLK0.n332 0 0.02fF $ **FLOATING
C6121 CLK0.n333 0 0.10fF $ **FLOATING
C6122 CLK0.n334 0 0.02fF $ **FLOATING
C6123 CLK0.n335 0 0.01fF $ **FLOATING
C6124 CLK0.n336 0 0.01fF $ **FLOATING
C6125 CLK0.n337 0 0.17fF $ **FLOATING
C6126 CLK0.t13 0 0.05fF
C6127 CLK0.n338 0 0.06fF $ **FLOATING
C6128 CLK0.n339 0 0.02fF $ **FLOATING
C6129 CLK0.n340 0 0.01fF $ **FLOATING
C6130 CLK0.n341 0 0.02fF $ **FLOATING
C6131 CLK0.n342 0 0.09fF $ **FLOATING
C6132 CLK0.n343 0 0.02fF $ **FLOATING
C6133 CLK0.n344 0 0.01fF $ **FLOATING
C6134 CLK0.n345 0 0.02fF $ **FLOATING
C6135 CLK0.t15 0 0.05fF
C6136 CLK0.n346 0 0.05fF $ **FLOATING
C6137 CLK0.n347 0 0.02fF $ **FLOATING
C6138 CLK0.n348 0 0.01fF $ **FLOATING
C6139 CLK0.n349 0 0.02fF $ **FLOATING
C6140 CLK3.n0 0 0.02fF $ **FLOATING
C6141 CLK3.n1 0 0.02fF $ **FLOATING
C6142 CLK3.n2 0 0.03fF $ **FLOATING
C6143 CLK3.n3 0 0.06fF $ **FLOATING
C6144 CLK3.n4 0 0.03fF $ **FLOATING
C6145 CLK3.n5 0 0.02fF $ **FLOATING
C6146 CLK3.t26 0 0.03fF
C6147 CLK3.t17 0 0.03fF
C6148 CLK3.n6 0 0.16fF $ **FLOATING
C6149 CLK3.n7 0 0.03fF $ **FLOATING
C6150 CLK3.n8 0 0.02fF $ **FLOATING
C6151 CLK3.n9 0 0.03fF $ **FLOATING
C6152 CLK3.n10 0 0.11fF $ **FLOATING
C6153 CLK3.n11 0 0.03fF $ **FLOATING
C6154 CLK3.n12 0 0.02fF $ **FLOATING
C6155 CLK3.t42 0 0.05fF
C6156 CLK3.n13 0 0.03fF $ **FLOATING
C6157 CLK3.n14 0 0.02fF $ **FLOATING
C6158 CLK3.n15 0 0.03fF $ **FLOATING
C6159 CLK3.t36 0 0.09fF
C6160 CLK3.n16 0 0.03fF $ **FLOATING
C6161 CLK3.n17 0 0.02fF $ **FLOATING
C6162 CLK3.t37 0 0.03fF
C6163 CLK3.t39 0 0.03fF
C6164 CLK3.n18 0 0.10fF $ **FLOATING
C6165 CLK3.n19 0 0.03fF $ **FLOATING
C6166 CLK3.n20 0 0.02fF $ **FLOATING
C6167 CLK3.n21 0 0.03fF $ **FLOATING
C6168 CLK3.n22 0 0.14fF $ **FLOATING
C6169 CLK3.n23 0 0.03fF $ **FLOATING
C6170 CLK3.n24 0 0.02fF $ **FLOATING
C6171 CLK3.n25 0 0.03fF $ **FLOATING
C6172 CLK3.n26 0 0.02fF $ **FLOATING
C6173 CLK3.n27 0 0.03fF $ **FLOATING
C6174 CLK3.n28 0 0.07fF $ **FLOATING
C6175 CLK3.n29 0 0.03fF $ **FLOATING
C6176 CLK3.n30 0 0.02fF $ **FLOATING
C6177 CLK3.t27 0 0.08fF
C6178 CLK3.n31 0 0.13fF $ **FLOATING
C6179 CLK3.n32 0 0.36fF $ **FLOATING
C6180 CLK3.n33 0 0.03fF $ **FLOATING
C6181 CLK3.n34 0 0.03fF $ **FLOATING
C6182 CLK3.n35 0 0.02fF $ **FLOATING
C6183 CLK3.n36 0 0.03fF $ **FLOATING
C6184 CLK3.n37 0 0.06fF $ **FLOATING
C6185 CLK3.n38 0 0.06fF $ **FLOATING
C6186 CLK3.n39 0 0.06fF $ **FLOATING
C6187 CLK3.n40 0 0.03fF $ **FLOATING
C6188 CLK3.n41 0 0.02fF $ **FLOATING
C6189 CLK3.n42 0 0.03fF $ **FLOATING
C6190 CLK3.n43 0 0.03fF $ **FLOATING
C6191 CLK3.t4 0 0.05fF
C6192 CLK3.n44 0 0.30fF $ **FLOATING
C6193 CLK3.n45 0 0.02fF $ **FLOATING
C6194 CLK3.n46 0 0.02fF $ **FLOATING
C6195 CLK3.n47 0 0.03fF $ **FLOATING
C6196 CLK3.n48 0 0.18fF $ **FLOATING
C6197 CLK3.n49 0 0.11fF $ **FLOATING
C6198 CLK3.t3 0 0.09fF
C6199 CLK3.n50 0 0.10fF $ **FLOATING
C6200 CLK3.n51 0 0.16fF $ **FLOATING
C6201 CLK3.n52 0 0.03fF $ **FLOATING
C6202 CLK3.n53 0 0.02fF $ **FLOATING
C6203 CLK3.n54 0 0.03fF $ **FLOATING
C6204 CLK3.n55 0 0.03fF $ **FLOATING
C6205 CLK3.n56 0 0.18fF $ **FLOATING
C6206 CLK3.n57 0 0.02fF $ **FLOATING
C6207 CLK3.n58 0 0.03fF $ **FLOATING
C6208 CLK3.n59 0 0.17fF $ **FLOATING
C6209 CLK3.t38 0 0.09fF
C6210 CLK3.n60 0 0.10fF $ **FLOATING
C6211 CLK3.t41 0 0.09fF
C6212 CLK3.n61 0 0.16fF $ **FLOATING
C6213 CLK3.n62 0 0.03fF $ **FLOATING
C6214 CLK3.n63 0 0.02fF $ **FLOATING
C6215 CLK3.n64 0 0.03fF $ **FLOATING
C6216 CLK3.n65 0 0.03fF $ **FLOATING
C6217 CLK3.n66 0 0.30fF $ **FLOATING
C6218 CLK3.n67 0 0.02fF $ **FLOATING
C6219 CLK3.n68 0 0.02fF $ **FLOATING
C6220 CLK3.n69 0 0.03fF $ **FLOATING
C6221 CLK3.n70 0 0.18fF $ **FLOATING
C6222 CLK3.n71 0 0.14fF $ **FLOATING
C6223 CLK3.n72 0 0.06fF $ **FLOATING
C6224 CLK3.n73 0 0.03fF $ **FLOATING
C6225 CLK3.n74 0 0.02fF $ **FLOATING
C6226 CLK3.n75 0 0.03fF $ **FLOATING
C6227 CLK3.n76 0 0.03fF $ **FLOATING
C6228 CLK3.n77 0 0.19fF $ **FLOATING
C6229 CLK3.n78 0 0.01fF $ **FLOATING
C6230 CLK3.n79 0 0.13fF $ **FLOATING
C6231 CLK3.t10 0 0.08fF
C6232 CLK3.n80 0 0.03fF $ **FLOATING
C6233 CLK3.n81 0 0.02fF $ **FLOATING
C6234 CLK3.n82 0 0.03fF $ **FLOATING
C6235 CLK3.n83 0 0.06fF $ **FLOATING
C6236 CLK3.n84 0 0.03fF $ **FLOATING
C6237 CLK3.n85 0 0.02fF $ **FLOATING
C6238 CLK3.t12 0 0.03fF
C6239 CLK3.t40 0 0.03fF
C6240 CLK3.n86 0 0.16fF $ **FLOATING
C6241 CLK3.n87 0 0.03fF $ **FLOATING
C6242 CLK3.n88 0 0.02fF $ **FLOATING
C6243 CLK3.n89 0 0.03fF $ **FLOATING
C6244 CLK3.n90 0 0.18fF $ **FLOATING
C6245 CLK3.n91 0 0.03fF $ **FLOATING
C6246 CLK3.n92 0 0.02fF $ **FLOATING
C6247 CLK3.t44 0 0.05fF
C6248 CLK3.n93 0 0.03fF $ **FLOATING
C6249 CLK3.n94 0 0.02fF $ **FLOATING
C6250 CLK3.n95 0 0.03fF $ **FLOATING
C6251 CLK3.t5 0 0.09fF
C6252 CLK3.n96 0 0.03fF $ **FLOATING
C6253 CLK3.n97 0 0.02fF $ **FLOATING
C6254 CLK3.t14 0 0.03fF
C6255 CLK3.t6 0 0.03fF
C6256 CLK3.n98 0 0.10fF $ **FLOATING
C6257 CLK3.n99 0 0.03fF $ **FLOATING
C6258 CLK3.n100 0 0.02fF $ **FLOATING
C6259 CLK3.n101 0 0.03fF $ **FLOATING
C6260 CLK3.n102 0 0.18fF $ **FLOATING
C6261 CLK3.n103 0 0.03fF $ **FLOATING
C6262 CLK3.n104 0 0.02fF $ **FLOATING
C6263 CLK3.t1 0 0.05fF
C6264 CLK3.n105 0 0.03fF $ **FLOATING
C6265 CLK3.n106 0 0.02fF $ **FLOATING
C6266 CLK3.n107 0 0.03fF $ **FLOATING
C6267 CLK3.n108 0 0.06fF $ **FLOATING
C6268 CLK3.n109 0 0.03fF $ **FLOATING
C6269 CLK3.n110 0 0.02fF $ **FLOATING
C6270 CLK3.n111 0 0.03fF $ **FLOATING
C6271 CLK3.n112 0 0.02fF $ **FLOATING
C6272 CLK3.n113 0 0.03fF $ **FLOATING
C6273 CLK3.n114 0 0.13fF $ **FLOATING
C6274 CLK3.n115 0 0.02fF $ **FLOATING
C6275 CLK3.n116 0 0.02fF $ **FLOATING
C6276 CLK3.n117 0 0.02fF $ **FLOATING
C6277 CLK3.t7 0 0.03fF
C6278 CLK3.n118 0 0.13fF $ **FLOATING
C6279 CLK3.n119 0 0.03fF $ **FLOATING
C6280 CLK3.n120 0 0.02fF $ **FLOATING
C6281 CLK3.n121 0 0.03fF $ **FLOATING
C6282 CLK3.n122 0 0.06fF $ **FLOATING
C6283 CLK3.n123 0 0.03fF $ **FLOATING
C6284 CLK3.n124 0 0.02fF $ **FLOATING
C6285 CLK3.n125 0 0.03fF $ **FLOATING
C6286 CLK3.n126 0 0.02fF $ **FLOATING
C6287 CLK3.n127 0 0.03fF $ **FLOATING
C6288 CLK3.n128 0 0.18fF $ **FLOATING
C6289 CLK3.n129 0 0.03fF $ **FLOATING
C6290 CLK3.n130 0 0.02fF $ **FLOATING
C6291 CLK3.t35 0 0.05fF
C6292 CLK3.n131 0 0.03fF $ **FLOATING
C6293 CLK3.n132 0 0.02fF $ **FLOATING
C6294 CLK3.n133 0 0.03fF $ **FLOATING
C6295 CLK3.t21 0 0.09fF
C6296 CLK3.n134 0 0.03fF $ **FLOATING
C6297 CLK3.n135 0 0.02fF $ **FLOATING
C6298 CLK3.t22 0 0.03fF
C6299 CLK3.t19 0 0.03fF
C6300 CLK3.n136 0 0.10fF $ **FLOATING
C6301 CLK3.n137 0 0.03fF $ **FLOATING
C6302 CLK3.n138 0 0.02fF $ **FLOATING
C6303 CLK3.n139 0 0.03fF $ **FLOATING
C6304 CLK3.n140 0 0.17fF $ **FLOATING
C6305 CLK3.t18 0 0.09fF
C6306 CLK3.n141 0 0.18fF $ **FLOATING
C6307 CLK3.n142 0 0.03fF $ **FLOATING
C6308 CLK3.n143 0 0.02fF $ **FLOATING
C6309 CLK3.t24 0 0.05fF
C6310 CLK3.n144 0 0.03fF $ **FLOATING
C6311 CLK3.n145 0 0.02fF $ **FLOATING
C6312 CLK3.n146 0 0.03fF $ **FLOATING
C6313 CLK3.n147 0 0.06fF $ **FLOATING
C6314 CLK3.n148 0 0.03fF $ **FLOATING
C6315 CLK3.n149 0 0.02fF $ **FLOATING
C6316 CLK3.t28 0 0.03fF
C6317 CLK3.t9 0 0.03fF
C6318 CLK3.n150 0 0.16fF $ **FLOATING
C6319 CLK3.n151 0 0.03fF $ **FLOATING
C6320 CLK3.n152 0 0.02fF $ **FLOATING
C6321 CLK3.n153 0 0.03fF $ **FLOATING
C6322 CLK3.n154 0 0.13fF $ **FLOATING
C6323 CLK3.n155 0 0.01fF $ **FLOATING
C6324 CLK3.n156 0 0.01fF $ **FLOATING
C6325 CLK3.n157 0 0.01fF $ **FLOATING
C6326 CLK3.n158 0 0.13fF $ **FLOATING
C6327 CLK3.t25 0 0.08fF
C6328 CLK3.n159 0 0.03fF $ **FLOATING
C6329 CLK3.n160 0 0.02fF $ **FLOATING
C6330 CLK3.n161 0 0.03fF $ **FLOATING
C6331 CLK3.n162 0 0.06fF $ **FLOATING
C6332 CLK3.n163 0 0.03fF $ **FLOATING
C6333 CLK3.n164 0 0.02fF $ **FLOATING
C6334 CLK3.t33 0 0.03fF
C6335 CLK3.t20 0 0.03fF
C6336 CLK3.n165 0 0.16fF $ **FLOATING
C6337 CLK3.n166 0 0.03fF $ **FLOATING
C6338 CLK3.n167 0 0.02fF $ **FLOATING
C6339 CLK3.n168 0 0.03fF $ **FLOATING
C6340 CLK3.n169 0 0.18fF $ **FLOATING
C6341 CLK3.n170 0 0.03fF $ **FLOATING
C6342 CLK3.n171 0 0.02fF $ **FLOATING
C6343 CLK3.t46 0 0.05fF
C6344 CLK3.n172 0 0.03fF $ **FLOATING
C6345 CLK3.n173 0 0.02fF $ **FLOATING
C6346 CLK3.n174 0 0.03fF $ **FLOATING
C6347 CLK3.t15 0 0.09fF
C6348 CLK3.n175 0 0.03fF $ **FLOATING
C6349 CLK3.n176 0 0.02fF $ **FLOATING
C6350 CLK3.t32 0 0.03fF
C6351 CLK3.t16 0 0.03fF
C6352 CLK3.n177 0 0.10fF $ **FLOATING
C6353 CLK3.n178 0 0.03fF $ **FLOATING
C6354 CLK3.n179 0 0.02fF $ **FLOATING
C6355 CLK3.n180 0 0.03fF $ **FLOATING
C6356 CLK3.n181 0 0.18fF $ **FLOATING
C6357 CLK3.n182 0 0.03fF $ **FLOATING
C6358 CLK3.n183 0 0.02fF $ **FLOATING
C6359 CLK3.t30 0 0.05fF
C6360 CLK3.n184 0 0.03fF $ **FLOATING
C6361 CLK3.n185 0 0.02fF $ **FLOATING
C6362 CLK3.n186 0 0.03fF $ **FLOATING
C6363 CLK3.n187 0 0.06fF $ **FLOATING
C6364 CLK3.n188 0 0.03fF $ **FLOATING
C6365 CLK3.n189 0 0.02fF $ **FLOATING
C6366 CLK3.n190 0 0.03fF $ **FLOATING
C6367 CLK3.n191 0 0.02fF $ **FLOATING
C6368 CLK3.n192 0 0.03fF $ **FLOATING
C6369 CLK3.n193 0 0.13fF $ **FLOATING
C6370 CLK3.t8 0 0.08fF
C6371 CLK3.n194 0 0.36fF $ **FLOATING
C6372 CLK3.n195 0 0.03fF $ **FLOATING
C6373 CLK3.n196 0 0.02fF $ **FLOATING
C6374 CLK3.n197 0 0.03fF $ **FLOATING
C6375 CLK3.n198 0 0.07fF $ **FLOATING
C6376 CLK3.n199 0 0.06fF $ **FLOATING
C6377 CLK3.n200 0 0.06fF $ **FLOATING
C6378 CLK3.n201 0 0.03fF $ **FLOATING
C6379 CLK3.n202 0 0.02fF $ **FLOATING
C6380 CLK3.n203 0 0.03fF $ **FLOATING
C6381 CLK3.n204 0 0.03fF $ **FLOATING
C6382 CLK3.n205 0 0.03fF $ **FLOATING
C6383 CLK3.n206 0 0.02fF $ **FLOATING
C6384 CLK3.n207 0 0.03fF $ **FLOATING
C6385 CLK3.n208 0 0.06fF $ **FLOATING
C6386 CLK3.n209 0 0.06fF $ **FLOATING
C6387 CLK3.n210 0 0.14fF $ **FLOATING
C6388 CLK3.n211 0 0.03fF $ **FLOATING
C6389 CLK3.n212 0 0.02fF $ **FLOATING
C6390 CLK3.n213 0 0.03fF $ **FLOATING
C6391 CLK3.n214 0 0.02fF $ **FLOATING
C6392 CLK3.n215 0 0.30fF $ **FLOATING
C6393 CLK3.n216 0 0.03fF $ **FLOATING
C6394 CLK3.n217 0 0.02fF $ **FLOATING
C6395 CLK3.n218 0 0.03fF $ **FLOATING
C6396 CLK3.n219 0 0.11fF $ **FLOATING
C6397 CLK3.t29 0 0.09fF
C6398 CLK3.n220 0 0.16fF $ **FLOATING
C6399 CLK3.n221 0 0.17fF $ **FLOATING
C6400 CLK3.t31 0 0.09fF
C6401 CLK3.n222 0 0.10fF $ **FLOATING
C6402 CLK3.n223 0 0.03fF $ **FLOATING
C6403 CLK3.n224 0 0.02fF $ **FLOATING
C6404 CLK3.n225 0 0.03fF $ **FLOATING
C6405 CLK3.n226 0 0.18fF $ **FLOATING
C6406 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/CLK 0 0.02fF $ **FLOATING
C6407 CLK3.n227 0 0.03fF $ **FLOATING
C6408 CLK3.n228 0 0.02fF $ **FLOATING
C6409 CLK3.n229 0 0.03fF $ **FLOATING
C6410 CLK3.n230 0 0.10fF $ **FLOATING
C6411 CLK3.n231 0 0.16fF $ **FLOATING
C6412 CLK3.t45 0 0.09fF
C6413 CLK3.n232 0 0.11fF $ **FLOATING
C6414 CLK3.n233 0 0.03fF $ **FLOATING
C6415 CLK3.n234 0 0.02fF $ **FLOATING
C6416 CLK3.n235 0 0.03fF $ **FLOATING
C6417 CLK3.n236 0 0.30fF $ **FLOATING
C6418 CLK3.n237 0 0.02fF $ **FLOATING
C6419 CLK3.n238 0 0.03fF $ **FLOATING
C6420 CLK3.n239 0 0.02fF $ **FLOATING
C6421 CLK3.n240 0 0.03fF $ **FLOATING
C6422 CLK3.n241 0 0.14fF $ **FLOATING
C6423 CLK3.n242 0 0.06fF $ **FLOATING
C6424 CLK3.n243 0 0.06fF $ **FLOATING
C6425 CLK3.n244 0 0.03fF $ **FLOATING
C6426 CLK3.n245 0 0.02fF $ **FLOATING
C6427 CLK3.n246 0 0.03fF $ **FLOATING
C6428 CLK3.n247 0 0.19fF $ **FLOATING
C6429 CLK3.n248 0 0.02fF $ **FLOATING
C6430 CLK3.n249 0 0.03fF $ **FLOATING
C6431 CLK3.n250 0 0.02fF $ **FLOATING
C6432 CLK3.n251 0 0.03fF $ **FLOATING
C6433 CLK3.n252 0 0.06fF $ **FLOATING
C6434 CLK3.n253 0 0.06fF $ **FLOATING
C6435 CLK3.n254 0 0.07fF $ **FLOATING
C6436 CLK3.n255 0 0.03fF $ **FLOATING
C6437 CLK3.n256 0 0.02fF $ **FLOATING
C6438 CLK3.n257 0 0.03fF $ **FLOATING
C6439 CLK3.n258 0 0.34fF $ **FLOATING
C6440 CLK3.n259 0 0.41fF $ **FLOATING
C6441 EESPFAL_Sbox_0/EESPFAL_s3_0/CLK3 0 0.61fF $ **FLOATING
C6442 EESPFAL_Sbox_0/EESPFAL_s2_0/CLK3 0 0.55fF $ **FLOATING
C6443 CLK3.n260 0 0.44fF $ **FLOATING
C6444 CLK3.n261 0 0.01fF $ **FLOATING
C6445 CLK3.n262 0 0.02fF $ **FLOATING
C6446 CLK3.n263 0 0.00fF $ **FLOATING
C6447 CLK3.t11 0 0.08fF
C6448 CLK3.n264 0 0.36fF $ **FLOATING
C6449 CLK3.n265 0 0.01fF $ **FLOATING
C6450 CLK3.n266 0 0.00fF $ **FLOATING
C6451 CLK3.n267 0 0.00fF $ **FLOATING
C6452 CLK3.n268 0 0.03fF $ **FLOATING
C6453 CLK3.n269 0 0.07fF $ **FLOATING
C6454 CLK3.n270 0 0.06fF $ **FLOATING
C6455 CLK3.n271 0 0.06fF $ **FLOATING
C6456 CLK3.n272 0 0.03fF $ **FLOATING
C6457 CLK3.n273 0 0.02fF $ **FLOATING
C6458 CLK3.n274 0 0.03fF $ **FLOATING
C6459 CLK3.n275 0 0.02fF $ **FLOATING
C6460 CLK3.n276 0 0.19fF $ **FLOATING
C6461 CLK3.n277 0 0.03fF $ **FLOATING
C6462 CLK3.n278 0 0.02fF $ **FLOATING
C6463 CLK3.n279 0 0.03fF $ **FLOATING
C6464 CLK3.n280 0 0.06fF $ **FLOATING
C6465 CLK3.n281 0 0.06fF $ **FLOATING
C6466 CLK3.n282 0 0.14fF $ **FLOATING
C6467 CLK3.n283 0 0.03fF $ **FLOATING
C6468 CLK3.n284 0 0.02fF $ **FLOATING
C6469 CLK3.n285 0 0.03fF $ **FLOATING
C6470 CLK3.n286 0 0.02fF $ **FLOATING
C6471 CLK3.n287 0 0.30fF $ **FLOATING
C6472 CLK3.n288 0 0.03fF $ **FLOATING
C6473 CLK3.n289 0 0.02fF $ **FLOATING
C6474 CLK3.n290 0 0.03fF $ **FLOATING
C6475 CLK3.n291 0 0.11fF $ **FLOATING
C6476 CLK3.t23 0 0.09fF
C6477 CLK3.n292 0 0.16fF $ **FLOATING
C6478 CLK3.n293 0 0.10fF $ **FLOATING
C6479 CLK3.n294 0 0.03fF $ **FLOATING
C6480 CLK3.n295 0 0.02fF $ **FLOATING
C6481 CLK3.n296 0 0.03fF $ **FLOATING
C6482 EESPFAL_Sbox_0/EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/CLK 0 0.02fF $ **FLOATING
C6483 CLK3.n297 0 0.18fF $ **FLOATING
C6484 CLK3.n298 0 0.03fF $ **FLOATING
C6485 CLK3.n299 0 0.02fF $ **FLOATING
C6486 CLK3.n300 0 0.03fF $ **FLOATING
C6487 CLK3.n301 0 0.10fF $ **FLOATING
C6488 CLK3.n302 0 0.16fF $ **FLOATING
C6489 CLK3.t34 0 0.09fF
C6490 CLK3.n303 0 0.11fF $ **FLOATING
C6491 CLK3.n304 0 0.03fF $ **FLOATING
C6492 CLK3.n305 0 0.02fF $ **FLOATING
C6493 CLK3.n306 0 0.03fF $ **FLOATING
C6494 CLK3.n307 0 0.30fF $ **FLOATING
C6495 CLK3.n308 0 0.02fF $ **FLOATING
C6496 CLK3.n309 0 0.03fF $ **FLOATING
C6497 CLK3.n310 0 0.02fF $ **FLOATING
C6498 CLK3.n311 0 0.03fF $ **FLOATING
C6499 CLK3.n312 0 0.14fF $ **FLOATING
C6500 CLK3.n313 0 0.06fF $ **FLOATING
C6501 CLK3.n314 0 0.06fF $ **FLOATING
C6502 CLK3.n315 0 0.03fF $ **FLOATING
C6503 CLK3.n316 0 0.02fF $ **FLOATING
C6504 CLK3.n317 0 0.03fF $ **FLOATING
C6505 CLK3.n318 0 0.03fF $ **FLOATING
C6506 CLK3.n319 0 0.03fF $ **FLOATING
C6507 CLK3.n320 0 0.02fF $ **FLOATING
C6508 CLK3.n321 0 0.03fF $ **FLOATING
C6509 CLK3.n322 0 0.06fF $ **FLOATING
C6510 CLK3.n323 0 0.06fF $ **FLOATING
C6511 CLK3.n324 0 0.07fF $ **FLOATING
C6512 CLK3.n325 0 0.03fF $ **FLOATING
C6513 CLK3.n326 0 0.02fF $ **FLOATING
C6514 CLK3.n327 0 0.03fF $ **FLOATING
C6515 CLK3.n328 0 0.09fF $ **FLOATING
C6516 CLK3.n329 0 0.08fF $ **FLOATING
C6517 CLK3.n330 0 0.03fF $ **FLOATING
C6518 CLK3.n331 0 0.10fF $ **FLOATING
C6519 CLK3.n332 0 0.01fF $ **FLOATING
C6520 CLK3.n333 0 0.12fF $ **FLOATING
C6521 CLK3.n334 0 0.10fF $ **FLOATING
C6522 CLK3.t2 0 0.03fF
C6523 CLK3.n335 0 0.10fF $ **FLOATING
C6524 CLK3.n336 0 0.02fF $ **FLOATING
C6525 CLK3.n337 0 0.02fF $ **FLOATING
C6526 CLK3.n338 0 0.02fF $ **FLOATING
C6527 CLK3.n339 0 0.09fF $ **FLOATING
C6528 CLK3.n340 0 0.09fF $ **FLOATING
C6529 CLK3.n341 0 0.03fF $ **FLOATING
C6530 CLK3.n342 0 0.02fF $ **FLOATING
C6531 CLK3.n343 0 0.03fF $ **FLOATING
C6532 CLK3.n344 0 0.07fF $ **FLOATING
C6533 CLK3.n345 0 0.06fF $ **FLOATING
C6534 CLK3.n346 0 0.06fF $ **FLOATING
C6535 CLK3.n347 0 0.03fF $ **FLOATING
C6536 CLK3.n348 0 0.02fF $ **FLOATING
C6537 CLK3.n349 0 0.03fF $ **FLOATING
C6538 CLK3.n350 0 0.03fF $ **FLOATING
C6539 CLK3.n351 0 0.03fF $ **FLOATING
C6540 CLK3.n352 0 0.02fF $ **FLOATING
C6541 CLK3.n353 0 0.03fF $ **FLOATING
C6542 CLK3.n354 0 0.06fF $ **FLOATING
C6543 CLK3.n355 0 0.06fF $ **FLOATING
C6544 CLK3.n356 0 0.14fF $ **FLOATING
C6545 CLK3.n357 0 0.03fF $ **FLOATING
C6546 CLK3.n358 0 0.02fF $ **FLOATING
C6547 CLK3.n359 0 0.03fF $ **FLOATING
C6548 CLK3.n360 0 0.02fF $ **FLOATING
C6549 CLK3.n361 0 0.30fF $ **FLOATING
C6550 CLK3.n362 0 0.03fF $ **FLOATING
C6551 CLK3.n363 0 0.02fF $ **FLOATING
C6552 CLK3.n364 0 0.03fF $ **FLOATING
C6553 CLK3.n365 0 0.11fF $ **FLOATING
C6554 CLK3.t0 0 0.09fF
C6555 CLK3.n366 0 0.16fF $ **FLOATING
C6556 CLK3.n367 0 0.17fF $ **FLOATING
C6557 CLK3.t13 0 0.09fF
C6558 CLK3.n368 0 0.10fF $ **FLOATING
C6559 CLK3.n369 0 0.03fF $ **FLOATING
C6560 CLK3.n370 0 0.02fF $ **FLOATING
C6561 CLK3.n371 0 0.03fF $ **FLOATING
C6562 CLK3.n372 0 0.18fF $ **FLOATING
C6563 EESPFAL_Sbox_0/EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/CLK 0 0.02fF $ **FLOATING
C6564 CLK3.n373 0 0.03fF $ **FLOATING
C6565 CLK3.n374 0 0.02fF $ **FLOATING
C6566 CLK3.n375 0 0.03fF $ **FLOATING
C6567 CLK3.n376 0 0.10fF $ **FLOATING
C6568 CLK3.n377 0 0.16fF $ **FLOATING
C6569 CLK3.t43 0 0.09fF
C6570 CLK3.n378 0 0.11fF $ **FLOATING
C6571 CLK3.n379 0 0.03fF $ **FLOATING
C6572 CLK3.n380 0 0.02fF $ **FLOATING
C6573 CLK3.n381 0 0.03fF $ **FLOATING
C6574 CLK3.n382 0 0.30fF $ **FLOATING
C6575 CLK3.n383 0 0.02fF $ **FLOATING
C6576 CLK3.n384 0 0.03fF $ **FLOATING
C6577 CLK3.n385 0 0.02fF $ **FLOATING
C6578 CLK3.n386 0 0.03fF $ **FLOATING
C6579 CLK3.n387 0 0.14fF $ **FLOATING
C6580 CLK3.n388 0 0.06fF $ **FLOATING
C6581 CLK3.n389 0 0.06fF $ **FLOATING
C6582 CLK3.n390 0 0.03fF $ **FLOATING
C6583 CLK3.n391 0 0.02fF $ **FLOATING
C6584 CLK3.n392 0 0.03fF $ **FLOATING
C6585 CLK3.n393 0 0.19fF $ **FLOATING
C6586 CLK3.n394 0 0.02fF $ **FLOATING
C6587 CLK3.n395 0 0.03fF $ **FLOATING
C6588 CLK3.n396 0 0.02fF $ **FLOATING
C6589 CLK3.n397 0 0.03fF $ **FLOATING
C6590 CLK3.n398 0 0.06fF $ **FLOATING
C6591 CLK3.n399 0 0.06fF $ **FLOATING
C6592 CLK3.n400 0 0.07fF $ **FLOATING
C6593 CLK3.n401 0 0.03fF $ **FLOATING
C6594 CLK3.n402 0 0.02fF $ **FLOATING
C6595 CLK3.n403 0 0.03fF $ **FLOATING
C6596 CLK3.n404 0 0.34fF $ **FLOATING
C6597 CLK3.n405 0 0.39fF $ **FLOATING
C6598 EESPFAL_Sbox_0/EESPFAL_s1_0/CLK3 0 0.03fF $ **FLOATING
C6599 CLK3.n406 0 0.58fF $ **FLOATING
C6600 CLK3.n407 0 0.34fF $ **FLOATING
C6601 CLK3.n408 0 0.02fF $ **FLOATING
C6602 CLK3.n409 0 0.02fF $ **FLOATING
C6603 CLK3.n410 0 0.01fF $ **FLOATING
C6604 CLK3.n411 0 0.02fF $ **FLOATING
C6605 CLK3.n412 0 0.03fF $ **FLOATING
C6606 CLK3.n413 0 0.06fF $ **FLOATING
C6607 CLK3.n414 0 0.07fF $ **FLOATING
C6608 CLK3.n415 0 0.13fF $ **FLOATING
C6609 CLK3.n416 0 0.25fF $ **FLOATING
C6610 EESPFAL_Sbox_0/CLK3 0 0.23fF $ **FLOATING
C6611 EESPFAL_Sbox_0/EESPFAL_s0_0/CLK3 0 0.01fF $ **FLOATING
.ends

