magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -240 -85 -110 45
<< l67d20 >>
rect -225 -10 -185 30
rect -165 -10 -125 30
rect -225 -70 -185 -30
rect -165 -70 -125 -30
<< l67d44 >>
rect -214 2 -197 19
rect -154 2 -137 19
rect -214 -59 -197 -42
rect -154 -59 -137 -42
<< l68d20 >>
rect -240 -85 -110 45
<< l69d20 >>
rect -240 -85 -110 45
<< l71d20 >>
rect -240 -85 -110 45
<< l70d20 >>
rect -240 -85 -110 45
<< l68d44 >>
rect -213 3 -198 18
rect -153 3 -138 18
rect -213 -58 -198 -43
rect -153 -58 -138 -43
<< l70d44 >>
rect -215 0 -195 20
rect -155 0 -135 20
rect -215 -60 -195 -40
rect -155 -60 -135 -40
<< end >>
