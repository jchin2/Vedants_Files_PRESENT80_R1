magic
tech sky130A
magscale 1 2
timestamp 1670967196
<< error_p >>
rect 17 -295 41 295
<< locali >>
rect -17 295 17 352
rect -17 -352 17 -295
<< rlocali >>
rect -17 -295 17 295
<< properties >>
string gencell sky130_fd_pr__res_generic_l1
string library sky130
string parameters w 0.170 l 2.95 m 1 nx 1 wmin 0.17 lmin 0.17 rho 12.8 val 222.117 dummy 0 dw 0.0 term 0.0 snake 0 roverlap 0
<< end >>
