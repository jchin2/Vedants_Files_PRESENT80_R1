magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -815 580 -125 630
<< l67d20 >>
rect -815 585 -125 625
<< l67d44 >>
rect -799 597 -782 614
rect -759 597 -742 614
rect -719 597 -702 614
rect -679 597 -662 614
rect -639 597 -622 614
rect -599 597 -582 614
rect -559 597 -542 614
rect -519 597 -502 614
rect -479 597 -462 614
rect -439 597 -422 614
rect -399 597 -382 614
rect -359 597 -342 614
rect -319 597 -302 614
rect -279 597 -262 614
rect -239 597 -222 614
rect -199 597 -182 614
rect -159 597 -142 614
<< l68d20 >>
rect -815 580 -125 630
<< end >>
