* NGSPICE file created from EESPFAL_NOR_v3.ext - technology: sky130A

.subckt EESPFAL_NOR_v3 A A_bar B B_bar OUT OUT_bar Dis GND CLK
X0 a_n1820_550# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=6e+12p ps=2.62e+07u w=1.5e+06u l=150000u
X1 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X2 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u M=2
X3 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X4 OUT_bar B_bar a_n1820_550# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X6 OUT A CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 CLK B OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

