magic
tech sky130A
timestamp 1667079175
<< nwell >>
rect -1170 735 -130 830
rect -855 540 -445 735
<< nmos >>
rect -1085 120 -1070 270
rect -1010 120 -995 270
rect -935 120 -920 270
rect -770 120 -755 270
rect -695 120 -680 270
rect -620 120 -605 270
rect -545 120 -530 270
rect -380 120 -365 270
rect -305 120 -290 270
rect -230 120 -215 270
<< pmos >>
rect -770 565 -755 715
rect -695 565 -680 715
rect -620 565 -605 715
rect -545 565 -530 715
<< ndiff >>
rect -1145 235 -1085 270
rect -1145 215 -1125 235
rect -1105 215 -1085 235
rect -1145 195 -1085 215
rect -1145 175 -1125 195
rect -1105 175 -1085 195
rect -1145 155 -1085 175
rect -1145 135 -1125 155
rect -1105 135 -1085 155
rect -1145 120 -1085 135
rect -1070 120 -1010 270
rect -995 120 -935 270
rect -920 235 -860 270
rect -920 215 -900 235
rect -880 215 -860 235
rect -920 195 -860 215
rect -920 175 -900 195
rect -880 175 -860 195
rect -920 155 -860 175
rect -920 135 -900 155
rect -880 135 -860 155
rect -920 120 -860 135
rect -830 235 -770 270
rect -830 215 -810 235
rect -790 215 -770 235
rect -830 195 -770 215
rect -830 175 -810 195
rect -790 175 -770 195
rect -830 155 -770 175
rect -830 135 -810 155
rect -790 135 -770 155
rect -830 120 -770 135
rect -755 235 -695 270
rect -755 215 -735 235
rect -715 215 -695 235
rect -755 195 -695 215
rect -755 175 -735 195
rect -715 175 -695 195
rect -755 155 -695 175
rect -755 135 -735 155
rect -715 135 -695 155
rect -755 120 -695 135
rect -680 235 -620 270
rect -680 215 -660 235
rect -640 215 -620 235
rect -680 195 -620 215
rect -680 175 -660 195
rect -640 175 -620 195
rect -680 155 -620 175
rect -680 135 -660 155
rect -640 135 -620 155
rect -680 120 -620 135
rect -605 235 -545 270
rect -605 215 -585 235
rect -565 215 -545 235
rect -605 195 -545 215
rect -605 175 -585 195
rect -565 175 -545 195
rect -605 155 -545 175
rect -605 135 -585 155
rect -565 135 -545 155
rect -605 120 -545 135
rect -530 235 -470 270
rect -530 215 -510 235
rect -490 215 -470 235
rect -530 195 -470 215
rect -530 175 -510 195
rect -490 175 -470 195
rect -530 155 -470 175
rect -530 135 -510 155
rect -490 135 -470 155
rect -530 120 -470 135
rect -440 235 -380 270
rect -440 215 -420 235
rect -400 215 -380 235
rect -440 195 -380 215
rect -440 175 -420 195
rect -400 175 -380 195
rect -440 155 -380 175
rect -440 135 -420 155
rect -400 135 -380 155
rect -440 120 -380 135
rect -365 235 -305 270
rect -365 215 -345 235
rect -325 215 -305 235
rect -365 195 -305 215
rect -365 175 -345 195
rect -325 175 -305 195
rect -365 155 -305 175
rect -365 135 -345 155
rect -325 135 -305 155
rect -365 120 -305 135
rect -290 235 -230 270
rect -290 215 -270 235
rect -250 215 -230 235
rect -290 195 -230 215
rect -290 175 -270 195
rect -250 175 -230 195
rect -290 155 -230 175
rect -290 135 -270 155
rect -250 135 -230 155
rect -290 120 -230 135
rect -215 235 -155 270
rect -215 215 -195 235
rect -175 215 -155 235
rect -215 195 -155 215
rect -215 175 -195 195
rect -175 175 -155 195
rect -215 155 -155 175
rect -215 135 -195 155
rect -175 135 -155 155
rect -215 120 -155 135
<< pdiff >>
rect -830 680 -770 715
rect -830 660 -810 680
rect -790 660 -770 680
rect -830 640 -770 660
rect -830 620 -810 640
rect -790 620 -770 640
rect -830 600 -770 620
rect -830 580 -810 600
rect -790 580 -770 600
rect -830 565 -770 580
rect -755 680 -695 715
rect -755 660 -735 680
rect -715 660 -695 680
rect -755 640 -695 660
rect -755 620 -735 640
rect -715 620 -695 640
rect -755 600 -695 620
rect -755 580 -735 600
rect -715 580 -695 600
rect -755 565 -695 580
rect -680 680 -620 715
rect -680 660 -660 680
rect -640 660 -620 680
rect -680 640 -620 660
rect -680 620 -660 640
rect -640 620 -620 640
rect -680 600 -620 620
rect -680 580 -660 600
rect -640 580 -620 600
rect -680 565 -620 580
rect -605 680 -545 715
rect -605 660 -585 680
rect -565 660 -545 680
rect -605 640 -545 660
rect -605 620 -585 640
rect -565 620 -545 640
rect -605 600 -545 620
rect -605 580 -585 600
rect -565 580 -545 600
rect -605 565 -545 580
rect -530 680 -470 715
rect -530 660 -510 680
rect -490 660 -470 680
rect -530 640 -470 660
rect -530 620 -510 640
rect -490 620 -470 640
rect -530 600 -470 620
rect -530 580 -510 600
rect -490 580 -470 600
rect -530 565 -470 580
<< ndiffc >>
rect -1125 215 -1105 235
rect -1125 175 -1105 195
rect -1125 135 -1105 155
rect -900 215 -880 235
rect -900 175 -880 195
rect -900 135 -880 155
rect -810 215 -790 235
rect -810 175 -790 195
rect -810 135 -790 155
rect -735 215 -715 235
rect -735 175 -715 195
rect -735 135 -715 155
rect -660 215 -640 235
rect -660 175 -640 195
rect -660 135 -640 155
rect -585 215 -565 235
rect -585 175 -565 195
rect -585 135 -565 155
rect -510 215 -490 235
rect -510 175 -490 195
rect -510 135 -490 155
rect -420 215 -400 235
rect -420 175 -400 195
rect -420 135 -400 155
rect -345 215 -325 235
rect -345 175 -325 195
rect -345 135 -325 155
rect -270 215 -250 235
rect -270 175 -250 195
rect -270 135 -250 155
rect -195 215 -175 235
rect -195 175 -175 195
rect -195 135 -175 155
<< pdiffc >>
rect -810 660 -790 680
rect -810 620 -790 640
rect -810 580 -790 600
rect -735 660 -715 680
rect -735 620 -715 640
rect -735 580 -715 600
rect -660 660 -640 680
rect -660 620 -640 640
rect -660 580 -640 600
rect -585 660 -565 680
rect -585 620 -565 640
rect -585 580 -565 600
rect -510 660 -490 680
rect -510 620 -490 640
rect -510 580 -490 600
<< psubdiff >>
rect -1150 35 -150 50
rect -1150 15 -1140 35
rect -1120 15 -1100 35
rect -1080 15 -1060 35
rect -1040 15 -1020 35
rect -1000 15 -980 35
rect -960 15 -940 35
rect -920 15 -900 35
rect -880 15 -860 35
rect -840 15 -820 35
rect -800 15 -780 35
rect -760 15 -740 35
rect -720 15 -700 35
rect -680 15 -660 35
rect -640 15 -620 35
rect -600 15 -580 35
rect -560 15 -540 35
rect -520 15 -500 35
rect -480 15 -460 35
rect -440 15 -420 35
rect -400 15 -380 35
rect -360 15 -340 35
rect -320 15 -300 35
rect -280 15 -260 35
rect -240 15 -220 35
rect -200 15 -180 35
rect -160 15 -150 35
rect -1150 0 -150 15
<< nsubdiff >>
rect -1150 790 -150 805
rect -1150 770 -1140 790
rect -1120 770 -1100 790
rect -1080 770 -1060 790
rect -1040 770 -1020 790
rect -1000 770 -980 790
rect -960 770 -940 790
rect -920 770 -900 790
rect -880 770 -860 790
rect -840 770 -820 790
rect -800 770 -780 790
rect -760 770 -740 790
rect -720 770 -700 790
rect -680 770 -660 790
rect -640 770 -620 790
rect -600 770 -580 790
rect -560 770 -540 790
rect -520 770 -500 790
rect -480 770 -460 790
rect -440 770 -420 790
rect -400 770 -380 790
rect -360 770 -340 790
rect -320 770 -300 790
rect -280 770 -260 790
rect -240 770 -220 790
rect -200 770 -180 790
rect -160 770 -150 790
rect -1150 755 -150 770
<< psubdiffcont >>
rect -1140 15 -1120 35
rect -1100 15 -1080 35
rect -1060 15 -1040 35
rect -1020 15 -1000 35
rect -980 15 -960 35
rect -940 15 -920 35
rect -900 15 -880 35
rect -860 15 -840 35
rect -820 15 -800 35
rect -780 15 -760 35
rect -740 15 -720 35
rect -700 15 -680 35
rect -660 15 -640 35
rect -620 15 -600 35
rect -580 15 -560 35
rect -540 15 -520 35
rect -500 15 -480 35
rect -460 15 -440 35
rect -420 15 -400 35
rect -380 15 -360 35
rect -340 15 -320 35
rect -300 15 -280 35
rect -260 15 -240 35
rect -220 15 -200 35
rect -180 15 -160 35
<< nsubdiffcont >>
rect -1140 770 -1120 790
rect -1100 770 -1080 790
rect -1060 770 -1040 790
rect -1020 770 -1000 790
rect -980 770 -960 790
rect -940 770 -920 790
rect -900 770 -880 790
rect -860 770 -840 790
rect -820 770 -800 790
rect -780 770 -760 790
rect -740 770 -720 790
rect -700 770 -680 790
rect -660 770 -640 790
rect -620 770 -600 790
rect -580 770 -560 790
rect -540 770 -520 790
rect -500 770 -480 790
rect -460 770 -440 790
rect -420 770 -400 790
rect -380 770 -360 790
rect -340 770 -320 790
rect -300 770 -280 790
rect -260 770 -240 790
rect -220 770 -200 790
rect -180 770 -160 790
<< poly >>
rect -770 730 -680 745
rect -770 715 -755 730
rect -695 715 -680 730
rect -620 730 -530 745
rect -620 715 -605 730
rect -545 715 -530 730
rect -770 550 -755 565
rect -695 490 -680 565
rect -620 550 -605 565
rect -545 550 -530 565
rect -645 540 -605 550
rect -645 520 -635 540
rect -615 520 -605 540
rect -645 510 -605 520
rect -695 480 -655 490
rect -695 460 -685 480
rect -665 460 -655 480
rect -695 450 -655 460
rect -1105 400 -1065 410
rect -1105 380 -1095 400
rect -1075 380 -1065 400
rect -1105 370 -1065 380
rect -1085 270 -1070 370
rect -1035 350 -995 360
rect -1035 330 -1025 350
rect -1005 330 -995 350
rect -1035 320 -995 330
rect -1010 270 -995 320
rect -960 310 -920 320
rect -960 290 -950 310
rect -930 290 -920 310
rect -960 280 -920 290
rect -935 270 -920 280
rect -770 270 -755 285
rect -695 270 -680 450
rect -620 270 -605 510
rect -255 430 -215 440
rect -255 410 -245 430
rect -225 410 -215 430
rect -255 400 -215 410
rect -330 380 -290 390
rect -330 360 -320 380
rect -300 360 -290 380
rect -330 350 -290 360
rect -405 330 -365 340
rect -405 310 -395 330
rect -375 310 -365 330
rect -405 300 -365 310
rect -545 270 -530 285
rect -380 270 -365 300
rect -305 270 -290 350
rect -230 270 -215 400
rect -1085 105 -1070 120
rect -1010 105 -995 120
rect -935 105 -920 120
rect -770 105 -755 120
rect -695 105 -680 120
rect -620 105 -605 120
rect -545 105 -530 120
rect -380 105 -365 120
rect -305 105 -290 120
rect -230 105 -215 120
rect -770 95 -730 105
rect -770 75 -760 95
rect -740 75 -730 95
rect -770 65 -730 75
rect -570 95 -530 105
rect -570 75 -560 95
rect -540 75 -530 95
rect -570 65 -530 75
<< polycont >>
rect -635 520 -615 540
rect -685 460 -665 480
rect -1095 380 -1075 400
rect -1025 330 -1005 350
rect -950 290 -930 310
rect -245 410 -225 430
rect -320 360 -300 380
rect -395 310 -375 330
rect -760 75 -740 95
rect -560 75 -540 95
<< locali >>
rect -1150 790 -150 800
rect -1150 770 -1140 790
rect -1120 770 -1100 790
rect -1080 770 -1060 790
rect -1040 770 -1020 790
rect -1000 770 -980 790
rect -960 770 -940 790
rect -920 770 -900 790
rect -880 770 -860 790
rect -840 770 -820 790
rect -800 770 -780 790
rect -760 770 -740 790
rect -720 770 -700 790
rect -680 770 -660 790
rect -640 770 -620 790
rect -600 770 -580 790
rect -560 770 -540 790
rect -520 770 -500 790
rect -480 770 -460 790
rect -440 770 -420 790
rect -400 770 -380 790
rect -360 770 -340 790
rect -320 770 -300 790
rect -280 770 -260 790
rect -240 770 -220 790
rect -200 770 -180 790
rect -160 770 -150 790
rect -1150 760 -150 770
rect -820 680 -780 695
rect -820 660 -810 680
rect -790 660 -780 680
rect -820 640 -780 660
rect -820 620 -810 640
rect -790 620 -780 640
rect -820 600 -780 620
rect -820 580 -810 600
rect -790 580 -780 600
rect -820 570 -780 580
rect -745 680 -705 695
rect -745 660 -735 680
rect -715 660 -705 680
rect -745 640 -705 660
rect -745 620 -735 640
rect -715 620 -705 640
rect -745 600 -705 620
rect -745 580 -735 600
rect -715 580 -705 600
rect -745 565 -705 580
rect -670 680 -630 695
rect -670 660 -660 680
rect -640 660 -630 680
rect -670 640 -630 660
rect -670 620 -660 640
rect -640 620 -630 640
rect -670 600 -630 620
rect -670 580 -660 600
rect -640 580 -630 600
rect -670 570 -630 580
rect -595 680 -555 695
rect -595 660 -585 680
rect -565 660 -555 680
rect -595 640 -555 660
rect -595 620 -585 640
rect -565 620 -555 640
rect -595 600 -555 620
rect -595 580 -585 600
rect -565 580 -555 600
rect -595 565 -555 580
rect -520 680 -480 695
rect -520 660 -510 680
rect -490 660 -480 680
rect -520 640 -480 660
rect -520 620 -510 640
rect -490 620 -480 640
rect -520 600 -480 620
rect -520 580 -510 600
rect -490 580 -480 600
rect -520 570 -480 580
rect -735 540 -715 565
rect -645 540 -605 550
rect -1145 520 -755 540
rect -795 510 -755 520
rect -855 490 -815 500
rect -1145 470 -845 490
rect -825 470 -815 490
rect -795 490 -785 510
rect -765 490 -755 510
rect -795 480 -755 490
rect -735 520 -635 540
rect -615 520 -605 540
rect -855 460 -815 470
rect -1145 440 -870 450
rect -1145 430 -900 440
rect -910 420 -900 430
rect -880 420 -870 440
rect -910 410 -870 420
rect -1145 400 -1065 410
rect -1145 390 -1095 400
rect -1105 380 -1095 390
rect -1075 380 -1065 400
rect -1105 370 -1065 380
rect -1035 350 -995 360
rect -1145 330 -1025 350
rect -1005 330 -995 350
rect -1035 320 -995 330
rect -960 310 -920 320
rect -960 300 -950 310
rect -1145 290 -950 300
rect -930 290 -920 310
rect -735 290 -715 520
rect -645 510 -605 520
rect -695 480 -655 490
rect -585 480 -565 565
rect -445 540 -405 550
rect -445 520 -435 540
rect -415 520 -155 540
rect -445 510 -405 520
rect -695 460 -685 480
rect -665 460 -155 480
rect -695 450 -655 460
rect -585 290 -565 460
rect -515 430 -475 440
rect -255 430 -215 440
rect -515 410 -505 430
rect -485 410 -245 430
rect -225 410 -215 430
rect -515 400 -475 410
rect -255 400 -215 410
rect -460 380 -420 390
rect -330 380 -290 390
rect -460 360 -450 380
rect -430 360 -320 380
rect -300 360 -290 380
rect -460 350 -420 360
rect -330 350 -290 360
rect -405 330 -365 340
rect -405 310 -395 330
rect -375 310 -365 330
rect -405 300 -365 310
rect -1145 280 -920 290
rect -890 270 -705 290
rect -890 250 -870 270
rect -1135 235 -1095 250
rect -1135 215 -1125 235
rect -1105 215 -1095 235
rect -1135 195 -1095 215
rect -1135 175 -1125 195
rect -1105 175 -1095 195
rect -1135 155 -1095 175
rect -1135 135 -1125 155
rect -1105 135 -1095 155
rect -1135 125 -1095 135
rect -910 235 -870 250
rect -910 215 -900 235
rect -880 215 -870 235
rect -910 195 -870 215
rect -910 175 -900 195
rect -880 175 -870 195
rect -910 155 -870 175
rect -910 135 -900 155
rect -880 135 -870 155
rect -910 125 -870 135
rect -820 235 -780 250
rect -820 215 -810 235
rect -790 215 -780 235
rect -820 195 -780 215
rect -820 175 -810 195
rect -790 175 -780 195
rect -820 155 -780 175
rect -820 135 -810 155
rect -790 135 -780 155
rect -820 125 -780 135
rect -745 235 -705 270
rect -595 270 -440 290
rect -745 215 -735 235
rect -715 215 -705 235
rect -745 195 -705 215
rect -745 175 -735 195
rect -715 175 -705 195
rect -745 155 -705 175
rect -745 135 -735 155
rect -715 135 -705 155
rect -745 125 -705 135
rect -670 235 -630 250
rect -670 215 -660 235
rect -640 215 -630 235
rect -670 195 -630 215
rect -670 175 -660 195
rect -640 175 -630 195
rect -670 155 -630 175
rect -670 135 -660 155
rect -640 135 -630 155
rect -670 125 -630 135
rect -595 235 -555 270
rect -460 250 -440 270
rect -595 215 -585 235
rect -565 215 -555 235
rect -595 195 -555 215
rect -595 175 -585 195
rect -565 175 -555 195
rect -595 155 -555 175
rect -595 135 -585 155
rect -565 135 -555 155
rect -595 125 -555 135
rect -520 235 -480 250
rect -520 215 -510 235
rect -490 215 -480 235
rect -460 235 -390 250
rect -460 225 -420 235
rect -520 195 -480 215
rect -520 175 -510 195
rect -490 175 -480 195
rect -520 155 -480 175
rect -520 135 -510 155
rect -490 135 -480 155
rect -520 125 -480 135
rect -430 215 -420 225
rect -400 215 -390 235
rect -430 195 -390 215
rect -430 175 -420 195
rect -400 175 -390 195
rect -430 155 -390 175
rect -430 135 -420 155
rect -400 135 -390 155
rect -430 125 -390 135
rect -355 235 -315 250
rect -355 215 -345 235
rect -325 215 -315 235
rect -355 195 -315 215
rect -355 175 -345 195
rect -325 175 -315 195
rect -355 155 -315 175
rect -355 135 -345 155
rect -325 135 -315 155
rect -355 125 -315 135
rect -280 235 -240 250
rect -280 215 -270 235
rect -250 215 -240 235
rect -280 195 -240 215
rect -280 175 -270 195
rect -250 175 -240 195
rect -280 155 -240 175
rect -280 135 -270 155
rect -250 135 -240 155
rect -280 125 -240 135
rect -205 235 -165 250
rect -205 215 -195 235
rect -175 215 -165 235
rect -205 195 -165 215
rect -205 175 -195 195
rect -175 175 -165 195
rect -205 155 -165 175
rect -205 135 -195 155
rect -175 135 -165 155
rect -205 125 -165 135
rect -420 105 -400 125
rect -270 105 -250 125
rect -770 95 -730 105
rect -570 95 -530 105
rect -1145 75 -760 95
rect -740 75 -560 95
rect -540 75 -530 95
rect -420 85 -250 105
rect -770 65 -730 75
rect -570 65 -530 75
rect -1150 35 -150 45
rect -1150 15 -1140 35
rect -1120 15 -1100 35
rect -1080 15 -1060 35
rect -1040 15 -1020 35
rect -1000 15 -980 35
rect -960 15 -940 35
rect -920 15 -900 35
rect -880 15 -860 35
rect -840 15 -820 35
rect -800 15 -780 35
rect -760 15 -740 35
rect -720 15 -700 35
rect -680 15 -660 35
rect -640 15 -620 35
rect -600 15 -580 35
rect -560 15 -540 35
rect -520 15 -500 35
rect -480 15 -460 35
rect -440 15 -420 35
rect -400 15 -380 35
rect -360 15 -340 35
rect -320 15 -300 35
rect -280 15 -260 35
rect -240 15 -220 35
rect -200 15 -180 35
rect -160 15 -150 35
rect -1150 5 -150 15
<< viali >>
rect -1140 770 -1120 790
rect -1100 770 -1080 790
rect -1060 770 -1040 790
rect -1020 770 -1000 790
rect -980 770 -960 790
rect -940 770 -920 790
rect -900 770 -880 790
rect -860 770 -840 790
rect -820 770 -800 790
rect -780 770 -760 790
rect -740 770 -720 790
rect -700 770 -680 790
rect -660 770 -640 790
rect -620 770 -600 790
rect -580 770 -560 790
rect -540 770 -520 790
rect -500 770 -480 790
rect -460 770 -440 790
rect -420 770 -400 790
rect -380 770 -360 790
rect -340 770 -320 790
rect -300 770 -280 790
rect -260 770 -240 790
rect -220 770 -200 790
rect -180 770 -160 790
rect -810 660 -790 680
rect -810 620 -790 640
rect -810 580 -790 600
rect -660 660 -640 680
rect -660 620 -640 640
rect -660 580 -640 600
rect -510 660 -490 680
rect -510 620 -490 640
rect -510 580 -490 600
rect -845 470 -825 490
rect -785 490 -765 510
rect -635 520 -615 540
rect -900 420 -880 440
rect -435 520 -415 540
rect -505 410 -485 430
rect -450 360 -430 380
rect -395 310 -375 330
rect -1125 215 -1105 235
rect -1125 175 -1105 195
rect -1125 135 -1105 155
rect -810 215 -790 235
rect -810 175 -790 195
rect -810 135 -790 155
rect -660 215 -640 235
rect -660 175 -640 195
rect -660 135 -640 155
rect -510 215 -490 235
rect -510 175 -490 195
rect -510 135 -490 155
rect -345 215 -325 235
rect -345 175 -325 195
rect -345 135 -325 155
rect -195 215 -175 235
rect -195 175 -175 195
rect -195 135 -175 155
rect -1140 15 -1120 35
rect -1100 15 -1080 35
rect -1060 15 -1040 35
rect -1020 15 -1000 35
rect -980 15 -960 35
rect -940 15 -920 35
rect -900 15 -880 35
rect -860 15 -840 35
rect -820 15 -800 35
rect -780 15 -760 35
rect -740 15 -720 35
rect -700 15 -680 35
rect -660 15 -640 35
rect -620 15 -600 35
rect -580 15 -560 35
rect -540 15 -520 35
rect -500 15 -480 35
rect -460 15 -440 35
rect -420 15 -400 35
rect -380 15 -360 35
rect -340 15 -320 35
rect -300 15 -280 35
rect -260 15 -240 35
rect -220 15 -200 35
rect -180 15 -160 35
<< metal1 >>
rect -1150 790 -150 805
rect -1150 770 -1140 790
rect -1120 770 -1100 790
rect -1080 770 -1060 790
rect -1040 770 -1020 790
rect -1000 770 -980 790
rect -960 770 -940 790
rect -920 770 -900 790
rect -880 770 -860 790
rect -840 770 -820 790
rect -800 770 -780 790
rect -760 770 -740 790
rect -720 770 -700 790
rect -680 770 -660 790
rect -640 770 -620 790
rect -600 770 -580 790
rect -560 770 -540 790
rect -520 770 -500 790
rect -480 770 -460 790
rect -440 770 -420 790
rect -400 770 -380 790
rect -360 770 -340 790
rect -320 770 -300 790
rect -280 770 -260 790
rect -240 770 -220 790
rect -200 770 -180 790
rect -160 770 -150 790
rect -1150 755 -150 770
rect -1125 250 -1105 755
rect -820 680 -780 755
rect -820 660 -810 680
rect -790 660 -780 680
rect -820 640 -780 660
rect -820 620 -810 640
rect -790 620 -780 640
rect -820 600 -780 620
rect -820 580 -810 600
rect -790 580 -780 600
rect -820 570 -780 580
rect -670 680 -630 755
rect -670 660 -660 680
rect -640 660 -630 680
rect -670 640 -630 660
rect -670 620 -660 640
rect -640 620 -630 640
rect -670 600 -630 620
rect -670 580 -660 600
rect -640 580 -630 600
rect -670 570 -630 580
rect -520 680 -480 755
rect -520 660 -510 680
rect -490 660 -480 680
rect -520 640 -480 660
rect -520 620 -510 640
rect -490 620 -480 640
rect -520 600 -480 620
rect -520 580 -510 600
rect -490 580 -480 600
rect -520 570 -480 580
rect -645 540 -605 550
rect -445 540 -405 550
rect -645 520 -635 540
rect -615 520 -435 540
rect -415 520 -405 540
rect -795 510 -755 520
rect -645 510 -605 520
rect -445 510 -405 520
rect -855 490 -815 500
rect -855 470 -845 490
rect -825 470 -815 490
rect -795 490 -785 510
rect -765 490 -755 510
rect -795 480 -755 490
rect -855 460 -815 470
rect -910 440 -870 450
rect -910 420 -900 440
rect -880 420 -870 440
rect -910 410 -870 420
rect -900 330 -880 410
rect -845 380 -825 460
rect -785 430 -765 480
rect -515 430 -475 440
rect -785 410 -505 430
rect -485 410 -475 430
rect -515 400 -475 410
rect -460 380 -420 390
rect -845 360 -450 380
rect -430 360 -420 380
rect -460 350 -420 360
rect -405 330 -365 340
rect -900 310 -395 330
rect -375 310 -365 330
rect -405 300 -365 310
rect -345 250 -325 755
rect -195 250 -175 755
rect -1135 235 -1095 250
rect -1135 215 -1125 235
rect -1105 215 -1095 235
rect -1135 195 -1095 215
rect -1135 175 -1125 195
rect -1105 175 -1095 195
rect -1135 155 -1095 175
rect -1135 135 -1125 155
rect -1105 135 -1095 155
rect -1135 125 -1095 135
rect -820 235 -780 250
rect -820 215 -810 235
rect -790 215 -780 235
rect -820 195 -780 215
rect -820 175 -810 195
rect -790 175 -780 195
rect -820 155 -780 175
rect -820 135 -810 155
rect -790 135 -780 155
rect -820 125 -780 135
rect -670 235 -630 250
rect -670 215 -660 235
rect -640 215 -630 235
rect -670 195 -630 215
rect -670 175 -660 195
rect -640 175 -630 195
rect -670 155 -630 175
rect -670 135 -660 155
rect -640 135 -630 155
rect -670 125 -630 135
rect -520 235 -480 250
rect -520 215 -510 235
rect -490 215 -480 235
rect -520 195 -480 215
rect -520 175 -510 195
rect -490 175 -480 195
rect -520 155 -480 175
rect -520 135 -510 155
rect -490 135 -480 155
rect -520 125 -480 135
rect -355 235 -315 250
rect -355 215 -345 235
rect -325 215 -315 235
rect -355 195 -315 215
rect -355 175 -345 195
rect -325 175 -315 195
rect -355 155 -315 175
rect -355 135 -345 155
rect -325 135 -315 155
rect -355 125 -315 135
rect -205 235 -165 250
rect -205 215 -195 235
rect -175 215 -165 235
rect -205 195 -165 215
rect -205 175 -195 195
rect -175 175 -165 195
rect -205 155 -165 175
rect -205 135 -195 155
rect -175 135 -165 155
rect -205 125 -165 135
rect -810 50 -790 125
rect -660 50 -640 125
rect -510 50 -490 125
rect -1150 35 -150 50
rect -1150 15 -1140 35
rect -1120 15 -1100 35
rect -1080 15 -1060 35
rect -1040 15 -1020 35
rect -1000 15 -980 35
rect -960 15 -940 35
rect -920 15 -900 35
rect -880 15 -860 35
rect -840 15 -820 35
rect -800 15 -780 35
rect -760 15 -740 35
rect -720 15 -700 35
rect -680 15 -660 35
rect -640 15 -620 35
rect -600 15 -580 35
rect -560 15 -540 35
rect -520 15 -500 35
rect -480 15 -460 35
rect -440 15 -420 35
rect -400 15 -380 35
rect -360 15 -340 35
rect -320 15 -300 35
rect -280 15 -260 35
rect -240 15 -220 35
rect -200 15 -180 35
rect -160 15 -150 35
rect -1150 0 -150 15
<< labels >>
rlabel viali -635 520 -615 540 7 OUT_bar
port 8 w
rlabel locali -685 460 -665 480 7 OUT
port 7 w
rlabel metal1 -660 770 -640 790 7 CLK
port 11 w
rlabel locali -1140 525 -1130 535 7 A
port 1 w
rlabel locali -1140 475 -1130 485 7 B
port 3 w
rlabel locali -760 75 -740 95 7 Dis
port 9 w
rlabel locali -1140 395 -1130 405 7 A_bar
port 2 w
rlabel locali -1140 435 -1130 445 7 C
port 5 w
rlabel locali -1140 285 -1130 295 7 C_bar
port 6 w
rlabel locali -1140 335 -1130 345 7 B_bar
port 4 w
rlabel metal1 -660 15 -640 35 7 GND!
port 10 w
<< end >>
