magic
tech sky130A
timestamp 1666645976
<< nwell >>
rect -370 185 -25 530
<< nmos >>
rect -500 -70 -485 80
rect -275 -70 -260 80
rect -200 -70 -185 80
rect -125 -70 -110 80
rect -50 -70 -35 80
rect 175 -70 190 80
<< pmos >>
rect -200 210 -185 510
rect -125 210 -110 510
<< ndiff >>
rect -560 45 -500 80
rect -560 25 -540 45
rect -520 25 -500 45
rect -560 5 -500 25
rect -560 -15 -540 5
rect -520 -15 -500 5
rect -560 -35 -500 -15
rect -560 -55 -540 -35
rect -520 -55 -500 -35
rect -560 -70 -500 -55
rect -485 45 -425 80
rect -485 25 -465 45
rect -445 25 -425 45
rect -485 5 -425 25
rect -485 -15 -465 5
rect -445 -15 -425 5
rect -485 -35 -425 -15
rect -485 -55 -465 -35
rect -445 -55 -425 -35
rect -485 -70 -425 -55
rect -335 45 -275 80
rect -335 25 -315 45
rect -295 25 -275 45
rect -335 5 -275 25
rect -335 -15 -315 5
rect -295 -15 -275 5
rect -335 -35 -275 -15
rect -335 -55 -315 -35
rect -295 -55 -275 -35
rect -335 -70 -275 -55
rect -260 45 -200 80
rect -260 25 -240 45
rect -220 25 -200 45
rect -260 5 -200 25
rect -260 -15 -240 5
rect -220 -15 -200 5
rect -260 -35 -200 -15
rect -260 -55 -240 -35
rect -220 -55 -200 -35
rect -260 -70 -200 -55
rect -185 45 -125 80
rect -185 25 -165 45
rect -145 25 -125 45
rect -185 5 -125 25
rect -185 -15 -165 5
rect -145 -15 -125 5
rect -185 -35 -125 -15
rect -185 -55 -165 -35
rect -145 -55 -125 -35
rect -185 -70 -125 -55
rect -110 45 -50 80
rect -110 25 -90 45
rect -70 25 -50 45
rect -110 5 -50 25
rect -110 -15 -90 5
rect -70 -15 -50 5
rect -110 -35 -50 -15
rect -110 -55 -90 -35
rect -70 -55 -50 -35
rect -110 -70 -50 -55
rect -35 45 25 80
rect -35 25 -15 45
rect 5 25 25 45
rect -35 5 25 25
rect -35 -15 -15 5
rect 5 -15 25 5
rect -35 -35 25 -15
rect -35 -55 -15 -35
rect 5 -55 25 -35
rect -35 -70 25 -55
rect 115 45 175 80
rect 115 25 135 45
rect 155 25 175 45
rect 115 5 175 25
rect 115 -15 135 5
rect 155 -15 175 5
rect 115 -35 175 -15
rect 115 -55 135 -35
rect 155 -55 175 -35
rect 115 -70 175 -55
rect 190 45 250 80
rect 190 25 210 45
rect 230 25 250 45
rect 190 5 250 25
rect 190 -15 210 5
rect 230 -15 250 5
rect 190 -35 250 -15
rect 190 -55 210 -35
rect 230 -55 250 -35
rect 190 -70 250 -55
<< pdiff >>
rect -260 485 -200 510
rect -260 465 -240 485
rect -220 465 -200 485
rect -260 445 -200 465
rect -260 425 -240 445
rect -220 425 -200 445
rect -260 405 -200 425
rect -260 385 -240 405
rect -220 385 -200 405
rect -260 365 -200 385
rect -260 345 -240 365
rect -220 345 -200 365
rect -260 325 -200 345
rect -260 305 -240 325
rect -220 305 -200 325
rect -260 285 -200 305
rect -260 265 -240 285
rect -220 265 -200 285
rect -260 245 -200 265
rect -260 225 -240 245
rect -220 225 -200 245
rect -260 210 -200 225
rect -185 485 -125 510
rect -185 465 -165 485
rect -145 465 -125 485
rect -185 445 -125 465
rect -185 425 -165 445
rect -145 425 -125 445
rect -185 405 -125 425
rect -185 385 -165 405
rect -145 385 -125 405
rect -185 365 -125 385
rect -185 345 -165 365
rect -145 345 -125 365
rect -185 325 -125 345
rect -185 305 -165 325
rect -145 305 -125 325
rect -185 285 -125 305
rect -185 265 -165 285
rect -145 265 -125 285
rect -185 245 -125 265
rect -185 225 -165 245
rect -145 225 -125 245
rect -185 210 -125 225
rect -110 485 -50 510
rect -110 465 -90 485
rect -70 465 -50 485
rect -110 445 -50 465
rect -110 425 -90 445
rect -70 425 -50 445
rect -110 405 -50 425
rect -110 385 -90 405
rect -70 385 -50 405
rect -110 365 -50 385
rect -110 345 -90 365
rect -70 345 -50 365
rect -110 325 -50 345
rect -110 305 -90 325
rect -70 305 -50 325
rect -110 285 -50 305
rect -110 265 -90 285
rect -70 265 -50 285
rect -110 245 -50 265
rect -110 225 -90 245
rect -70 225 -50 245
rect -110 210 -50 225
<< ndiffc >>
rect -540 25 -520 45
rect -540 -15 -520 5
rect -540 -55 -520 -35
rect -465 25 -445 45
rect -465 -15 -445 5
rect -465 -55 -445 -35
rect -315 25 -295 45
rect -315 -15 -295 5
rect -315 -55 -295 -35
rect -240 25 -220 45
rect -240 -15 -220 5
rect -240 -55 -220 -35
rect -165 25 -145 45
rect -165 -15 -145 5
rect -165 -55 -145 -35
rect -90 25 -70 45
rect -90 -15 -70 5
rect -90 -55 -70 -35
rect -15 25 5 45
rect -15 -15 5 5
rect -15 -55 5 -35
rect 135 25 155 45
rect 135 -15 155 5
rect 135 -55 155 -35
rect 210 25 230 45
rect 210 -15 230 5
rect 210 -55 230 -35
<< pdiffc >>
rect -240 465 -220 485
rect -240 425 -220 445
rect -240 385 -220 405
rect -240 345 -220 365
rect -240 305 -220 325
rect -240 265 -220 285
rect -240 225 -220 245
rect -165 465 -145 485
rect -165 425 -145 445
rect -165 385 -145 405
rect -165 345 -145 365
rect -165 305 -145 325
rect -165 265 -145 285
rect -165 225 -145 245
rect -90 465 -70 485
rect -90 425 -70 445
rect -90 385 -70 405
rect -90 345 -70 365
rect -90 305 -70 325
rect -90 265 -70 285
rect -90 225 -70 245
<< psubdiff >>
rect -620 45 -560 80
rect -620 25 -600 45
rect -580 25 -560 45
rect -620 5 -560 25
rect -620 -15 -600 5
rect -580 -15 -560 5
rect -620 -35 -560 -15
rect -620 -55 -600 -35
rect -580 -55 -560 -35
rect -620 -70 -560 -55
rect -395 45 -335 80
rect -395 25 -375 45
rect -355 25 -335 45
rect -395 5 -335 25
rect -395 -15 -375 5
rect -355 -15 -335 5
rect -395 -35 -335 -15
rect -395 -55 -375 -35
rect -355 -55 -335 -35
rect -395 -70 -335 -55
rect 55 45 115 80
rect 55 25 75 45
rect 95 25 115 45
rect 55 5 115 25
rect 55 -15 75 5
rect 95 -15 115 5
rect 55 -35 115 -15
rect 55 -55 75 -35
rect 95 -55 115 -35
rect 55 -70 115 -55
<< nsubdiff >>
rect -350 485 -290 510
rect -350 465 -330 485
rect -310 465 -290 485
rect -350 445 -290 465
rect -350 425 -330 445
rect -310 425 -290 445
rect -350 405 -290 425
rect -350 385 -330 405
rect -310 385 -290 405
rect -350 365 -290 385
rect -350 345 -330 365
rect -310 345 -290 365
rect -350 325 -290 345
rect -350 305 -330 325
rect -310 305 -290 325
rect -350 285 -290 305
rect -350 265 -330 285
rect -310 265 -290 285
rect -350 245 -290 265
rect -350 225 -330 245
rect -310 225 -290 245
rect -350 210 -290 225
<< psubdiffcont >>
rect -600 25 -580 45
rect -600 -15 -580 5
rect -600 -55 -580 -35
rect -375 25 -355 45
rect -375 -15 -355 5
rect -375 -55 -355 -35
rect 75 25 95 45
rect 75 -15 95 5
rect 75 -55 95 -35
<< nsubdiffcont >>
rect -330 465 -310 485
rect -330 425 -310 445
rect -330 385 -310 405
rect -330 345 -310 365
rect -330 305 -310 325
rect -330 265 -310 285
rect -330 225 -310 245
<< poly >>
rect 160 675 200 685
rect 160 655 170 675
rect 190 655 200 675
rect 160 645 200 655
rect -515 620 -475 630
rect -515 600 -505 620
rect -485 600 -475 620
rect -515 590 -475 600
rect -500 80 -485 590
rect -200 510 -185 525
rect -125 510 -110 525
rect -200 135 -185 210
rect -125 195 -110 210
rect -150 185 -110 195
rect -150 165 -140 185
rect -120 165 -110 185
rect -150 155 -110 165
rect -200 125 -160 135
rect -200 105 -190 125
rect -170 105 -160 125
rect -200 95 -160 105
rect -275 80 -260 95
rect -200 80 -185 95
rect -125 80 -110 155
rect -50 80 -35 95
rect 175 80 190 645
rect -500 -250 -485 -70
rect -275 -110 -260 -70
rect -200 -85 -185 -70
rect -125 -85 -110 -70
rect -50 -110 -35 -70
rect -275 -125 -35 -110
rect -275 -200 -255 -125
rect -285 -210 -245 -200
rect -285 -230 -275 -210
rect -255 -230 -245 -210
rect -285 -240 -245 -230
rect -515 -260 -475 -250
rect -515 -280 -505 -260
rect -485 -280 -475 -260
rect -515 -290 -475 -280
rect 175 -300 190 -70
rect 160 -310 200 -300
rect 160 -330 170 -310
rect 190 -330 200 -310
rect 160 -340 200 -330
<< polycont >>
rect 170 655 190 675
rect -505 600 -485 620
rect -140 165 -120 185
rect -190 105 -170 125
rect -275 -230 -255 -210
rect -505 -280 -485 -260
rect 170 -330 190 -310
<< locali >>
rect -90 775 -50 785
rect -620 755 -80 775
rect -60 755 250 775
rect -90 745 -50 755
rect -260 725 -220 735
rect -620 705 -250 725
rect -230 705 250 725
rect -260 695 -220 705
rect 160 675 200 685
rect -620 655 170 675
rect 190 655 250 675
rect 160 645 200 655
rect -515 620 -475 630
rect -620 600 -505 620
rect -485 600 250 620
rect -515 590 -475 600
rect -340 485 -300 495
rect -340 465 -330 485
rect -310 465 -300 485
rect -340 445 -300 465
rect -340 425 -330 445
rect -310 425 -300 445
rect -340 405 -300 425
rect -340 385 -330 405
rect -310 385 -300 405
rect -340 365 -300 385
rect -340 345 -330 365
rect -310 345 -300 365
rect -340 325 -300 345
rect -340 305 -330 325
rect -310 305 -300 325
rect -340 285 -300 305
rect -340 265 -330 285
rect -310 265 -300 285
rect -340 245 -300 265
rect -340 225 -330 245
rect -310 225 -300 245
rect -340 215 -300 225
rect -250 485 -210 495
rect -250 465 -240 485
rect -220 465 -210 485
rect -250 445 -210 465
rect -250 425 -240 445
rect -220 425 -210 445
rect -250 405 -210 425
rect -250 385 -240 405
rect -220 385 -210 405
rect -250 365 -210 385
rect -250 345 -240 365
rect -220 345 -210 365
rect -250 325 -210 345
rect -250 305 -240 325
rect -220 305 -210 325
rect -250 285 -210 305
rect -250 265 -240 285
rect -220 265 -210 285
rect -250 245 -210 265
rect -250 225 -240 245
rect -220 225 -210 245
rect -250 210 -210 225
rect -175 485 -135 495
rect -175 465 -165 485
rect -145 465 -135 485
rect -175 445 -135 465
rect -175 425 -165 445
rect -145 425 -135 445
rect -175 405 -135 425
rect -175 385 -165 405
rect -145 385 -135 405
rect -175 365 -135 385
rect -175 345 -165 365
rect -145 345 -135 365
rect -175 325 -135 345
rect -175 305 -165 325
rect -145 305 -135 325
rect -175 285 -135 305
rect -175 265 -165 285
rect -145 265 -135 285
rect -175 245 -135 265
rect -175 225 -165 245
rect -145 225 -135 245
rect -175 215 -135 225
rect -100 485 -60 495
rect -100 465 -90 485
rect -70 465 -60 485
rect -100 445 -60 465
rect -100 425 -90 445
rect -70 425 -60 445
rect -100 405 -60 425
rect -100 385 -90 405
rect -70 385 -60 405
rect -100 365 -60 385
rect -100 345 -90 365
rect -70 345 -60 365
rect -100 325 -60 345
rect -100 305 -90 325
rect -70 305 -60 325
rect -100 285 -60 305
rect -100 265 -90 285
rect -70 265 -60 285
rect -100 245 -60 265
rect -100 225 -90 245
rect -70 225 -60 245
rect -100 210 -60 225
rect -250 185 -220 210
rect -150 185 -110 195
rect -250 165 -140 185
rect -120 165 -110 185
rect -250 140 -220 165
rect -150 155 -110 165
rect -465 130 -220 140
rect -90 145 -60 210
rect -90 135 230 145
rect -465 110 -250 130
rect -230 110 -220 130
rect -465 100 -220 110
rect -465 60 -435 100
rect -240 80 -220 100
rect -200 125 -160 135
rect -90 125 -80 135
rect -200 105 -190 125
rect -170 115 -80 125
rect -60 115 230 135
rect -170 105 230 115
rect -200 95 -160 105
rect -90 80 -70 105
rect -610 45 -570 60
rect -610 25 -600 45
rect -580 25 -570 45
rect -610 5 -570 25
rect -610 -15 -600 5
rect -580 -15 -570 5
rect -610 -35 -570 -15
rect -610 -55 -600 -35
rect -580 -55 -570 -35
rect -610 -65 -570 -55
rect -550 45 -510 60
rect -550 25 -540 45
rect -520 25 -510 45
rect -550 5 -510 25
rect -550 -15 -540 5
rect -520 -15 -510 5
rect -550 -35 -510 -15
rect -550 -55 -540 -35
rect -520 -55 -510 -35
rect -550 -65 -510 -55
rect -475 45 -435 60
rect -475 25 -465 45
rect -445 25 -435 45
rect -475 5 -435 25
rect -475 -15 -465 5
rect -445 -15 -435 5
rect -475 -35 -435 -15
rect -475 -55 -465 -35
rect -445 -55 -435 -35
rect -475 -65 -435 -55
rect -385 45 -345 60
rect -385 25 -375 45
rect -355 25 -345 45
rect -385 5 -345 25
rect -385 -15 -375 5
rect -355 -15 -345 5
rect -385 -35 -345 -15
rect -385 -55 -375 -35
rect -355 -55 -345 -35
rect -385 -65 -345 -55
rect -325 45 -285 60
rect -325 25 -315 45
rect -295 25 -285 45
rect -325 5 -285 25
rect -325 -15 -315 5
rect -295 -15 -285 5
rect -325 -35 -285 -15
rect -325 -55 -315 -35
rect -295 -55 -285 -35
rect -325 -65 -285 -55
rect -250 45 -210 80
rect -250 25 -240 45
rect -220 25 -210 45
rect -250 5 -210 25
rect -250 -15 -240 5
rect -220 -15 -210 5
rect -250 -35 -210 -15
rect -250 -55 -240 -35
rect -220 -55 -210 -35
rect -250 -65 -210 -55
rect -175 45 -135 60
rect -175 25 -165 45
rect -145 25 -135 45
rect -175 5 -135 25
rect -175 -15 -165 5
rect -145 -15 -135 5
rect -175 -35 -135 -15
rect -175 -55 -165 -35
rect -145 -55 -135 -35
rect -175 -65 -135 -55
rect -100 45 -60 80
rect 200 60 230 105
rect -100 25 -90 45
rect -70 25 -60 45
rect -100 5 -60 25
rect -100 -15 -90 5
rect -70 -15 -60 5
rect -100 -35 -60 -15
rect -100 -55 -90 -35
rect -70 -55 -60 -35
rect -100 -65 -60 -55
rect -25 45 15 60
rect -25 25 -15 45
rect 5 25 15 45
rect -25 5 15 25
rect -25 -15 -15 5
rect 5 -15 15 5
rect -25 -35 15 -15
rect -25 -55 -15 -35
rect 5 -55 15 -35
rect -25 -65 15 -55
rect 65 45 105 60
rect 65 25 75 45
rect 95 25 105 45
rect 65 5 105 25
rect 65 -15 75 5
rect 95 -15 105 5
rect 65 -35 105 -15
rect 65 -55 75 -35
rect 95 -55 105 -35
rect 65 -65 105 -55
rect 125 45 165 60
rect 125 25 135 45
rect 155 25 165 45
rect 125 5 165 25
rect 125 -15 135 5
rect 155 -15 165 5
rect 125 -35 165 -15
rect 125 -55 135 -35
rect 155 -55 165 -35
rect 125 -65 165 -55
rect 200 45 240 60
rect 200 25 210 45
rect 230 25 240 45
rect 200 5 240 25
rect 200 -15 210 5
rect 230 -15 240 5
rect 200 -35 240 -15
rect 200 -55 210 -35
rect 230 -55 240 -35
rect 200 -65 240 -55
rect -285 -210 -245 -200
rect -620 -230 -275 -210
rect -255 -230 250 -210
rect -285 -240 -245 -230
rect -515 -260 -475 -250
rect -620 -280 -505 -260
rect -485 -280 250 -260
rect -515 -290 -475 -280
rect 160 -310 200 -300
rect -620 -330 170 -310
rect 190 -330 250 -310
rect 160 -340 200 -330
rect -260 -360 -220 -350
rect -620 -380 -250 -360
rect -230 -380 250 -360
rect -260 -390 -220 -380
rect -90 -410 -50 -400
rect -620 -430 -80 -410
rect -60 -430 250 -410
rect -90 -440 -50 -430
<< viali >>
rect -80 755 -60 775
rect -250 705 -230 725
rect -330 465 -310 485
rect -330 425 -310 445
rect -330 385 -310 405
rect -330 345 -310 365
rect -330 305 -310 325
rect -330 265 -310 285
rect -330 225 -310 245
rect -165 465 -145 485
rect -165 425 -145 445
rect -165 385 -145 405
rect -165 345 -145 365
rect -165 305 -145 325
rect -165 265 -145 285
rect -165 225 -145 245
rect -250 110 -230 130
rect -80 115 -60 135
rect -600 25 -580 45
rect -600 -15 -580 5
rect -600 -55 -580 -35
rect -540 25 -520 45
rect -540 -15 -520 5
rect -540 -55 -520 -35
rect -375 25 -355 45
rect -375 -15 -355 5
rect -375 -55 -355 -35
rect -315 25 -295 45
rect -315 -15 -295 5
rect -315 -55 -295 -35
rect -165 25 -145 45
rect -165 -15 -145 5
rect -165 -55 -145 -35
rect -15 25 5 45
rect -15 -15 5 5
rect -15 -55 5 -35
rect 75 25 95 45
rect 75 -15 95 5
rect 75 -55 95 -35
rect 135 25 155 45
rect 135 -15 155 5
rect 135 -55 155 -35
rect -250 -380 -230 -360
rect -80 -430 -60 -410
<< metal1 >>
rect -90 780 -50 785
rect -90 750 -85 780
rect -55 750 -50 780
rect -90 745 -50 750
rect -260 730 -220 735
rect -260 700 -255 730
rect -225 700 -220 730
rect -260 695 -220 700
rect -620 540 250 590
rect -340 485 -300 540
rect -340 465 -330 485
rect -310 465 -300 485
rect -340 445 -300 465
rect -340 425 -330 445
rect -310 425 -300 445
rect -340 405 -300 425
rect -340 385 -330 405
rect -310 385 -300 405
rect -340 365 -300 385
rect -340 345 -330 365
rect -310 345 -300 365
rect -340 325 -300 345
rect -340 305 -330 325
rect -310 305 -300 325
rect -340 285 -300 305
rect -340 265 -330 285
rect -310 265 -300 285
rect -340 245 -300 265
rect -340 225 -330 245
rect -310 225 -300 245
rect -340 215 -300 225
rect -175 485 -135 540
rect -175 465 -165 485
rect -145 465 -135 485
rect -175 445 -135 465
rect -175 425 -165 445
rect -145 425 -135 445
rect -175 405 -135 425
rect -175 385 -165 405
rect -145 385 -135 405
rect -175 365 -135 385
rect -175 345 -165 365
rect -145 345 -135 365
rect -175 325 -135 345
rect -175 305 -165 325
rect -145 305 -135 325
rect -175 285 -135 305
rect -175 265 -165 285
rect -145 265 -135 285
rect -175 245 -135 265
rect -175 225 -165 245
rect -145 225 -135 245
rect -175 215 -135 225
rect -90 140 -50 145
rect -260 135 -220 140
rect -260 105 -255 135
rect -225 105 -220 135
rect -90 110 -85 140
rect -55 110 -50 140
rect -90 105 -50 110
rect -260 100 -220 105
rect -610 45 -510 60
rect -610 25 -600 45
rect -580 25 -540 45
rect -520 25 -510 45
rect -610 5 -510 25
rect -610 -15 -600 5
rect -580 -15 -540 5
rect -520 -15 -510 5
rect -610 -35 -510 -15
rect -610 -55 -600 -35
rect -580 -55 -540 -35
rect -520 -55 -510 -35
rect -610 -135 -510 -55
rect -385 45 -285 60
rect -385 25 -375 45
rect -355 25 -315 45
rect -295 25 -285 45
rect -385 5 -285 25
rect -385 -15 -375 5
rect -355 -15 -315 5
rect -295 -15 -285 5
rect -385 -35 -285 -15
rect -385 -55 -375 -35
rect -355 -55 -315 -35
rect -295 -55 -285 -35
rect -385 -135 -285 -55
rect -175 45 -135 60
rect -175 25 -165 45
rect -145 25 -135 45
rect -175 5 -135 25
rect -175 -15 -165 5
rect -145 -15 -135 5
rect -175 -35 -135 -15
rect -175 -55 -165 -35
rect -145 -55 -135 -35
rect -175 -135 -135 -55
rect -25 45 15 60
rect -25 25 -15 45
rect 5 25 15 45
rect -25 5 15 25
rect -25 -15 -15 5
rect 5 -15 15 5
rect -25 -35 15 -15
rect -25 -55 -15 -35
rect 5 -55 15 -35
rect -25 -135 15 -55
rect 65 45 165 60
rect 65 25 75 45
rect 95 25 135 45
rect 155 25 165 45
rect 65 5 165 25
rect 65 -15 75 5
rect 95 -15 135 5
rect 155 -15 165 5
rect 65 -35 165 -15
rect 65 -55 75 -35
rect 95 -55 135 -35
rect 155 -55 165 -35
rect 65 -135 165 -55
rect -620 -185 250 -135
rect -260 -355 -220 -350
rect -260 -385 -255 -355
rect -225 -385 -220 -355
rect -260 -390 -220 -385
rect -90 -405 -50 -400
rect -90 -435 -85 -405
rect -55 -435 -50 -405
rect -90 -440 -50 -435
<< via1 >>
rect -85 775 -55 780
rect -85 755 -80 775
rect -80 755 -60 775
rect -60 755 -55 775
rect -85 750 -55 755
rect -255 725 -225 730
rect -255 705 -250 725
rect -250 705 -230 725
rect -230 705 -225 725
rect -255 700 -225 705
rect -255 130 -225 135
rect -255 110 -250 130
rect -250 110 -230 130
rect -230 110 -225 130
rect -255 105 -225 110
rect -85 135 -55 140
rect -85 115 -80 135
rect -80 115 -60 135
rect -60 115 -55 135
rect -85 110 -55 115
rect -255 -360 -225 -355
rect -255 -380 -250 -360
rect -250 -380 -230 -360
rect -230 -380 -225 -360
rect -255 -385 -225 -380
rect -85 -410 -55 -405
rect -85 -430 -80 -410
rect -80 -430 -60 -410
rect -60 -430 -55 -410
rect -85 -435 -55 -430
<< metal2 >>
rect -90 780 -50 785
rect -90 750 -85 780
rect -55 750 -50 780
rect -260 730 -220 735
rect -260 700 -255 730
rect -225 700 -220 730
rect -260 135 -220 700
rect -260 105 -255 135
rect -225 105 -220 135
rect -260 -355 -220 105
rect -260 -385 -255 -355
rect -225 -385 -220 -355
rect -260 -390 -220 -385
rect -90 140 -50 750
rect -90 110 -85 140
rect -55 110 -50 140
rect -90 -405 -50 110
rect -90 -435 -85 -405
rect -55 -435 -50 -405
rect -90 -440 -50 -435
<< labels >>
rlabel metal1 -165 -170 -145 -150 7 GND
rlabel metal1 -165 550 -145 570 7 CLK
rlabel metal2 -250 110 -230 130 7 OUT
rlabel metal2 -80 115 -60 135 7 OUT_bar
rlabel locali -505 -280 -485 -260 7 A_bar
rlabel locali 170 -330 190 -310 7 A
<< end >>
