magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -302 -271 302 271
<< l67d20 >>
rect -256 35 -221 251
rect -97 35 -62 251
rect 62 35 97 251
rect 221 35 256 251
rect -256 -251 -221 -35
rect -97 -251 -62 -35
rect 62 -251 97 -35
rect 221 -251 256 -35
<< l66d20 >>
rect -256 -251 -221 251
rect -97 -251 -62 251
rect 62 -251 97 251
rect 221 -251 256 251
<< l66d44 >>
rect -247 44 -230 61
rect -247 44 -230 61
rect 230 224 247 241
rect 230 188 247 205
rect -247 -241 -230 -224
rect -247 -241 -230 -224
rect 230 -61 247 -44
rect 230 -97 247 -80
rect -247 -205 -230 -188
rect -247 -169 -230 -152
rect -247 -133 -230 -116
rect -247 -97 -230 -80
rect -247 -61 -230 -44
rect -247 -205 -230 -188
rect -247 -169 -230 -152
rect -247 -133 -230 -116
rect -247 -97 -230 -80
rect -247 -61 -230 -44
rect -88 -61 -71 -44
rect -88 -97 -71 -80
rect -88 -133 -71 -116
rect -88 -169 -71 -152
rect -88 -205 -71 -188
rect -88 -61 -71 -44
rect -88 -97 -71 -80
rect -88 -133 -71 -116
rect -88 -169 -71 -152
rect -88 -205 -71 -188
rect -88 -241 -71 -224
rect -88 -241 -71 -224
rect 71 -61 88 -44
rect 71 -97 88 -80
rect 71 -133 88 -116
rect 71 -169 88 -152
rect 71 -205 88 -188
rect 71 -61 88 -44
rect 71 -97 88 -80
rect 71 -133 88 -116
rect 71 -169 88 -152
rect 71 -205 88 -188
rect 71 -241 88 -224
rect 71 -241 88 -224
rect 230 -133 247 -116
rect 230 -169 247 -152
rect 230 -205 247 -188
rect 230 -61 247 -44
rect 230 -97 247 -80
rect 230 -133 247 -116
rect 230 -169 247 -152
rect 230 -205 247 -188
rect 230 -241 247 -224
rect 230 -241 247 -224
rect -247 80 -230 97
rect -247 116 -230 133
rect -247 152 -230 169
rect -247 188 -230 205
rect -247 224 -230 241
rect -247 80 -230 97
rect -247 116 -230 133
rect -247 152 -230 169
rect -247 188 -230 205
rect -247 224 -230 241
rect -88 224 -71 241
rect -88 188 -71 205
rect -88 152 -71 169
rect -88 116 -71 133
rect -88 80 -71 97
rect -88 224 -71 241
rect -88 188 -71 205
rect -88 152 -71 169
rect -88 116 -71 133
rect -88 80 -71 97
rect -88 44 -71 61
rect -88 44 -71 61
rect 71 224 88 241
rect 71 188 88 205
rect 71 152 88 169
rect 71 116 88 133
rect 71 80 88 97
rect 71 224 88 241
rect 71 188 88 205
rect 71 152 88 169
rect 71 116 88 133
rect 71 80 88 97
rect 71 44 88 61
rect 71 44 88 61
rect 230 152 247 169
rect 230 116 247 133
rect 230 80 247 97
rect 230 224 247 241
rect 230 188 247 205
rect 230 152 247 169
rect 230 116 247 133
rect 230 80 247 97
rect 230 44 247 61
rect 230 44 247 61
<< l94d20 >>
rect -267 -262 -210 262
rect -108 -262 -51 262
rect 51 -262 108 262
rect 210 -262 267 262
<< l67d44 >>
rect 71 224 88 241
rect 230 224 247 241
rect 71 188 88 205
rect 230 188 247 205
rect 71 152 88 169
rect 230 152 247 169
rect 71 116 88 133
rect 230 116 247 133
rect 71 80 88 97
rect 230 80 247 97
rect 71 44 88 61
rect 230 44 247 61
rect 71 224 88 241
rect 230 224 247 241
rect 71 188 88 205
rect 230 188 247 205
rect 71 152 88 169
rect 230 152 247 169
rect 71 116 88 133
rect 230 116 247 133
rect 71 80 88 97
rect 230 80 247 97
rect 71 44 88 61
rect 230 44 247 61
rect 71 44 88 61
rect 71 44 88 61
rect 71 80 88 97
rect 71 80 88 97
rect 71 116 88 133
rect 71 116 88 133
rect 71 152 88 169
rect 71 152 88 169
rect 71 188 88 205
rect 71 188 88 205
rect 71 224 88 241
rect 71 224 88 241
rect 230 224 247 241
rect 230 188 247 205
rect 230 152 247 169
rect 230 116 247 133
rect 230 80 247 97
rect 230 44 247 61
rect 230 44 247 61
rect 230 44 247 61
rect 230 80 247 97
rect 230 80 247 97
rect 230 116 247 133
rect 230 116 247 133
rect 230 152 247 169
rect 230 152 247 169
rect 230 188 247 205
rect 230 188 247 205
rect 230 224 247 241
rect 230 224 247 241
rect -88 152 -71 169
rect -88 152 -71 169
rect -88 188 -71 205
rect -88 188 -71 205
rect -88 224 -71 241
rect -88 224 -71 241
rect -247 224 -230 241
rect -247 224 -230 241
rect -247 116 -230 133
rect -88 116 -71 133
rect -247 188 -230 205
rect -247 188 -230 205
rect -247 224 -230 241
rect -88 224 -71 241
rect -247 152 -230 169
rect -247 152 -230 169
rect -247 80 -230 97
rect -88 80 -71 97
rect -247 116 -230 133
rect -247 116 -230 133
rect -247 152 -230 169
rect -88 152 -71 169
rect -247 80 -230 97
rect -247 80 -230 97
rect -247 44 -230 61
rect -88 44 -71 61
rect -247 44 -230 61
rect -247 44 -230 61
rect -247 188 -230 205
rect -88 188 -71 205
rect -88 44 -71 61
rect -88 44 -71 61
rect -88 80 -71 97
rect -88 80 -71 97
rect -88 116 -71 133
rect -88 116 -71 133
rect -88 -133 -71 -116
rect -88 -133 -71 -116
rect -88 -97 -71 -80
rect -88 -97 -71 -80
rect -88 -61 -71 -44
rect -88 -61 -71 -44
rect -247 -61 -230 -44
rect -247 -61 -230 -44
rect -247 -97 -230 -80
rect -247 -97 -230 -80
rect -247 -133 -230 -116
rect -247 -133 -230 -116
rect -247 -169 -230 -152
rect -247 -169 -230 -152
rect -247 -205 -230 -188
rect -247 -205 -230 -188
rect -247 -241 -230 -224
rect -247 -241 -230 -224
rect -88 -241 -71 -224
rect -88 -241 -71 -224
rect -88 -205 -71 -188
rect -88 -205 -71 -188
rect -88 -169 -71 -152
rect -88 -169 -71 -152
rect 230 -61 247 -44
rect 230 -97 247 -80
rect 230 -133 247 -116
rect 230 -169 247 -152
rect 230 -205 247 -188
rect 230 -241 247 -224
rect 230 -241 247 -224
rect 230 -241 247 -224
rect 230 -205 247 -188
rect 230 -205 247 -188
rect 230 -169 247 -152
rect 230 -169 247 -152
rect 230 -133 247 -116
rect 230 -133 247 -116
rect 230 -97 247 -80
rect 230 -97 247 -80
rect 230 -61 247 -44
rect 230 -61 247 -44
rect 71 -97 88 -80
rect 230 -97 247 -80
rect 71 -169 88 -152
rect 230 -169 247 -152
rect 71 -61 88 -44
rect 230 -61 247 -44
rect 71 -205 88 -188
rect 230 -205 247 -188
rect 71 -133 88 -116
rect 230 -133 247 -116
rect 71 -241 88 -224
rect 230 -241 247 -224
rect 71 -241 88 -224
rect 71 -241 88 -224
rect 71 -205 88 -188
rect 71 -205 88 -188
rect 71 -169 88 -152
rect 71 -169 88 -152
rect 71 -133 88 -116
rect 71 -133 88 -116
rect 71 -97 88 -80
rect 71 -97 88 -80
rect 71 -61 88 -44
rect 71 -61 88 -44
<< l68d20 >>
rect -251 37 -226 248
rect -92 37 -67 248
rect 67 37 92 248
rect 226 37 251 248
rect -251 -248 -226 -37
rect -92 -248 -67 -37
rect 67 -248 92 -37
rect 226 -248 251 -37
<< l79d20 >>
rect -302 -271 302 271
<< l95d20 >>
rect -266 -260 -212 260
rect -107 -260 -53 260
rect 53 -260 107 260
rect 212 -260 266 260
<< l66d13 >>
rect -256 -41 -221 41
rect -97 -41 -62 41
rect 62 -41 97 41
rect 221 -41 256 41
<< end >>
