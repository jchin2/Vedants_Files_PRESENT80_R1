magic
tech sky130A
magscale 1 2
timestamp 1673474122
<< locali >>
rect -446 3710 290 3750
rect 2570 3650 2650 3670
rect -445 3610 290 3650
rect 2570 3647 2910 3650
rect 2570 3613 2593 3647
rect 2627 3613 2910 3647
rect 2570 3610 2910 3613
rect 4578 3620 4658 3640
rect 4578 3617 4930 3620
rect 2570 3590 2650 3610
rect 4578 3583 4601 3617
rect 4635 3583 4930 3617
rect 4578 3580 4930 3583
rect 4578 3560 4658 3580
rect -446 3510 290 3550
rect 2780 3530 2860 3550
rect 2780 3527 2910 3530
rect 2780 3493 2803 3527
rect 2837 3493 2910 3527
rect 2780 3490 2910 3493
rect 4692 3504 4772 3527
rect 2780 3470 2860 3490
rect 4692 3470 4715 3504
rect 4749 3500 4772 3504
rect 4749 3470 4930 3500
rect 4692 3460 4930 3470
rect -445 3410 290 3450
rect 2660 3430 2740 3450
rect 4692 3447 4772 3460
rect 2530 3427 2910 3430
rect 2530 3393 2683 3427
rect 2717 3393 2910 3427
rect 2530 3390 2910 3393
rect 4820 3400 4900 3420
rect 4820 3397 4930 3400
rect 2530 3310 2570 3390
rect 2660 3370 2740 3390
rect 4590 3340 4732 3380
rect 4820 3363 4843 3397
rect 4877 3363 4930 3397
rect 4820 3360 4930 3363
rect 4820 3340 4900 3360
rect 6579 3349 6601 3372
rect 2740 3307 2820 3330
rect 2740 3273 2763 3307
rect 2797 3273 2820 3307
rect 2570 3247 2650 3270
rect 2570 3213 2593 3247
rect 2627 3213 2650 3247
rect 2570 3190 2650 3213
rect 2740 3250 2820 3273
rect 2860 3290 2910 3330
rect 4692 3300 4732 3340
rect 2740 3150 2780 3250
rect 2860 3210 2900 3290
rect 2610 3110 2780 3150
rect 2850 3170 2900 3210
rect 4578 3257 4658 3280
rect 4692 3260 4933 3300
rect 4578 3223 4601 3257
rect 4635 3223 4658 3257
rect 6580 3230 6600 3250
rect 4578 3200 4658 3223
rect 290 2817 370 2840
rect 290 2783 313 2817
rect 347 2783 370 2817
rect 290 2760 370 2783
rect 10 2697 290 2720
rect 10 2663 43 2697
rect 77 2663 290 2697
rect 10 2640 290 2663
rect 290 2580 370 2600
rect 2610 2580 2650 3110
rect 2850 3070 2890 3170
rect 290 2577 590 2580
rect 290 2543 313 2577
rect 347 2543 590 2577
rect 290 2540 590 2543
rect 2290 2540 2650 2580
rect 2750 3030 2890 3070
rect 4652 3123 4772 3146
rect 4652 3089 4715 3123
rect 4749 3089 4772 3123
rect 4652 3066 4772 3089
rect 290 2520 370 2540
rect 2290 2140 2330 2540
rect 2750 2500 2790 3030
rect 2910 2817 2990 2840
rect 2910 2783 2933 2817
rect 2967 2783 2990 2817
rect 2910 2760 2990 2783
rect 2910 2577 2990 2600
rect 2910 2543 2933 2577
rect 2967 2543 2990 2577
rect 2910 2520 2990 2543
rect 2270 2100 2330 2140
rect 2370 2460 2790 2500
rect -446 2060 -218 2100
rect -138 2060 590 2100
rect 2370 2020 2410 2460
rect 4652 2140 4692 3066
rect 4820 3001 4900 3021
rect 4590 2100 4692 2140
rect 4726 2998 4900 3001
rect 4726 2964 4843 2998
rect 4877 2964 4900 2998
rect 4726 2961 4900 2964
rect -446 1960 -104 2000
rect -24 1960 590 2000
rect 2270 1980 2410 2020
rect 2450 2030 2910 2070
rect -446 1860 -331 1900
rect -252 1860 590 1900
rect -367 1740 590 1780
rect -24 1250 590 1290
rect -138 1130 590 1170
rect -252 1030 590 1070
rect 2450 1020 2490 2030
rect 4726 2020 4766 2961
rect 4820 2941 4900 2961
rect 4930 2817 5010 2840
rect 4930 2783 4953 2817
rect 4987 2783 5010 2817
rect 4930 2760 5010 2783
rect 2570 1970 2650 1990
rect 4590 1980 4766 2020
rect 2570 1967 2910 1970
rect 2570 1933 2593 1967
rect 2627 1933 2910 1967
rect 2570 1930 2910 1933
rect 2570 1910 2650 1930
rect 2270 980 2490 1020
rect 2530 1830 2910 1870
rect -366 930 590 970
rect 2530 900 2570 1830
rect 2660 1750 2740 1770
rect 2660 1747 2910 1750
rect 2660 1713 2683 1747
rect 2717 1713 2910 1747
rect 2660 1710 2910 1713
rect 2660 1690 2740 1710
rect 2270 860 2570 900
rect 290 460 370 480
rect 290 457 590 460
rect 290 423 313 457
rect 347 423 590 457
rect 290 420 590 423
rect 290 400 370 420
<< viali >>
rect 2593 3613 2627 3647
rect 4601 3583 4635 3617
rect 2803 3493 2837 3527
rect 4715 3470 4749 3504
rect 2683 3393 2717 3427
rect 4843 3363 4877 3397
rect 2763 3273 2797 3307
rect 2593 3213 2627 3247
rect 4601 3223 4635 3257
rect 313 2783 347 2817
rect 43 2663 77 2697
rect 313 2543 347 2577
rect 4715 3089 4749 3123
rect 2933 2783 2967 2817
rect 2933 2543 2967 2577
rect 4843 2964 4877 2998
rect 4953 2783 4987 2817
rect 2593 1933 2627 1967
rect 2683 1713 2717 1747
rect 313 423 347 457
<< metal1 >>
rect 150 3810 290 3910
rect 4530 3840 4570 3880
rect 4950 3840 4990 3880
rect 10 2697 110 2720
rect 10 2663 43 2697
rect 77 2663 110 2697
rect -426 990 -386 1720
rect -312 1090 -272 1840
rect -198 1190 -158 2041
rect -84 1310 -44 1940
rect 10 370 110 2663
rect 150 1550 250 3810
rect 2570 3647 2650 3670
rect 2570 3613 2593 3647
rect 2627 3613 2650 3647
rect 2570 3590 2650 3613
rect 4578 3617 4658 3640
rect 2590 3270 2630 3590
rect 4578 3583 4601 3617
rect 4635 3583 4658 3617
rect 4578 3560 4658 3583
rect 2780 3527 2860 3550
rect 2780 3493 2803 3527
rect 2837 3493 2860 3527
rect 2780 3470 2860 3493
rect 2660 3436 2740 3450
rect 2660 3384 2674 3436
rect 2726 3384 2740 3436
rect 2660 3370 2740 3384
rect 2780 3330 2820 3470
rect 2740 3307 2820 3330
rect 2740 3273 2763 3307
rect 2797 3273 2820 3307
rect 4598 3280 4638 3560
rect 4692 3504 4772 3527
rect 4692 3470 4715 3504
rect 4749 3470 4772 3504
rect 4692 3447 4772 3470
rect 2570 3256 2650 3270
rect 2570 3204 2584 3256
rect 2636 3204 2650 3256
rect 2740 3250 2820 3273
rect 4578 3257 4658 3280
rect 2570 3190 2650 3204
rect 4578 3223 4601 3257
rect 4635 3223 4658 3257
rect 4578 3200 4658 3223
rect 4711 3146 4751 3447
rect 4820 3397 4900 3420
rect 4820 3363 4843 3397
rect 4877 3363 4900 3397
rect 4820 3340 4900 3363
rect 4692 3123 4772 3146
rect 4692 3089 4715 3123
rect 4749 3089 4772 3123
rect 4692 3066 4772 3089
rect 4840 3021 4880 3340
rect 4820 2998 4900 3021
rect 4820 2964 4843 2998
rect 4877 2964 4900 2998
rect 4820 2941 4900 2964
rect 290 2826 370 2840
rect 290 2774 304 2826
rect 356 2774 370 2826
rect 290 2760 370 2774
rect 2910 2826 2990 2840
rect 2910 2774 2924 2826
rect 2976 2774 2990 2826
rect 2910 2760 2990 2774
rect 4930 2826 5010 2840
rect 4930 2774 4944 2826
rect 4996 2774 5010 2826
rect 4930 2760 5010 2774
rect 2570 2630 2910 2730
rect 4590 2630 4930 2730
rect 290 2586 370 2600
rect 290 2534 304 2586
rect 356 2534 370 2586
rect 290 2520 370 2534
rect 2910 2586 2990 2600
rect 2910 2534 2924 2586
rect 2976 2534 2990 2586
rect 2910 2520 2990 2534
rect 2570 1976 2650 1990
rect 2570 1924 2584 1976
rect 2636 1924 2650 1976
rect 2570 1910 2650 1924
rect 2660 1756 2740 1770
rect 2660 1704 2674 1756
rect 2726 1704 2740 1756
rect 2660 1690 2740 1704
rect 150 1450 590 1550
rect 290 466 370 480
rect 290 414 304 466
rect 356 414 370 466
rect 290 400 370 414
rect 10 270 590 370
<< via1 >>
rect 2674 3427 2726 3436
rect 2674 3393 2683 3427
rect 2683 3393 2717 3427
rect 2717 3393 2726 3427
rect 2674 3384 2726 3393
rect 2584 3247 2636 3256
rect 2584 3213 2593 3247
rect 2593 3213 2627 3247
rect 2627 3213 2636 3247
rect 2584 3204 2636 3213
rect 4504 2894 4556 2946
rect 304 2817 356 2826
rect 304 2783 313 2817
rect 313 2783 347 2817
rect 347 2783 356 2817
rect 304 2774 356 2783
rect 2924 2817 2976 2826
rect 2924 2783 2933 2817
rect 2933 2783 2967 2817
rect 2967 2783 2976 2817
rect 2924 2774 2976 2783
rect 4944 2817 4996 2826
rect 4944 2783 4953 2817
rect 4953 2783 4987 2817
rect 4987 2783 4996 2817
rect 4944 2774 4996 2783
rect 304 2577 356 2586
rect 304 2543 313 2577
rect 313 2543 347 2577
rect 347 2543 356 2577
rect 304 2534 356 2543
rect 2924 2577 2976 2586
rect 2924 2543 2933 2577
rect 2933 2543 2967 2577
rect 2967 2543 2976 2577
rect 2924 2534 2976 2543
rect 4504 2414 4556 2466
rect 2584 1967 2636 1976
rect 2584 1933 2593 1967
rect 2593 1933 2627 1967
rect 2627 1933 2636 1967
rect 2584 1924 2636 1933
rect 2674 1747 2726 1756
rect 2674 1713 2683 1747
rect 2683 1713 2717 1747
rect 2717 1713 2726 1747
rect 2674 1704 2726 1713
rect 304 457 356 466
rect 304 423 313 457
rect 313 423 347 457
rect 347 423 356 457
rect 304 414 356 423
<< metal2 >>
rect 310 2840 350 4000
rect 2660 3436 2740 3450
rect 2660 3384 2674 3436
rect 2726 3384 2740 3436
rect 2660 3370 2740 3384
rect 2570 3256 2650 3270
rect 2570 3204 2584 3256
rect 2636 3204 2650 3256
rect 2570 3190 2650 3204
rect 290 2826 370 2840
rect 290 2774 304 2826
rect 356 2774 370 2826
rect 290 2760 370 2774
rect 310 2600 350 2760
rect 290 2586 370 2600
rect 290 2534 304 2586
rect 356 2534 370 2586
rect 290 2520 370 2534
rect 310 480 350 2520
rect 2590 1990 2630 3190
rect 2570 1976 2650 1990
rect 2570 1924 2584 1976
rect 2636 1924 2650 1976
rect 2570 1910 2650 1924
rect 2680 1770 2720 3370
rect 2930 2840 2970 4000
rect 4490 2946 4570 2960
rect 4490 2894 4504 2946
rect 4556 2894 4570 2946
rect 2910 2826 2990 2840
rect 2910 2774 2924 2826
rect 2976 2774 2990 2826
rect 2910 2760 2990 2774
rect 2930 2600 2970 2760
rect 2910 2586 2990 2600
rect 2910 2534 2924 2586
rect 2976 2534 2990 2586
rect 2910 2520 2990 2534
rect 4490 2466 4570 2894
rect 4950 2840 4990 4000
rect 4930 2826 5010 2840
rect 4930 2774 4944 2826
rect 4996 2774 5010 2826
rect 4930 2760 5010 2774
rect 4490 2414 4504 2466
rect 4556 2414 4570 2466
rect 4490 2400 4570 2414
rect 2660 1756 2740 1770
rect 2660 1704 2674 1756
rect 2726 1704 2740 1756
rect 2660 1690 2740 1704
rect 290 466 370 480
rect 290 414 304 466
rect 356 414 370 466
rect 290 400 370 414
use EESPFAL_NAND_v3  EESPFAL_NAND_v3_0
timestamp 1673383081
transform 1 0 7260 0 1 2550
box -4390 54 -2630 1410
use EESPFAL_NAND_v3  EESPFAL_NAND_v3_1
timestamp 1673383081
transform 1 0 4940 0 1 190
box -4390 54 -2630 1410
use EESPFAL_NAND_v3  EESPFAL_NAND_v3_2
timestamp 1673383081
transform 1 0 7260 0 -1 2810
box -4390 54 -2630 1410
use EESPFAL_NOR_v3  EESPFAL_NOR_v3_0
timestamp 1673383081
transform 1 0 6900 0 1 2320
box -2010 284 -250 1640
use EESPFAL_NOR_v3  EESPFAL_NOR_v3_1
timestamp 1673383081
transform 1 0 2560 0 -1 3040
box -2010 284 -250 1640
use EESPFAL_XOR_v3  EESPFAL_XOR_v3_0
timestamp 1673383081
transform 1 0 1580 0 1 2460
box -1330 144 1030 1500
use Li_mcon_M1  Li_mcon_M1_0
timestamp 1673383081
transform 1 0 -84 0 1 1960
box -20 -20 60 60
use Li_mcon_M1  Li_mcon_M1_1
timestamp 1673383081
transform 1 0 -198 0 1 2060
box -20 -20 60 60
use Li_mcon_M1  Li_mcon_M1_2
timestamp 1673383081
transform 1 0 -312 0 1 1860
box -20 -20 60 60
use Li_mcon_M1  Li_mcon_M1_3
timestamp 1673383081
transform 1 0 -426 0 1 1740
box -20 -20 60 60
use Li_mcon_M1  Li_mcon_M1_4
timestamp 1673383081
transform 1 0 -426 0 -1 970
box -20 -20 60 60
use Li_mcon_M1  Li_mcon_M1_5
timestamp 1673383081
transform 1 0 -312 0 -1 1070
box -20 -20 60 60
use Li_mcon_M1  Li_mcon_M1_6
timestamp 1673383081
transform 1 0 -198 0 -1 1170
box -20 -20 60 60
use Li_mcon_M1  Li_mcon_M1_7
timestamp 1673383081
transform 1 0 -84 0 -1 1290
box -20 -20 60 60
<< labels >>
flabel locali s 20 3720 40 3740 2 FreeSans 2000 0 0 0 x0 
port 1 nsew
flabel locali s 20 3620 40 3640 2 FreeSans 2000 0 0 0 x0_bar
port 2 nsew
flabel locali s 20 3520 40 3540 2 FreeSans 2000 0 0 0 x3
port 3 nsew
flabel locali s 20 3420 40 3440 2 FreeSans 2000 0 0 0 x3_bar
port 4 nsew
flabel locali s 20 2070 40 2090 2 FreeSans 2000 0 0 0 x1_bar
port 5 nsew
flabel locali s 20 1969 40 1989 2 FreeSans 2000 0 0 0 x2
port 6 nsew
flabel locali s 20 1870 40 1890 2 FreeSans 2000 0 0 0 x2_bar
port 7 nsew
flabel locali s 20 1750 40 1770 2 FreeSans 2000 0 0 0 x1
port 8 nsew
flabel locali s 6579 3349 6601 3372 2 FreeSans 2000 0 0 0 s0_bar
port 9 nsew
flabel locali s 6580 3230 6600 3250 2 FreeSans 2000 0 0 0 s0
port 10 nsew
flabel metal1 s 180 3840 220 3880 2 FreeSans 2000 0 0 0 CLK1
port 11 nsew
flabel metal1 s 40 2660 80 2700 2 FreeSans 2000 0 0 0 GND
port 12 nsew
flabel metal1 s 4530 3840 4570 3880 2 FreeSans 2000 0 0 0 CLK2
port 13 nsew
flabel metal1 s 4950 3840 4990 3880 2 FreeSans 2000 0 0 0 CLK3
port 14 nsew
flabel metal2 s 4960 3972 4981 3993 2 FreeSans 2000 0 0 0 Dis3
port 15 nsew
flabel metal2 s 2940 3973 2960 3994 2 FreeSans 2000 0 0 0 Dis2
port 16 nsew
flabel metal2 s 321 3974 341 3993 2 FreeSans 2000 0 0 0 Dis1
port 17 nsew
<< properties >>
string path 24.850 14.200 24.850 20.000 
<< end >>
