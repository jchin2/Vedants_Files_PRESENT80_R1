magic
tech sky130A
magscale 1 2
timestamp 1670967604
<< locali >>
rect -1610 67 -230 90
rect -1610 33 -1549 67
rect -1515 33 -1477 67
rect -1443 33 -1405 67
rect -1371 33 -1333 67
rect -1299 33 -1261 67
rect -1227 33 -1189 67
rect -1155 33 -1117 67
rect -1083 33 -1045 67
rect -1011 33 -973 67
rect -939 33 -901 67
rect -867 33 -829 67
rect -795 33 -757 67
rect -723 33 -685 67
rect -651 33 -613 67
rect -579 33 -541 67
rect -507 33 -469 67
rect -435 33 -397 67
rect -363 33 -325 67
rect -291 33 -230 67
rect -1610 10 -230 33
<< viali >>
rect -1549 33 -1515 67
rect -1477 33 -1443 67
rect -1405 33 -1371 67
rect -1333 33 -1299 67
rect -1261 33 -1227 67
rect -1189 33 -1155 67
rect -1117 33 -1083 67
rect -1045 33 -1011 67
rect -973 33 -939 67
rect -901 33 -867 67
rect -829 33 -795 67
rect -757 33 -723 67
rect -685 33 -651 67
rect -613 33 -579 67
rect -541 33 -507 67
rect -469 33 -435 67
rect -397 33 -363 67
rect -325 33 -291 67
<< metal1 >>
rect -1610 67 -230 100
rect -1610 33 -1549 67
rect -1515 33 -1477 67
rect -1443 33 -1405 67
rect -1371 33 -1333 67
rect -1299 33 -1261 67
rect -1227 33 -1189 67
rect -1155 33 -1117 67
rect -1083 33 -1045 67
rect -1011 33 -973 67
rect -939 33 -901 67
rect -867 33 -829 67
rect -795 33 -757 67
rect -723 33 -685 67
rect -651 33 -613 67
rect -579 33 -541 67
rect -507 33 -469 67
rect -435 33 -397 67
rect -363 33 -325 67
rect -291 33 -230 67
rect -1610 0 -230 33
<< end >>
