* NGSPICE file created from CMOS_s0_flat.ext - technology: sky130A

.subckt CMOS_s0_flat GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar s0 VDD
X0 VDD.t12 CMOS_AND_0/A a_425_640# VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X1 VDD.t3 x0.t0 a_n1990_n1548# VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X2 VDD.t17 x2.t0 a_n787_n1548# VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X3 CMOS_AND_0/AND a_425_640# VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X4 CMOS_AND_1/B a_n2140_n1548# GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n787_n1548# x1_bar.t0 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X6 a_n787_640# x1.t0 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X7 a_n787_30# x1.t1 GND.t5 GND.t0 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 CMOS_AND_1/A a_n787_n1548# GND.t20 GND.t14 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X9 CMOS_AND_0/A x0.t1 a_n2290_640# VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X10 a_1637_640# CMOS_AND_0/AND VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X11 CMOS_AND_1/A a_n787_n1548# VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X12 a_n1990_n638# x0_bar.t0 a_n2140_n1548# GND.t2 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X13 a_1637_30# CMOS_AND_0/AND GND.t19 GND.t18 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X14 VDD.t8 x3.t0 a_n1990_640# VDD.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X15 CMOS_AND_0/A x3.t1 a_n2290_30# GND.t7 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X16 a_425_640# CMOS_AND_0/B VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X17 a_425_30# CMOS_AND_0/B GND.t23 GND.t21 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X18 CMOS_AND_0/B a_n787_30# VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X19 s0.t1 a_1637_30# VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X20 a_n787_30# x2_bar.t0 a_n787_640# VDD.t9 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X21 a_n2140_n1548# x0.t2 a_n2290_n638# GND.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X22 a_n2290_n638# x3.t2 GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X23 a_n787_n638# x1_bar.t1 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X24 a_n787_n1548# x2.t1 a_n787_n638# GND.t3 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X25 GND.t4 x2_bar.t1 a_n787_30# GND.t3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X26 a_1637_30# CMOS_AND_1/AND a_1637_640# VDD.t18 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X27 a_n2140_n1548# x3.t3 a_n2290_n1548# VDD.t13 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X28 a_n1990_30# x3_bar.t0 CMOS_AND_0/A GND.t2 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X29 a_425_n638# CMOS_AND_1/B GND.t22 GND.t21 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X30 a_425_n1548# CMOS_AND_1/A a_425_n638# GND.t6 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X31 a_n2290_n1548# x0_bar.t1 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X32 CMOS_AND_1/B a_n2140_n1548# VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X33 a_n1990_640# x0_bar.t2 CMOS_AND_0/A VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X34 CMOS_AND_0/AND a_425_640# GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X35 CMOS_AND_0/B a_n787_30# GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X36 GND.t29 x0_bar.t3 a_n1990_30# GND.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X37 a_n2290_640# x3_bar.t1 VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X38 CMOS_AND_1/AND a_425_n1548# VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X39 GND.t30 x3_bar.t2 a_n1990_n638# GND.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X40 a_n2290_30# x0.t3 GND.t24 GND.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X41 GND.t13 CMOS_AND_1/AND a_1637_30# GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X42 a_425_n1548# CMOS_AND_1/B VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X43 VDD.t36 CMOS_AND_1/A a_425_n1548# VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X44 a_425_640# CMOS_AND_0/A a_425_30# GND.t6 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X45 s0.t0 a_1637_30# GND.t26 GND.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X46 a_n1990_n1548# x3_bar.t3 a_n2140_n1548# VDD.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X47 CMOS_AND_1/AND a_425_n1548# GND.t27 GND.t8 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
R0 VDD.n261 VDD.t13 38.206
R1 VDD.n119 VDD.t6 36.141
R2 VDD.n288 VDD.t39 32.01
R3 VDD.n269 VDD.t0 32.01
R4 VDD.n306 VDD.t10 29.945
R5 VDD.n249 VDD.t41 29.945
R6 VDD.n331 VDD.t37 24.782
R7 VDD.n80 VDD.t29 24.782
R8 VDD.n33 VDD.t23 24.782
R9 VDD.n155 VDD.t27 24.782
R10 VDD.n202 VDD.t4 24.782
R11 VDD.n314 VDD.t7 23.75
R12 VDD.n241 VDD.t2 23.75
R13 VDD.n287 VDD.t40 22.029
R14 VDD.n318 VDD.t8 22.029
R15 VDD.n326 VDD.t38 22.029
R16 VDD.n101 VDD.t20 22.029
R17 VDD.n88 VDD.t30 22.029
R18 VDD.n67 VDD.t12 22.029
R19 VDD.n54 VDD.t15 22.029
R20 VDD.n41 VDD.t24 22.029
R21 VDD.n8 VDD.t32 22.029
R22 VDD.n129 VDD.t34 22.029
R23 VDD.n142 VDD.t36 22.029
R24 VDD.n163 VDD.t28 22.029
R25 VDD.n176 VDD.t26 22.029
R26 VDD.n189 VDD.t17 22.029
R27 VDD.n210 VDD.t5 22.029
R28 VDD.n223 VDD.t22 22.029
R29 VDD.n240 VDD.t3 22.029
R30 VDD.n273 VDD.t1 22.029
R31 VDD.n339 VDD.t9 18.586
R32 VDD.n72 VDD.t11 18.586
R33 VDD.n25 VDD.t18 18.586
R34 VDD.n147 VDD.t35 18.586
R35 VDD.n194 VDD.t16 18.586
R36 VDD.n219 VDD.t21 18.586
R37 VDD.n97 VDD.t19 12.391
R38 VDD.n50 VDD.t14 12.391
R39 VDD.n4 VDD.t31 12.391
R40 VDD.n125 VDD.t33 12.391
R41 VDD.n172 VDD.t25 12.391
R42 VDD.n300 VDD.n299 11.52
R43 VDD.n74 VDD.n71 11.52
R44 VDD.n27 VDD.n24 11.52
R45 VDD.n149 VDD.n146 11.52
R46 VDD.n196 VDD.n193 11.52
R47 VDD.n263 VDD.n260 11.52
R48 VDD.n123 VDD.n122 8.855
R49 VDD.n170 VDD.n169 8.855
R50 VDD.n217 VDD.n216 8.855
R51 VDD.n221 VDD.n220 8.855
R52 VDD.n220 VDD.n219 8.855
R53 VDD.n226 VDD.n225 8.855
R54 VDD.n225 VDD.n224 8.855
R55 VDD.n230 VDD.n229 8.855
R56 VDD.n229 VDD.n228 8.855
R57 VDD.n234 VDD.n233 8.855
R58 VDD.n233 VDD.n232 8.855
R59 VDD.n238 VDD.n237 8.855
R60 VDD.n237 VDD.n236 8.855
R61 VDD.n243 VDD.n242 8.855
R62 VDD.n242 VDD.n241 8.855
R63 VDD.n247 VDD.n246 8.855
R64 VDD.n246 VDD.n245 8.855
R65 VDD.n251 VDD.n250 8.855
R66 VDD.n250 VDD.n249 8.855
R67 VDD.n255 VDD.n254 8.855
R68 VDD.n254 VDD.n253 8.855
R69 VDD.n260 VDD.n259 8.855
R70 VDD.n259 VDD.n258 8.855
R71 VDD.n263 VDD.n262 8.855
R72 VDD.n262 VDD.n261 8.855
R73 VDD.n267 VDD.n266 8.855
R74 VDD.n266 VDD.n265 8.855
R75 VDD.n271 VDD.n270 8.855
R76 VDD.n270 VDD.n269 8.855
R77 VDD.n276 VDD.n275 8.855
R78 VDD.n174 VDD.n173 8.855
R79 VDD.n173 VDD.n172 8.855
R80 VDD.n179 VDD.n178 8.855
R81 VDD.n178 VDD.n177 8.855
R82 VDD.n183 VDD.n182 8.855
R83 VDD.n182 VDD.n181 8.855
R84 VDD.n187 VDD.n186 8.855
R85 VDD.n186 VDD.n185 8.855
R86 VDD.n193 VDD.n192 8.855
R87 VDD.n192 VDD.n191 8.855
R88 VDD.n196 VDD.n195 8.855
R89 VDD.n195 VDD.n194 8.855
R90 VDD.n200 VDD.n199 8.855
R91 VDD.n199 VDD.n198 8.855
R92 VDD.n204 VDD.n203 8.855
R93 VDD.n203 VDD.n202 8.855
R94 VDD.n208 VDD.n207 8.855
R95 VDD.n127 VDD.n126 8.855
R96 VDD.n126 VDD.n125 8.855
R97 VDD.n132 VDD.n131 8.855
R98 VDD.n131 VDD.n130 8.855
R99 VDD.n136 VDD.n135 8.855
R100 VDD.n135 VDD.n134 8.855
R101 VDD.n140 VDD.n139 8.855
R102 VDD.n139 VDD.n138 8.855
R103 VDD.n146 VDD.n145 8.855
R104 VDD.n145 VDD.n144 8.855
R105 VDD.n149 VDD.n148 8.855
R106 VDD.n148 VDD.n147 8.855
R107 VDD.n153 VDD.n152 8.855
R108 VDD.n152 VDD.n151 8.855
R109 VDD.n157 VDD.n156 8.855
R110 VDD.n156 VDD.n155 8.855
R111 VDD.n161 VDD.n160 8.855
R112 VDD.n2 VDD.n1 8.855
R113 VDD.n6 VDD.n5 8.855
R114 VDD.n5 VDD.n4 8.855
R115 VDD.n11 VDD.n10 8.855
R116 VDD.n10 VDD.n9 8.855
R117 VDD.n15 VDD.n14 8.855
R118 VDD.n14 VDD.n13 8.855
R119 VDD.n19 VDD.n18 8.855
R120 VDD.n18 VDD.n17 8.855
R121 VDD.n24 VDD.n23 8.855
R122 VDD.n23 VDD.n22 8.855
R123 VDD.n27 VDD.n26 8.855
R124 VDD.n26 VDD.n25 8.855
R125 VDD.n31 VDD.n30 8.855
R126 VDD.n30 VDD.n29 8.855
R127 VDD.n35 VDD.n34 8.855
R128 VDD.n34 VDD.n33 8.855
R129 VDD.n39 VDD.n38 8.855
R130 VDD.n48 VDD.n47 8.855
R131 VDD.n52 VDD.n51 8.855
R132 VDD.n51 VDD.n50 8.855
R133 VDD.n57 VDD.n56 8.855
R134 VDD.n56 VDD.n55 8.855
R135 VDD.n61 VDD.n60 8.855
R136 VDD.n60 VDD.n59 8.855
R137 VDD.n65 VDD.n64 8.855
R138 VDD.n64 VDD.n63 8.855
R139 VDD.n71 VDD.n70 8.855
R140 VDD.n70 VDD.n69 8.855
R141 VDD.n74 VDD.n73 8.855
R142 VDD.n73 VDD.n72 8.855
R143 VDD.n78 VDD.n77 8.855
R144 VDD.n77 VDD.n76 8.855
R145 VDD.n82 VDD.n81 8.855
R146 VDD.n81 VDD.n80 8.855
R147 VDD.n86 VDD.n85 8.855
R148 VDD.n95 VDD.n94 8.855
R149 VDD.n99 VDD.n98 8.855
R150 VDD.n98 VDD.n97 8.855
R151 VDD.n104 VDD.n103 8.855
R152 VDD.n103 VDD.n102 8.855
R153 VDD.n108 VDD.n107 8.855
R154 VDD.n107 VDD.n106 8.855
R155 VDD.n112 VDD.n111 8.855
R156 VDD.n111 VDD.n110 8.855
R157 VDD.n116 VDD.n115 8.855
R158 VDD.n115 VDD.n114 8.855
R159 VDD.n341 VDD.n340 8.855
R160 VDD.n340 VDD.n339 8.855
R161 VDD.n337 VDD.n336 8.855
R162 VDD.n336 VDD.n335 8.855
R163 VDD.n333 VDD.n332 8.855
R164 VDD.n332 VDD.n331 8.855
R165 VDD.n329 VDD.n328 8.855
R166 VDD.n321 VDD.n320 8.855
R167 VDD.n316 VDD.n315 8.855
R168 VDD.n315 VDD.n314 8.855
R169 VDD.n312 VDD.n311 8.855
R170 VDD.n311 VDD.n310 8.855
R171 VDD.n308 VDD.n307 8.855
R172 VDD.n307 VDD.n306 8.855
R173 VDD.n304 VDD.n303 8.855
R174 VDD.n303 VDD.n302 8.855
R175 VDD.n300 VDD.n120 8.855
R176 VDD.n120 VDD.n119 8.855
R177 VDD.n299 VDD.n298 8.855
R178 VDD.n298 VDD.n297 8.855
R179 VDD.n294 VDD.n293 8.855
R180 VDD.n293 VDD.n292 8.855
R181 VDD.n290 VDD.n289 8.855
R182 VDD.n289 VDD.n288 8.855
R183 VDD.n285 VDD.n284 8.855
R184 VDD.n280 VDD.n279 4.91
R185 VDD.n279 VDD.n278 4.65
R186 VDD.n218 VDD.n217 4.65
R187 VDD.n222 VDD.n221 4.65
R188 VDD.n227 VDD.n226 4.65
R189 VDD.n231 VDD.n230 4.65
R190 VDD.n235 VDD.n234 4.65
R191 VDD.n239 VDD.n238 4.65
R192 VDD.n244 VDD.n243 4.65
R193 VDD.n248 VDD.n247 4.65
R194 VDD.n252 VDD.n251 4.65
R195 VDD.n256 VDD.n255 4.65
R196 VDD.n260 VDD.n257 4.65
R197 VDD.n264 VDD.n263 4.65
R198 VDD.n268 VDD.n267 4.65
R199 VDD.n272 VDD.n271 4.65
R200 VDD.n277 VDD.n276 4.65
R201 VDD.n214 VDD.n213 4.65
R202 VDD.n212 VDD.n211 4.65
R203 VDD.n171 VDD.n170 4.65
R204 VDD.n175 VDD.n174 4.65
R205 VDD.n180 VDD.n179 4.65
R206 VDD.n184 VDD.n183 4.65
R207 VDD.n188 VDD.n187 4.65
R208 VDD.n193 VDD.n190 4.65
R209 VDD.n197 VDD.n196 4.65
R210 VDD.n201 VDD.n200 4.65
R211 VDD.n205 VDD.n204 4.65
R212 VDD.n209 VDD.n208 4.65
R213 VDD.n167 VDD.n166 4.65
R214 VDD.n165 VDD.n164 4.65
R215 VDD.n128 VDD.n127 4.65
R216 VDD.n133 VDD.n132 4.65
R217 VDD.n137 VDD.n136 4.65
R218 VDD.n141 VDD.n140 4.65
R219 VDD.n146 VDD.n143 4.65
R220 VDD.n150 VDD.n149 4.65
R221 VDD.n154 VDD.n153 4.65
R222 VDD.n158 VDD.n157 4.65
R223 VDD.n162 VDD.n161 4.65
R224 VDD.n7 VDD.n6 4.65
R225 VDD.n12 VDD.n11 4.65
R226 VDD.n16 VDD.n15 4.65
R227 VDD.n20 VDD.n19 4.65
R228 VDD.n24 VDD.n21 4.65
R229 VDD.n28 VDD.n27 4.65
R230 VDD.n32 VDD.n31 4.65
R231 VDD.n36 VDD.n35 4.65
R232 VDD.n40 VDD.n39 4.65
R233 VDD.n43 VDD.n42 4.65
R234 VDD.n45 VDD.n44 4.65
R235 VDD.n49 VDD.n48 4.65
R236 VDD.n53 VDD.n52 4.65
R237 VDD.n58 VDD.n57 4.65
R238 VDD.n62 VDD.n61 4.65
R239 VDD.n66 VDD.n65 4.65
R240 VDD.n71 VDD.n68 4.65
R241 VDD.n75 VDD.n74 4.65
R242 VDD.n79 VDD.n78 4.65
R243 VDD.n83 VDD.n82 4.65
R244 VDD.n87 VDD.n86 4.65
R245 VDD.n90 VDD.n89 4.65
R246 VDD.n92 VDD.n91 4.65
R247 VDD.n96 VDD.n95 4.65
R248 VDD.n100 VDD.n99 4.65
R249 VDD.n105 VDD.n104 4.65
R250 VDD.n109 VDD.n108 4.65
R251 VDD.n113 VDD.n112 4.65
R252 VDD.n117 VDD.n116 4.65
R253 VDD.n342 VDD.n341 4.65
R254 VDD.n338 VDD.n337 4.65
R255 VDD.n334 VDD.n333 4.65
R256 VDD.n330 VDD.n329 4.65
R257 VDD.n325 VDD.n324 4.65
R258 VDD.n323 VDD.n118 4.65
R259 VDD.n322 VDD.n321 4.65
R260 VDD.n317 VDD.n316 4.65
R261 VDD.n313 VDD.n312 4.65
R262 VDD.n309 VDD.n308 4.65
R263 VDD.n305 VDD.n304 4.65
R264 VDD.n301 VDD.n300 4.65
R265 VDD.n299 VDD.n296 4.65
R266 VDD.n295 VDD.n294 4.65
R267 VDD.n291 VDD.n290 4.65
R268 VDD.n286 VDD.n285 4.65
R269 VDD.n282 VDD.n281 4.65
R270 VDD.n1 VDD.n0 4.288
R271 VDD.n47 VDD.n46 4.288
R272 VDD.n94 VDD.n93 4.288
R273 VDD.n320 VDD.n319 4.288
R274 VDD.n122 VDD.n121 4.288
R275 VDD.n169 VDD.n168 4.288
R276 VDD.n216 VDD.n215 4.288
R277 VDD.n275 VDD.n274 4.288
R278 VDD.n207 VDD.n206 4.288
R279 VDD.n160 VDD.n159 4.288
R280 VDD.n38 VDD.n37 4.288
R281 VDD.n85 VDD.n84 4.288
R282 VDD.n328 VDD.n327 4.288
R283 VDD.n284 VDD.n283 4.288
R284 VDD.n3 VDD.n2 2.562
R285 VDD.n124 VDD.n123 2.562
R286 VDD.n7 VDD.n3 1.145
R287 VDD.n128 VDD.n124 1.145
R288 VDD.n325 VDD.n323 0.957
R289 VDD.n167 VDD.n165 0.525
R290 VDD.n45 VDD.n43 0.525
R291 VDD.n92 VDD.n90 0.525
R292 VDD.n214 VDD.n212 0.507
R293 VDD.n282 VDD.n280 0.135
R294 VDD.n137 VDD.n133 0.09
R295 VDD.n141 VDD.n137 0.09
R296 VDD.n143 VDD.n141 0.09
R297 VDD.n154 VDD.n150 0.09
R298 VDD.n158 VDD.n154 0.09
R299 VDD.n162 VDD.n158 0.09
R300 VDD.n171 VDD.n167 0.09
R301 VDD.n175 VDD.n171 0.09
R302 VDD.n184 VDD.n180 0.09
R303 VDD.n188 VDD.n184 0.09
R304 VDD.n190 VDD.n188 0.09
R305 VDD.n201 VDD.n197 0.09
R306 VDD.n205 VDD.n201 0.09
R307 VDD.n209 VDD.n205 0.09
R308 VDD.n218 VDD.n214 0.09
R309 VDD.n222 VDD.n218 0.09
R310 VDD.n231 VDD.n227 0.09
R311 VDD.n235 VDD.n231 0.09
R312 VDD.n239 VDD.n235 0.09
R313 VDD.n248 VDD.n244 0.09
R314 VDD.n252 VDD.n248 0.09
R315 VDD.n256 VDD.n252 0.09
R316 VDD.n257 VDD.n256 0.09
R317 VDD.n268 VDD.n264 0.09
R318 VDD.n272 VDD.n268 0.09
R319 VDD.n279 VDD.n277 0.09
R320 VDD.n16 VDD.n12 0.09
R321 VDD.n20 VDD.n16 0.09
R322 VDD.n21 VDD.n20 0.09
R323 VDD.n32 VDD.n28 0.09
R324 VDD.n36 VDD.n32 0.09
R325 VDD.n40 VDD.n36 0.09
R326 VDD.n49 VDD.n45 0.09
R327 VDD.n53 VDD.n49 0.09
R328 VDD.n62 VDD.n58 0.09
R329 VDD.n66 VDD.n62 0.09
R330 VDD.n68 VDD.n66 0.09
R331 VDD.n79 VDD.n75 0.09
R332 VDD.n83 VDD.n79 0.09
R333 VDD.n87 VDD.n83 0.09
R334 VDD.n96 VDD.n92 0.09
R335 VDD.n100 VDD.n96 0.09
R336 VDD.n109 VDD.n105 0.09
R337 VDD.n113 VDD.n109 0.09
R338 VDD.n117 VDD.n113 0.09
R339 VDD.n342 VDD.n338 0.09
R340 VDD.n338 VDD.n334 0.09
R341 VDD.n334 VDD.n330 0.09
R342 VDD.n323 VDD.n322 0.09
R343 VDD.n317 VDD.n313 0.09
R344 VDD.n313 VDD.n309 0.09
R345 VDD.n309 VDD.n305 0.09
R346 VDD.n305 VDD.n301 0.09
R347 VDD.n296 VDD.n295 0.09
R348 VDD.n295 VDD.n291 0.09
R349 VDD.n286 VDD.n282 0.09
R350 VDD.n129 VDD.n128 0.078
R351 VDD.n176 VDD.n175 0.078
R352 VDD.n8 VDD.n7 0.078
R353 VDD.n54 VDD.n53 0.078
R354 VDD.n101 VDD.n100 0.078
R355 VDD.n223 VDD.n222 0.071
R356 VDD.n150 CMOS_AND_1/VDD 0.065
R357 VDD.n197 CMOS_AND_2/VDD 0.065
R358 VDD.n244 VDD.n240 0.065
R359 VDD.n264 CMOS_XNOR_0/VDD 0.065
R360 VDD.n28 CMOS_OR_0/VDD 0.065
R361 VDD.n75 CMOS_AND_0/VDD 0.065
R362 CMOS_OR_1/VDD VDD.n342 0.065
R363 VDD.n318 VDD.n317 0.065
R364 VDD.n296 VDD 0.065
R365 VDD.n165 VDD.n163 0.056
R366 VDD.n212 VDD.n210 0.056
R367 VDD.n43 VDD.n41 0.056
R368 VDD.n90 VDD.n88 0.056
R369 VDD.n326 VDD.n325 0.056
R370 VDD.n273 VDD.n272 0.055
R371 VDD.n291 VDD.n287 0.055
R372 VDD.n277 VDD.n273 0.035
R373 VDD.n287 VDD.n286 0.035
R374 VDD.n163 VDD.n162 0.033
R375 VDD.n210 VDD.n209 0.033
R376 VDD.n41 VDD.n40 0.033
R377 VDD.n88 VDD.n87 0.033
R378 VDD.n330 VDD.n326 0.033
R379 VDD.n280 VDD 0.027
R380 VDD.n240 VDD.n239 0.025
R381 VDD.n257 CMOS_XNOR_0/VDD 0.025
R382 VDD.n21 CMOS_OR_0/VDD 0.025
R383 CMOS_OR_1/VDD VDD.n117 0.025
R384 VDD.n322 VDD.n318 0.025
R385 VDD.n301 VDD 0.025
R386 VDD.n227 VDD.n223 0.018
R387 VDD.n143 VDD.n142 0.017
R388 VDD.n190 VDD.n189 0.017
R389 VDD.n68 VDD.n67 0.017
R390 VDD.n133 VDD.n129 0.011
R391 VDD.n180 VDD.n176 0.011
R392 VDD.n12 VDD.n8 0.011
R393 VDD.n58 VDD.n54 0.011
R394 VDD.n105 VDD.n101 0.011
R395 VDD.n142 CMOS_AND_1/VDD 0.007
R396 VDD.n189 CMOS_AND_2/VDD 0.007
R397 VDD.n67 CMOS_AND_0/VDD 0.007
R398 x0.n0 x0.t1 993.097
R399 x0.t0 x0.t2 923.343
R400 CMOS_XNOR_0/B x0.t0 633.02
R401 x0.n1 CMOS_XNOR_0/B 539.008
R402 x0 x0.n1 391.88
R403 x0.n0 x0.t3 356.59
R404 x0 x0.n0 78.72
R405 x0.n1 x0 1.597
R406 x2.t1 x2.t0 1221.07
R407 x2 x2.t1 392.02
R408 GND.n69 GND.t16 1283.79
R409 GND.n70 GND.n69 284.705
R410 GND.n192 GND.t18 180.204
R411 GND.n48 GND.t7 150.98
R412 GND.n200 GND.t12 135.153
R413 GND.n36 GND.t10 133.725
R414 GND.n56 GND.t2 125.098
R415 GND.n147 GND.t21 103.529
R416 GND.n102 GND.t0 103.529
R417 GND.n64 GND.t28 99.215
R418 GND.n4 GND.t25 90.102
R419 GND.n156 GND.t6 77.647
R420 GND.n111 GND.t3 77.647
R421 GND.n176 GND.t8 51.764
R422 GND.n131 GND.t14 51.764
R423 GND.n30 GND 37.93
R424 GND.n35 GND.t24 30.21
R425 GND.n175 GND.t27 30.21
R426 GND.n142 GND.t22 30.21
R427 GND.n130 GND.t20 30.21
R428 GND.n97 GND.t1 30.21
R429 GND.n68 GND.t30 30.21
R430 GND.n35 GND.t11 30.21
R431 GND.n84 GND.t17 30.21
R432 GND.n8 GND.t26 30.21
R433 GND.n25 GND.t13 30.21
R434 GND.n187 GND.t19 30.21
R435 GND.n175 GND.t9 30.21
R436 GND.n142 GND.t23 30.21
R437 GND.n130 GND.t15 30.21
R438 GND.n28 GND.t4 30.21
R439 GND.n97 GND.t5 30.21
R440 GND.n68 GND.t29 30.21
R441 GND.n94 GND.n93 17.263
R442 GND.n161 GND.n158 11.52
R443 GND.n116 GND.n113 11.52
R444 GND.n50 GND.n47 11.52
R445 GND.n2 GND.n1 9.154
R446 GND.n182 GND.n181 9.154
R447 GND.n137 GND.n136 9.154
R448 GND.n133 GND.n132 9.154
R449 GND.n132 GND.n131 9.154
R450 GND.n128 GND.n127 9.154
R451 GND.n127 GND.n126 9.154
R452 GND.n124 GND.n123 9.154
R453 GND.n123 GND.n122 9.154
R454 GND.n120 GND.n119 9.154
R455 GND.n119 GND.n118 9.154
R456 GND.n116 GND.n115 9.154
R457 GND.n115 GND.n114 9.154
R458 GND.n113 GND.n112 9.154
R459 GND.n112 GND.n111 9.154
R460 GND.n108 GND.n107 9.154
R461 GND.n107 GND.n106 9.154
R462 GND.n104 GND.n103 9.154
R463 GND.n103 GND.n102 9.154
R464 GND.n100 GND.n99 9.154
R465 GND.n178 GND.n177 9.154
R466 GND.n177 GND.n176 9.154
R467 GND.n173 GND.n172 9.154
R468 GND.n172 GND.n171 9.154
R469 GND.n169 GND.n168 9.154
R470 GND.n168 GND.n167 9.154
R471 GND.n165 GND.n164 9.154
R472 GND.n164 GND.n163 9.154
R473 GND.n161 GND.n160 9.154
R474 GND.n160 GND.n159 9.154
R475 GND.n158 GND.n157 9.154
R476 GND.n157 GND.n156 9.154
R477 GND.n153 GND.n152 9.154
R478 GND.n152 GND.n151 9.154
R479 GND.n149 GND.n148 9.154
R480 GND.n148 GND.n147 9.154
R481 GND.n145 GND.n144 9.154
R482 GND.n6 GND.n5 9.154
R483 GND.n5 GND.n4 9.154
R484 GND.n11 GND.n10 9.154
R485 GND.n10 GND.n9 9.154
R486 GND.n15 GND.n14 9.154
R487 GND.n14 GND.n13 9.154
R488 GND.n19 GND.n18 9.154
R489 GND.n18 GND.n17 9.154
R490 GND.n23 GND.n22 9.154
R491 GND.n22 GND.n21 9.154
R492 GND.n202 GND.n201 9.154
R493 GND.n201 GND.n200 9.154
R494 GND.n198 GND.n197 9.154
R495 GND.n197 GND.n196 9.154
R496 GND.n194 GND.n193 9.154
R497 GND.n193 GND.n192 9.154
R498 GND.n190 GND.n189 9.154
R499 GND.n90 GND.n89 9.154
R500 GND.n87 GND.n86 9.154
R501 GND.n82 GND.n81 9.154
R502 GND.n79 GND.n78 9.154
R503 GND.n75 GND.n74 9.154
R504 GND.n72 GND.n71 9.154
R505 GND.n71 GND.n70 9.154
R506 GND.n66 GND.n65 9.154
R507 GND.n65 GND.n64 9.154
R508 GND.n62 GND.n61 9.154
R509 GND.n61 GND.n60 9.154
R510 GND.n58 GND.n57 9.154
R511 GND.n57 GND.n56 9.154
R512 GND.n54 GND.n53 9.154
R513 GND.n53 GND.n52 9.154
R514 GND.n50 GND.n49 9.154
R515 GND.n49 GND.n48 9.154
R516 GND.n47 GND.n46 9.154
R517 GND.n46 GND.n45 9.154
R518 GND.n42 GND.n41 9.154
R519 GND.n41 GND.n40 9.154
R520 GND.n38 GND.n37 9.154
R521 GND.n37 GND.n36 9.154
R522 GND.n33 GND.n32 9.154
R523 GND.n86 GND.n85 8.108
R524 GND.n78 GND.n77 8.108
R525 GND.n96 GND.n29 4.65
R526 GND.n138 GND.n137 4.65
R527 GND.n134 GND.n133 4.65
R528 GND.n129 GND.n128 4.65
R529 GND.n125 GND.n124 4.65
R530 GND.n121 GND.n120 4.65
R531 GND.n117 GND.n116 4.65
R532 GND.n113 GND.n110 4.65
R533 GND.n109 GND.n108 4.65
R534 GND.n105 GND.n104 4.65
R535 GND.n101 GND.n100 4.65
R536 GND.n140 GND.n139 4.65
R537 GND.n141 GND.n27 4.65
R538 GND.n183 GND.n182 4.65
R539 GND.n179 GND.n178 4.65
R540 GND.n174 GND.n173 4.65
R541 GND.n170 GND.n169 4.65
R542 GND.n166 GND.n165 4.65
R543 GND.n162 GND.n161 4.65
R544 GND.n158 GND.n155 4.65
R545 GND.n154 GND.n153 4.65
R546 GND.n150 GND.n149 4.65
R547 GND.n146 GND.n145 4.65
R548 GND.n185 GND.n184 4.65
R549 GND.n186 GND.n26 4.65
R550 GND.n7 GND.n6 4.65
R551 GND.n12 GND.n11 4.65
R552 GND.n16 GND.n15 4.65
R553 GND.n20 GND.n19 4.65
R554 GND.n24 GND.n23 4.65
R555 GND.n203 GND.n202 4.65
R556 GND.n199 GND.n198 4.65
R557 GND.n195 GND.n194 4.65
R558 GND.n191 GND.n190 4.65
R559 GND.n91 GND.n90 4.65
R560 GND.n88 GND.n87 4.65
R561 GND.n83 GND.n82 4.65
R562 GND.n80 GND.n79 4.65
R563 GND.n76 GND.n75 4.65
R564 GND.n73 GND.n72 4.65
R565 GND.n67 GND.n66 4.65
R566 GND.n63 GND.n62 4.65
R567 GND.n59 GND.n58 4.65
R568 GND.n55 GND.n54 4.65
R569 GND.n51 GND.n50 4.65
R570 GND.n47 GND.n44 4.65
R571 GND.n43 GND.n42 4.65
R572 GND.n39 GND.n38 4.65
R573 GND.n95 GND.n94 4.65
R574 GND.n181 GND.n180 2.759
R575 GND.n136 GND.n135 2.759
R576 GND.n99 GND.n98 2.759
R577 GND.n144 GND.n143 2.759
R578 GND.n34 GND.n30 2.612
R579 GND.n3 GND.n2 2.562
R580 GND.n34 GND.n33 2.562
R581 GND.n1 GND.n0 1.853
R582 GND.n189 GND.n188 1.853
R583 GND.n32 GND.n31 1.593
R584 GND.n7 GND.n3 1.145
R585 GND.n35 GND.n34 1.09
R586 GND.n186 GND.n185 0.525
R587 GND.n141 GND.n140 0.525
R588 GND.n93 GND.n92 0.524
R589 GND.n96 GND.n95 0.507
R590 GND.n16 GND.n12 0.09
R591 GND.n20 GND.n16 0.09
R592 GND.n24 GND.n20 0.09
R593 GND.n203 GND.n199 0.09
R594 GND.n199 GND.n195 0.09
R595 GND.n195 GND.n191 0.09
R596 GND.n185 GND.n183 0.09
R597 GND.n183 GND.n179 0.09
R598 GND.n174 GND.n170 0.09
R599 GND.n170 GND.n166 0.09
R600 GND.n166 GND.n162 0.09
R601 GND.n155 GND.n154 0.09
R602 GND.n154 GND.n150 0.09
R603 GND.n150 GND.n146 0.09
R604 GND.n140 GND.n138 0.09
R605 GND.n138 GND.n134 0.09
R606 GND.n129 GND.n125 0.09
R607 GND.n125 GND.n121 0.09
R608 GND.n121 GND.n117 0.09
R609 GND.n110 GND.n109 0.09
R610 GND.n109 GND.n105 0.09
R611 GND.n105 GND.n101 0.09
R612 GND.n95 GND.n91 0.09
R613 GND.n91 GND.n88 0.09
R614 GND.n83 GND.n80 0.09
R615 GND.n80 GND.n76 0.09
R616 GND.n76 GND.n73 0.09
R617 GND.n67 GND.n63 0.09
R618 GND.n63 GND.n59 0.09
R619 GND.n59 GND.n55 0.09
R620 GND.n55 GND.n51 0.09
R621 GND.n44 GND.n43 0.09
R622 GND.n43 GND.n39 0.09
R623 GND.n8 GND.n7 0.078
R624 GND.n179 GND.n175 0.078
R625 GND.n134 GND.n130 0.078
R626 GND.n88 GND.n84 0.071
R627 CMOS_OR_0/GND GND.n203 0.065
R628 GND.n155 CMOS_AND_0/GND 0.065
R629 GND.n110 CMOS_AND_2/GND 0.065
R630 GND.n68 GND.n67 0.065
R631 GND.n44 GND 0.065
R632 GND.n187 GND.n186 0.056
R633 GND.n142 GND.n141 0.056
R634 GND.n97 GND.n96 0.056
R635 GND.n39 GND.n35 0.055
R636 GND.n191 GND.n187 0.033
R637 GND.n146 GND.n142 0.033
R638 GND.n101 GND.n97 0.033
R639 GND.n162 CMOS_AND_0/GND 0.025
R640 GND.n73 GND.n68 0.025
R641 GND.n51 GND 0.025
R642 GND.n25 GND.n24 0.018
R643 GND.n117 GND.n28 0.018
R644 GND.n84 GND.n83 0.018
R645 GND.n12 GND.n8 0.011
R646 GND.n175 GND.n174 0.011
R647 GND.n130 GND.n129 0.011
R648 CMOS_OR_0/GND GND.n25 0.006
R649 CMOS_AND_2/GND GND.n28 0.006
R650 x1_bar.n0 x1_bar.t1 579.86
R651 x1_bar.n0 x1_bar.t0 547.727
R652 x1_bar x1_bar.n0 78.72
R653 x1.n0 x1.t1 579.86
R654 x1.n0 x1.t0 547.727
R655 x1 x1.n0 78.72
R656 x0_bar.t3 x0_bar.t2 1345.61
R657 x0_bar.n0 x0_bar.t1 681.713
R658 x0_bar.n0 x0_bar.t0 528.72
R659 x0_bar x0_bar.n1 507.08
R660 x0_bar x0_bar.t3 392.02
R661 x0_bar.n1 CMOS_XNOR_0/B_bar 346.157
R662 CMOS_XNOR_0/B_bar x0_bar.n0 3.68
R663 x0_bar.n1 x0_bar 2.166
R664 x3.n0 x3.t3 993.097
R665 x3.t0 x3.t1 924.95
R666 x3 x3.t0 633.02
R667 x3.n0 x3.t2 356.59
R668 x3 x3.n1 317
R669 x3.n1 CMOS_XNOR_0/A 176.128
R670 CMOS_XNOR_0/A x3.n0 78.72
R671 x3.n1 x3 0.154
R672 s0 s0.t1 117.353
R673 s0.n0 s0.t0 95.65
R674 s0 s0.n0 10.009
R675 s0.n0 s0 0.913
R676 x2_bar.t1 x2_bar.t0 1221.07
R677 x2_bar x2_bar.t1 392.02
R678 x3_bar.t2 x3_bar.t3 1345.61
R679 x3_bar.n0 x3_bar.t1 683.32
R680 x3_bar.n0 x3_bar.t0 528.72
R681 CMOS_XNOR_0/A_bar x3_bar.t2 392.02
R682 x3_bar.n1 CMOS_XNOR_0/A_bar 287.515
R683 x3_bar x3_bar.n1 125.96
R684 x3_bar x3_bar.n0 3.68
R685 x3_bar.n1 x3_bar 1.205
C0 x1_bar CMOS_AND_1/A 0.00fF
C1 a_n787_n1548# x0_bar 0.00fF
C2 a_n1990_n1548# CMOS_AND_1/B 0.00fF
C3 CMOS_AND_1/B a_n787_640# 0.00fF
C4 a_n787_n1548# CMOS_AND_1/B 0.09fF
C5 CMOS_AND_0/A a_n1990_30# 0.01fF
C6 x2 a_n2290_30# 0.00fF
C7 CMOS_AND_0/AND a_n787_30# 0.00fF
C8 a_n2290_640# x1 0.01fF
C9 a_425_640# a_n787_640# 0.00fF
C10 a_n787_n1548# a_n2290_n1548# 0.00fF
C11 a_n2290_n638# a_n787_n1548# 0.00fF
C12 a_n787_30# a_n2290_30# 0.00fF
C13 x2 CMOS_AND_0/A 0.05fF
C14 x0 x1 0.06fF
C15 a_n2290_640# VDD 0.04fF
C16 a_n2140_n1548# x1 0.01fF
C17 CMOS_AND_0/B x1 0.00fF
C18 a_n2290_640# x3 0.02fF
C19 a_n787_30# CMOS_AND_0/A 0.07fF
C20 x1 x0_bar 2.42fF
C21 a_n787_n638# VDD 0.01fF
C22 CMOS_AND_1/A a_425_n638# 0.01fF
C23 CMOS_AND_0/AND a_425_30# 0.00fF
C24 x1 CMOS_AND_1/B 0.01fF
C25 x0 VDD 1.06fF
C26 a_n2140_n1548# VDD 1.01fF
C27 CMOS_AND_0/B VDD 0.58fF
C28 CMOS_AND_1/AND VDD 0.44fF
C29 x3 x0 0.31fF
C30 a_425_n1548# a_n787_n1548# 0.01fF
C31 a_425_640# x1 0.00fF
C32 a_n2140_n1548# x3 0.06fF
C33 x0_bar VDD 0.38fF
C34 x1 a_n2290_n1548# 0.00fF
C35 a_n2290_n638# x1 0.00fF
C36 CMOS_AND_0/B x3 0.00fF
C37 x3 x0_bar 0.36fF
C38 CMOS_AND_1/B VDD 0.78fF
C39 x2 a_n1990_30# 0.00fF
C40 x0 a_n1990_n638# 0.01fF
C41 a_n2140_n1548# a_n1990_n638# 0.01fF
C42 x3 CMOS_AND_1/B 0.00fF
C43 a_425_30# CMOS_AND_0/A 0.01fF
C44 a_425_640# VDD 0.81fF
C45 a_n787_30# a_n1990_30# 0.00fF
C46 x0_bar a_n1990_n638# 0.00fF
C47 a_n2290_n1548# VDD 0.03fF
C48 a_n2290_n638# VDD 0.00fF
C49 x3 a_n2290_n1548# 0.00fF
C50 CMOS_AND_1/B a_n1990_n638# 0.00fF
C51 a_n2290_n638# x3 0.00fF
C52 a_n2290_30# x3_bar 0.00fF
C53 a_n1990_n1548# a_n787_n1548# 0.00fF
C54 CMOS_AND_1/AND s0 0.00fF
C55 a_n787_n1548# a_n787_640# 0.00fF
C56 x1_bar a_n2290_640# 0.00fF
C57 x2_bar a_n2290_640# 0.00fF
C58 a_1637_30# VDD 0.50fF
C59 a_n787_30# x2 0.00fF
C60 CMOS_AND_0/A x3_bar 0.16fF
C61 x2_bar a_n787_n638# 0.00fF
C62 a_n1990_640# x0 0.00fF
C63 a_425_640# s0 0.00fF
C64 a_n1990_640# a_n2140_n1548# 0.00fF
C65 x1_bar x0 0.13fF
C66 x1_bar a_n2140_n1548# 0.21fF
C67 x2_bar x0 0.07fF
C68 x2_bar a_n2140_n1548# 0.04fF
C69 a_425_n1548# VDD 0.79fF
C70 x2_bar CMOS_AND_0/B 0.00fF
C71 a_n1990_640# x0_bar 0.01fF
C72 x1_bar x0_bar 0.08fF
C73 CMOS_AND_1/A CMOS_AND_0/A 0.07fF
C74 x2_bar x0_bar 0.13fF
C75 x1_bar CMOS_AND_1/B 0.42fF
C76 x2_bar CMOS_AND_1/B 0.01fF
C77 a_n1990_n1548# x1 0.00fF
C78 a_1637_30# s0 0.06fF
C79 x1 a_n787_640# 0.01fF
C80 x1_bar a_n2290_n1548# 0.01fF
C81 x2_bar a_425_640# 0.00fF
C82 a_n2290_n638# x1_bar 0.00fF
C83 a_n1990_30# x3_bar 0.00fF
C84 x2_bar a_n2290_n1548# 0.00fF
C85 x2_bar a_n2290_n638# 0.00fF
C86 a_n787_30# a_425_30# 0.00fF
C87 a_n1990_n1548# VDD 0.04fF
C88 a_n787_640# VDD 0.05fF
C89 a_n787_n1548# VDD 0.79fF
C90 x3 a_n1990_n1548# 0.00fF
C91 x3 a_n787_n1548# 0.00fF
C92 x2 x3_bar 0.14fF
C93 a_425_n638# CMOS_AND_1/AND 0.00fF
C94 a_n787_n1548# a_n1990_n638# 0.00fF
C95 a_n787_30# x3_bar 0.00fF
C96 a_425_n1548# x1_bar 0.00fF
C97 CMOS_AND_1/A x2 0.01fF
C98 a_425_n638# a_425_640# 0.00fF
C99 x1 VDD 1.09fF
C100 x3 x1 0.14fF
C101 a_1637_640# CMOS_AND_1/AND 0.01fF
C102 CMOS_AND_0/AND CMOS_AND_0/B 0.01fF
C103 x1_bar a_n1990_n1548# 0.01fF
C104 x2_bar a_n1990_n1548# 0.00fF
C105 x1 a_n1990_n638# 0.00fF
C106 CMOS_AND_0/AND CMOS_AND_1/AND 0.09fF
C107 x1_bar a_n787_n1548# 0.04fF
C108 x2_bar a_n787_640# 0.01fF
C109 x2_bar a_n787_n1548# 0.00fF
C110 a_n2290_640# CMOS_AND_0/A 0.02fF
C111 x0 a_n2290_30# 0.00fF
C112 x3 VDD 1.08fF
C113 a_425_30# CMOS_AND_1/A 0.00fF
C114 a_425_n1548# a_425_n638# 0.01fF
C115 a_n2290_30# x0_bar 0.01fF
C116 a_1637_640# a_425_640# 0.00fF
C117 a_n787_n638# CMOS_AND_0/A 0.00fF
C118 a_n1990_n638# VDD 0.00fF
C119 CMOS_AND_0/AND a_425_640# 0.07fF
C120 x0 CMOS_AND_0/A 0.03fF
C121 a_n2140_n1548# CMOS_AND_0/A 0.03fF
C122 x3 a_n1990_n638# 0.00fF
C123 CMOS_AND_0/B CMOS_AND_0/A 0.32fF
C124 CMOS_AND_0/A CMOS_AND_1/AND 0.01fF
C125 CMOS_AND_0/A x0_bar 0.11fF
C126 s0 VDD 0.37fF
C127 CMOS_AND_0/A CMOS_AND_1/B 0.01fF
C128 a_1637_640# a_1637_30# 0.01fF
C129 a_n1990_640# x1 0.01fF
C130 CMOS_AND_0/AND a_1637_30# 0.05fF
C131 x1_bar x1 3.44fF
C132 x2_bar x1 0.17fF
C133 a_425_640# CMOS_AND_0/A 0.06fF
C134 a_425_n638# a_n787_n1548# 0.00fF
C135 x0 a_n1990_30# 0.00fF
C136 a_n2140_n1548# a_n1990_30# 0.00fF
C137 a_n1990_640# VDD 0.05fF
C138 x1_bar VDD 1.43fF
C139 a_n2290_640# x2 0.00fF
C140 x2_bar VDD 0.24fF
C141 a_n1990_30# x0_bar 0.01fF
C142 a_n1990_640# x3 0.03fF
C143 x1_bar x3 0.07fF
C144 CMOS_AND_0/A a_1637_30# 0.00fF
C145 x2_bar x3 2.86fF
C146 a_n787_30# a_n2290_640# 0.00fF
C147 a_n787_n638# x2 0.01fF
C148 x0 x2 0.09fF
C149 x1_bar a_n1990_n638# 0.00fF
C150 a_n2140_n1548# x2 0.20fF
C151 x2_bar a_n1990_n638# 0.00fF
C152 a_n787_30# a_n787_n638# 0.00fF
C153 x2 x0_bar 0.09fF
C154 a_425_n1548# CMOS_AND_0/A 0.00fF
C155 a_n787_30# x0 0.00fF
C156 CMOS_AND_0/B a_n787_30# 0.07fF
C157 x2 CMOS_AND_1/B 0.17fF
C158 a_n787_30# x0_bar 0.00fF
C159 x2 a_n2290_n1548# 0.01fF
C160 a_n2290_n638# x2 0.01fF
C161 a_n787_30# CMOS_AND_1/B 0.01fF
C162 a_425_n638# VDD 0.01fF
C163 a_n787_30# a_425_640# 0.01fF
C164 CMOS_AND_0/A a_n1990_n1548# 0.00fF
C165 a_n1990_640# x1_bar 0.00fF
C166 a_n1990_640# x2_bar 0.00fF
C167 CMOS_AND_0/A a_n787_640# 0.02fF
C168 x2_bar x1_bar 0.05fF
C169 CMOS_AND_0/A a_n787_n1548# 0.01fF
C170 CMOS_AND_0/B a_425_30# 0.00fF
C171 a_n2290_640# x3_bar 0.01fF
C172 a_425_n1548# x2 0.00fF
C173 a_425_30# a_425_640# 0.01fF
C174 x1 a_n2290_30# 0.00fF
C175 x0 x3_bar 0.32fF
C176 a_1637_640# VDD 0.06fF
C177 a_n2140_n1548# x3_bar 0.14fF
C178 CMOS_AND_0/AND VDD 0.58fF
C179 x0_bar x3_bar 0.31fF
C180 a_n787_n638# CMOS_AND_1/A 0.00fF
C181 CMOS_AND_0/A x1 0.21fF
C182 a_n2290_30# VDD 0.01fF
C183 CMOS_AND_1/B x3_bar 0.00fF
C184 CMOS_AND_1/A x0 0.00fF
C185 a_n2140_n1548# CMOS_AND_1/A 0.00fF
C186 a_425_30# a_1637_30# 0.00fF
C187 CMOS_AND_0/B CMOS_AND_1/A 0.01fF
C188 CMOS_AND_1/A CMOS_AND_1/AND 0.01fF
C189 x3 a_n2290_30# 0.01fF
C190 x2 a_n1990_n1548# 0.01fF
C191 a_n2290_n1548# x3_bar 0.01fF
C192 a_n2290_n638# x3_bar 0.01fF
C193 x2 a_n787_640# 0.00fF
C194 x2 a_n787_n1548# 0.05fF
C195 CMOS_AND_0/A VDD 1.15fF
C196 CMOS_AND_1/A CMOS_AND_1/B 0.18fF
C197 a_1637_640# s0 0.00fF
C198 a_425_n1548# a_425_30# 0.00fF
C199 x3 CMOS_AND_0/A 0.32fF
C200 CMOS_AND_0/AND s0 0.01fF
C201 a_n787_30# a_n787_640# 0.01fF
C202 a_n787_30# a_n787_n1548# 0.01fF
C203 CMOS_AND_1/A a_425_640# 0.00fF
C204 CMOS_AND_0/A a_n1990_n638# 0.00fF
C205 a_n1990_30# x1 0.00fF
C206 a_n1990_30# VDD 0.01fF
C207 x2 x1 0.05fF
C208 x3 a_n1990_30# 0.01fF
C209 x1_bar a_n2290_30# 0.00fF
C210 x2_bar a_n2290_30# 0.00fF
C211 a_n787_30# x1 0.04fF
C212 a_425_n1548# CMOS_AND_1/A 0.07fF
C213 x2 VDD 0.38fF
C214 a_n1990_640# CMOS_AND_0/A 0.03fF
C215 x1_bar CMOS_AND_0/A 0.02fF
C216 x2_bar CMOS_AND_0/A 0.21fF
C217 x3 x2 0.10fF
C218 a_n1990_n1548# x3_bar 0.01fF
C219 a_n787_30# VDD 0.51fF
C220 a_n787_n1548# x3_bar 0.00fF
C221 x2 a_n1990_n638# 0.01fF
C222 a_n787_30# x3 0.01fF
C223 a_n2290_640# x0 0.00fF
C224 CMOS_AND_1/A a_n787_n1548# 0.05fF
C225 a_n2290_640# x0_bar 0.01fF
C226 a_n2140_n1548# a_n787_n638# 0.00fF
C227 x1_bar a_n1990_30# 0.00fF
C228 x2_bar a_n1990_30# 0.00fF
C229 a_n2140_n1548# x0 0.37fF
C230 a_425_30# VDD 0.01fF
C231 CMOS_AND_0/B CMOS_AND_1/AND 0.00fF
C232 x0 x0_bar 2.88fF
C233 a_425_n638# CMOS_AND_0/A 0.00fF
C234 a_n2140_n1548# x0_bar 0.15fF
C235 a_n787_n638# CMOS_AND_1/B 0.01fF
C236 x1 x3_bar 0.07fF
C237 x0 CMOS_AND_1/B 0.01fF
C238 a_n2140_n1548# CMOS_AND_1/B 0.12fF
C239 a_n1990_640# x2 0.00fF
C240 CMOS_AND_0/B CMOS_AND_1/B 0.01fF
C241 x1_bar x2 2.97fF
C242 x2_bar x2 3.89fF
C243 CMOS_AND_1/AND CMOS_AND_1/B 0.00fF
C244 x0_bar CMOS_AND_1/B 0.01fF
C245 x0 a_n2290_n1548# 0.02fF
C246 a_n2290_n638# x0 0.01fF
C247 a_n2140_n1548# a_n2290_n1548# 0.02fF
C248 a_n2290_n638# a_n2140_n1548# 0.01fF
C249 CMOS_AND_0/B a_425_640# 0.04fF
C250 a_1637_640# CMOS_AND_0/AND 0.01fF
C251 a_n1990_640# a_n787_30# 0.00fF
C252 a_425_640# CMOS_AND_1/AND 0.00fF
C253 x3_bar VDD 0.40fF
C254 x2_bar a_n787_30# 0.08fF
C255 a_n2290_n1548# x0_bar 0.01fF
C256 a_n2290_n638# x0_bar 0.00fF
C257 x3 x3_bar 3.47fF
C258 a_n2290_n1548# CMOS_AND_1/B 0.00fF
C259 a_n2290_n638# CMOS_AND_1/B 0.00fF
C260 CMOS_AND_1/A VDD 0.53fF
C261 CMOS_AND_0/B a_1637_30# 0.00fF
C262 x3_bar a_n1990_n638# 0.01fF
C263 CMOS_AND_1/AND a_1637_30# 0.08fF
C264 CMOS_AND_0/AND CMOS_AND_0/A 0.00fF
C265 a_425_n1548# a_n787_n638# 0.00fF
C266 CMOS_AND_0/A a_n2290_30# 0.01fF
C267 a_425_n1548# CMOS_AND_1/AND 0.05fF
C268 a_425_640# a_1637_30# 0.01fF
C269 a_425_n1548# CMOS_AND_1/B 0.04fF
C270 a_n1990_640# x3_bar 0.01fF
C271 a_425_n1548# a_425_640# 0.01fF
C272 x1_bar x3_bar 0.07fF
C273 x2_bar x3_bar 0.06fF
C274 a_n787_n638# a_n787_n1548# 0.01fF
C275 x0 a_n1990_n1548# 0.02fF
C276 a_n2140_n1548# a_n1990_n1548# 0.03fF
C277 x0 a_n787_n1548# 0.00fF
C278 a_n2140_n1548# a_n787_n1548# 0.02fF
C279 CMOS_AND_0/B a_n787_640# 0.00fF
C280 a_n1990_n1548# x0_bar 0.00fF
C281 CMOS_AND_1/AND a_n787_n1548# 0.00fF
C282 a_n1990_n1548# GND 0.00fF
C283 a_n2290_n1548# GND 0.00fF
C284 a_425_n638# GND 0.03fF
C285 a_n787_n638# GND 0.03fF
C286 a_n1990_n638# GND 0.02fF
C287 a_n2290_n638# GND 0.01fF
C288 a_425_n1548# GND 0.55fF
C289 CMOS_AND_1/B GND 0.93fF
C290 a_n787_n1548# GND 0.50fF
C291 x1_bar GND 6.70fF
C292 a_n2140_n1548# GND 0.59fF
C293 CMOS_AND_1/A GND 0.96fF
C294 x2 GND 8.05fF
C295 a_425_30# GND 0.03fF
C296 a_n1990_30# GND 0.02fF
C297 a_n2290_30# GND 0.01fF
C298 s0 GND 0.58fF
C299 a_1637_640# GND 0.02fF
C300 a_n787_640# GND 0.01fF
C301 a_n1990_640# GND 0.00fF
C302 a_n2290_640# GND 0.00fF
C303 a_1637_30# GND 0.67fF
C304 CMOS_AND_1/AND GND 1.29fF
C305 CMOS_AND_0/AND GND 0.64fF
C306 a_425_640# GND 0.50fF
C307 CMOS_AND_0/A GND 1.60fF
C308 CMOS_AND_0/B GND 0.57fF
C309 a_n787_30# GND 0.61fF
C310 x2_bar GND 8.02fF
C311 x1 GND 6.48fF
C312 x0_bar GND 3.60fF
C313 x0 GND 2.82fF
C314 x3_bar GND 5.55fF
C315 x3 GND 1.80fF
C316 VDD GND 26.54fF
C317 x3_bar.t0 GND 0.26fF
C318 x3_bar.t1 GND 0.26fF
C319 x3_bar.n0 GND 0.70fF $ **FLOATING
C320 x3_bar.t3 GND 0.36fF
C321 x3_bar.t2 GND 0.32fF
C322 CMOS_XNOR_0/A_bar GND 0.55fF $ **FLOATING
C323 x3_bar.n1 GND 4.79fF $ **FLOATING
C324 x2_bar.t0 GND 0.29fF
C325 x2_bar.t1 GND 0.24fF
C326 x3.t1 GND 0.63fF
C327 x3.t0 GND 0.43fF
C328 x3.t2 GND 0.09fF
C329 x3.t3 GND 0.22fF
C330 x3.n0 GND 0.25fF $ **FLOATING
C331 CMOS_XNOR_0/A GND 0.25fF $ **FLOATING
C332 x3.n1 GND 3.86fF $ **FLOATING
C333 x0_bar.t2 GND 0.29fF
C334 x0_bar.t3 GND 0.26fF
C335 x0_bar.t0 GND 0.21fF
C336 x0_bar.t1 GND 0.21fF
C337 x0_bar.n0 GND 0.57fF $ **FLOATING
C338 CMOS_XNOR_0/B_bar GND 0.33fF $ **FLOATING
C339 x0_bar.n1 GND 3.92fF $ **FLOATING
C340 x1.t0 GND 0.16fF
C341 x1.t1 GND 0.11fF
C342 x1.n0 GND 0.23fF $ **FLOATING
C343 x1_bar.t1 GND 0.12fF
C344 x1_bar.t0 GND 0.18fF
C345 x1_bar.n0 GND 0.25fF $ **FLOATING
C346 x2.t0 GND 0.30fF
C347 x2.t1 GND 0.25fF
C348 x0.t1 GND 0.16fF
C349 x0.t3 GND 0.06fF
C350 x0.n0 GND 0.18fF $ **FLOATING
C351 x0.t2 GND 0.45fF
C352 x0.t0 GND 0.30fF
C353 CMOS_XNOR_0/B GND 0.45fF $ **FLOATING
C354 x0.n1 GND 2.73fF $ **FLOATING
C355 VDD.t20 GND 0.07fF
C356 VDD.t30 GND 0.07fF
C357 CMOS_AND_0/VDD GND 0.01fF $ **FLOATING
C358 VDD.t15 GND 0.07fF
C359 VDD.t24 GND 0.07fF
C360 CMOS_OR_0/VDD GND 0.01fF $ **FLOATING
C361 VDD.t32 GND 0.07fF
C362 VDD.n0 GND 0.18fF $ **FLOATING
C363 VDD.n1 GND 0.02fF $ **FLOATING
C364 VDD.n2 GND 0.01fF $ **FLOATING
C365 VDD.n3 GND 0.14fF $ **FLOATING
C366 VDD.t31 GND 0.09fF
C367 VDD.n4 GND 0.09fF $ **FLOATING
C368 VDD.n5 GND 0.02fF $ **FLOATING
C369 VDD.n6 GND 0.01fF $ **FLOATING
C370 VDD.n7 GND 0.05fF $ **FLOATING
C371 VDD.n8 GND 0.34fF $ **FLOATING
C372 VDD.n9 GND 0.16fF $ **FLOATING
C373 VDD.n10 GND 0.02fF $ **FLOATING
C374 VDD.n11 GND 0.01fF $ **FLOATING
C375 VDD.n12 GND 0.01fF $ **FLOATING
C376 VDD.n13 GND 0.16fF $ **FLOATING
C377 VDD.n14 GND 0.02fF $ **FLOATING
C378 VDD.n15 GND 0.01fF $ **FLOATING
C379 VDD.n16 GND 0.02fF $ **FLOATING
C380 VDD.n17 GND 0.16fF $ **FLOATING
C381 VDD.n18 GND 0.02fF $ **FLOATING
C382 VDD.n19 GND 0.01fF $ **FLOATING
C383 VDD.n20 GND 0.02fF $ **FLOATING
C384 VDD.n21 GND 0.01fF $ **FLOATING
C385 VDD.n22 GND 0.16fF $ **FLOATING
C386 VDD.n23 GND 0.02fF $ **FLOATING
C387 VDD.n24 GND 0.01fF $ **FLOATING
C388 VDD.t18 GND 0.08fF
C389 VDD.n25 GND 0.10fF $ **FLOATING
C390 VDD.n26 GND 0.02fF $ **FLOATING
C391 VDD.n27 GND 0.01fF $ **FLOATING
C392 VDD.n28 GND 0.01fF $ **FLOATING
C393 VDD.n29 GND 0.14fF $ **FLOATING
C394 VDD.n30 GND 0.02fF $ **FLOATING
C395 VDD.n31 GND 0.01fF $ **FLOATING
C396 VDD.n32 GND 0.02fF $ **FLOATING
C397 VDD.t23 GND 0.09fF
C398 VDD.n33 GND 0.10fF $ **FLOATING
C399 VDD.n34 GND 0.02fF $ **FLOATING
C400 VDD.n35 GND 0.01fF $ **FLOATING
C401 VDD.n36 GND 0.02fF $ **FLOATING
C402 VDD.n37 GND 0.17fF $ **FLOATING
C403 VDD.n38 GND 0.02fF $ **FLOATING
C404 VDD.n39 GND 0.01fF $ **FLOATING
C405 VDD.n40 GND 0.01fF $ **FLOATING
C406 VDD.n41 GND 0.34fF $ **FLOATING
C407 VDD.n42 GND 0.17fF $ **FLOATING
C408 VDD.n43 GND 0.06fF $ **FLOATING
C409 VDD.n44 GND 0.14fF $ **FLOATING
C410 VDD.n45 GND 0.06fF $ **FLOATING
C411 VDD.n46 GND 0.18fF $ **FLOATING
C412 VDD.n47 GND 0.02fF $ **FLOATING
C413 VDD.n48 GND 0.01fF $ **FLOATING
C414 VDD.n49 GND 0.02fF $ **FLOATING
C415 VDD.t14 GND 0.09fF
C416 VDD.n50 GND 0.09fF $ **FLOATING
C417 VDD.n51 GND 0.02fF $ **FLOATING
C418 VDD.n52 GND 0.01fF $ **FLOATING
C419 VDD.n53 GND 0.02fF $ **FLOATING
C420 VDD.n54 GND 0.34fF $ **FLOATING
C421 VDD.n55 GND 0.16fF $ **FLOATING
C422 VDD.n56 GND 0.02fF $ **FLOATING
C423 VDD.n57 GND 0.01fF $ **FLOATING
C424 VDD.n58 GND 0.01fF $ **FLOATING
C425 VDD.n59 GND 0.16fF $ **FLOATING
C426 VDD.n60 GND 0.02fF $ **FLOATING
C427 VDD.n61 GND 0.01fF $ **FLOATING
C428 VDD.n62 GND 0.02fF $ **FLOATING
C429 VDD.n63 GND 0.16fF $ **FLOATING
C430 VDD.n64 GND 0.02fF $ **FLOATING
C431 VDD.n65 GND 0.01fF $ **FLOATING
C432 VDD.n66 GND 0.02fF $ **FLOATING
C433 VDD.t12 GND 0.07fF
C434 VDD.n67 GND 0.33fF $ **FLOATING
C435 VDD.n68 GND 0.01fF $ **FLOATING
C436 VDD.n69 GND 0.16fF $ **FLOATING
C437 VDD.n70 GND 0.02fF $ **FLOATING
C438 VDD.n71 GND 0.01fF $ **FLOATING
C439 VDD.t11 GND 0.08fF
C440 VDD.n72 GND 0.10fF $ **FLOATING
C441 VDD.n73 GND 0.02fF $ **FLOATING
C442 VDD.n74 GND 0.01fF $ **FLOATING
C443 VDD.n75 GND 0.01fF $ **FLOATING
C444 VDD.n76 GND 0.14fF $ **FLOATING
C445 VDD.n77 GND 0.02fF $ **FLOATING
C446 VDD.n78 GND 0.01fF $ **FLOATING
C447 VDD.n79 GND 0.02fF $ **FLOATING
C448 VDD.t29 GND 0.09fF
C449 VDD.n80 GND 0.10fF $ **FLOATING
C450 VDD.n81 GND 0.02fF $ **FLOATING
C451 VDD.n82 GND 0.01fF $ **FLOATING
C452 VDD.n83 GND 0.02fF $ **FLOATING
C453 VDD.n84 GND 0.17fF $ **FLOATING
C454 VDD.n85 GND 0.02fF $ **FLOATING
C455 VDD.n86 GND 0.01fF $ **FLOATING
C456 VDD.n87 GND 0.01fF $ **FLOATING
C457 VDD.n88 GND 0.34fF $ **FLOATING
C458 VDD.n89 GND 0.17fF $ **FLOATING
C459 VDD.n90 GND 0.06fF $ **FLOATING
C460 VDD.n91 GND 0.14fF $ **FLOATING
C461 VDD.n92 GND 0.06fF $ **FLOATING
C462 VDD.n93 GND 0.18fF $ **FLOATING
C463 VDD.n94 GND 0.02fF $ **FLOATING
C464 VDD.n95 GND 0.01fF $ **FLOATING
C465 VDD.n96 GND 0.02fF $ **FLOATING
C466 VDD.t19 GND 0.09fF
C467 VDD.n97 GND 0.09fF $ **FLOATING
C468 VDD.n98 GND 0.02fF $ **FLOATING
C469 VDD.n99 GND 0.01fF $ **FLOATING
C470 VDD.n100 GND 0.02fF $ **FLOATING
C471 VDD.n101 GND 0.34fF $ **FLOATING
C472 VDD.n102 GND 0.16fF $ **FLOATING
C473 VDD.n103 GND 0.02fF $ **FLOATING
C474 VDD.n104 GND 0.01fF $ **FLOATING
C475 VDD.n105 GND 0.01fF $ **FLOATING
C476 VDD.n106 GND 0.16fF $ **FLOATING
C477 VDD.n107 GND 0.02fF $ **FLOATING
C478 VDD.n108 GND 0.01fF $ **FLOATING
C479 VDD.n109 GND 0.02fF $ **FLOATING
C480 VDD.n110 GND 0.16fF $ **FLOATING
C481 VDD.n111 GND 0.02fF $ **FLOATING
C482 VDD.n112 GND 0.01fF $ **FLOATING
C483 VDD.n113 GND 0.02fF $ **FLOATING
C484 VDD.n114 GND 0.16fF $ **FLOATING
C485 VDD.n115 GND 0.02fF $ **FLOATING
C486 VDD.n116 GND 0.01fF $ **FLOATING
C487 VDD.n117 GND 0.01fF $ **FLOATING
C488 VDD.t38 GND 0.07fF
C489 VDD.n118 GND 0.13fF $ **FLOATING
C490 VDD.t8 GND 0.07fF
C491 VDD.t6 GND 0.08fF
C492 VDD.n119 GND 0.12fF $ **FLOATING
C493 VDD.n120 GND 0.02fF $ **FLOATING
C494 VDD.t40 GND 0.07fF
C495 VDD.t1 GND 0.07fF
C496 CMOS_XNOR_0/VDD GND 0.01fF $ **FLOATING
C497 VDD.t3 GND 0.07fF
C498 VDD.t22 GND 0.07fF
C499 VDD.t5 GND 0.07fF
C500 CMOS_AND_2/VDD GND 0.01fF $ **FLOATING
C501 VDD.t26 GND 0.07fF
C502 VDD.t28 GND 0.07fF
C503 CMOS_AND_1/VDD GND 0.01fF $ **FLOATING
C504 VDD.t34 GND 0.07fF
C505 VDD.n121 GND 0.18fF $ **FLOATING
C506 VDD.n122 GND 0.02fF $ **FLOATING
C507 VDD.n123 GND 0.01fF $ **FLOATING
C508 VDD.n124 GND 0.14fF $ **FLOATING
C509 VDD.t33 GND 0.09fF
C510 VDD.n125 GND 0.09fF $ **FLOATING
C511 VDD.n126 GND 0.02fF $ **FLOATING
C512 VDD.n127 GND 0.01fF $ **FLOATING
C513 VDD.n128 GND 0.05fF $ **FLOATING
C514 VDD.n129 GND 0.34fF $ **FLOATING
C515 VDD.n130 GND 0.16fF $ **FLOATING
C516 VDD.n131 GND 0.02fF $ **FLOATING
C517 VDD.n132 GND 0.01fF $ **FLOATING
C518 VDD.n133 GND 0.01fF $ **FLOATING
C519 VDD.n134 GND 0.16fF $ **FLOATING
C520 VDD.n135 GND 0.02fF $ **FLOATING
C521 VDD.n136 GND 0.01fF $ **FLOATING
C522 VDD.n137 GND 0.02fF $ **FLOATING
C523 VDD.n138 GND 0.16fF $ **FLOATING
C524 VDD.n139 GND 0.02fF $ **FLOATING
C525 VDD.n140 GND 0.01fF $ **FLOATING
C526 VDD.n141 GND 0.02fF $ **FLOATING
C527 VDD.t36 GND 0.07fF
C528 VDD.n142 GND 0.33fF $ **FLOATING
C529 VDD.n143 GND 0.01fF $ **FLOATING
C530 VDD.n144 GND 0.16fF $ **FLOATING
C531 VDD.n145 GND 0.02fF $ **FLOATING
C532 VDD.n146 GND 0.01fF $ **FLOATING
C533 VDD.t35 GND 0.08fF
C534 VDD.n147 GND 0.10fF $ **FLOATING
C535 VDD.n148 GND 0.02fF $ **FLOATING
C536 VDD.n149 GND 0.01fF $ **FLOATING
C537 VDD.n150 GND 0.01fF $ **FLOATING
C538 VDD.n151 GND 0.14fF $ **FLOATING
C539 VDD.n152 GND 0.02fF $ **FLOATING
C540 VDD.n153 GND 0.01fF $ **FLOATING
C541 VDD.n154 GND 0.02fF $ **FLOATING
C542 VDD.t27 GND 0.09fF
C543 VDD.n155 GND 0.10fF $ **FLOATING
C544 VDD.n156 GND 0.02fF $ **FLOATING
C545 VDD.n157 GND 0.01fF $ **FLOATING
C546 VDD.n158 GND 0.02fF $ **FLOATING
C547 VDD.n159 GND 0.17fF $ **FLOATING
C548 VDD.n160 GND 0.02fF $ **FLOATING
C549 VDD.n161 GND 0.01fF $ **FLOATING
C550 VDD.n162 GND 0.01fF $ **FLOATING
C551 VDD.n163 GND 0.34fF $ **FLOATING
C552 VDD.n164 GND 0.17fF $ **FLOATING
C553 VDD.n165 GND 0.06fF $ **FLOATING
C554 VDD.n166 GND 0.14fF $ **FLOATING
C555 VDD.n167 GND 0.06fF $ **FLOATING
C556 VDD.n168 GND 0.18fF $ **FLOATING
C557 VDD.n169 GND 0.02fF $ **FLOATING
C558 VDD.n170 GND 0.01fF $ **FLOATING
C559 VDD.n171 GND 0.02fF $ **FLOATING
C560 VDD.t25 GND 0.09fF
C561 VDD.n172 GND 0.09fF $ **FLOATING
C562 VDD.n173 GND 0.02fF $ **FLOATING
C563 VDD.n174 GND 0.01fF $ **FLOATING
C564 VDD.n175 GND 0.02fF $ **FLOATING
C565 VDD.n176 GND 0.34fF $ **FLOATING
C566 VDD.n177 GND 0.16fF $ **FLOATING
C567 VDD.n178 GND 0.02fF $ **FLOATING
C568 VDD.n179 GND 0.01fF $ **FLOATING
C569 VDD.n180 GND 0.01fF $ **FLOATING
C570 VDD.n181 GND 0.16fF $ **FLOATING
C571 VDD.n182 GND 0.02fF $ **FLOATING
C572 VDD.n183 GND 0.01fF $ **FLOATING
C573 VDD.n184 GND 0.02fF $ **FLOATING
C574 VDD.n185 GND 0.16fF $ **FLOATING
C575 VDD.n186 GND 0.02fF $ **FLOATING
C576 VDD.n187 GND 0.01fF $ **FLOATING
C577 VDD.n188 GND 0.02fF $ **FLOATING
C578 VDD.t17 GND 0.07fF
C579 VDD.n189 GND 0.33fF $ **FLOATING
C580 VDD.n190 GND 0.01fF $ **FLOATING
C581 VDD.n191 GND 0.16fF $ **FLOATING
C582 VDD.n192 GND 0.02fF $ **FLOATING
C583 VDD.n193 GND 0.01fF $ **FLOATING
C584 VDD.t16 GND 0.08fF
C585 VDD.n194 GND 0.10fF $ **FLOATING
C586 VDD.n195 GND 0.02fF $ **FLOATING
C587 VDD.n196 GND 0.01fF $ **FLOATING
C588 VDD.n197 GND 0.01fF $ **FLOATING
C589 VDD.n198 GND 0.14fF $ **FLOATING
C590 VDD.n199 GND 0.02fF $ **FLOATING
C591 VDD.n200 GND 0.01fF $ **FLOATING
C592 VDD.n201 GND 0.02fF $ **FLOATING
C593 VDD.t4 GND 0.09fF
C594 VDD.n202 GND 0.10fF $ **FLOATING
C595 VDD.n203 GND 0.02fF $ **FLOATING
C596 VDD.n204 GND 0.01fF $ **FLOATING
C597 VDD.n205 GND 0.02fF $ **FLOATING
C598 VDD.n206 GND 0.17fF $ **FLOATING
C599 VDD.n207 GND 0.02fF $ **FLOATING
C600 VDD.n208 GND 0.01fF $ **FLOATING
C601 VDD.n209 GND 0.01fF $ **FLOATING
C602 VDD.n210 GND 0.34fF $ **FLOATING
C603 VDD.n211 GND 0.17fF $ **FLOATING
C604 VDD.n212 GND 0.05fF $ **FLOATING
C605 VDD.n213 GND 0.15fF $ **FLOATING
C606 VDD.n214 GND 0.06fF $ **FLOATING
C607 VDD.n215 GND 0.18fF $ **FLOATING
C608 VDD.n216 GND 0.02fF $ **FLOATING
C609 VDD.n217 GND 0.01fF $ **FLOATING
C610 VDD.n218 GND 0.02fF $ **FLOATING
C611 VDD.t21 GND 0.09fF
C612 VDD.n219 GND 0.10fF $ **FLOATING
C613 VDD.n220 GND 0.02fF $ **FLOATING
C614 VDD.n221 GND 0.01fF $ **FLOATING
C615 VDD.n222 GND 0.02fF $ **FLOATING
C616 VDD.n223 GND 0.34fF $ **FLOATING
C617 VDD.n224 GND 0.16fF $ **FLOATING
C618 VDD.n225 GND 0.02fF $ **FLOATING
C619 VDD.n226 GND 0.01fF $ **FLOATING
C620 VDD.n227 GND 0.01fF $ **FLOATING
C621 VDD.n228 GND 0.16fF $ **FLOATING
C622 VDD.n229 GND 0.02fF $ **FLOATING
C623 VDD.n230 GND 0.01fF $ **FLOATING
C624 VDD.n231 GND 0.02fF $ **FLOATING
C625 VDD.n232 GND 0.16fF $ **FLOATING
C626 VDD.n233 GND 0.02fF $ **FLOATING
C627 VDD.n234 GND 0.01fF $ **FLOATING
C628 VDD.n235 GND 0.02fF $ **FLOATING
C629 VDD.n236 GND 0.16fF $ **FLOATING
C630 VDD.n237 GND 0.02fF $ **FLOATING
C631 VDD.n238 GND 0.01fF $ **FLOATING
C632 VDD.n239 GND 0.01fF $ **FLOATING
C633 VDD.n240 GND 0.34fF $ **FLOATING
C634 VDD.t2 GND 0.08fF
C635 VDD.n241 GND 0.10fF $ **FLOATING
C636 VDD.n242 GND 0.02fF $ **FLOATING
C637 VDD.n243 GND 0.01fF $ **FLOATING
C638 VDD.n244 GND 0.01fF $ **FLOATING
C639 VDD.n245 GND 0.13fF $ **FLOATING
C640 VDD.n246 GND 0.02fF $ **FLOATING
C641 VDD.n247 GND 0.01fF $ **FLOATING
C642 VDD.n248 GND 0.02fF $ **FLOATING
C643 VDD.t41 GND 0.08fF
C644 VDD.n249 GND 0.11fF $ **FLOATING
C645 VDD.n250 GND 0.02fF $ **FLOATING
C646 VDD.n251 GND 0.01fF $ **FLOATING
C647 VDD.n252 GND 0.02fF $ **FLOATING
C648 VDD.n253 GND 0.13fF $ **FLOATING
C649 VDD.n254 GND 0.02fF $ **FLOATING
C650 VDD.n255 GND 0.01fF $ **FLOATING
C651 VDD.n256 GND 0.02fF $ **FLOATING
C652 VDD.n257 GND 0.01fF $ **FLOATING
C653 VDD.n258 GND 0.12fF $ **FLOATING
C654 VDD.n259 GND 0.02fF $ **FLOATING
C655 VDD.n260 GND 0.01fF $ **FLOATING
C656 VDD.t13 GND 0.08fF
C657 VDD.n261 GND 0.12fF $ **FLOATING
C658 VDD.n262 GND 0.02fF $ **FLOATING
C659 VDD.n263 GND 0.01fF $ **FLOATING
C660 VDD.n264 GND 0.01fF $ **FLOATING
C661 VDD.n265 GND 0.12fF $ **FLOATING
C662 VDD.n266 GND 0.02fF $ **FLOATING
C663 VDD.n267 GND 0.01fF $ **FLOATING
C664 VDD.n268 GND 0.02fF $ **FLOATING
C665 VDD.t0 GND 0.08fF
C666 VDD.n269 GND 0.12fF $ **FLOATING
C667 VDD.n270 GND 0.02fF $ **FLOATING
C668 VDD.n271 GND 0.01fF $ **FLOATING
C669 VDD.n272 GND 0.01fF $ **FLOATING
C670 VDD.n273 GND 0.34fF $ **FLOATING
C671 VDD.n274 GND 0.18fF $ **FLOATING
C672 VDD.n275 GND 0.02fF $ **FLOATING
C673 VDD.n276 GND 0.01fF $ **FLOATING
C674 VDD.n277 GND 0.01fF $ **FLOATING
C675 VDD.n278 GND 0.10fF $ **FLOATING
C676 VDD.n279 GND 0.32fF $ **FLOATING
C677 VDD.n280 GND 0.31fF $ **FLOATING
C678 VDD.n281 GND 0.10fF $ **FLOATING
C679 VDD.n282 GND 0.02fF $ **FLOATING
C680 VDD.n283 GND 0.18fF $ **FLOATING
C681 VDD.n284 GND 0.02fF $ **FLOATING
C682 VDD.n285 GND 0.01fF $ **FLOATING
C683 VDD.n286 GND 0.01fF $ **FLOATING
C684 VDD.n287 GND 0.34fF $ **FLOATING
C685 VDD.t39 GND 0.08fF
C686 VDD.n288 GND 0.12fF $ **FLOATING
C687 VDD.n289 GND 0.02fF $ **FLOATING
C688 VDD.n290 GND 0.01fF $ **FLOATING
C689 VDD.n291 GND 0.01fF $ **FLOATING
C690 VDD.n292 GND 0.12fF $ **FLOATING
C691 VDD.n293 GND 0.02fF $ **FLOATING
C692 VDD.n294 GND 0.01fF $ **FLOATING
C693 VDD.n295 GND 0.02fF $ **FLOATING
C694 VDD.n296 GND 0.01fF $ **FLOATING
C695 VDD.n297 GND 0.12fF $ **FLOATING
C696 VDD.n298 GND 0.02fF $ **FLOATING
C697 VDD.n299 GND 0.01fF $ **FLOATING
C698 VDD.n300 GND 0.01fF $ **FLOATING
C699 VDD.n301 GND 0.01fF $ **FLOATING
C700 VDD.n302 GND 0.13fF $ **FLOATING
C701 VDD.n303 GND 0.02fF $ **FLOATING
C702 VDD.n304 GND 0.01fF $ **FLOATING
C703 VDD.n305 GND 0.02fF $ **FLOATING
C704 VDD.t10 GND 0.08fF
C705 VDD.n306 GND 0.11fF $ **FLOATING
C706 VDD.n307 GND 0.02fF $ **FLOATING
C707 VDD.n308 GND 0.01fF $ **FLOATING
C708 VDD.n309 GND 0.02fF $ **FLOATING
C709 VDD.n310 GND 0.13fF $ **FLOATING
C710 VDD.n311 GND 0.02fF $ **FLOATING
C711 VDD.n312 GND 0.01fF $ **FLOATING
C712 VDD.n313 GND 0.02fF $ **FLOATING
C713 VDD.t7 GND 0.08fF
C714 VDD.n314 GND 0.11fF $ **FLOATING
C715 VDD.n315 GND 0.02fF $ **FLOATING
C716 VDD.n316 GND 0.01fF $ **FLOATING
C717 VDD.n317 GND 0.01fF $ **FLOATING
C718 VDD.n318 GND 0.34fF $ **FLOATING
C719 VDD.n319 GND 0.19fF $ **FLOATING
C720 VDD.n320 GND 0.02fF $ **FLOATING
C721 VDD.n321 GND 0.01fF $ **FLOATING
C722 VDD.n322 GND 0.01fF $ **FLOATING
C723 VDD.n323 GND 0.10fF $ **FLOATING
C724 VDD.n324 GND 0.17fF $ **FLOATING
C725 VDD.n325 GND 0.10fF $ **FLOATING
C726 VDD.n326 GND 0.34fF $ **FLOATING
C727 VDD.n327 GND 0.17fF $ **FLOATING
C728 VDD.n328 GND 0.02fF $ **FLOATING
C729 VDD.n329 GND 0.01fF $ **FLOATING
C730 VDD.n330 GND 0.01fF $ **FLOATING
C731 VDD.t37 GND 0.09fF
C732 VDD.n331 GND 0.10fF $ **FLOATING
C733 VDD.n332 GND 0.02fF $ **FLOATING
C734 VDD.n333 GND 0.01fF $ **FLOATING
C735 VDD.n334 GND 0.02fF $ **FLOATING
C736 VDD.n335 GND 0.14fF $ **FLOATING
C737 VDD.n336 GND 0.02fF $ **FLOATING
C738 VDD.n337 GND 0.01fF $ **FLOATING
C739 VDD.n338 GND 0.02fF $ **FLOATING
C740 VDD.t9 GND 0.08fF
C741 VDD.n339 GND 0.10fF $ **FLOATING
C742 VDD.n340 GND 0.02fF $ **FLOATING
C743 VDD.n341 GND 0.01fF $ **FLOATING
C744 VDD.n342 GND 0.01fF $ **FLOATING
C745 CMOS_OR_1/VDD GND 0.01fF $ **FLOATING
.ends

