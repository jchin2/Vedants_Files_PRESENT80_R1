.subckt Buffer A VP VN OUT
*.PININFO A:I VP:B VN:B OUT:O
x1 VP A net1 VN INV_VP_VN
x2 VP net1 OUT VN INV_VP_VN
.ends

* expanding   symbol:  INV_VP_VN.sym # of pins=4
* sym_path: /home/jchin2/skywater_stuff/INV_VP_VN.sym
* sch_path: /home/jchin2/skywater_stuff/INV_VP_VN.sch
.subckt INV_VP_VN  VP A INV VN
*.PININFO A:I INV:O VP:B VN:B
XM1 INV A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 INV A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

** flattened .save nodes
.end
