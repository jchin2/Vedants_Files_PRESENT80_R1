magic
tech sky130A
magscale 1 2
timestamp 1674172301
<< locali >>
rect -4582 907 -3870 947
rect -4468 807 -3870 847
rect -1591 839 -1303 879
rect -4810 707 -3870 747
rect -4696 607 -3870 647
rect -1591 507 -1551 839
rect 272 692 661 732
rect 150 537 158 577
rect -1284 417 -1230 457
rect -1576 249 -1496 268
rect -1284 249 -1244 417
rect 272 407 312 692
rect 2180 537 2337 577
rect 2180 417 2183 457
rect 150 367 312 407
rect -1576 246 -1244 249
rect -1576 212 -1553 246
rect -1519 212 -1244 246
rect -1576 209 -1244 212
rect -1576 188 -1496 209
rect -2490 -23 -1230 17
rect -3910 -163 -3847 -83
rect -2490 -263 -1230 -223
rect -1576 -446 -1496 -427
rect -1576 -449 -1244 -446
rect -1576 -483 -1553 -449
rect -1519 -483 -1244 -449
rect -1576 -486 -1244 -483
rect -1576 -507 -1496 -486
rect -1284 -663 -1244 -486
rect 150 -653 158 -613
rect -1590 -703 -1385 -663
rect -1284 -703 -1230 -663
rect 2180 -703 2183 -663
rect -4012 -893 -3870 -853
rect -4126 -993 -3870 -953
rect -4240 -1093 -3870 -1053
rect -1425 -1085 -1385 -703
rect 130 -773 500 -733
rect 130 -823 170 -773
rect 2180 -823 2254 -783
rect 272 -873 500 -833
rect 272 -941 312 -873
rect 238 -981 312 -941
rect -1425 -1125 -1318 -1085
rect -4354 -1193 -3870 -1153
rect 134 -1557 508 -1517
rect -4240 -1903 -3719 -1863
rect 134 -1930 174 -1557
rect 2214 -1644 2254 -823
rect 2297 -1551 2337 537
rect 2297 -1591 2453 -1551
rect 2214 -1684 2539 -1644
rect -4810 -2023 -3719 -1983
rect -4126 -2133 -3719 -2093
rect -1377 -2163 -1369 -2123
rect -4354 -2213 -3719 -2173
rect 176 -2186 290 -2146
rect 176 -2243 216 -2186
rect 2351 -2214 2385 -2174
rect -4696 -2293 -3719 -2253
rect -1739 -2283 -1536 -2243
rect 11 -2283 216 -2243
rect -4012 -2393 -3719 -2353
rect -1576 -2363 -1536 -2283
rect 2499 -2294 2539 -1684
rect 2351 -2334 2539 -2294
rect -1576 -2403 -1369 -2363
rect 11 -2453 25 -2413
rect 128 -2803 168 -2587
rect -439 -2843 168 -2803
rect 279 -2844 1121 -2804
rect -3898 -2983 -3729 -2903
<< viali >>
rect -1553 212 -1519 246
rect -1553 -483 -1519 -449
<< metal1 >>
rect -1590 1007 -1230 1107
rect -4890 -3000 -4810 947
rect -4776 -3000 -4696 947
rect -4662 -3000 -4582 947
rect -4548 -3000 -4468 947
rect -4434 -3000 -4354 947
rect -4320 -3000 -4240 947
rect -4206 -3000 -4126 947
rect -4092 -2999 -4012 947
rect -1010 717 -970 889
rect 238 812 420 852
rect 238 711 480 751
rect -1299 452 -1259 710
rect 440 647 480 711
rect 158 471 420 511
rect -1510 412 -1259 452
rect -3960 -146 -3916 -100
rect -3978 -2983 -3898 -163
rect -1590 -173 -1230 -73
rect 150 -173 661 -73
rect 238 -653 480 -613
rect -1510 -793 -1259 -753
rect -1299 -954 -1259 -793
rect 440 -913 480 -653
rect -1010 -1135 -970 -963
rect 238 -1088 420 -1048
rect -1591 -1353 -1230 -1253
rect 280 -1353 500 -1253
rect 280 -1483 380 -1353
rect -89 -1583 380 -1483
rect -89 -1713 11 -1583
rect -3835 -1813 -3729 -1713
rect 45 -2078 290 -2038
rect -1718 -2163 -1457 -2123
rect -1718 -2342 -1678 -2163
rect 45 -2393 85 -2078
rect 1921 -2354 1961 -2232
rect -1729 -2993 -1369 -2893
rect 11 -2993 361 -2893
<< metal2 >>
rect -3835 -1724 -3755 1200
rect -3699 -2783 -3659 1200
rect -1238 821 158 861
rect -1238 750 106 790
rect 66 749 106 750
rect 66 709 159 749
rect 10 -981 158 -941
rect 10 -994 50 -981
rect -1238 -1034 50 -994
rect -1238 -1107 158 -1067
rect 266 -1160 306 1200
rect 222 -1200 306 -1160
rect 133 -2507 173 -2010
rect 222 -2785 262 -1200
rect 381 -1724 421 1200
rect 528 -1497 568 1200
rect 2100 1097 2180 1200
rect 2263 417 2379 457
rect 2080 -323 2160 77
rect 2183 -1964 2223 -723
rect 2339 -1854 2379 417
rect 370 -2076 463 -2036
rect 423 -2084 463 -2076
rect 423 -2124 791 -2084
rect 290 -2212 1901 -2172
rect 2493 -2174 2533 -1610
rect 2448 -2214 2533 -2174
rect 371 -2300 2401 -2260
rect 371 -2404 2401 -2364
<< metal3 >>
rect -4002 899 -1040 959
rect -4116 198 -1586 258
rect -4458 -496 -1486 -436
rect -4572 -1205 -1040 -1145
use EESPFAL_3in_NAND_v2  EESPFAL_3in_NAND_v2_0
timestamp 1502773982
transform 1 0 -1099 0 1 -3393
box -2670 374 -590 1730
use EESPFAL_3in_NOR_v2  EESPFAL_3in_NOR_v2_0
timestamp 1502773982
transform -1 0 61 0 1 -3324
box -2340 304 -260 1660
use EESPFAL_INV4  EESPFAL_INV4_0
timestamp 1502773982
transform 1 0 1961 0 1 -3613
box -3390 594 -1900 1950
use EESPFAL_INV4  EESPFAL_INV4_1
timestamp 1502773982
transform 1 0 2100 0 -1 547
box -3390 594 -1900 1950
use EESPFAL_INV4  EESPFAL_INV4_2
timestamp 1502773982
transform 1 0 2100 0 1 -793
box -3390 594 -1900 1950
use EESPFAL_NAND_v3  EESPFAL_NAND_v3_0
timestamp 1502773982
transform 1 0 1409 0 1 481
box -949 -680 811 676
use EESPFAL_NAND_v3  EESPFAL_NAND_v3_1
timestamp 1502773982
transform 1 0 1409 0 -1 -727
box -949 -680 811 676
use EESPFAL_XOR_v3  EESPFAL_XOR_v3_0
timestamp 1502773982
transform 1 0 -2580 0 1 -343
box -1330 144 1030 1500
use EESPFAL_XOR_v3  EESPFAL_XOR_v3_1
timestamp 1502773982
transform 1 0 -2580 0 -1 97
box -1330 144 1030 1500
use Li_via_M1  Li_via_M1_0
timestamp 1502773982
transform 1 0 -4280 0 1 -1075
box -40 -38 40 42
use Li_via_M1  Li_via_M1_1
timestamp 1502773982
transform 1 0 198 0 1 -635
box -40 -38 40 42
use Li_via_M1  Li_via_M1_2
timestamp 1502773982
transform 1 0 460 0 1 -1076
box -40 -38 40 42
use Li_via_M1  Li_via_M1_3
timestamp 1502773982
transform 1 0 1941 0 1 -2396
box -40 -38 40 42
use Li_via_M1  Li_via_M1_4
timestamp 1502773982
transform 1 0 65 0 1 -2435
box -40 -38 40 42
use Li_via_M1  Li_via_M1_5
timestamp 1502773982
transform 1 0 -1417 0 1 -2145
box -40 -38 40 42
use Li_via_M1  Li_via_M1_6
timestamp 1502773982
transform 1 0 -1699 0 1 -2384
box -40 -38 40 42
use Li_via_M1  Li_via_M1_7
timestamp 1502773982
transform 1 0 -3938 0 1 -2945
box -40 -38 40 42
use Li_via_M1  Li_via_M1_8
timestamp 1502773982
transform 1 0 -4280 0 1 -1885
box -40 -38 40 42
use Li_via_M1  Li_via_M1_9
timestamp 1502773982
transform 1 0 -4394 0 1 -2181
box -40 -38 40 42
use Li_via_M1  Li_via_M1_10
timestamp 1502773982
transform 1 0 -4052 0 1 -2375
box -40 -38 40 42
use Li_via_M1  Li_via_M1_11
timestamp 1502773982
transform 1 0 -4394 0 1 -1175
box -40 -38 40 42
use Li_via_M1  Li_via_M1_12
timestamp 1502773982
transform 1 0 -4850 0 1 -2005
box -40 -38 40 42
use Li_via_M1  Li_via_M1_13
timestamp 1502773982
transform 1 0 -4736 0 1 -2275
box -40 -38 40 42
use Li_via_M1  Li_via_M1_14
timestamp 1502773982
transform 1 0 -4166 0 1 -2101
box -40 -38 40 42
use Li_via_M1  Li_via_M1_15
timestamp 1502773982
transform 1 0 -4736 0 1 625
box -40 -38 40 42
use Li_via_M1  Li_via_M1_16
timestamp 1502773982
transform 1 0 -4850 0 1 725
box -40 -38 40 42
use Li_via_M1  Li_via_M1_17
timestamp 1502773982
transform -1 0 -1550 0 1 -795
box -40 -38 40 42
use Li_via_M1  Li_via_M1_18
timestamp 1502773982
transform 1 0 -4622 0 1 925
box -40 -38 40 42
use Li_via_M1  Li_via_M1_19
timestamp 1502773982
transform 1 0 -4052 0 1 -875
box -40 -38 40 42
use Li_via_M1  Li_via_M1_20
timestamp 1502773982
transform 1 0 -4508 0 1 825
box -40 -38 40 42
use Li_via_M1  Li_via_M1_21
timestamp 1502773982
transform -1 0 -1550 0 -1 435
box -40 -38 40 42
use Li_via_M1  Li_via_M1_22
timestamp 1502773982
transform 1 0 -3938 0 1 -125
box -40 -38 40 42
use Li_via_M1  Li_via_M1_23
timestamp 1502773982
transform 1 0 460 0 1 -955
box -40 -38 40 42
use Li_via_M1  Li_via_M1_24
timestamp 1502773982
transform 1 0 460 0 1 485
box -40 -38 40 42
use Li_via_M1  Li_via_M1_25
timestamp 1502773982
transform 1 0 198 0 1 549
box -40 -38 40 42
use Li_via_M1  Li_via_M1_26
timestamp 1502773982
transform 1 0 460 0 1 605
box -40 -38 40 42
use Li_via_M1  Li_via_M1_27
timestamp 1502773982
transform 1 0 460 0 1 825
box -40 -38 40 42
use Li_via_M1  Li_via_M1_28
timestamp 1502773982
transform 1 0 -4166 0 1 -975
box -40 -38 40 42
use Li_via_M2  Li_via_M2_0
timestamp 1502773982
transform 1 0 2379 0 1 -1896
box -40 -38 40 42
use Li_via_M2  Li_via_M2_1
timestamp 1502773982
transform 1 0 2379 0 1 -1896
box -40 -38 40 42
use Li_via_M2  Li_via_M2_2
timestamp 1502773982
transform 1 0 2183 0 1 -2006
box -40 -38 40 42
use Li_via_M2  Li_via_M2_3
timestamp 1502773982
transform 1 0 2183 0 1 -2006
box -40 -38 40 42
use Li_via_M2  Li_via_M2_4
timestamp 1502773982
transform 1 0 401 0 1 -1766
box -40 -38 40 42
use Li_via_M2  Li_via_M2_5
timestamp 1502773982
transform 1 0 242 0 1 -2827
box -40 -38 40 42
use Li_via_M2  Li_via_M2_6
timestamp 1502773982
transform 1 0 2425 0 1 -2194
box -40 -38 40 42
use Li_via_M2  Li_via_M2_7
timestamp 1502773982
transform 1 0 2425 0 1 -2194
box -40 -38 40 42
use Li_via_M2  Li_via_M2_8
timestamp 1502773982
transform 1 0 2493 0 1 -1572
box -40 -38 40 42
use Li_via_M2  Li_via_M2_9
timestamp 1502773982
transform 1 0 2493 0 1 -1572
box -40 -38 40 42
use Li_via_M2  Li_via_M2_10
timestamp 1502773982
transform 1 0 331 0 1 -2396
box -40 -38 40 42
use Li_via_M2  Li_via_M2_11
timestamp 1502773982
transform 1 0 331 0 1 -2282
box -40 -38 40 42
use Li_via_M2  Li_via_M2_12
timestamp 1502773982
transform 1 0 330 0 1 -2168
box -40 -38 40 42
use Li_via_M2  Li_via_M2_13
timestamp 1502773982
transform 1 0 548 0 1 -1539
box -40 -38 40 42
use Li_via_M2  Li_via_M2_14
timestamp 1502773982
transform 1 0 154 0 1 -1972
box -40 -38 40 42
use Li_via_M2  Li_via_M2_15
timestamp 1502773982
transform 1 0 148 0 1 -2549
box -40 -38 40 42
use Li_via_M2  Li_via_M2_16
timestamp 1502773982
transform 1 0 -3679 0 1 -2825
box -40 -38 40 42
use Li_via_M2  Li_via_M2_17
timestamp 1502773982
transform 1 0 -1278 0 1 -1109
box -40 -38 40 42
use Li_via_M2  Li_via_M2_18
timestamp 1502773982
transform 1 0 -3679 0 1 -5
box -40 -38 40 42
use Li_via_M2  Li_via_M2_19
timestamp 1502773982
transform 1 0 -3679 0 1 -245
box -40 -38 40 42
use Li_via_M2  Li_via_M2_20
timestamp 1502773982
transform 1 0 -1278 0 -1 863
box -40 -38 40 42
use Li_via_M2  Li_via_M2_21
timestamp 1502773982
transform 1 0 2223 0 1 435
box -40 -38 40 42
use Li_via_M2  Li_via_M2_22
timestamp 1502773982
transform 1 0 2223 0 1 435
box -40 -38 40 42
use Li_via_M2  Li_via_M2_23
timestamp 1502773982
transform 1 0 2223 0 1 -685
box -40 -38 40 42
use Li_via_M2  Li_via_M2_24
timestamp 1502773982
transform 1 0 2223 0 1 -685
box -40 -38 40 42
use Li_via_M2  Li_via_M2_25
timestamp 1502773982
transform 1 0 2120 0 1 115
box -40 -38 40 42
use Li_via_M2  Li_via_M2_26
timestamp 1502773982
transform 1 0 2120 0 1 115
box -40 -38 40 42
use Li_via_M2  Li_via_M2_27
timestamp 1502773982
transform 1 0 2120 0 1 -365
box -40 -38 40 42
use Li_via_M2  Li_via_M2_28
timestamp 1502773982
transform 1 0 2120 0 1 -365
box -40 -38 40 42
use Li_via_M2  Li_via_M2_29
timestamp 1502773982
transform 1 0 548 0 1 -5
box -40 -38 40 42
use Li_via_M2  Li_via_M2_30
timestamp 1502773982
transform 1 0 2140 0 1 1055
box -40 -38 40 42
use Li_via_M2  Li_via_M2_31
timestamp 1502773982
transform 1 0 548 0 1 -244
box -40 -38 40 42
use Li_via_M2  Li_via_M2_32
timestamp 1502773982
transform 1 0 198 0 1 -963
box -40 -38 40 42
use M1_M3  M1_M3_0
timestamp 1502773982
transform 1 0 -930 0 1 -1135
box -110 -90 -10 10
use M1_M3  M1_M3_1
timestamp 1502773982
transform 1 0 -4562 0 1 -1135
box -110 -90 -10 10
use M1_M3  M1_M3_2
timestamp 1502773982
transform 1 0 -4448 0 1 -428
box -110 -90 -10 10
use M1_M3  M1_M3_3
timestamp 1502773982
transform 1 0 -1476 0 1 -427
box -110 -90 -10 10
use M1_M3  M1_M3_4
timestamp 1502773982
transform 1 0 -1476 0 1 268
box -110 -90 -10 10
use M1_M3  M1_M3_5
timestamp 1502773982
transform 1 0 -4106 0 1 268
box -110 -90 -10 10
use M1_M3  M1_M3_6
timestamp 1502773982
transform 1 0 -3992 0 1 968
box -110 -90 -10 10
use M1_M3  M1_M3_7
timestamp 1502773982
transform 1 0 -930 0 1 969
box -110 -90 -10 10
use M1_via_M2  M1_via_M2_0
timestamp 1502773982
transform 1 0 198 0 1 -1071
box -40 -38 40 42
use M1_via_M2  M1_via_M2_1
timestamp 1502773982
transform 1 0 1941 0 1 -2194
box -40 -38 40 42
use M1_via_M2  M1_via_M2_2
timestamp 1502773982
transform 1 0 330 0 1 -2058
box -40 -38 40 42
use M1_via_M2  M1_via_M2_3
timestamp 1502773982
transform 1 0 -1278 0 1 -996
box -40 -38 40 42
use M1_via_M2  M1_via_M2_4
timestamp 1502773982
transform 1 0 -3795 0 1 -1305
box -40 -38 40 42
use M1_via_M2  M1_via_M2_5
timestamp 1502773982
transform 1 0 -3795 0 1 -1766
box -40 -38 40 42
use M1_via_M2  M1_via_M2_6
timestamp 1502773982
transform 1 0 -1278 0 -1 752
box -40 -38 40 42
use M1_via_M2  M1_via_M2_7
timestamp 1502773982
transform 1 0 -3794 0 1 1055
box -40 -38 40 42
use M1_via_M2  M1_via_M2_8
timestamp 1502773982
transform 1 0 198 0 1 729
box -40 -38 40 42
use M1_via_M2  M1_via_M2_9
timestamp 1502773982
transform 1 0 198 0 1 838
box -40 -38 40 42
<< labels >>
flabel metal1 s -3960 -146 -3916 -100 2 FreeSans 2000 0 0 0 GND
port 1 nsew
flabel metal1 s -4880 873 -4819 933 2 FreeSans 2500 0 0 0 x0
port 2 nsew
flabel metal1 s -4767 812 -4706 872 2 FreeSans 2500 0 0 0 x0_bar
port 3 nsew
flabel metal1 s -4652 873 -4591 933 2 FreeSans 2500 0 0 0 x1
port 4 nsew
flabel metal1 s -4538 812 -4477 872 2 FreeSans 2500 0 0 0 x1_bar
port 5 nsew
flabel metal1 s -4423 877 -4362 937 2 FreeSans 2500 0 0 0 x2
port 6 nsew
flabel metal1 s -4311 813 -4250 873 2 FreeSans 2500 0 0 0 x2_bar
port 7 nsew
flabel metal1 s -4196 874 -4135 934 2 FreeSans 2500 0 0 0 x3
port 8 nsew
flabel metal1 s -4082 813 -4021 873 2 FreeSans 2500 0 0 0 x3_bar
port 9 nsew
flabel metal2 s 2370 -2290 2390 -2270 2 FreeSans 2000 0 0 0 s3_bar
port 10 nsew
flabel metal2 s 2381 -2281 2381 -2281 2 FreeSans 2000 0 0 0 s1_bar
port 11 nsew
flabel metal2 s 2381 -2281 2381 -2281 2 FreeSans 2000 0 0 0 s1_bar
port 11 nsew
flabel metal2 s -3810 1159 -3779 1190 2 FreeSans 2000 0 0 0 CLK1
port 12 nsew
flabel metal2 s -3690 1165 -3667 1189 2 FreeSans 2000 0 0 0 Dis1
port 13 nsew
flabel metal2 s 277 1172 296 1193 2 FreeSans 2000 0 0 0 Dis3
port 14 nsew
flabel metal2 s 388 1169 413 1194 2 FreeSans 2000 0 0 0 CLK3
port 15 nsew
flabel metal2 s 536 1171 561 1195 2 FreeSans 2000 0 0 0 Dis2
port 16 nsew
flabel metal2 s 2124 1161 2158 1195 2 FreeSans 2000 0 0 0 CLK2
port 17 nsew
flabel metal2 s 2381 -2281 2381 -2281 2 FreeSans 2000 0 0 0 s1_bar
port 11 nsew
<< properties >>
string path -102.900 5.700 -39.650 5.700 
<< end >>
