**.subckt INV_VP_VN_sim
x1 VDD A OUT GND INV_VP_VN
Vdd VDD GND 1.8
Vin1 A GND pulse(0,1.8,1ns,1ns,1ns,1us,2us)
**** begin user architecture code

.lib /research/pdk/open_pdks/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include ~/magic_layout_stuff/INV_VP_VN.spice
.control
tran 0.1n 10u
plot v(A)
plot v(OUT)
.endc
.save all

**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
