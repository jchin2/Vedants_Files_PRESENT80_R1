magic
tech sky130A
magscale 1 2
timestamp 1671058898
<< error_p >>
rect 80 30 200 930
rect 230 30 350 930
rect 380 30 500 930
rect 530 30 650 930
rect 680 30 800 930
rect 830 30 950 930
rect 980 30 1100 930
rect 1130 30 1250 930
rect 1280 30 1400 930
rect 1430 30 1550 930
rect 1580 30 1700 930
<< pwell >>
rect 54 4 1726 956
<< nmoslvt >>
rect 200 30 230 930
rect 350 30 380 930
rect 500 30 530 930
rect 650 30 680 930
rect 800 30 830 930
rect 950 30 980 930
rect 1100 30 1130 930
rect 1250 30 1280 930
rect 1400 30 1430 930
rect 1550 30 1580 930
<< ndiff >>
rect 80 871 200 930
rect 80 837 123 871
rect 157 837 200 871
rect 80 803 200 837
rect 80 769 123 803
rect 157 769 200 803
rect 80 735 200 769
rect 80 701 123 735
rect 157 701 200 735
rect 80 667 200 701
rect 80 633 123 667
rect 157 633 200 667
rect 80 599 200 633
rect 80 565 123 599
rect 157 565 200 599
rect 80 531 200 565
rect 80 497 123 531
rect 157 497 200 531
rect 80 463 200 497
rect 80 429 123 463
rect 157 429 200 463
rect 80 395 200 429
rect 80 361 123 395
rect 157 361 200 395
rect 80 327 200 361
rect 80 293 123 327
rect 157 293 200 327
rect 80 259 200 293
rect 80 225 123 259
rect 157 225 200 259
rect 80 191 200 225
rect 80 157 123 191
rect 157 157 200 191
rect 80 123 200 157
rect 80 89 123 123
rect 157 89 200 123
rect 80 30 200 89
rect 230 871 350 930
rect 230 837 273 871
rect 307 837 350 871
rect 230 803 350 837
rect 230 769 273 803
rect 307 769 350 803
rect 230 735 350 769
rect 230 701 273 735
rect 307 701 350 735
rect 230 667 350 701
rect 230 633 273 667
rect 307 633 350 667
rect 230 599 350 633
rect 230 565 273 599
rect 307 565 350 599
rect 230 531 350 565
rect 230 497 273 531
rect 307 497 350 531
rect 230 463 350 497
rect 230 429 273 463
rect 307 429 350 463
rect 230 395 350 429
rect 230 361 273 395
rect 307 361 350 395
rect 230 327 350 361
rect 230 293 273 327
rect 307 293 350 327
rect 230 259 350 293
rect 230 225 273 259
rect 307 225 350 259
rect 230 191 350 225
rect 230 157 273 191
rect 307 157 350 191
rect 230 123 350 157
rect 230 89 273 123
rect 307 89 350 123
rect 230 30 350 89
rect 380 871 500 930
rect 380 837 423 871
rect 457 837 500 871
rect 380 803 500 837
rect 380 769 423 803
rect 457 769 500 803
rect 380 735 500 769
rect 380 701 423 735
rect 457 701 500 735
rect 380 667 500 701
rect 380 633 423 667
rect 457 633 500 667
rect 380 599 500 633
rect 380 565 423 599
rect 457 565 500 599
rect 380 531 500 565
rect 380 497 423 531
rect 457 497 500 531
rect 380 463 500 497
rect 380 429 423 463
rect 457 429 500 463
rect 380 395 500 429
rect 380 361 423 395
rect 457 361 500 395
rect 380 327 500 361
rect 380 293 423 327
rect 457 293 500 327
rect 380 259 500 293
rect 380 225 423 259
rect 457 225 500 259
rect 380 191 500 225
rect 380 157 423 191
rect 457 157 500 191
rect 380 123 500 157
rect 380 89 423 123
rect 457 89 500 123
rect 380 30 500 89
rect 530 871 650 930
rect 530 837 573 871
rect 607 837 650 871
rect 530 803 650 837
rect 530 769 573 803
rect 607 769 650 803
rect 530 735 650 769
rect 530 701 573 735
rect 607 701 650 735
rect 530 667 650 701
rect 530 633 573 667
rect 607 633 650 667
rect 530 599 650 633
rect 530 565 573 599
rect 607 565 650 599
rect 530 531 650 565
rect 530 497 573 531
rect 607 497 650 531
rect 530 463 650 497
rect 530 429 573 463
rect 607 429 650 463
rect 530 395 650 429
rect 530 361 573 395
rect 607 361 650 395
rect 530 327 650 361
rect 530 293 573 327
rect 607 293 650 327
rect 530 259 650 293
rect 530 225 573 259
rect 607 225 650 259
rect 530 191 650 225
rect 530 157 573 191
rect 607 157 650 191
rect 530 123 650 157
rect 530 89 573 123
rect 607 89 650 123
rect 530 30 650 89
rect 680 871 800 930
rect 680 837 723 871
rect 757 837 800 871
rect 680 803 800 837
rect 680 769 723 803
rect 757 769 800 803
rect 680 735 800 769
rect 680 701 723 735
rect 757 701 800 735
rect 680 667 800 701
rect 680 633 723 667
rect 757 633 800 667
rect 680 599 800 633
rect 680 565 723 599
rect 757 565 800 599
rect 680 531 800 565
rect 680 497 723 531
rect 757 497 800 531
rect 680 463 800 497
rect 680 429 723 463
rect 757 429 800 463
rect 680 395 800 429
rect 680 361 723 395
rect 757 361 800 395
rect 680 327 800 361
rect 680 293 723 327
rect 757 293 800 327
rect 680 259 800 293
rect 680 225 723 259
rect 757 225 800 259
rect 680 191 800 225
rect 680 157 723 191
rect 757 157 800 191
rect 680 123 800 157
rect 680 89 723 123
rect 757 89 800 123
rect 680 30 800 89
rect 830 871 950 930
rect 830 837 873 871
rect 907 837 950 871
rect 830 803 950 837
rect 830 769 873 803
rect 907 769 950 803
rect 830 735 950 769
rect 830 701 873 735
rect 907 701 950 735
rect 830 667 950 701
rect 830 633 873 667
rect 907 633 950 667
rect 830 599 950 633
rect 830 565 873 599
rect 907 565 950 599
rect 830 531 950 565
rect 830 497 873 531
rect 907 497 950 531
rect 830 463 950 497
rect 830 429 873 463
rect 907 429 950 463
rect 830 395 950 429
rect 830 361 873 395
rect 907 361 950 395
rect 830 327 950 361
rect 830 293 873 327
rect 907 293 950 327
rect 830 259 950 293
rect 830 225 873 259
rect 907 225 950 259
rect 830 191 950 225
rect 830 157 873 191
rect 907 157 950 191
rect 830 123 950 157
rect 830 89 873 123
rect 907 89 950 123
rect 830 30 950 89
rect 980 871 1100 930
rect 980 837 1023 871
rect 1057 837 1100 871
rect 980 803 1100 837
rect 980 769 1023 803
rect 1057 769 1100 803
rect 980 735 1100 769
rect 980 701 1023 735
rect 1057 701 1100 735
rect 980 667 1100 701
rect 980 633 1023 667
rect 1057 633 1100 667
rect 980 599 1100 633
rect 980 565 1023 599
rect 1057 565 1100 599
rect 980 531 1100 565
rect 980 497 1023 531
rect 1057 497 1100 531
rect 980 463 1100 497
rect 980 429 1023 463
rect 1057 429 1100 463
rect 980 395 1100 429
rect 980 361 1023 395
rect 1057 361 1100 395
rect 980 327 1100 361
rect 980 293 1023 327
rect 1057 293 1100 327
rect 980 259 1100 293
rect 980 225 1023 259
rect 1057 225 1100 259
rect 980 191 1100 225
rect 980 157 1023 191
rect 1057 157 1100 191
rect 980 123 1100 157
rect 980 89 1023 123
rect 1057 89 1100 123
rect 980 30 1100 89
rect 1130 871 1250 930
rect 1130 837 1173 871
rect 1207 837 1250 871
rect 1130 803 1250 837
rect 1130 769 1173 803
rect 1207 769 1250 803
rect 1130 735 1250 769
rect 1130 701 1173 735
rect 1207 701 1250 735
rect 1130 667 1250 701
rect 1130 633 1173 667
rect 1207 633 1250 667
rect 1130 599 1250 633
rect 1130 565 1173 599
rect 1207 565 1250 599
rect 1130 531 1250 565
rect 1130 497 1173 531
rect 1207 497 1250 531
rect 1130 463 1250 497
rect 1130 429 1173 463
rect 1207 429 1250 463
rect 1130 395 1250 429
rect 1130 361 1173 395
rect 1207 361 1250 395
rect 1130 327 1250 361
rect 1130 293 1173 327
rect 1207 293 1250 327
rect 1130 259 1250 293
rect 1130 225 1173 259
rect 1207 225 1250 259
rect 1130 191 1250 225
rect 1130 157 1173 191
rect 1207 157 1250 191
rect 1130 123 1250 157
rect 1130 89 1173 123
rect 1207 89 1250 123
rect 1130 30 1250 89
rect 1280 871 1400 930
rect 1280 837 1323 871
rect 1357 837 1400 871
rect 1280 803 1400 837
rect 1280 769 1323 803
rect 1357 769 1400 803
rect 1280 735 1400 769
rect 1280 701 1323 735
rect 1357 701 1400 735
rect 1280 667 1400 701
rect 1280 633 1323 667
rect 1357 633 1400 667
rect 1280 599 1400 633
rect 1280 565 1323 599
rect 1357 565 1400 599
rect 1280 531 1400 565
rect 1280 497 1323 531
rect 1357 497 1400 531
rect 1280 463 1400 497
rect 1280 429 1323 463
rect 1357 429 1400 463
rect 1280 395 1400 429
rect 1280 361 1323 395
rect 1357 361 1400 395
rect 1280 327 1400 361
rect 1280 293 1323 327
rect 1357 293 1400 327
rect 1280 259 1400 293
rect 1280 225 1323 259
rect 1357 225 1400 259
rect 1280 191 1400 225
rect 1280 157 1323 191
rect 1357 157 1400 191
rect 1280 123 1400 157
rect 1280 89 1323 123
rect 1357 89 1400 123
rect 1280 30 1400 89
rect 1430 861 1550 930
rect 1430 827 1473 861
rect 1507 827 1550 861
rect 1430 793 1550 827
rect 1430 759 1473 793
rect 1507 759 1550 793
rect 1430 725 1550 759
rect 1430 691 1473 725
rect 1507 691 1550 725
rect 1430 657 1550 691
rect 1430 623 1473 657
rect 1507 623 1550 657
rect 1430 589 1550 623
rect 1430 555 1473 589
rect 1507 555 1550 589
rect 1430 521 1550 555
rect 1430 487 1473 521
rect 1507 487 1550 521
rect 1430 453 1550 487
rect 1430 419 1473 453
rect 1507 419 1550 453
rect 1430 385 1550 419
rect 1430 351 1473 385
rect 1507 351 1550 385
rect 1430 317 1550 351
rect 1430 283 1473 317
rect 1507 283 1550 317
rect 1430 249 1550 283
rect 1430 215 1473 249
rect 1507 215 1550 249
rect 1430 181 1550 215
rect 1430 147 1473 181
rect 1507 147 1550 181
rect 1430 113 1550 147
rect 1430 79 1473 113
rect 1507 79 1550 113
rect 1430 30 1550 79
rect 1580 871 1700 930
rect 1580 837 1623 871
rect 1657 837 1700 871
rect 1580 803 1700 837
rect 1580 769 1623 803
rect 1657 769 1700 803
rect 1580 735 1700 769
rect 1580 701 1623 735
rect 1657 701 1700 735
rect 1580 667 1700 701
rect 1580 633 1623 667
rect 1657 633 1700 667
rect 1580 599 1700 633
rect 1580 565 1623 599
rect 1657 565 1700 599
rect 1580 531 1700 565
rect 1580 497 1623 531
rect 1657 497 1700 531
rect 1580 463 1700 497
rect 1580 429 1623 463
rect 1657 429 1700 463
rect 1580 395 1700 429
rect 1580 361 1623 395
rect 1657 361 1700 395
rect 1580 327 1700 361
rect 1580 293 1623 327
rect 1657 293 1700 327
rect 1580 259 1700 293
rect 1580 225 1623 259
rect 1657 225 1700 259
rect 1580 191 1700 225
rect 1580 157 1623 191
rect 1657 157 1700 191
rect 1580 123 1700 157
rect 1580 89 1623 123
rect 1657 89 1700 123
rect 1580 30 1700 89
<< ndiffc >>
rect 123 837 157 871
rect 123 769 157 803
rect 123 701 157 735
rect 123 633 157 667
rect 123 565 157 599
rect 123 497 157 531
rect 123 429 157 463
rect 123 361 157 395
rect 123 293 157 327
rect 123 225 157 259
rect 123 157 157 191
rect 123 89 157 123
rect 273 837 307 871
rect 273 769 307 803
rect 273 701 307 735
rect 273 633 307 667
rect 273 565 307 599
rect 273 497 307 531
rect 273 429 307 463
rect 273 361 307 395
rect 273 293 307 327
rect 273 225 307 259
rect 273 157 307 191
rect 273 89 307 123
rect 423 837 457 871
rect 423 769 457 803
rect 423 701 457 735
rect 423 633 457 667
rect 423 565 457 599
rect 423 497 457 531
rect 423 429 457 463
rect 423 361 457 395
rect 423 293 457 327
rect 423 225 457 259
rect 423 157 457 191
rect 423 89 457 123
rect 573 837 607 871
rect 573 769 607 803
rect 573 701 607 735
rect 573 633 607 667
rect 573 565 607 599
rect 573 497 607 531
rect 573 429 607 463
rect 573 361 607 395
rect 573 293 607 327
rect 573 225 607 259
rect 573 157 607 191
rect 573 89 607 123
rect 723 837 757 871
rect 723 769 757 803
rect 723 701 757 735
rect 723 633 757 667
rect 723 565 757 599
rect 723 497 757 531
rect 723 429 757 463
rect 723 361 757 395
rect 723 293 757 327
rect 723 225 757 259
rect 723 157 757 191
rect 723 89 757 123
rect 873 837 907 871
rect 873 769 907 803
rect 873 701 907 735
rect 873 633 907 667
rect 873 565 907 599
rect 873 497 907 531
rect 873 429 907 463
rect 873 361 907 395
rect 873 293 907 327
rect 873 225 907 259
rect 873 157 907 191
rect 873 89 907 123
rect 1023 837 1057 871
rect 1023 769 1057 803
rect 1023 701 1057 735
rect 1023 633 1057 667
rect 1023 565 1057 599
rect 1023 497 1057 531
rect 1023 429 1057 463
rect 1023 361 1057 395
rect 1023 293 1057 327
rect 1023 225 1057 259
rect 1023 157 1057 191
rect 1023 89 1057 123
rect 1173 837 1207 871
rect 1173 769 1207 803
rect 1173 701 1207 735
rect 1173 633 1207 667
rect 1173 565 1207 599
rect 1173 497 1207 531
rect 1173 429 1207 463
rect 1173 361 1207 395
rect 1173 293 1207 327
rect 1173 225 1207 259
rect 1173 157 1207 191
rect 1173 89 1207 123
rect 1323 837 1357 871
rect 1323 769 1357 803
rect 1323 701 1357 735
rect 1323 633 1357 667
rect 1323 565 1357 599
rect 1323 497 1357 531
rect 1323 429 1357 463
rect 1323 361 1357 395
rect 1323 293 1357 327
rect 1323 225 1357 259
rect 1323 157 1357 191
rect 1323 89 1357 123
rect 1473 827 1507 861
rect 1473 759 1507 793
rect 1473 691 1507 725
rect 1473 623 1507 657
rect 1473 555 1507 589
rect 1473 487 1507 521
rect 1473 419 1507 453
rect 1473 351 1507 385
rect 1473 283 1507 317
rect 1473 215 1507 249
rect 1473 147 1507 181
rect 1473 79 1507 113
rect 1623 837 1657 871
rect 1623 769 1657 803
rect 1623 701 1657 735
rect 1623 633 1657 667
rect 1623 565 1657 599
rect 1623 497 1657 531
rect 1623 429 1657 463
rect 1623 361 1657 395
rect 1623 293 1657 327
rect 1623 225 1657 259
rect 1623 157 1657 191
rect 1623 89 1657 123
<< poly >>
rect 200 930 230 980
rect 350 930 380 980
rect 500 930 530 980
rect 650 930 680 980
rect 800 930 830 980
rect 950 930 980 980
rect 1100 930 1130 980
rect 1250 930 1280 980
rect 1400 930 1430 980
rect 1550 930 1580 980
rect 200 0 230 30
rect 350 0 380 30
rect 500 0 530 30
rect 650 0 680 30
rect 800 0 830 30
rect 950 0 980 30
rect 1100 0 1130 30
rect 1250 0 1280 30
rect 1400 0 1430 30
rect 1550 0 1580 30
<< locali >>
rect 100 871 180 910
rect 100 837 123 871
rect 157 837 180 871
rect 100 803 180 837
rect 100 769 123 803
rect 157 769 180 803
rect 100 735 180 769
rect 100 701 123 735
rect 157 701 180 735
rect 100 667 180 701
rect 100 633 123 667
rect 157 633 180 667
rect 100 599 180 633
rect 100 565 123 599
rect 157 565 180 599
rect 100 531 180 565
rect 100 497 123 531
rect 157 497 180 531
rect 100 463 180 497
rect 100 429 123 463
rect 157 429 180 463
rect 100 395 180 429
rect 100 361 123 395
rect 157 361 180 395
rect 100 327 180 361
rect 100 293 123 327
rect 157 293 180 327
rect 100 259 180 293
rect 100 225 123 259
rect 157 225 180 259
rect 100 191 180 225
rect 100 157 123 191
rect 157 157 180 191
rect 100 123 180 157
rect 100 89 123 123
rect 157 89 180 123
rect 100 50 180 89
rect 250 871 330 910
rect 250 837 273 871
rect 307 837 330 871
rect 250 803 330 837
rect 250 769 273 803
rect 307 769 330 803
rect 250 735 330 769
rect 250 701 273 735
rect 307 701 330 735
rect 250 667 330 701
rect 250 633 273 667
rect 307 633 330 667
rect 250 599 330 633
rect 250 565 273 599
rect 307 565 330 599
rect 250 531 330 565
rect 250 497 273 531
rect 307 497 330 531
rect 250 463 330 497
rect 250 429 273 463
rect 307 429 330 463
rect 250 395 330 429
rect 250 361 273 395
rect 307 361 330 395
rect 250 327 330 361
rect 250 293 273 327
rect 307 293 330 327
rect 250 259 330 293
rect 250 225 273 259
rect 307 225 330 259
rect 250 191 330 225
rect 250 157 273 191
rect 307 157 330 191
rect 250 123 330 157
rect 250 89 273 123
rect 307 89 330 123
rect 250 50 330 89
rect 400 871 480 910
rect 400 837 423 871
rect 457 837 480 871
rect 400 803 480 837
rect 400 769 423 803
rect 457 769 480 803
rect 400 735 480 769
rect 400 701 423 735
rect 457 701 480 735
rect 400 667 480 701
rect 400 633 423 667
rect 457 633 480 667
rect 400 599 480 633
rect 400 565 423 599
rect 457 565 480 599
rect 400 531 480 565
rect 400 497 423 531
rect 457 497 480 531
rect 400 463 480 497
rect 400 429 423 463
rect 457 429 480 463
rect 400 395 480 429
rect 400 361 423 395
rect 457 361 480 395
rect 400 327 480 361
rect 400 293 423 327
rect 457 293 480 327
rect 400 259 480 293
rect 400 225 423 259
rect 457 225 480 259
rect 400 191 480 225
rect 400 157 423 191
rect 457 157 480 191
rect 400 123 480 157
rect 400 89 423 123
rect 457 89 480 123
rect 400 50 480 89
rect 550 871 630 910
rect 550 837 573 871
rect 607 837 630 871
rect 550 803 630 837
rect 550 769 573 803
rect 607 769 630 803
rect 550 735 630 769
rect 550 701 573 735
rect 607 701 630 735
rect 550 667 630 701
rect 550 633 573 667
rect 607 633 630 667
rect 550 599 630 633
rect 550 565 573 599
rect 607 565 630 599
rect 550 531 630 565
rect 550 497 573 531
rect 607 497 630 531
rect 550 463 630 497
rect 550 429 573 463
rect 607 429 630 463
rect 550 395 630 429
rect 550 361 573 395
rect 607 361 630 395
rect 550 327 630 361
rect 550 293 573 327
rect 607 293 630 327
rect 550 259 630 293
rect 550 225 573 259
rect 607 225 630 259
rect 550 191 630 225
rect 550 157 573 191
rect 607 157 630 191
rect 550 123 630 157
rect 550 89 573 123
rect 607 89 630 123
rect 550 50 630 89
rect 700 871 780 910
rect 700 837 723 871
rect 757 837 780 871
rect 700 803 780 837
rect 700 769 723 803
rect 757 769 780 803
rect 700 735 780 769
rect 700 701 723 735
rect 757 701 780 735
rect 700 667 780 701
rect 700 633 723 667
rect 757 633 780 667
rect 700 599 780 633
rect 700 565 723 599
rect 757 565 780 599
rect 700 531 780 565
rect 700 497 723 531
rect 757 497 780 531
rect 700 463 780 497
rect 700 429 723 463
rect 757 429 780 463
rect 700 395 780 429
rect 700 361 723 395
rect 757 361 780 395
rect 700 327 780 361
rect 700 293 723 327
rect 757 293 780 327
rect 700 259 780 293
rect 700 225 723 259
rect 757 225 780 259
rect 700 191 780 225
rect 700 157 723 191
rect 757 157 780 191
rect 700 123 780 157
rect 700 89 723 123
rect 757 89 780 123
rect 700 50 780 89
rect 850 871 930 910
rect 850 837 873 871
rect 907 837 930 871
rect 850 803 930 837
rect 850 769 873 803
rect 907 769 930 803
rect 850 735 930 769
rect 850 701 873 735
rect 907 701 930 735
rect 850 667 930 701
rect 850 633 873 667
rect 907 633 930 667
rect 850 599 930 633
rect 850 565 873 599
rect 907 565 930 599
rect 850 531 930 565
rect 850 497 873 531
rect 907 497 930 531
rect 850 463 930 497
rect 850 429 873 463
rect 907 429 930 463
rect 850 395 930 429
rect 850 361 873 395
rect 907 361 930 395
rect 850 327 930 361
rect 850 293 873 327
rect 907 293 930 327
rect 850 259 930 293
rect 850 225 873 259
rect 907 225 930 259
rect 850 191 930 225
rect 850 157 873 191
rect 907 157 930 191
rect 850 123 930 157
rect 850 89 873 123
rect 907 89 930 123
rect 850 50 930 89
rect 1000 871 1080 910
rect 1000 837 1023 871
rect 1057 837 1080 871
rect 1000 803 1080 837
rect 1000 769 1023 803
rect 1057 769 1080 803
rect 1000 735 1080 769
rect 1000 701 1023 735
rect 1057 701 1080 735
rect 1000 667 1080 701
rect 1000 633 1023 667
rect 1057 633 1080 667
rect 1000 599 1080 633
rect 1000 565 1023 599
rect 1057 565 1080 599
rect 1000 531 1080 565
rect 1000 497 1023 531
rect 1057 497 1080 531
rect 1000 463 1080 497
rect 1000 429 1023 463
rect 1057 429 1080 463
rect 1000 395 1080 429
rect 1000 361 1023 395
rect 1057 361 1080 395
rect 1000 327 1080 361
rect 1000 293 1023 327
rect 1057 293 1080 327
rect 1000 259 1080 293
rect 1000 225 1023 259
rect 1057 225 1080 259
rect 1000 191 1080 225
rect 1000 157 1023 191
rect 1057 157 1080 191
rect 1000 123 1080 157
rect 1000 89 1023 123
rect 1057 89 1080 123
rect 1000 50 1080 89
rect 1150 871 1230 910
rect 1150 837 1173 871
rect 1207 837 1230 871
rect 1150 803 1230 837
rect 1150 769 1173 803
rect 1207 769 1230 803
rect 1150 735 1230 769
rect 1150 701 1173 735
rect 1207 701 1230 735
rect 1150 667 1230 701
rect 1150 633 1173 667
rect 1207 633 1230 667
rect 1150 599 1230 633
rect 1150 565 1173 599
rect 1207 565 1230 599
rect 1150 531 1230 565
rect 1150 497 1173 531
rect 1207 497 1230 531
rect 1150 463 1230 497
rect 1150 429 1173 463
rect 1207 429 1230 463
rect 1150 395 1230 429
rect 1150 361 1173 395
rect 1207 361 1230 395
rect 1150 327 1230 361
rect 1150 293 1173 327
rect 1207 293 1230 327
rect 1150 259 1230 293
rect 1150 225 1173 259
rect 1207 225 1230 259
rect 1150 191 1230 225
rect 1150 157 1173 191
rect 1207 157 1230 191
rect 1150 123 1230 157
rect 1150 89 1173 123
rect 1207 89 1230 123
rect 1150 50 1230 89
rect 1300 871 1380 910
rect 1300 837 1323 871
rect 1357 837 1380 871
rect 1300 803 1380 837
rect 1300 769 1323 803
rect 1357 769 1380 803
rect 1300 735 1380 769
rect 1300 701 1323 735
rect 1357 701 1380 735
rect 1300 667 1380 701
rect 1300 633 1323 667
rect 1357 633 1380 667
rect 1300 599 1380 633
rect 1300 565 1323 599
rect 1357 565 1380 599
rect 1300 531 1380 565
rect 1300 497 1323 531
rect 1357 497 1380 531
rect 1300 463 1380 497
rect 1300 429 1323 463
rect 1357 429 1380 463
rect 1300 395 1380 429
rect 1300 361 1323 395
rect 1357 361 1380 395
rect 1300 327 1380 361
rect 1300 293 1323 327
rect 1357 293 1380 327
rect 1300 259 1380 293
rect 1300 225 1323 259
rect 1357 225 1380 259
rect 1300 191 1380 225
rect 1300 157 1323 191
rect 1357 157 1380 191
rect 1300 123 1380 157
rect 1300 89 1323 123
rect 1357 89 1380 123
rect 1300 50 1380 89
rect 1450 861 1530 910
rect 1450 827 1473 861
rect 1507 827 1530 861
rect 1450 793 1530 827
rect 1450 759 1473 793
rect 1507 759 1530 793
rect 1450 725 1530 759
rect 1450 691 1473 725
rect 1507 691 1530 725
rect 1450 657 1530 691
rect 1450 623 1473 657
rect 1507 623 1530 657
rect 1450 589 1530 623
rect 1450 555 1473 589
rect 1507 555 1530 589
rect 1450 521 1530 555
rect 1450 487 1473 521
rect 1507 487 1530 521
rect 1450 453 1530 487
rect 1450 419 1473 453
rect 1507 419 1530 453
rect 1450 385 1530 419
rect 1450 351 1473 385
rect 1507 351 1530 385
rect 1450 317 1530 351
rect 1450 283 1473 317
rect 1507 283 1530 317
rect 1450 249 1530 283
rect 1450 215 1473 249
rect 1507 215 1530 249
rect 1450 181 1530 215
rect 1450 147 1473 181
rect 1507 147 1530 181
rect 1450 113 1530 147
rect 1450 79 1473 113
rect 1507 79 1530 113
rect 1450 50 1530 79
rect 1600 871 1680 910
rect 1600 837 1623 871
rect 1657 837 1680 871
rect 1600 803 1680 837
rect 1600 769 1623 803
rect 1657 769 1680 803
rect 1600 735 1680 769
rect 1600 701 1623 735
rect 1657 701 1680 735
rect 1600 667 1680 701
rect 1600 633 1623 667
rect 1657 633 1680 667
rect 1600 599 1680 633
rect 1600 565 1623 599
rect 1657 565 1680 599
rect 1600 531 1680 565
rect 1600 497 1623 531
rect 1657 497 1680 531
rect 1600 463 1680 497
rect 1600 429 1623 463
rect 1657 429 1680 463
rect 1600 395 1680 429
rect 1600 361 1623 395
rect 1657 361 1680 395
rect 1600 327 1680 361
rect 1600 293 1623 327
rect 1657 293 1680 327
rect 1600 259 1680 293
rect 1600 225 1623 259
rect 1657 225 1680 259
rect 1600 191 1680 225
rect 1600 157 1623 191
rect 1657 157 1680 191
rect 1600 123 1680 157
rect 1600 89 1623 123
rect 1657 89 1680 123
rect 1600 50 1680 89
<< end >>
