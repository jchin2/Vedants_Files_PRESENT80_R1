magic
tech sky130A
timestamp 1670902135
<< locali >>
rect -225 20 -185 30
rect -225 0 -215 20
rect -195 0 -185 20
rect -225 -10 -185 0
rect -165 20 -125 30
rect -165 0 -155 20
rect -135 0 -125 20
rect -165 -10 -125 0
rect -225 -40 -185 -30
rect -225 -60 -215 -40
rect -195 -60 -185 -40
rect -225 -70 -185 -60
rect -165 -40 -125 -30
rect -165 -60 -155 -40
rect -135 -60 -125 -40
rect -165 -70 -125 -60
<< viali >>
rect -215 0 -195 20
rect -155 0 -135 20
rect -215 -60 -195 -40
rect -155 -60 -135 -40
<< metal1 >>
rect -240 25 -110 45
rect -240 -5 -220 25
rect -190 -5 -160 25
rect -130 -5 -110 25
rect -240 -35 -110 -5
rect -240 -65 -220 -35
rect -190 -65 -160 -35
rect -130 -65 -110 -35
rect -240 -85 -110 -65
<< via1 >>
rect -220 20 -190 25
rect -220 0 -215 20
rect -215 0 -195 20
rect -195 0 -190 20
rect -220 -5 -190 0
rect -160 20 -130 25
rect -160 0 -155 20
rect -155 0 -135 20
rect -135 0 -130 20
rect -160 -5 -130 0
rect -220 -40 -190 -35
rect -220 -60 -215 -40
rect -215 -60 -195 -40
rect -195 -60 -190 -40
rect -220 -65 -190 -60
rect -160 -40 -130 -35
rect -160 -60 -155 -40
rect -155 -60 -135 -40
rect -135 -60 -130 -40
rect -160 -65 -130 -60
<< metal2 >>
rect -240 25 -110 45
rect -240 -5 -220 25
rect -190 -5 -160 25
rect -130 -5 -110 25
rect -240 -35 -110 -5
rect -240 -65 -220 -35
rect -190 -65 -160 -35
rect -130 -65 -110 -35
rect -240 -85 -110 -65
<< metal3 >>
rect -240 30 -110 45
rect -240 -10 -225 30
rect -185 -10 -165 30
rect -125 -10 -110 30
rect -240 -30 -110 -10
rect -240 -70 -225 -30
rect -185 -70 -165 -30
rect -125 -70 -110 -30
rect -240 -85 -110 -70
<< via3 >>
rect -225 -10 -185 30
rect -165 -10 -125 30
rect -225 -70 -185 -30
rect -165 -70 -125 -30
<< metal4 >>
rect -240 30 -110 45
rect -240 -10 -225 30
rect -185 -10 -165 30
rect -125 -10 -110 30
rect -240 -30 -110 -10
rect -240 -70 -225 -30
rect -185 -70 -165 -30
rect -125 -70 -110 -30
rect -240 -85 -110 -70
<< end >>
