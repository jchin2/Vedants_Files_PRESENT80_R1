magic
tech sky130A
magscale 1 2
timestamp 1670986233
<< metal3 >>
rect -7369 7572 -2470 7600
rect -7369 2628 -2554 7572
rect -2490 2628 -2470 7572
rect -7369 2600 -2470 2628
rect -2390 7572 2509 7600
rect -2390 2628 2425 7572
rect 2489 2628 2509 7572
rect -2390 2600 2509 2628
rect 2589 7572 7488 7600
rect 2589 2628 7404 7572
rect 7468 2628 7488 7572
rect 2589 2600 7488 2628
rect -7369 2472 -2470 2500
rect -7369 -2472 -2554 2472
rect -2490 -2472 -2470 2472
rect -7369 -2500 -2470 -2472
rect -2390 2472 2509 2500
rect -2390 -2472 2425 2472
rect 2489 -2472 2509 2472
rect -2390 -2500 2509 -2472
rect 2589 2472 7488 2500
rect 2589 -2472 7404 2472
rect 7468 -2472 7488 2472
rect 2589 -2500 7488 -2472
rect -7369 -2628 -2470 -2600
rect -7369 -7572 -2554 -2628
rect -2490 -7572 -2470 -2628
rect -7369 -7600 -2470 -7572
rect -2390 -2628 2509 -2600
rect -2390 -7572 2425 -2628
rect 2489 -7572 2509 -2628
rect -2390 -7600 2509 -7572
rect 2589 -2628 7488 -2600
rect 2589 -7572 7404 -2628
rect 7468 -7572 7488 -2628
rect 2589 -7600 7488 -7572
<< via3 >>
rect -2554 2628 -2490 7572
rect 2425 2628 2489 7572
rect 7404 2628 7468 7572
rect -2554 -2472 -2490 2472
rect 2425 -2472 2489 2472
rect 7404 -2472 7468 2472
rect -2554 -7572 -2490 -2628
rect 2425 -7572 2489 -2628
rect 7404 -7572 7468 -2628
<< mimcap >>
rect -7269 7460 -2669 7500
rect -7269 2740 -7229 7460
rect -2709 2740 -2669 7460
rect -7269 2700 -2669 2740
rect -2290 7460 2310 7500
rect -2290 2740 -2250 7460
rect 2270 2740 2310 7460
rect -2290 2700 2310 2740
rect 2689 7460 7289 7500
rect 2689 2740 2729 7460
rect 7249 2740 7289 7460
rect 2689 2700 7289 2740
rect -7269 2360 -2669 2400
rect -7269 -2360 -7229 2360
rect -2709 -2360 -2669 2360
rect -7269 -2400 -2669 -2360
rect -2290 2360 2310 2400
rect -2290 -2360 -2250 2360
rect 2270 -2360 2310 2360
rect -2290 -2400 2310 -2360
rect 2689 2360 7289 2400
rect 2689 -2360 2729 2360
rect 7249 -2360 7289 2360
rect 2689 -2400 7289 -2360
rect -7269 -2740 -2669 -2700
rect -7269 -7460 -7229 -2740
rect -2709 -7460 -2669 -2740
rect -7269 -7500 -2669 -7460
rect -2290 -2740 2310 -2700
rect -2290 -7460 -2250 -2740
rect 2270 -7460 2310 -2740
rect -2290 -7500 2310 -7460
rect 2689 -2740 7289 -2700
rect 2689 -7460 2729 -2740
rect 7249 -7460 7289 -2740
rect 2689 -7500 7289 -7460
<< mimcapcontact >>
rect -7229 2740 -2709 7460
rect -2250 2740 2270 7460
rect 2729 2740 7249 7460
rect -7229 -2360 -2709 2360
rect -2250 -2360 2270 2360
rect 2729 -2360 7249 2360
rect -7229 -7460 -2709 -2740
rect -2250 -7460 2270 -2740
rect 2729 -7460 7249 -2740
<< metal4 >>
rect -5021 7461 -4917 7650
rect -2601 7588 -2497 7650
rect -2601 7572 -2474 7588
rect -7230 7460 -2708 7461
rect -7230 2740 -7229 7460
rect -2709 2740 -2708 7460
rect -7230 2739 -2708 2740
rect -5021 2361 -4917 2739
rect -2601 2628 -2554 7572
rect -2490 2628 -2474 7572
rect -42 7461 62 7650
rect 2378 7588 2482 7650
rect 2378 7572 2505 7588
rect -2251 7460 2271 7461
rect -2251 2740 -2250 7460
rect 2270 2740 2271 7460
rect -2251 2739 2271 2740
rect -2601 2612 -2474 2628
rect -2601 2488 -2497 2612
rect -2601 2472 -2474 2488
rect -7230 2360 -2708 2361
rect -7230 -2360 -7229 2360
rect -2709 -2360 -2708 2360
rect -7230 -2361 -2708 -2360
rect -5021 -2739 -4917 -2361
rect -2601 -2472 -2554 2472
rect -2490 -2472 -2474 2472
rect -42 2361 62 2739
rect 2378 2628 2425 7572
rect 2489 2628 2505 7572
rect 4937 7461 5041 7650
rect 7357 7588 7461 7650
rect 7357 7572 7484 7588
rect 2728 7460 7250 7461
rect 2728 2740 2729 7460
rect 7249 2740 7250 7460
rect 2728 2739 7250 2740
rect 2378 2612 2505 2628
rect 2378 2488 2482 2612
rect 2378 2472 2505 2488
rect -2251 2360 2271 2361
rect -2251 -2360 -2250 2360
rect 2270 -2360 2271 2360
rect -2251 -2361 2271 -2360
rect -2601 -2488 -2474 -2472
rect -2601 -2612 -2497 -2488
rect -2601 -2628 -2474 -2612
rect -7230 -2740 -2708 -2739
rect -7230 -7460 -7229 -2740
rect -2709 -7460 -2708 -2740
rect -7230 -7461 -2708 -7460
rect -5021 -7650 -4917 -7461
rect -2601 -7572 -2554 -2628
rect -2490 -7572 -2474 -2628
rect -42 -2739 62 -2361
rect 2378 -2472 2425 2472
rect 2489 -2472 2505 2472
rect 4937 2361 5041 2739
rect 7357 2628 7404 7572
rect 7468 2628 7484 7572
rect 7357 2612 7484 2628
rect 7357 2488 7461 2612
rect 7357 2472 7484 2488
rect 2728 2360 7250 2361
rect 2728 -2360 2729 2360
rect 7249 -2360 7250 2360
rect 2728 -2361 7250 -2360
rect 2378 -2488 2505 -2472
rect 2378 -2612 2482 -2488
rect 2378 -2628 2505 -2612
rect -2251 -2740 2271 -2739
rect -2251 -7460 -2250 -2740
rect 2270 -7460 2271 -2740
rect -2251 -7461 2271 -7460
rect -2601 -7588 -2474 -7572
rect -2601 -7650 -2497 -7588
rect -42 -7650 62 -7461
rect 2378 -7572 2425 -2628
rect 2489 -7572 2505 -2628
rect 4937 -2739 5041 -2361
rect 7357 -2472 7404 2472
rect 7468 -2472 7484 2472
rect 7357 -2488 7484 -2472
rect 7357 -2612 7461 -2488
rect 7357 -2628 7484 -2612
rect 2728 -2740 7250 -2739
rect 2728 -7460 2729 -2740
rect 7249 -7460 7250 -2740
rect 2728 -7461 7250 -7460
rect 2378 -7588 2505 -7572
rect 2378 -7650 2482 -7588
rect 4937 -7650 5041 -7461
rect 7357 -7572 7404 -2628
rect 7468 -7572 7484 -2628
rect 7357 -7588 7484 -7572
rect 7357 -7650 7461 -7588
<< properties >>
string FIXED_BBOX 2469 2600 7269 7600
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 23 l 24 val 1.121k carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
