magic
tech sky130A
timestamp 1671245489
<< pwell >>
rect -628 -3 268 1003
<< nmoslvt >>
rect -495 10 -480 990
rect -420 10 -405 990
rect -345 10 -330 990
rect -270 10 -255 990
rect -195 10 -180 990
rect -120 10 -105 990
rect -45 10 -30 990
rect 30 10 45 990
rect 105 10 120 990
rect 180 10 195 990
<< ndiff >>
rect -555 970 -495 990
rect -555 30 -535 970
rect -515 30 -495 970
rect -555 10 -495 30
rect -480 970 -420 990
rect -480 30 -460 970
rect -440 30 -420 970
rect -480 10 -420 30
rect -405 970 -345 990
rect -405 30 -385 970
rect -365 30 -345 970
rect -405 10 -345 30
rect -330 970 -270 990
rect -330 30 -310 970
rect -290 30 -270 970
rect -330 10 -270 30
rect -255 970 -195 990
rect -255 30 -235 970
rect -215 30 -195 970
rect -255 10 -195 30
rect -180 970 -120 990
rect -180 30 -160 970
rect -140 30 -120 970
rect -180 10 -120 30
rect -105 970 -45 990
rect -105 30 -85 970
rect -65 30 -45 970
rect -105 10 -45 30
rect -30 970 30 990
rect -30 30 -10 970
rect 10 30 30 970
rect -30 10 30 30
rect 45 970 105 990
rect 45 30 65 970
rect 85 30 105 970
rect 45 10 105 30
rect 120 970 180 990
rect 120 30 140 970
rect 160 30 180 970
rect 120 10 180 30
rect 195 970 255 990
rect 195 30 215 970
rect 235 30 255 970
rect 195 10 255 30
<< ndiffc >>
rect -535 30 -515 970
rect -460 30 -440 970
rect -385 30 -365 970
rect -310 30 -290 970
rect -235 30 -215 970
rect -160 30 -140 970
rect -85 30 -65 970
rect -10 30 10 970
rect 65 30 85 970
rect 140 30 160 970
rect 215 30 235 970
<< psubdiff >>
rect -615 970 -555 990
rect -615 30 -595 970
rect -575 30 -555 970
rect -615 10 -555 30
<< psubdiffcont >>
rect -595 30 -575 970
<< poly >>
rect -495 990 -480 1005
rect -420 990 -405 1005
rect -345 990 -330 1005
rect -270 990 -255 1005
rect -195 990 -180 1005
rect -120 990 -105 1005
rect -45 990 -30 1005
rect 30 990 45 1005
rect 105 990 120 1005
rect 180 990 195 1005
rect -495 -5 -480 10
rect -420 -5 -405 10
rect -345 -5 -330 10
rect -270 -5 -255 10
rect -195 -5 -180 10
rect -120 -5 -105 10
rect -45 -5 -30 10
rect 30 -5 45 10
rect 105 -5 120 10
rect 180 -5 195 10
<< locali >>
rect -605 970 -505 980
rect -605 30 -595 970
rect -575 30 -535 970
rect -515 30 -505 970
rect -605 20 -505 30
rect -470 970 -430 980
rect -470 30 -460 970
rect -440 30 -430 970
rect -470 20 -430 30
rect -395 970 -355 980
rect -395 30 -385 970
rect -365 30 -355 970
rect -395 20 -355 30
rect -320 970 -280 980
rect -320 30 -310 970
rect -290 30 -280 970
rect -320 20 -280 30
rect -245 970 -205 980
rect -245 30 -235 970
rect -215 30 -205 970
rect -245 20 -205 30
rect -170 970 -130 980
rect -170 30 -160 970
rect -140 30 -130 970
rect -170 20 -130 30
rect -95 970 -55 980
rect -95 30 -85 970
rect -65 30 -55 970
rect -95 20 -55 30
rect -20 970 20 980
rect -20 30 -10 970
rect 10 30 20 970
rect -20 20 20 30
rect 55 970 95 980
rect 55 30 65 970
rect 85 30 95 970
rect 55 20 95 30
rect 130 970 170 980
rect 130 30 140 970
rect 160 30 170 970
rect 130 20 170 30
rect 205 970 245 980
rect 205 30 215 970
rect 235 30 245 970
rect 205 20 245 30
<< end >>
