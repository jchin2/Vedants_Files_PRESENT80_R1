magic
tech sky130A
magscale 1 2
timestamp 1672688233
<< nwell >>
rect 0 1170 1760 1356
rect 470 780 1290 1170
<< pwell >>
rect 14 4 1746 596
<< nmos >>
rect 160 270 190 570
rect 310 270 340 570
rect 640 270 670 570
rect 790 270 820 570
rect 940 270 970 570
rect 1090 270 1120 570
rect 1420 270 1450 570
rect 1570 270 1600 570
<< pmos >>
rect 640 830 670 1130
rect 790 830 820 1130
rect 940 830 970 1130
rect 1090 830 1120 1130
<< ndiff >>
rect 40 497 160 570
rect 40 463 83 497
rect 117 463 160 497
rect 40 417 160 463
rect 40 383 83 417
rect 117 383 160 417
rect 40 337 160 383
rect 40 303 83 337
rect 117 303 160 337
rect 40 270 160 303
rect 190 497 310 570
rect 190 463 233 497
rect 267 463 310 497
rect 190 417 310 463
rect 190 383 233 417
rect 267 383 310 417
rect 190 337 310 383
rect 190 303 233 337
rect 267 303 310 337
rect 190 270 310 303
rect 340 497 460 570
rect 340 463 383 497
rect 417 463 460 497
rect 340 417 460 463
rect 340 383 383 417
rect 417 383 460 417
rect 340 337 460 383
rect 340 303 383 337
rect 417 303 460 337
rect 340 270 460 303
rect 520 497 640 570
rect 520 463 563 497
rect 597 463 640 497
rect 520 417 640 463
rect 520 383 563 417
rect 597 383 640 417
rect 520 337 640 383
rect 520 303 563 337
rect 597 303 640 337
rect 520 270 640 303
rect 670 497 790 570
rect 670 463 713 497
rect 747 463 790 497
rect 670 417 790 463
rect 670 383 713 417
rect 747 383 790 417
rect 670 337 790 383
rect 670 303 713 337
rect 747 303 790 337
rect 670 270 790 303
rect 820 497 940 570
rect 820 463 863 497
rect 897 463 940 497
rect 820 417 940 463
rect 820 383 863 417
rect 897 383 940 417
rect 820 337 940 383
rect 820 303 863 337
rect 897 303 940 337
rect 820 270 940 303
rect 970 497 1090 570
rect 970 463 1013 497
rect 1047 463 1090 497
rect 970 417 1090 463
rect 970 383 1013 417
rect 1047 383 1090 417
rect 970 337 1090 383
rect 970 303 1013 337
rect 1047 303 1090 337
rect 970 270 1090 303
rect 1120 497 1240 570
rect 1120 463 1163 497
rect 1197 463 1240 497
rect 1120 417 1240 463
rect 1120 383 1163 417
rect 1197 383 1240 417
rect 1120 337 1240 383
rect 1120 303 1163 337
rect 1197 303 1240 337
rect 1120 270 1240 303
rect 1300 497 1420 570
rect 1300 463 1343 497
rect 1377 463 1420 497
rect 1300 417 1420 463
rect 1300 383 1343 417
rect 1377 383 1420 417
rect 1300 337 1420 383
rect 1300 303 1343 337
rect 1377 303 1420 337
rect 1300 270 1420 303
rect 1450 270 1570 570
rect 1600 497 1720 570
rect 1600 463 1643 497
rect 1677 463 1720 497
rect 1600 417 1720 463
rect 1600 383 1643 417
rect 1677 383 1720 417
rect 1600 337 1720 383
rect 1600 303 1643 337
rect 1677 303 1720 337
rect 1600 270 1720 303
<< pdiff >>
rect 520 1057 640 1130
rect 520 1023 563 1057
rect 597 1023 640 1057
rect 520 977 640 1023
rect 520 943 563 977
rect 597 943 640 977
rect 520 897 640 943
rect 520 863 563 897
rect 597 863 640 897
rect 520 830 640 863
rect 670 1057 790 1130
rect 670 1023 713 1057
rect 747 1023 790 1057
rect 670 977 790 1023
rect 670 943 713 977
rect 747 943 790 977
rect 670 897 790 943
rect 670 863 713 897
rect 747 863 790 897
rect 670 830 790 863
rect 820 1057 940 1130
rect 820 1023 863 1057
rect 897 1023 940 1057
rect 820 977 940 1023
rect 820 943 863 977
rect 897 943 940 977
rect 820 897 940 943
rect 820 863 863 897
rect 897 863 940 897
rect 820 830 940 863
rect 970 1057 1090 1130
rect 970 1023 1013 1057
rect 1047 1023 1090 1057
rect 970 977 1090 1023
rect 970 943 1013 977
rect 1047 943 1090 977
rect 970 897 1090 943
rect 970 863 1013 897
rect 1047 863 1090 897
rect 970 830 1090 863
rect 1120 1057 1240 1130
rect 1120 1023 1163 1057
rect 1197 1023 1240 1057
rect 1120 977 1240 1023
rect 1120 943 1163 977
rect 1197 943 1240 977
rect 1120 897 1240 943
rect 1120 863 1163 897
rect 1197 863 1240 897
rect 1120 830 1240 863
<< ndiffc >>
rect 83 463 117 497
rect 83 383 117 417
rect 83 303 117 337
rect 233 463 267 497
rect 233 383 267 417
rect 233 303 267 337
rect 383 463 417 497
rect 383 383 417 417
rect 383 303 417 337
rect 563 463 597 497
rect 563 383 597 417
rect 563 303 597 337
rect 713 463 747 497
rect 713 383 747 417
rect 713 303 747 337
rect 863 463 897 497
rect 863 383 897 417
rect 863 303 897 337
rect 1013 463 1047 497
rect 1013 383 1047 417
rect 1013 303 1047 337
rect 1163 463 1197 497
rect 1163 383 1197 417
rect 1163 303 1197 337
rect 1343 463 1377 497
rect 1343 383 1377 417
rect 1343 303 1377 337
rect 1643 463 1677 497
rect 1643 383 1677 417
rect 1643 303 1677 337
<< pdiffc >>
rect 563 1023 597 1057
rect 563 943 597 977
rect 563 863 597 897
rect 713 1023 747 1057
rect 713 943 747 977
rect 713 863 747 897
rect 863 1023 897 1057
rect 863 943 897 977
rect 863 863 897 897
rect 1013 1023 1047 1057
rect 1013 943 1047 977
rect 1013 863 1047 897
rect 1163 1023 1197 1057
rect 1163 943 1197 977
rect 1163 863 1197 897
<< psubdiff >>
rect 40 97 1720 130
rect 40 63 63 97
rect 97 63 143 97
rect 177 63 223 97
rect 257 63 303 97
rect 337 63 383 97
rect 417 63 463 97
rect 497 63 543 97
rect 577 63 623 97
rect 657 63 703 97
rect 737 63 783 97
rect 817 63 863 97
rect 897 63 943 97
rect 977 63 1023 97
rect 1057 63 1103 97
rect 1137 63 1183 97
rect 1217 63 1263 97
rect 1297 63 1343 97
rect 1377 63 1423 97
rect 1457 63 1503 97
rect 1537 63 1583 97
rect 1617 63 1663 97
rect 1697 63 1720 97
rect 40 30 1720 63
<< nsubdiff >>
rect 40 1277 1720 1310
rect 40 1243 63 1277
rect 97 1243 143 1277
rect 177 1243 223 1277
rect 257 1243 303 1277
rect 337 1243 383 1277
rect 417 1243 463 1277
rect 497 1243 543 1277
rect 577 1243 623 1277
rect 657 1243 703 1277
rect 737 1243 783 1277
rect 817 1243 863 1277
rect 897 1243 943 1277
rect 977 1243 1023 1277
rect 1057 1243 1103 1277
rect 1137 1243 1183 1277
rect 1217 1243 1263 1277
rect 1297 1243 1343 1277
rect 1377 1243 1423 1277
rect 1457 1243 1503 1277
rect 1537 1243 1583 1277
rect 1617 1243 1663 1277
rect 1697 1243 1720 1277
rect 40 1210 1720 1243
<< psubdiffcont >>
rect 63 63 97 97
rect 143 63 177 97
rect 223 63 257 97
rect 303 63 337 97
rect 383 63 417 97
rect 463 63 497 97
rect 543 63 577 97
rect 623 63 657 97
rect 703 63 737 97
rect 783 63 817 97
rect 863 63 897 97
rect 943 63 977 97
rect 1023 63 1057 97
rect 1103 63 1137 97
rect 1183 63 1217 97
rect 1263 63 1297 97
rect 1343 63 1377 97
rect 1423 63 1457 97
rect 1503 63 1537 97
rect 1583 63 1617 97
rect 1663 63 1697 97
<< nsubdiffcont >>
rect 63 1243 97 1277
rect 143 1243 177 1277
rect 223 1243 257 1277
rect 303 1243 337 1277
rect 383 1243 417 1277
rect 463 1243 497 1277
rect 543 1243 577 1277
rect 623 1243 657 1277
rect 703 1243 737 1277
rect 783 1243 817 1277
rect 863 1243 897 1277
rect 943 1243 977 1277
rect 1023 1243 1057 1277
rect 1103 1243 1137 1277
rect 1183 1243 1217 1277
rect 1263 1243 1297 1277
rect 1343 1243 1377 1277
rect 1423 1243 1457 1277
rect 1503 1243 1537 1277
rect 1583 1243 1617 1277
rect 1663 1243 1697 1277
<< poly >>
rect 640 1160 820 1190
rect 640 1130 670 1160
rect 790 1130 820 1160
rect 940 1160 1120 1190
rect 940 1130 970 1160
rect 1090 1130 1120 1160
rect 260 827 340 850
rect 1520 1047 1600 1070
rect 1520 1013 1543 1047
rect 1577 1013 1600 1047
rect 1520 990 1600 1013
rect 1370 927 1450 950
rect 1370 893 1393 927
rect 1427 893 1450 927
rect 1370 870 1450 893
rect 260 793 283 827
rect 317 793 340 827
rect 640 800 670 830
rect 260 770 340 793
rect 110 727 190 750
rect 110 693 133 727
rect 167 693 190 727
rect 110 670 190 693
rect 160 570 190 670
rect 310 570 340 770
rect 790 675 820 830
rect 940 800 970 830
rect 1090 800 1120 830
rect 890 777 970 800
rect 890 743 913 777
rect 947 743 970 777
rect 890 720 970 743
rect 790 652 870 675
rect 790 618 813 652
rect 847 618 870 652
rect 640 570 670 600
rect 790 595 870 618
rect 790 570 820 595
rect 940 570 970 720
rect 1090 570 1120 600
rect 1420 570 1450 870
rect 1570 570 1600 990
rect 160 240 190 270
rect 310 240 340 270
rect 640 240 670 270
rect 790 240 820 270
rect 940 240 970 270
rect 1090 240 1120 270
rect 1420 240 1450 270
rect 1570 240 1600 270
rect 640 217 720 240
rect 640 183 663 217
rect 697 183 720 217
rect 640 160 720 183
rect 1040 217 1120 240
rect 1040 183 1063 217
rect 1097 183 1120 217
rect 1040 160 1120 183
<< polycont >>
rect 1543 1013 1577 1047
rect 1393 893 1427 927
rect 283 793 317 827
rect 133 693 167 727
rect 913 743 947 777
rect 813 618 847 652
rect 663 183 697 217
rect 1063 183 1097 217
<< locali >>
rect 40 1277 1720 1300
rect 40 1243 63 1277
rect 97 1243 143 1277
rect 177 1243 223 1277
rect 257 1243 303 1277
rect 337 1243 383 1277
rect 417 1243 463 1277
rect 497 1243 543 1277
rect 577 1243 623 1277
rect 657 1243 703 1277
rect 737 1243 783 1277
rect 817 1243 863 1277
rect 897 1243 943 1277
rect 977 1243 1023 1277
rect 1057 1243 1103 1277
rect 1137 1243 1183 1277
rect 1217 1243 1263 1277
rect 1297 1243 1343 1277
rect 1377 1243 1423 1277
rect 1457 1243 1503 1277
rect 1537 1243 1583 1277
rect 1617 1243 1663 1277
rect 1697 1243 1720 1277
rect 40 1220 1720 1243
rect 390 1050 470 1070
rect 40 1047 470 1050
rect 40 1013 413 1047
rect 447 1013 470 1047
rect 40 1010 470 1013
rect 390 990 470 1010
rect 540 1057 620 1090
rect 540 1023 563 1057
rect 597 1023 620 1057
rect 540 977 620 1023
rect 390 930 470 950
rect 40 927 470 930
rect 40 893 413 927
rect 447 893 470 927
rect 40 890 470 893
rect 390 870 470 890
rect 540 943 563 977
rect 597 943 620 977
rect 540 897 620 943
rect 540 863 563 897
rect 597 863 620 897
rect 260 830 340 850
rect 540 840 620 863
rect 690 1057 770 1090
rect 690 1023 713 1057
rect 747 1023 770 1057
rect 690 977 770 1023
rect 690 943 713 977
rect 747 943 770 977
rect 690 897 770 943
rect 690 863 713 897
rect 747 863 770 897
rect 690 830 770 863
rect 840 1057 920 1090
rect 840 1023 863 1057
rect 897 1023 920 1057
rect 840 977 920 1023
rect 840 943 863 977
rect 897 943 920 977
rect 840 897 920 943
rect 840 863 863 897
rect 897 863 920 897
rect 840 840 920 863
rect 990 1057 1070 1090
rect 990 1023 1013 1057
rect 1047 1023 1070 1057
rect 990 977 1070 1023
rect 990 943 1013 977
rect 1047 943 1070 977
rect 990 897 1070 943
rect 990 863 1013 897
rect 1047 863 1070 897
rect 990 830 1070 863
rect 1140 1057 1220 1090
rect 1140 1023 1163 1057
rect 1197 1023 1220 1057
rect 1140 977 1220 1023
rect 1520 1047 1600 1070
rect 1520 1013 1543 1047
rect 1577 1013 1600 1047
rect 1520 990 1600 1013
rect 1140 943 1163 977
rect 1197 943 1220 977
rect 1140 897 1220 943
rect 1140 863 1163 897
rect 1197 863 1220 897
rect 1370 927 1450 950
rect 1370 893 1393 927
rect 1427 893 1450 927
rect 1370 870 1450 893
rect 1140 840 1220 863
rect 40 827 340 830
rect 40 793 283 827
rect 317 793 340 827
rect 40 790 340 793
rect 260 770 340 790
rect 710 780 750 830
rect 890 780 970 800
rect 710 777 970 780
rect 110 730 190 750
rect 40 727 190 730
rect 40 693 133 727
rect 167 693 190 727
rect 40 690 190 693
rect 110 670 190 690
rect 710 743 913 777
rect 947 743 970 777
rect 710 740 970 743
rect 710 610 750 740
rect 890 720 970 740
rect 80 570 750 610
rect 790 660 870 675
rect 1010 660 1050 830
rect 1290 780 1370 800
rect 1290 777 1720 780
rect 1290 743 1313 777
rect 1347 743 1720 777
rect 1290 740 1720 743
rect 1290 720 1370 740
rect 790 652 1720 660
rect 790 618 813 652
rect 847 620 1720 652
rect 847 618 870 620
rect 790 595 870 618
rect 80 530 120 570
rect 380 530 420 570
rect 711 530 750 570
rect 1010 530 1050 620
rect 1340 530 1380 620
rect 60 497 140 530
rect 60 463 83 497
rect 117 463 140 497
rect 60 417 140 463
rect 60 383 83 417
rect 117 383 140 417
rect 60 337 140 383
rect 60 303 83 337
rect 117 303 140 337
rect 60 280 140 303
rect 210 497 290 530
rect 210 463 233 497
rect 267 463 290 497
rect 210 417 290 463
rect 210 383 233 417
rect 267 383 290 417
rect 210 337 290 383
rect 210 303 233 337
rect 267 303 290 337
rect 210 280 290 303
rect 360 497 440 530
rect 360 463 383 497
rect 417 463 440 497
rect 360 417 440 463
rect 360 383 383 417
rect 417 383 440 417
rect 360 337 440 383
rect 360 303 383 337
rect 417 303 440 337
rect 360 280 440 303
rect 540 497 620 530
rect 540 463 563 497
rect 597 463 620 497
rect 540 417 620 463
rect 540 383 563 417
rect 597 383 620 417
rect 540 337 620 383
rect 540 303 563 337
rect 597 303 620 337
rect 540 280 620 303
rect 690 497 770 530
rect 690 463 713 497
rect 747 463 770 497
rect 690 417 770 463
rect 690 383 713 417
rect 747 383 770 417
rect 690 337 770 383
rect 690 303 713 337
rect 747 303 770 337
rect 690 280 770 303
rect 840 497 920 530
rect 840 463 863 497
rect 897 463 920 497
rect 840 417 920 463
rect 840 383 863 417
rect 897 383 920 417
rect 840 337 920 383
rect 840 303 863 337
rect 897 303 920 337
rect 840 280 920 303
rect 990 497 1070 530
rect 990 463 1013 497
rect 1047 463 1070 497
rect 990 417 1070 463
rect 990 383 1013 417
rect 1047 383 1070 417
rect 990 337 1070 383
rect 990 303 1013 337
rect 1047 303 1070 337
rect 990 280 1070 303
rect 1140 497 1220 530
rect 1140 463 1163 497
rect 1197 463 1220 497
rect 1140 417 1220 463
rect 1140 383 1163 417
rect 1197 383 1220 417
rect 1140 337 1220 383
rect 1140 303 1163 337
rect 1197 303 1220 337
rect 1140 280 1220 303
rect 1320 497 1400 530
rect 1320 463 1343 497
rect 1377 463 1400 497
rect 1320 417 1400 463
rect 1320 383 1343 417
rect 1377 383 1400 417
rect 1320 337 1400 383
rect 1320 303 1343 337
rect 1377 303 1400 337
rect 1320 280 1400 303
rect 1620 497 1700 530
rect 1620 463 1643 497
rect 1677 463 1700 497
rect 1620 417 1700 463
rect 1620 383 1643 417
rect 1677 383 1700 417
rect 1620 337 1700 383
rect 1620 303 1643 337
rect 1677 303 1700 337
rect 1620 280 1700 303
rect 640 220 720 240
rect 1040 220 1120 240
rect 40 217 1120 220
rect 40 183 663 217
rect 697 183 1063 217
rect 1097 183 1120 217
rect 40 180 1120 183
rect 640 160 720 180
rect 1040 160 1120 180
rect 40 97 1720 120
rect 40 63 63 97
rect 97 63 143 97
rect 177 63 223 97
rect 257 63 303 97
rect 337 63 383 97
rect 417 63 463 97
rect 497 63 543 97
rect 577 63 623 97
rect 657 63 703 97
rect 737 63 783 97
rect 817 63 863 97
rect 897 63 943 97
rect 977 63 1023 97
rect 1057 63 1103 97
rect 1137 63 1183 97
rect 1217 63 1263 97
rect 1297 63 1343 97
rect 1377 63 1423 97
rect 1457 63 1503 97
rect 1537 63 1583 97
rect 1617 63 1663 97
rect 1697 63 1720 97
rect 40 40 1720 63
<< viali >>
rect 63 1243 97 1277
rect 143 1243 177 1277
rect 223 1243 257 1277
rect 303 1243 337 1277
rect 383 1243 417 1277
rect 463 1243 497 1277
rect 543 1243 577 1277
rect 623 1243 657 1277
rect 703 1243 737 1277
rect 783 1243 817 1277
rect 863 1243 897 1277
rect 943 1243 977 1277
rect 1023 1243 1057 1277
rect 1103 1243 1137 1277
rect 1183 1243 1217 1277
rect 1263 1243 1297 1277
rect 1343 1243 1377 1277
rect 1423 1243 1457 1277
rect 1503 1243 1537 1277
rect 1583 1243 1617 1277
rect 1663 1243 1697 1277
rect 413 1013 447 1047
rect 563 1023 597 1057
rect 413 893 447 927
rect 563 943 597 977
rect 563 863 597 897
rect 863 1023 897 1057
rect 863 943 897 977
rect 863 863 897 897
rect 1163 1023 1197 1057
rect 1543 1013 1577 1047
rect 1163 943 1197 977
rect 1163 863 1197 897
rect 1393 893 1427 927
rect 913 743 947 777
rect 1313 743 1347 777
rect 233 463 267 497
rect 233 383 267 417
rect 233 303 267 337
rect 563 463 597 497
rect 563 383 597 417
rect 563 303 597 337
rect 863 463 897 497
rect 863 383 897 417
rect 863 303 897 337
rect 1163 463 1197 497
rect 1163 383 1197 417
rect 1163 303 1197 337
rect 1643 463 1677 497
rect 1643 383 1677 417
rect 1643 303 1677 337
rect 63 63 97 97
rect 143 63 177 97
rect 223 63 257 97
rect 303 63 337 97
rect 383 63 417 97
rect 463 63 497 97
rect 543 63 577 97
rect 623 63 657 97
rect 703 63 737 97
rect 783 63 817 97
rect 863 63 897 97
rect 943 63 977 97
rect 1023 63 1057 97
rect 1103 63 1137 97
rect 1183 63 1217 97
rect 1263 63 1297 97
rect 1343 63 1377 97
rect 1423 63 1457 97
rect 1503 63 1537 97
rect 1583 63 1617 97
rect 1663 63 1697 97
<< metal1 >>
rect 40 1277 1720 1310
rect 40 1243 63 1277
rect 97 1243 143 1277
rect 177 1243 223 1277
rect 257 1243 303 1277
rect 337 1243 383 1277
rect 417 1243 463 1277
rect 497 1243 543 1277
rect 577 1243 623 1277
rect 657 1243 703 1277
rect 737 1243 783 1277
rect 817 1243 863 1277
rect 897 1243 943 1277
rect 977 1243 1023 1277
rect 1057 1243 1103 1277
rect 1137 1243 1183 1277
rect 1217 1243 1263 1277
rect 1297 1243 1343 1277
rect 1377 1243 1423 1277
rect 1457 1243 1503 1277
rect 1537 1243 1583 1277
rect 1617 1243 1663 1277
rect 1697 1243 1720 1277
rect 40 1210 1720 1243
rect 230 530 270 1210
rect 390 1056 470 1070
rect 390 1004 404 1056
rect 456 1004 470 1056
rect 390 990 470 1004
rect 540 1057 620 1210
rect 540 1023 563 1057
rect 597 1023 620 1057
rect 540 977 620 1023
rect 390 936 470 950
rect 390 884 404 936
rect 456 884 470 936
rect 390 870 470 884
rect 540 943 563 977
rect 597 943 620 977
rect 540 897 620 943
rect 540 863 563 897
rect 597 863 620 897
rect 540 840 620 863
rect 840 1057 920 1210
rect 840 1023 863 1057
rect 897 1023 920 1057
rect 840 977 920 1023
rect 840 943 863 977
rect 897 943 920 977
rect 840 897 920 943
rect 840 863 863 897
rect 897 863 920 897
rect 840 840 920 863
rect 1140 1057 1220 1210
rect 1140 1023 1163 1057
rect 1197 1023 1220 1057
rect 1140 977 1220 1023
rect 1520 1056 1600 1070
rect 1520 1004 1534 1056
rect 1586 1004 1600 1056
rect 1520 990 1600 1004
rect 1140 943 1163 977
rect 1197 943 1220 977
rect 1140 897 1220 943
rect 1140 863 1163 897
rect 1197 863 1220 897
rect 1370 936 1450 950
rect 1370 884 1384 936
rect 1436 884 1450 936
rect 1370 870 1450 884
rect 1140 840 1220 863
rect 890 780 970 800
rect 1290 780 1370 800
rect 890 777 1370 780
rect 890 743 913 777
rect 947 743 1313 777
rect 1347 743 1370 777
rect 890 740 1370 743
rect 890 720 970 740
rect 1290 720 1370 740
rect 1640 530 1680 1210
rect 210 497 290 530
rect 210 463 233 497
rect 267 463 290 497
rect 210 417 290 463
rect 210 383 233 417
rect 267 383 290 417
rect 210 337 290 383
rect 210 303 233 337
rect 267 303 290 337
rect 210 280 290 303
rect 540 497 620 530
rect 540 463 563 497
rect 597 463 620 497
rect 540 417 620 463
rect 540 383 563 417
rect 597 383 620 417
rect 540 337 620 383
rect 540 303 563 337
rect 597 303 620 337
rect 540 280 620 303
rect 840 497 920 530
rect 840 463 863 497
rect 897 463 920 497
rect 840 417 920 463
rect 840 383 863 417
rect 897 383 920 417
rect 840 337 920 383
rect 840 303 863 337
rect 897 303 920 337
rect 840 280 920 303
rect 1140 497 1220 530
rect 1140 463 1163 497
rect 1197 463 1220 497
rect 1140 417 1220 463
rect 1140 383 1163 417
rect 1197 383 1220 417
rect 1140 337 1220 383
rect 1140 303 1163 337
rect 1197 303 1220 337
rect 1140 280 1220 303
rect 1620 497 1700 530
rect 1620 463 1643 497
rect 1677 463 1700 497
rect 1620 417 1700 463
rect 1620 383 1643 417
rect 1677 383 1700 417
rect 1620 337 1700 383
rect 1620 303 1643 337
rect 1677 303 1700 337
rect 1620 280 1700 303
rect 560 130 600 280
rect 860 130 900 280
rect 1160 130 1200 280
rect 40 97 1720 130
rect 40 63 63 97
rect 97 63 143 97
rect 177 63 223 97
rect 257 63 303 97
rect 337 63 383 97
rect 417 63 463 97
rect 497 63 543 97
rect 577 63 623 97
rect 657 63 703 97
rect 737 63 783 97
rect 817 63 863 97
rect 897 63 943 97
rect 977 63 1023 97
rect 1057 63 1103 97
rect 1137 63 1183 97
rect 1217 63 1263 97
rect 1297 63 1343 97
rect 1377 63 1423 97
rect 1457 63 1503 97
rect 1537 63 1583 97
rect 1617 63 1663 97
rect 1697 63 1720 97
rect 40 30 1720 63
<< via1 >>
rect 404 1047 456 1056
rect 404 1013 413 1047
rect 413 1013 447 1047
rect 447 1013 456 1047
rect 404 1004 456 1013
rect 404 927 456 936
rect 404 893 413 927
rect 413 893 447 927
rect 447 893 456 927
rect 404 884 456 893
rect 1534 1047 1586 1056
rect 1534 1013 1543 1047
rect 1543 1013 1577 1047
rect 1577 1013 1586 1047
rect 1534 1004 1586 1013
rect 1384 927 1436 936
rect 1384 893 1393 927
rect 1393 893 1427 927
rect 1427 893 1436 927
rect 1384 884 1436 893
<< metal2 >>
rect 390 1056 470 1070
rect 390 1004 404 1056
rect 456 1050 470 1056
rect 1520 1056 1600 1070
rect 1520 1050 1534 1056
rect 456 1010 1534 1050
rect 456 1004 470 1010
rect 390 990 470 1004
rect 1520 1004 1534 1010
rect 1586 1004 1600 1056
rect 1520 990 1600 1004
rect 390 936 470 950
rect 390 884 404 936
rect 456 930 470 936
rect 1370 936 1450 950
rect 1370 930 1384 936
rect 456 890 1384 930
rect 456 884 470 890
rect 390 870 470 884
rect 1370 884 1384 890
rect 1436 884 1450 936
rect 1370 870 1450 884
<< labels >>
rlabel locali s 810 615 850 655 4 OUT
port 1 nsew
rlabel locali s 50 1020 70 1040 4 A
port 2 nsew
rlabel locali s 50 800 70 820 4 A_bar
port 3 nsew
rlabel locali s 50 900 70 920 4 B
port 4 nsew
rlabel locali s 50 700 70 720 4 B_bar
port 5 nsew
rlabel locali s 660 180 700 220 4 Dis
port 6 nsew
rlabel metal1 s 910 740 950 780 4 OUT_bar
port 7 nsew
rlabel metal1 s 860 60 900 100 4 GND!
port 8 nsew
rlabel metal1 s 860 1240 900 1280 4 CLK
port 9 nsew
<< end >>
