magic
tech sky130A
timestamp 1665783531
<< nwell >>
rect -1080 910 -175 1000
rect -770 545 -500 910
<< nmos >>
rect -990 290 -975 440
rect -915 290 -900 440
rect -750 290 -735 440
rect -675 290 -660 440
rect -600 290 -585 440
rect -525 290 -510 440
rect -360 290 -345 440
rect -285 290 -270 440
<< pmos >>
rect -675 570 -660 870
rect -600 570 -585 870
<< ndiff >>
rect -1050 405 -990 440
rect -1050 385 -1030 405
rect -1010 385 -990 405
rect -1050 365 -990 385
rect -1050 345 -1030 365
rect -1010 345 -990 365
rect -1050 325 -990 345
rect -1050 305 -1030 325
rect -1010 305 -990 325
rect -1050 290 -990 305
rect -975 405 -915 440
rect -975 385 -955 405
rect -935 385 -915 405
rect -975 365 -915 385
rect -975 345 -955 365
rect -935 345 -915 365
rect -975 325 -915 345
rect -975 305 -955 325
rect -935 305 -915 325
rect -975 290 -915 305
rect -900 405 -840 440
rect -900 385 -880 405
rect -860 385 -840 405
rect -900 365 -840 385
rect -900 345 -880 365
rect -860 345 -840 365
rect -900 325 -840 345
rect -900 305 -880 325
rect -860 305 -840 325
rect -900 290 -840 305
rect -810 405 -750 440
rect -810 385 -790 405
rect -770 385 -750 405
rect -810 365 -750 385
rect -810 345 -790 365
rect -770 345 -750 365
rect -810 325 -750 345
rect -810 305 -790 325
rect -770 305 -750 325
rect -810 290 -750 305
rect -735 405 -675 440
rect -735 385 -715 405
rect -695 385 -675 405
rect -735 365 -675 385
rect -735 345 -715 365
rect -695 345 -675 365
rect -735 325 -675 345
rect -735 305 -715 325
rect -695 305 -675 325
rect -735 290 -675 305
rect -660 405 -600 440
rect -660 385 -640 405
rect -620 385 -600 405
rect -660 365 -600 385
rect -660 345 -640 365
rect -620 345 -600 365
rect -660 325 -600 345
rect -660 305 -640 325
rect -620 305 -600 325
rect -660 290 -600 305
rect -585 405 -525 440
rect -585 385 -565 405
rect -545 385 -525 405
rect -585 365 -525 385
rect -585 345 -565 365
rect -545 345 -525 365
rect -585 325 -525 345
rect -585 305 -565 325
rect -545 305 -525 325
rect -585 290 -525 305
rect -510 405 -450 440
rect -510 385 -490 405
rect -470 385 -450 405
rect -510 365 -450 385
rect -510 345 -490 365
rect -470 345 -450 365
rect -510 325 -450 345
rect -510 305 -490 325
rect -470 305 -450 325
rect -510 290 -450 305
rect -420 405 -360 440
rect -420 385 -400 405
rect -380 385 -360 405
rect -420 365 -360 385
rect -420 345 -400 365
rect -380 345 -360 365
rect -420 325 -360 345
rect -420 305 -400 325
rect -380 305 -360 325
rect -420 290 -360 305
rect -345 290 -285 440
rect -270 405 -210 440
rect -270 385 -250 405
rect -230 385 -210 405
rect -270 365 -210 385
rect -270 345 -250 365
rect -230 345 -210 365
rect -270 325 -210 345
rect -270 305 -250 325
rect -230 305 -210 325
rect -270 290 -210 305
<< pdiff >>
rect -735 845 -675 870
rect -735 825 -715 845
rect -695 825 -675 845
rect -735 805 -675 825
rect -735 785 -715 805
rect -695 785 -675 805
rect -735 765 -675 785
rect -735 745 -715 765
rect -695 745 -675 765
rect -735 725 -675 745
rect -735 705 -715 725
rect -695 705 -675 725
rect -735 685 -675 705
rect -735 665 -715 685
rect -695 665 -675 685
rect -735 645 -675 665
rect -735 625 -715 645
rect -695 625 -675 645
rect -735 605 -675 625
rect -735 585 -715 605
rect -695 585 -675 605
rect -735 570 -675 585
rect -660 845 -600 870
rect -660 825 -640 845
rect -620 825 -600 845
rect -660 805 -600 825
rect -660 785 -640 805
rect -620 785 -600 805
rect -660 765 -600 785
rect -660 745 -640 765
rect -620 745 -600 765
rect -660 725 -600 745
rect -660 705 -640 725
rect -620 705 -600 725
rect -660 685 -600 705
rect -660 665 -640 685
rect -620 665 -600 685
rect -660 645 -600 665
rect -660 625 -640 645
rect -620 625 -600 645
rect -660 605 -600 625
rect -660 585 -640 605
rect -620 585 -600 605
rect -660 570 -600 585
rect -585 845 -525 870
rect -585 825 -565 845
rect -545 825 -525 845
rect -585 805 -525 825
rect -585 785 -565 805
rect -545 785 -525 805
rect -585 765 -525 785
rect -585 745 -565 765
rect -545 745 -525 765
rect -585 725 -525 745
rect -585 705 -565 725
rect -545 705 -525 725
rect -585 685 -525 705
rect -585 665 -565 685
rect -545 665 -525 685
rect -585 645 -525 665
rect -585 625 -565 645
rect -545 625 -525 645
rect -585 605 -525 625
rect -585 585 -565 605
rect -545 585 -525 605
rect -585 570 -525 585
<< ndiffc >>
rect -1030 385 -1010 405
rect -1030 345 -1010 365
rect -1030 305 -1010 325
rect -955 385 -935 405
rect -955 345 -935 365
rect -955 305 -935 325
rect -880 385 -860 405
rect -880 345 -860 365
rect -880 305 -860 325
rect -790 385 -770 405
rect -790 345 -770 365
rect -790 305 -770 325
rect -715 385 -695 405
rect -715 345 -695 365
rect -715 305 -695 325
rect -640 385 -620 405
rect -640 345 -620 365
rect -640 305 -620 325
rect -565 385 -545 405
rect -565 345 -545 365
rect -565 305 -545 325
rect -490 385 -470 405
rect -490 345 -470 365
rect -490 305 -470 325
rect -400 385 -380 405
rect -400 345 -380 365
rect -400 305 -380 325
rect -250 385 -230 405
rect -250 345 -230 365
rect -250 305 -230 325
<< pdiffc >>
rect -715 825 -695 845
rect -715 785 -695 805
rect -715 745 -695 765
rect -715 705 -695 725
rect -715 665 -695 685
rect -715 625 -695 645
rect -715 585 -695 605
rect -640 825 -620 845
rect -640 785 -620 805
rect -640 745 -620 765
rect -640 705 -620 725
rect -640 665 -620 685
rect -640 625 -620 645
rect -640 585 -620 605
rect -565 825 -545 845
rect -565 785 -545 805
rect -565 745 -545 765
rect -565 705 -545 725
rect -565 665 -545 685
rect -565 625 -545 645
rect -565 585 -545 605
<< psubdiff >>
rect -1065 -15 -200 0
rect -1065 -35 -1045 -15
rect -1025 -35 -1005 -15
rect -985 -35 -965 -15
rect -945 -35 -925 -15
rect -905 -35 -885 -15
rect -865 -35 -845 -15
rect -825 -35 -805 -15
rect -785 -35 -765 -15
rect -745 -35 -725 -15
rect -705 -35 -685 -15
rect -665 -35 -645 -15
rect -625 -35 -605 -15
rect -585 -35 -565 -15
rect -545 -35 -525 -15
rect -505 -35 -485 -15
rect -465 -35 -445 -15
rect -425 -35 -400 -15
rect -380 -35 -360 -15
rect -340 -35 -320 -15
rect -300 -35 -280 -15
rect -260 -35 -240 -15
rect -220 -35 -200 -15
rect -1065 -50 -200 -35
<< nsubdiff >>
rect -1060 965 -195 980
rect -1060 945 -1040 965
rect -1020 945 -1000 965
rect -980 945 -960 965
rect -940 945 -920 965
rect -900 945 -880 965
rect -860 945 -840 965
rect -820 945 -800 965
rect -780 945 -760 965
rect -740 945 -720 965
rect -700 945 -680 965
rect -660 945 -640 965
rect -620 945 -600 965
rect -580 945 -560 965
rect -540 945 -520 965
rect -500 945 -480 965
rect -460 945 -440 965
rect -420 945 -400 965
rect -380 945 -355 965
rect -335 945 -315 965
rect -295 945 -275 965
rect -255 945 -235 965
rect -215 945 -195 965
rect -1060 930 -195 945
<< psubdiffcont >>
rect -1045 -35 -1025 -15
rect -1005 -35 -985 -15
rect -965 -35 -945 -15
rect -925 -35 -905 -15
rect -885 -35 -865 -15
rect -845 -35 -825 -15
rect -805 -35 -785 -15
rect -765 -35 -745 -15
rect -725 -35 -705 -15
rect -685 -35 -665 -15
rect -645 -35 -625 -15
rect -605 -35 -585 -15
rect -565 -35 -545 -15
rect -525 -35 -505 -15
rect -485 -35 -465 -15
rect -445 -35 -425 -15
rect -400 -35 -380 -15
rect -360 -35 -340 -15
rect -320 -35 -300 -15
rect -280 -35 -260 -15
rect -240 -35 -220 -15
<< nsubdiffcont >>
rect -1040 945 -1020 965
rect -1000 945 -980 965
rect -960 945 -940 965
rect -920 945 -900 965
rect -880 945 -860 965
rect -840 945 -820 965
rect -800 945 -780 965
rect -760 945 -740 965
rect -720 945 -700 965
rect -680 945 -660 965
rect -640 945 -620 965
rect -600 945 -580 965
rect -560 945 -540 965
rect -520 945 -500 965
rect -480 945 -460 965
rect -440 945 -420 965
rect -400 945 -380 965
rect -355 945 -335 965
rect -315 945 -295 965
rect -275 945 -255 965
rect -235 945 -215 965
<< poly >>
rect -675 870 -660 885
rect -600 870 -585 885
rect -675 495 -660 570
rect -600 555 -585 570
rect -625 545 -585 555
rect -625 525 -615 545
rect -595 525 -585 545
rect -625 515 -585 525
rect -675 485 -635 495
rect -675 465 -665 485
rect -645 465 -635 485
rect -675 455 -635 465
rect -990 440 -975 455
rect -915 440 -900 455
rect -750 440 -735 455
rect -675 440 -660 455
rect -600 440 -585 515
rect -525 440 -510 455
rect -360 440 -345 455
rect -285 440 -270 455
rect -990 225 -975 290
rect -990 215 -950 225
rect -990 195 -980 215
rect -960 195 -950 215
rect -990 185 -950 195
rect -915 175 -900 290
rect -750 275 -735 290
rect -675 275 -660 290
rect -600 275 -585 290
rect -525 275 -510 290
rect -750 265 -710 275
rect -750 245 -740 265
rect -720 245 -710 265
rect -750 235 -710 245
rect -550 265 -510 275
rect -550 245 -540 265
rect -520 245 -510 265
rect -550 235 -510 245
rect -915 165 -875 175
rect -915 145 -905 165
rect -885 145 -875 165
rect -915 135 -875 145
rect -360 115 -345 290
rect -360 105 -320 115
rect -360 85 -350 105
rect -330 85 -320 105
rect -360 75 -320 85
rect -285 65 -270 290
rect -285 55 -245 65
rect -285 35 -275 55
rect -255 35 -245 55
rect -285 25 -245 35
<< polycont >>
rect -615 525 -595 545
rect -665 465 -645 485
rect -980 195 -960 215
rect -740 245 -720 265
rect -540 245 -520 265
rect -905 145 -885 165
rect -350 85 -330 105
rect -275 35 -255 55
<< locali >>
rect -1060 965 -195 975
rect -1060 945 -1040 965
rect -1020 945 -1000 965
rect -980 945 -960 965
rect -940 945 -920 965
rect -900 945 -880 965
rect -860 945 -840 965
rect -820 945 -800 965
rect -780 945 -760 965
rect -740 945 -720 965
rect -700 945 -680 965
rect -660 945 -640 965
rect -620 945 -600 965
rect -580 945 -560 965
rect -540 945 -520 965
rect -500 945 -480 965
rect -460 945 -440 965
rect -420 945 -400 965
rect -380 945 -355 965
rect -335 945 -315 965
rect -295 945 -275 965
rect -255 945 -235 965
rect -215 945 -195 965
rect -1060 935 -195 945
rect -725 845 -685 855
rect -725 825 -715 845
rect -695 825 -685 845
rect -725 805 -685 825
rect -725 785 -715 805
rect -695 785 -685 805
rect -725 765 -685 785
rect -725 745 -715 765
rect -695 745 -685 765
rect -725 725 -685 745
rect -725 705 -715 725
rect -695 705 -685 725
rect -725 685 -685 705
rect -725 665 -715 685
rect -695 665 -685 685
rect -725 645 -685 665
rect -725 625 -715 645
rect -695 625 -685 645
rect -725 605 -685 625
rect -725 585 -715 605
rect -695 585 -685 605
rect -725 570 -685 585
rect -650 845 -610 855
rect -650 825 -640 845
rect -620 825 -610 845
rect -650 805 -610 825
rect -650 785 -640 805
rect -620 785 -610 805
rect -650 765 -610 785
rect -650 745 -640 765
rect -620 745 -610 765
rect -650 725 -610 745
rect -650 705 -640 725
rect -620 705 -610 725
rect -650 685 -610 705
rect -650 665 -640 685
rect -620 665 -610 685
rect -650 645 -610 665
rect -650 625 -640 645
rect -620 625 -610 645
rect -650 605 -610 625
rect -650 585 -640 605
rect -620 585 -610 605
rect -650 575 -610 585
rect -575 845 -535 855
rect -575 825 -565 845
rect -545 825 -535 845
rect -575 805 -535 825
rect -575 785 -565 805
rect -545 785 -535 805
rect -575 765 -535 785
rect -575 745 -565 765
rect -545 745 -535 765
rect -575 725 -535 745
rect -575 705 -565 725
rect -545 705 -535 725
rect -575 685 -535 705
rect -575 665 -565 685
rect -545 665 -535 685
rect -575 645 -535 665
rect -575 625 -565 645
rect -545 625 -535 645
rect -575 605 -535 625
rect -575 585 -565 605
rect -545 585 -535 605
rect -575 570 -535 585
rect -715 545 -695 570
rect -625 545 -585 555
rect -715 525 -615 545
rect -595 525 -585 545
rect -715 480 -695 525
rect -625 515 -585 525
rect -1030 460 -695 480
rect -1030 420 -1010 460
rect -880 420 -860 460
rect -715 440 -695 460
rect -675 485 -635 495
rect -565 485 -545 570
rect -675 465 -665 485
rect -645 465 -230 485
rect -675 455 -635 465
rect -565 440 -545 465
rect -1040 405 -1000 420
rect -1040 385 -1030 405
rect -1010 385 -1000 405
rect -1040 365 -1000 385
rect -1040 345 -1030 365
rect -1010 345 -1000 365
rect -1040 325 -1000 345
rect -1040 305 -1030 325
rect -1010 305 -1000 325
rect -1040 295 -1000 305
rect -965 405 -925 420
rect -965 385 -955 405
rect -935 385 -925 405
rect -965 365 -925 385
rect -965 345 -955 365
rect -935 345 -925 365
rect -965 325 -925 345
rect -965 305 -955 325
rect -935 305 -925 325
rect -965 295 -925 305
rect -890 405 -850 420
rect -890 385 -880 405
rect -860 385 -850 405
rect -890 365 -850 385
rect -890 345 -880 365
rect -860 345 -850 365
rect -890 325 -850 345
rect -890 305 -880 325
rect -860 305 -850 325
rect -890 295 -850 305
rect -800 405 -760 420
rect -800 385 -790 405
rect -770 385 -760 405
rect -800 365 -760 385
rect -800 345 -790 365
rect -770 345 -760 365
rect -800 325 -760 345
rect -800 305 -790 325
rect -770 305 -760 325
rect -800 295 -760 305
rect -725 405 -685 440
rect -725 385 -715 405
rect -695 385 -685 405
rect -725 365 -685 385
rect -725 345 -715 365
rect -695 345 -685 365
rect -725 325 -685 345
rect -725 305 -715 325
rect -695 305 -685 325
rect -725 295 -685 305
rect -650 405 -610 420
rect -650 385 -640 405
rect -620 385 -610 405
rect -650 365 -610 385
rect -650 345 -640 365
rect -620 345 -610 365
rect -650 325 -610 345
rect -650 305 -640 325
rect -620 305 -610 325
rect -650 295 -610 305
rect -575 405 -535 440
rect -250 420 -230 465
rect -575 385 -565 405
rect -545 385 -535 405
rect -575 365 -535 385
rect -575 345 -565 365
rect -545 345 -535 365
rect -575 325 -535 345
rect -575 305 -565 325
rect -545 305 -535 325
rect -575 295 -535 305
rect -500 405 -460 420
rect -500 385 -490 405
rect -470 385 -460 405
rect -500 365 -460 385
rect -500 345 -490 365
rect -470 345 -460 365
rect -500 325 -460 345
rect -500 305 -490 325
rect -470 305 -460 325
rect -500 295 -460 305
rect -410 405 -370 420
rect -410 385 -400 405
rect -380 385 -370 405
rect -410 365 -370 385
rect -410 345 -400 365
rect -380 345 -370 365
rect -410 325 -370 345
rect -410 305 -400 325
rect -380 305 -370 325
rect -410 295 -370 305
rect -260 405 -220 420
rect -260 385 -250 405
rect -230 385 -220 405
rect -260 365 -220 385
rect -260 345 -250 365
rect -230 345 -220 365
rect -260 325 -220 345
rect -260 305 -250 325
rect -230 305 -220 325
rect -260 295 -220 305
rect -750 265 -710 275
rect -550 265 -510 275
rect -1050 245 -740 265
rect -720 245 -540 265
rect -520 245 -510 265
rect -750 235 -710 245
rect -550 235 -510 245
rect -990 215 -950 225
rect -1050 195 -980 215
rect -960 195 -950 215
rect -990 185 -950 195
rect -915 165 -875 175
rect -1050 145 -905 165
rect -885 145 -875 165
rect -915 135 -875 145
rect -360 105 -320 115
rect -1050 85 -350 105
rect -330 85 -320 105
rect -360 75 -320 85
rect -285 55 -245 65
rect -1050 35 -275 55
rect -255 35 -245 55
rect -285 25 -245 35
rect -1065 -15 -200 -5
rect -1065 -35 -1045 -15
rect -1025 -35 -1005 -15
rect -985 -35 -965 -15
rect -945 -35 -925 -15
rect -905 -35 -885 -15
rect -865 -35 -845 -15
rect -825 -35 -805 -15
rect -785 -35 -765 -15
rect -745 -35 -725 -15
rect -705 -35 -685 -15
rect -665 -35 -645 -15
rect -625 -35 -605 -15
rect -585 -35 -565 -15
rect -545 -35 -525 -15
rect -505 -35 -485 -15
rect -465 -35 -445 -15
rect -425 -35 -400 -15
rect -380 -35 -360 -15
rect -340 -35 -320 -15
rect -300 -35 -280 -15
rect -260 -35 -240 -15
rect -220 -35 -200 -15
rect -1065 -45 -200 -35
<< viali >>
rect -1040 945 -1020 965
rect -1000 945 -980 965
rect -960 945 -940 965
rect -920 945 -900 965
rect -880 945 -860 965
rect -840 945 -820 965
rect -800 945 -780 965
rect -760 945 -740 965
rect -720 945 -700 965
rect -680 945 -660 965
rect -640 945 -620 965
rect -600 945 -580 965
rect -560 945 -540 965
rect -520 945 -500 965
rect -480 945 -460 965
rect -440 945 -420 965
rect -400 945 -380 965
rect -355 945 -335 965
rect -315 945 -295 965
rect -275 945 -255 965
rect -235 945 -215 965
rect -640 825 -620 845
rect -640 785 -620 805
rect -640 745 -620 765
rect -640 705 -620 725
rect -640 665 -620 685
rect -640 625 -620 645
rect -640 585 -620 605
rect -955 385 -935 405
rect -955 345 -935 365
rect -955 305 -935 325
rect -790 385 -770 405
rect -790 345 -770 365
rect -790 305 -770 325
rect -640 385 -620 405
rect -640 345 -620 365
rect -640 305 -620 325
rect -490 385 -470 405
rect -490 345 -470 365
rect -490 305 -470 325
rect -400 385 -380 405
rect -400 345 -380 365
rect -400 305 -380 325
rect -1045 -35 -1025 -15
rect -1005 -35 -985 -15
rect -965 -35 -945 -15
rect -925 -35 -905 -15
rect -885 -35 -865 -15
rect -845 -35 -825 -15
rect -805 -35 -785 -15
rect -765 -35 -745 -15
rect -725 -35 -705 -15
rect -685 -35 -665 -15
rect -645 -35 -625 -15
rect -605 -35 -585 -15
rect -565 -35 -545 -15
rect -525 -35 -505 -15
rect -485 -35 -465 -15
rect -445 -35 -425 -15
rect -400 -35 -380 -15
rect -360 -35 -340 -15
rect -320 -35 -300 -15
rect -280 -35 -260 -15
rect -240 -35 -220 -15
<< metal1 >>
rect -1060 965 -195 980
rect -1060 945 -1040 965
rect -1020 945 -1000 965
rect -980 945 -960 965
rect -940 945 -920 965
rect -900 945 -880 965
rect -860 945 -840 965
rect -820 945 -800 965
rect -780 945 -760 965
rect -740 945 -720 965
rect -700 945 -680 965
rect -660 945 -640 965
rect -620 945 -600 965
rect -580 945 -560 965
rect -540 945 -520 965
rect -500 945 -480 965
rect -460 945 -440 965
rect -420 945 -400 965
rect -380 945 -355 965
rect -335 945 -315 965
rect -295 945 -275 965
rect -255 945 -235 965
rect -215 945 -195 965
rect -1060 930 -195 945
rect -955 420 -935 930
rect -640 855 -620 930
rect -650 845 -610 855
rect -650 825 -640 845
rect -620 825 -610 845
rect -650 805 -610 825
rect -650 785 -640 805
rect -620 785 -610 805
rect -650 765 -610 785
rect -650 745 -640 765
rect -620 745 -610 765
rect -650 725 -610 745
rect -650 705 -640 725
rect -620 705 -610 725
rect -650 685 -610 705
rect -650 665 -640 685
rect -620 665 -610 685
rect -650 645 -610 665
rect -650 625 -640 645
rect -620 625 -610 645
rect -650 605 -610 625
rect -650 585 -640 605
rect -620 585 -610 605
rect -650 575 -610 585
rect -400 420 -380 930
rect -965 405 -925 420
rect -965 385 -955 405
rect -935 385 -925 405
rect -965 365 -925 385
rect -965 345 -955 365
rect -935 345 -925 365
rect -965 325 -925 345
rect -965 305 -955 325
rect -935 305 -925 325
rect -965 295 -925 305
rect -800 405 -760 420
rect -800 385 -790 405
rect -770 385 -760 405
rect -800 365 -760 385
rect -800 345 -790 365
rect -770 345 -760 365
rect -800 325 -760 345
rect -800 305 -790 325
rect -770 305 -760 325
rect -800 295 -760 305
rect -650 405 -610 420
rect -650 385 -640 405
rect -620 385 -610 405
rect -650 365 -610 385
rect -650 345 -640 365
rect -620 345 -610 365
rect -650 325 -610 345
rect -650 305 -640 325
rect -620 305 -610 325
rect -650 295 -610 305
rect -500 405 -460 420
rect -500 385 -490 405
rect -470 385 -460 405
rect -500 365 -460 385
rect -500 345 -490 365
rect -470 345 -460 365
rect -500 325 -460 345
rect -500 305 -490 325
rect -470 305 -460 325
rect -500 295 -460 305
rect -410 405 -370 420
rect -410 385 -400 405
rect -380 385 -370 405
rect -410 365 -370 385
rect -410 345 -400 365
rect -380 345 -370 365
rect -410 325 -370 345
rect -410 305 -400 325
rect -380 305 -370 325
rect -410 295 -370 305
rect -790 0 -770 295
rect -640 0 -620 295
rect -490 0 -470 295
rect -1065 -15 -200 0
rect -1065 -35 -1045 -15
rect -1025 -35 -1005 -15
rect -985 -35 -965 -15
rect -945 -35 -925 -15
rect -905 -35 -885 -15
rect -865 -35 -845 -15
rect -825 -35 -805 -15
rect -785 -35 -765 -15
rect -745 -35 -725 -15
rect -705 -35 -685 -15
rect -665 -35 -645 -15
rect -625 -35 -605 -15
rect -585 -35 -565 -15
rect -545 -35 -525 -15
rect -505 -35 -485 -15
rect -465 -35 -445 -15
rect -425 -35 -400 -15
rect -380 -35 -360 -15
rect -340 -35 -320 -15
rect -300 -35 -280 -15
rect -260 -35 -240 -15
rect -220 -35 -200 -15
rect -1065 -50 -200 -35
<< labels >>
rlabel locali -440 90 -430 100 7 A
port 1 w
rlabel locali -1045 200 -1035 210 7 A_bar
port 2 w
rlabel locali -440 40 -430 50 7 B
port 3 w
rlabel locali -1045 150 -1035 160 7 B_bar
port 4 w
rlabel locali -490 470 -480 480 3 OUT
port 5 e
rlabel locali -790 465 -780 475 7 OUT_bar
port 6 w
rlabel locali -805 250 -795 260 7 Dis
port 7 w
rlabel metal1 -640 945 -620 965 1 CLK
port 8 n
rlabel metal1 -645 -35 -625 -15 5 GND!
port 9 s
<< end >>
