* NGSPICE file created from EESPFAL_s0.ext - technology: sky130A

.subckt EESPFAL_XOR_v3 OUT A A_bar B B_bar Dis OUT_bar GND CLK
X0 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X2 a_n840_410# A CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=7.5e+12p ps=3.22e+07u w=1.5e+06u l=150000u
X3 a_n1140_410# B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_420_410# B_bar OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X5 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X7 a_720_410# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar B a_n840_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 CLK A_bar a_n1140_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK A a_420_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 OUT B a_720_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_NOR_v3 OUT A A_bar B B_bar Dis OUT_bar GND CLK
X0 a_n1820_550# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=6e+12p ps=2.62e+07u w=1.5e+06u l=150000u
X1 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X2 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u M=2
X3 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X4 OUT_bar B_bar a_n1820_550# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X6 OUT A CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 CLK B OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_NAND_v3 OUT A A_bar B B_bar Dis OUT_bar GND CLK
X0 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X2 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X3 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X5 OUT_bar A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6e+12p ps=2.62e+07u w=1.5e+06u l=150000u
X6 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_501_n414# B OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 CLK A a_501_n414# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 CLK B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_s0 GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar CLK1 Dis1 CLK3 Dis2
+ CLK2 Dis3 s0 s0_bar
XEESPFAL_XOR_v3_0 EESPFAL_NAND_v3_0/A x0 x0_bar x3 x3_bar Dis1 EESPFAL_NAND_v3_1/A
+ GND CLK1 EESPFAL_XOR_v3
XEESPFAL_NOR_v3_0 s0 EESPFAL_NOR_v3_0/A EESPFAL_NOR_v3_0/A_bar EESPFAL_NOR_v3_0/B
+ EESPFAL_NOR_v3_0/B_bar Dis3 s0_bar GND CLK3 EESPFAL_NOR_v3
XEESPFAL_NOR_v3_1 EESPFAL_NAND_v3_0/B x1 x1_bar x2_bar x2 Dis1 EESPFAL_NAND_v3_0/B_bar
+ GND CLK1 EESPFAL_NOR_v3
XEESPFAL_NAND_v3_0 EESPFAL_NOR_v3_0/A EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_0/B
+ EESPFAL_NAND_v3_0/B_bar Dis2 EESPFAL_NOR_v3_0/A_bar GND CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_1 EESPFAL_NOR_v3_0/B EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/B
+ EESPFAL_NAND_v3_1/B_bar Dis2 EESPFAL_NOR_v3_0/B_bar GND CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_2 EESPFAL_NAND_v3_1/B x2 x2_bar x1_bar x1 Dis1 EESPFAL_NAND_v3_1/B_bar
+ GND CLK1 EESPFAL_NAND_v3
.ends

