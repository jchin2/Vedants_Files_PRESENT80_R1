* NGSPICE file created from EESPFAL_s2_draft2.ext - technology: sky130A

.subckt EESPFAL_4in_NAND OUT A A_bar B B_bar C C_bar D D_bar Dis OUT_bar GND CLK
X0 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=3.6e+12p pd=1.68e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X1 CLK B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=8.5e+12p pd=3.68e+07u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n1040_180# B a_n1190_180# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 OUT_bar OUT CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u M=2
X4 CLK D_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n1340_180# D OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT_bar A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar C_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X11 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK A a_n1040_180# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_n1190_180# C a_n1340_180# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_INV4 OUT_bar A A_bar Dis OUT GND CLK
X0 OUT A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=5.25e+12p ps=2.32e+07u w=1.5e+06u l=150000u
X1 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X2 GND Dis OUT_bar GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X3 GND OUT_bar OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X5 OUT_bar OUT GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 CLK A OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT Dis GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_XOR_v3 OUT A A_bar B B_bar Dis OUT_bar GND CLK
X0 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X2 a_n840_410# A CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=7.5e+12p ps=3.22e+07u w=1.5e+06u l=150000u
X3 a_n1140_410# B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_420_410# B_bar OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X5 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X7 a_720_410# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar B a_n840_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 CLK A_bar a_n1140_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK A a_420_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 OUT B a_720_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_3in_NOR_v2 OUT A A_bar B B_bar C C_bar Dis OUT_bar GND CLK
X0 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 OUT B CLK GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=7.7e+12p ps=3.36e+07u w=1.5e+06u l=150000u
X2 OUT_bar OUT CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X3 a_n1990_570# B_bar a_n2140_570# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X4 CLK A OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X6 CLK C OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n2140_570# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 OUT_bar C_bar a_n1990_570# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_NAND_v3 OUT A A_bar B B_bar Dis OUT_bar GND CLK
X0 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 CLK A a_n2940_320# GND sky130_fd_pr__nfet_01v8 ad=6e+12p pd=2.62e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X2 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X3 CLK B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X4 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X5 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 OUT_bar A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n2940_320# B OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_s2_draft2 GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar CLK1 Dis1 Dis3
+ Dis2 CLK3 CLK2 s2_bar s2
XEESPFAL_4in_NAND_0 EESPFAL_INV4_2/A x3_bar x3 x1 x1_bar x0 x0_bar x2 x2_bar Dis1
+ EESPFAL_INV4_2/A_bar GND CLK1 EESPFAL_4in_NAND
XEESPFAL_INV4_1 EESPFAL_NAND_v3_1/B x1 x1_bar Dis1 EESPFAL_INV4_1/OUT GND CLK1 EESPFAL_INV4
XEESPFAL_INV4_0 EESPFAL_NAND_v3_0/B x2_bar x2 Dis1 EESPFAL_INV4_0/OUT GND CLK1 EESPFAL_INV4
XEESPFAL_INV4_2 EESPFAL_INV4_2/OUT_bar EESPFAL_INV4_2/A EESPFAL_INV4_2/A_bar Dis2
+ EESPFAL_INV4_2/OUT GND CLK2 EESPFAL_INV4
XEESPFAL_XOR_v3_0 EESPFAL_XOR_v3_0/OUT x3 x3_bar x2 x2_bar Dis1 EESPFAL_NAND_v3_1/A
+ GND CLK1 EESPFAL_XOR_v3
XEESPFAL_XOR_v3_1 EESPFAL_NAND_v3_0/A x1 x1_bar x0 x0_bar Dis1 EESPFAL_NAND_v3_0/A_bar
+ GND CLK1 EESPFAL_XOR_v3
XEESPFAL_3in_NOR_v2_0 s2 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_0/OUT
+ EESPFAL_NAND_v3_0/OUT_bar EESPFAL_INV4_2/OUT_bar EESPFAL_INV4_2/OUT Dis3 s2_bar
+ GND CLK3 EESPFAL_3in_NOR_v2
XEESPFAL_NAND_v3_0 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/A_bar
+ EESPFAL_NAND_v3_0/B EESPFAL_INV4_0/OUT Dis2 EESPFAL_NAND_v3_0/OUT_bar GND CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_1 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/A EESPFAL_XOR_v3_0/OUT
+ EESPFAL_NAND_v3_1/B EESPFAL_INV4_1/OUT Dis2 EESPFAL_NAND_v3_1/OUT_bar GND CLK2 EESPFAL_NAND_v3
.ends

