* NGSPICE file created from Mixer_LVS_test1.ext - technology: sky130A

.subckt Mixer_LVS_test1 v_bias_p RFP RFN LOP LON VoutP VoutN Ground VDD
X0 VDD v_bias_p a_2038_n6423# VDD sky130_fd_pr__pfet_01v8_lvt ad=1.425e+13p pd=5.35e+07u as=5.7e+12p ps=2.14e+07u w=4.75e+06u l=500000u M=4
X1 a_2038_n6423# LON VoutN Ground sky130_fd_pr__nfet_01v8_lvt ad=1.83e+13p pd=6.94e+07u as=1.008e+13p ps=3.84e+07u w=4.2e+06u l=500000u M=4
X2 VDD v_bias_p a_5592_n6455# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.7e+12p ps=2.14e+07u w=4.75e+06u l=500000u M=4
X3 Ground RFP a_2038_n6423# Ground sky130_fd_pr__nfet_01v8_lvt ad=1.425e+13p pd=5.35e+07u as=0p ps=0u w=4.75e+06u l=500000u M=4
X4 Ground RFN a_5592_n6455# Ground sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.83e+13p ps=6.94e+07u w=4.75e+06u l=500000u M=4
X5 VoutP LOP a_2038_n6423# Ground sky130_fd_pr__nfet_01v8_lvt ad=1.008e+13p pd=3.84e+07u as=0p ps=0u w=4.2e+06u l=500000u M=4
X6 VoutN LOP a_5592_n6455# Ground sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.2e+06u l=500000u M=4
X7 VoutP VDD Ground sky130_fd_pr__res_xhigh_po w=350000u l=690000u
X8 VoutP LON a_5592_n6455# Ground sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.2e+06u l=500000u M=4
X9 VoutN VDD Ground sky130_fd_pr__res_xhigh_po w=350000u l=690000u
.ends

