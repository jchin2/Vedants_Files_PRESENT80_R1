* NGSPICE file created from CMOS_PRESENT80_SB.ext - technology: sky130A

.subckt CMOS_XOR GND B A_bar A B_bar XOR VDD
X0 a_90_0# A_bar XOR VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X1 VDD B a_90_0# VDD sky130_fd_pr__pfet_01v8 ad=3.6e+12p pd=1.44e+07u as=0p ps=0u w=3e+06u l=150000u
X2 a_n210_n610# A GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X3 GND A_bar a_90_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X4 XOR A a_n210_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X5 a_n210_0# B_bar VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X6 a_90_n610# B_bar XOR GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X7 XOR B a_n210_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt CMOS_INV OUT A VDD GND
X0 OUT A GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X1 OUT A VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
.ends

.subckt CMOS_4in_XOR VDD x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar x2 x2_bar k2 k2_bar
+ x3 x3_bar k3 k3_bar XOR1 XOR0 XOR2 XOR3 XOR0_bar XOR1_bar XOR2_bar XOR3_bar CMOS_XOR_3/GND
XCMOS_XOR_1 CMOS_XOR_3/GND k3 x3_bar x3 k3_bar XOR3 VDD CMOS_XOR
XCMOS_XOR_2 CMOS_XOR_3/GND k1 x1_bar x1 k1_bar XOR1 VDD CMOS_XOR
XCMOS_XOR_3 CMOS_XOR_3/GND k0 x0_bar x0 k0_bar XOR0 VDD CMOS_XOR
XCMOS_INV_0 XOR3_bar XOR3 VDD CMOS_XOR_3/GND CMOS_INV
XCMOS_INV_1 XOR1_bar XOR1 VDD CMOS_XOR_3/GND CMOS_INV
XCMOS_INV_2 XOR0_bar XOR0 VDD CMOS_XOR_3/GND CMOS_INV
XCMOS_INV_3 XOR2_bar XOR2 VDD CMOS_XOR_3/GND CMOS_INV
XCMOS_XOR_0 CMOS_XOR_3/GND k2 x2_bar x2 k2_bar XOR2 VDD CMOS_XOR
.ends

.subckt CMOS_AND GND AND A B VDD
X0 a_n265_0# B VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=5.4e+12p ps=2.16e+07u w=3e+06u l=150000u
X1 VDD A a_n265_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2 a_n265_0# A a_n265_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 AND a_n265_0# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X4 a_n265_n610# B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X5 AND a_n265_0# GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt CMOS_3in_OR GND A B C OR VDD
X0 a_n480_n610# B GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X1 OR a_n480_n610# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X2 a_n480_n610# C a_n180_0# VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X3 GND A a_n480_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 OR a_n480_n610# GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n330_0# A VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X6 a_n180_0# B a_n330_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X7 GND C a_n480_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt CMOS_XNOR GND XNOR B A_bar A B_bar a_n233_n610# VDD
X0 XNOR a_n233_n610# GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X1 a_n383_n610# A GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n233_n610# B a_n383_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n383_0# B_bar VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=5.4e+12p ps=2.16e+07u w=3e+06u l=150000u
X4 a_n233_n610# A a_n383_0# VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X5 a_n83_0# A_bar a_n233_n610# VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X6 a_n83_n610# B_bar a_n233_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 GND A_bar a_n83_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 XNOR a_n233_n610# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X9 VDD B a_n83_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
.ends

.subckt CMOS_3in_AND GND A B C OUT VDD
X0 a_n180_n610# B a_n330_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X1 OUT a_n480_0# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=5.4e+12p ps=2.16e+07u w=3e+06u l=150000u
X2 VDD A a_n480_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X3 a_n330_n610# C GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X4 OUT a_n480_0# GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 VDD C a_n480_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X6 a_n480_0# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X7 a_n480_0# A a_n180_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt CMOS_s3 CMOS_XOR_0/GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar s3 VDD
XCMOS_AND_0 CMOS_XOR_0/GND CMOS_AND_0/AND CMOS_AND_0/A x1 VDD CMOS_AND
XCMOS_AND_1 CMOS_XOR_0/GND CMOS_AND_1/AND CMOS_AND_1/A x3_bar VDD CMOS_AND
XCMOS_3in_OR_0 CMOS_XOR_0/GND CMOS_AND_1/AND CMOS_AND_0/AND CMOS_3in_OR_0/C s3 VDD
+ CMOS_3in_OR
XCMOS_XNOR_0 CMOS_XOR_0/GND CMOS_AND_1/A x0 x1_bar x1 x0_bar CMOS_XNOR_0/a_n233_n610#
+ VDD CMOS_XNOR
XCMOS_3in_AND_0 CMOS_XOR_0/GND x2_bar x0 x3 CMOS_3in_OR_0/C VDD CMOS_3in_AND
XCMOS_XOR_0 CMOS_XOR_0/GND x3 x2_bar x2 x3_bar CMOS_AND_0/A VDD CMOS_XOR
.ends

.subckt CMOS_s1 CMOS_XOR_0/GND x0 x0_bar x1 x1_bar x2 x2_bar x3 s1 x3_bar VDD
XCMOS_AND_0 CMOS_XOR_0/GND CMOS_AND_0/AND CMOS_AND_0/A x2_bar VDD CMOS_AND
XCMOS_AND_1 CMOS_XOR_0/GND CMOS_AND_1/AND CMOS_AND_1/A x3 VDD CMOS_AND
XCMOS_3in_OR_0 CMOS_XOR_0/GND CMOS_AND_1/AND CMOS_AND_0/AND CMOS_3in_OR_0/C s1 VDD
+ CMOS_3in_OR
XCMOS_XNOR_0 CMOS_XOR_0/GND CMOS_AND_1/A x2 x0_bar x0 x2_bar CMOS_XNOR_0/a_n233_n610#
+ VDD CMOS_XNOR
XCMOS_3in_AND_0 CMOS_XOR_0/GND x3_bar x1 x0_bar CMOS_3in_OR_0/C VDD CMOS_3in_AND
XCMOS_XOR_0 CMOS_XOR_0/GND x3 x1_bar x1 x3_bar CMOS_AND_0/A VDD CMOS_XOR
.ends

.subckt CMOS_4in_AND GND OUT A B C D VDD
X0 a_n405_0# A a_n105_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X1 VDD C a_n405_0# VDD sky130_fd_pr__pfet_01v8 ad=7.2e+12p pd=2.88e+07u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X2 a_n405_0# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 a_n405_0# D VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4 VDD A a_n405_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X5 a_n105_n610# B a_n255_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X6 OUT a_n405_0# GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X7 a_n255_n610# C a_n405_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X8 OUT a_n405_0# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X9 a_n405_n610# D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt CMOS_s2 CMOS_XOR_0/GND x0 x0_bar x1 x2 x2_bar x3 s2 x3_bar x1_bar VDD
XCMOS_AND_0 CMOS_XOR_0/GND CMOS_AND_0/AND CMOS_AND_0/A x2_bar VDD CMOS_AND
XCMOS_AND_1 CMOS_XOR_0/GND CMOS_AND_1/AND CMOS_AND_1/A x1_bar VDD CMOS_AND
XCMOS_3in_OR_0 CMOS_XOR_0/GND CMOS_AND_1/AND CMOS_AND_0/AND CMOS_3in_OR_0/C s2 VDD
+ CMOS_3in_OR
XCMOS_4in_AND_0 CMOS_XOR_0/GND CMOS_3in_OR_0/C x3_bar x1 x0 x2 VDD CMOS_4in_AND
XCMOS_XNOR_0 CMOS_XOR_0/GND CMOS_AND_1/A x2 x3_bar x3 x2_bar CMOS_XNOR_0/a_n233_n610#
+ VDD CMOS_XNOR
XCMOS_XOR_0 CMOS_XOR_0/GND x0 x1_bar x1 x0_bar CMOS_AND_0/A VDD CMOS_XOR
.ends

.subckt CMOS_OR GND OR B A VDD
X0 a_n265_0# A VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X1 a_n265_n610# B a_n265_0# VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X2 GND B a_n265_n610# GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 OR a_n265_n610# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X4 a_n265_n610# A GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 OR a_n265_n610# GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt CMOS_s0 x3 x2_bar x2 x1_bar x1 x0 CMOS_OR_1/GND s0 x3_bar x0_bar VDD
XCMOS_AND_0 CMOS_OR_1/GND CMOS_OR_0/A CMOS_AND_0/A CMOS_OR_1/OR VDD CMOS_AND
XCMOS_AND_1 CMOS_OR_1/GND CMOS_OR_0/B CMOS_AND_1/A CMOS_AND_1/B VDD CMOS_AND
XCMOS_AND_2 CMOS_OR_1/GND CMOS_AND_1/A x2 x1_bar VDD CMOS_AND
XCMOS_XNOR_0 CMOS_OR_1/GND CMOS_AND_1/B x0 x3_bar x3 x0_bar li_n1053_n744# VDD CMOS_XNOR
XCMOS_OR_0 CMOS_OR_1/GND s0 CMOS_OR_0/B CMOS_OR_0/A VDD CMOS_OR
XCMOS_OR_1 CMOS_OR_1/GND CMOS_OR_1/OR x2_bar x1 VDD CMOS_OR
XCMOS_XOR_0 CMOS_OR_1/GND x3 x0_bar x0 x3_bar CMOS_AND_0/A VDD CMOS_XOR
.ends

.subckt CMOS_sbox x3 x2 x1_bar x1 x0_bar x0 CMOS_s0_0/CMOS_OR_1/GND s0 s1 s2 s3 x2_bar
+ x3_bar VDD
XCMOS_s3_0 CMOS_s0_0/CMOS_OR_1/GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar s3 VDD
+ CMOS_s3
XCMOS_s1_0 CMOS_s0_0/CMOS_OR_1/GND x0 x0_bar x1 x1_bar x2 x2_bar x3 s1 x3_bar VDD
+ CMOS_s1
XCMOS_s2_0 CMOS_s0_0/CMOS_OR_1/GND x0 x0_bar x1 x2 x2_bar x3 s2 x3_bar x1_bar VDD
+ CMOS_s2
XCMOS_s0_0 x3 x2_bar x2 x1_bar x1 x0 CMOS_s0_0/CMOS_OR_1/GND s0 x3_bar x0_bar VDD
+ CMOS_s0
.ends

.subckt CMOS_PRESENT80_R1 k0 k0_bar x0 x0_bar x1_bar x1 k1_bar k1 k2 k2_bar x2 x2_bar
+ x3_bar x3 k3_bar k3 s2 s1 s0 s3 CMOS_4in_XOR_0/CMOS_XOR_3/GND VDD
XCMOS_4in_XOR_0 VDD x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar x2 x2_bar k2 k2_bar x3
+ x3_bar k3 k3_bar CMOS_sbox_0/x1 CMOS_sbox_0/x0 CMOS_sbox_0/x2 CMOS_sbox_0/x3 CMOS_sbox_0/x0_bar
+ CMOS_sbox_0/x1_bar CMOS_sbox_0/x2_bar CMOS_sbox_0/x3_bar CMOS_4in_XOR_0/CMOS_XOR_3/GND
+ CMOS_4in_XOR
XCMOS_sbox_0 CMOS_sbox_0/x3 CMOS_sbox_0/x2 CMOS_sbox_0/x1_bar CMOS_sbox_0/x1 CMOS_sbox_0/x0_bar
+ CMOS_sbox_0/x0 CMOS_4in_XOR_0/CMOS_XOR_3/GND s0 s1 s2 s3 CMOS_sbox_0/x2_bar CMOS_sbox_0/x3_bar
+ VDD CMOS_sbox
.ends

.subckt CMOS_PRESENT80_SB8andSB11 CMOS_PRESENT80_R1_1/s3 CMOS_PRESENT80_R1_2/k2_bar
+ CMOS_PRESENT80_R1_1/s2 CMOS_PRESENT80_R1_2/x2_bar CMOS_PRESENT80_R1_1/s1 CMOS_PRESENT80_R1_0/k1_bar
+ CMOS_PRESENT80_R1_1/s0 CMOS_PRESENT80_R1_0/x1_bar CMOS_PRESENT80_R1_3/k3 CMOS_PRESENT80_R1_0/k3
+ CMOS_PRESENT80_R1_3/k2 CMOS_PRESENT80_R1_1/x3 CMOS_PRESENT80_R1_0/k2 CMOS_PRESENT80_R1_3/k3_bar
+ CMOS_PRESENT80_R1_3/k1 CMOS_PRESENT80_R1_3/x3_bar CMOS_PRESENT80_R1_1/x2 CMOS_PRESENT80_R1_0/k1
+ CMOS_PRESENT80_R1_3/k0 CMOS_PRESENT80_R1_1/x1 CMOS_PRESENT80_R1_0/k0 CMOS_PRESENT80_R1_1/k2_bar
+ CMOS_PRESENT80_R1_1/x2_bar CMOS_PRESENT80_R1_1/x0 CMOS_PRESENT80_R1_3/k0_bar CMOS_PRESENT80_R1_3/x0_bar
+ CMOS_PRESENT80_R1_3/s3 CMOS_PRESENT80_R1_2/k3_bar CMOS_PRESENT80_R1_0/s3 CMOS_PRESENT80_R1_2/x3_bar
+ CMOS_PRESENT80_R1_3/s2 CMOS_PRESENT80_R1_0/s2 CMOS_PRESENT80_R1_3/s1 CMOS_PRESENT80_R1_0/k2_bar
+ CMOS_PRESENT80_R1_0/x2_bar CMOS_PRESENT80_R1_0/s1 CMOS_PRESENT80_R1_3/s0 CMOS_PRESENT80_R1_2/k0_bar
+ CMOS_PRESENT80_R1_2/x0_bar CMOS_PRESENT80_R1_0/s0 CMOS_PRESENT80_R1_2/k3 CMOS_PRESENT80_R1_3/x3
+ CMOS_PRESENT80_R1_2/k2 CMOS_PRESENT80_R1_0/x3 CMOS_PRESENT80_R1_3/x2 CMOS_PRESENT80_R1_2/k1
+ CMOS_PRESENT80_R1_0/x2 CMOS_PRESENT80_R1_1/k3_bar CMOS_PRESENT80_R1_3/x1 CMOS_PRESENT80_R1_1/x3_bar
+ CMOS_PRESENT80_R1_2/k0 CMOS_PRESENT80_R1_0/x1 CMOS_PRESENT80_R1_3/k1_bar CMOS_PRESENT80_R1_3/x0
+ CMOS_PRESENT80_R1_3/x1_bar CMOS_PRESENT80_R1_0/x0 CMOS_PRESENT80_R1_1/k0_bar CMOS_PRESENT80_R1_1/x0_bar
+ CMOS_PRESENT80_R1_2/s3 CMOS_PRESENT80_R1_2/s2 CMOS_PRESENT80_R1_0/k3_bar CMOS_PRESENT80_R1_0/x3_bar
+ CMOS_PRESENT80_R1_2/s1 CMOS_PRESENT80_R1_2/k1_bar CMOS_PRESENT80_R1_2/x1_bar CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1_2/s0 CMOS_PRESENT80_R1_0/k0_bar CMOS_PRESENT80_R1_0/x0_bar CMOS_PRESENT80_R1_1/k3
+ CMOS_PRESENT80_R1_2/x3 CMOS_PRESENT80_R1_1/k2 CMOS_PRESENT80_R1_2/x2 CMOS_PRESENT80_R1_1/k1
+ CMOS_PRESENT80_R1_3/k2_bar CMOS_PRESENT80_R1_2/x1 CMOS_PRESENT80_R1_3/x2_bar CMOS_PRESENT80_R1_1/k0
+ CMOS_PRESENT80_R1_2/x0 CMOS_PRESENT80_R1_1/k1_bar CMOS_PRESENT80_R1_1/x1_bar CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND
XCMOS_PRESENT80_R1_0 CMOS_PRESENT80_R1_0/k0 CMOS_PRESENT80_R1_0/k0_bar CMOS_PRESENT80_R1_0/x0
+ CMOS_PRESENT80_R1_0/x0_bar CMOS_PRESENT80_R1_0/x1_bar CMOS_PRESENT80_R1_0/x1 CMOS_PRESENT80_R1_0/k1_bar
+ CMOS_PRESENT80_R1_0/k1 CMOS_PRESENT80_R1_0/k2 CMOS_PRESENT80_R1_0/k2_bar CMOS_PRESENT80_R1_0/x2
+ CMOS_PRESENT80_R1_0/x2_bar CMOS_PRESENT80_R1_0/x3_bar CMOS_PRESENT80_R1_0/x3 CMOS_PRESENT80_R1_0/k3_bar
+ CMOS_PRESENT80_R1_0/k3 CMOS_PRESENT80_R1_0/s2 CMOS_PRESENT80_R1_0/s1 CMOS_PRESENT80_R1_0/s0
+ CMOS_PRESENT80_R1_0/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_2 CMOS_PRESENT80_R1_2/k0 CMOS_PRESENT80_R1_2/k0_bar CMOS_PRESENT80_R1_2/x0
+ CMOS_PRESENT80_R1_2/x0_bar CMOS_PRESENT80_R1_2/x1_bar CMOS_PRESENT80_R1_2/x1 CMOS_PRESENT80_R1_2/k1_bar
+ CMOS_PRESENT80_R1_2/k1 CMOS_PRESENT80_R1_2/k2 CMOS_PRESENT80_R1_2/k2_bar CMOS_PRESENT80_R1_2/x2
+ CMOS_PRESENT80_R1_2/x2_bar CMOS_PRESENT80_R1_2/x3_bar CMOS_PRESENT80_R1_2/x3 CMOS_PRESENT80_R1_2/k3_bar
+ CMOS_PRESENT80_R1_2/k3 CMOS_PRESENT80_R1_2/s2 CMOS_PRESENT80_R1_2/s1 CMOS_PRESENT80_R1_2/s0
+ CMOS_PRESENT80_R1_2/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_1 CMOS_PRESENT80_R1_1/k0 CMOS_PRESENT80_R1_1/k0_bar CMOS_PRESENT80_R1_1/x0
+ CMOS_PRESENT80_R1_1/x0_bar CMOS_PRESENT80_R1_1/x1_bar CMOS_PRESENT80_R1_1/x1 CMOS_PRESENT80_R1_1/k1_bar
+ CMOS_PRESENT80_R1_1/k1 CMOS_PRESENT80_R1_1/k2 CMOS_PRESENT80_R1_1/k2_bar CMOS_PRESENT80_R1_1/x2
+ CMOS_PRESENT80_R1_1/x2_bar CMOS_PRESENT80_R1_1/x3_bar CMOS_PRESENT80_R1_1/x3 CMOS_PRESENT80_R1_1/k3_bar
+ CMOS_PRESENT80_R1_1/k3 CMOS_PRESENT80_R1_1/s2 CMOS_PRESENT80_R1_1/s1 CMOS_PRESENT80_R1_1/s0
+ CMOS_PRESENT80_R1_1/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_3 CMOS_PRESENT80_R1_3/k0 CMOS_PRESENT80_R1_3/k0_bar CMOS_PRESENT80_R1_3/x0
+ CMOS_PRESENT80_R1_3/x0_bar CMOS_PRESENT80_R1_3/x1_bar CMOS_PRESENT80_R1_3/x1 CMOS_PRESENT80_R1_3/k1_bar
+ CMOS_PRESENT80_R1_3/k1 CMOS_PRESENT80_R1_3/k2 CMOS_PRESENT80_R1_3/k2_bar CMOS_PRESENT80_R1_3/x2
+ CMOS_PRESENT80_R1_3/x2_bar CMOS_PRESENT80_R1_3/x3_bar CMOS_PRESENT80_R1_3/x3 CMOS_PRESENT80_R1_3/k3_bar
+ CMOS_PRESENT80_R1_3/k3 CMOS_PRESENT80_R1_3/s2 CMOS_PRESENT80_R1_3/s1 CMOS_PRESENT80_R1_3/s0
+ CMOS_PRESENT80_R1_3/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
.ends

.subckt CMOS_PRESENT80_SB12andSB15 CMOS_PRESENT80_R1_1/s3 CMOS_PRESENT80_R1_2/x2_bar
+ CMOS_PRESENT80_R1_1/s2 CMOS_PRESENT80_R1_2/k2_bar CMOS_PRESENT80_R1_1/s1 CMOS_PRESENT80_R1_0/k1_bar
+ CMOS_PRESENT80_R1_0/x1_bar CMOS_PRESENT80_R1_1/s0 CMOS_PRESENT80_R1_3/k3 CMOS_PRESENT80_R1_0/k3
+ CMOS_PRESENT80_R1_3/k2 CMOS_PRESENT80_R1_3/k3_bar CMOS_PRESENT80_R1_1/x3 CMOS_PRESENT80_R1_0/k2
+ CMOS_PRESENT80_R1_3/k1 CMOS_PRESENT80_R1_3/x3_bar CMOS_PRESENT80_R1_1/x2 CMOS_PRESENT80_R1_0/k1
+ CMOS_PRESENT80_R1_3/k0 CMOS_PRESENT80_R1_1/x1 CMOS_PRESENT80_R1_1/k2_bar CMOS_PRESENT80_R1_1/x2_bar
+ CMOS_PRESENT80_R1_0/k0 CMOS_PRESENT80_R1_1/x0 CMOS_PRESENT80_R1_3/k0_bar CMOS_PRESENT80_R1_3/x0_bar
+ CMOS_PRESENT80_R1_0/s3 CMOS_PRESENT80_R1_3/s3 CMOS_PRESENT80_R1_3/s2 CMOS_PRESENT80_R1_2/k3_bar
+ CMOS_PRESENT80_R1_2/x3_bar CMOS_PRESENT80_R1_3/s1 CMOS_PRESENT80_R1_0/s2 CMOS_PRESENT80_R1_2/k0_bar
+ CMOS_PRESENT80_R1_0/k2_bar CMOS_PRESENT80_R1_3/s0 CMOS_PRESENT80_R1_0/s1 CMOS_PRESENT80_R1_0/x2_bar
+ CMOS_PRESENT80_R1_2/k3 CMOS_PRESENT80_R1_0/s0 CMOS_PRESENT80_R1_2/x0_bar CMOS_PRESENT80_R1_2/k2
+ CMOS_PRESENT80_R1_3/x3 CMOS_PRESENT80_R1_2/k1 CMOS_PRESENT80_R1_0/x3 CMOS_PRESENT80_R1_0/x2
+ CMOS_PRESENT80_R1_3/x2 CMOS_PRESENT80_R1_1/k3_bar CMOS_PRESENT80_R1_3/x1 CMOS_PRESENT80_R1_2/k0
+ CMOS_PRESENT80_R1_0/x1 CMOS_PRESENT80_R1_1/x3_bar CMOS_PRESENT80_R1_3/x0 CMOS_PRESENT80_R1_3/x1_bar
+ CMOS_PRESENT80_R1_0/x0 CMOS_PRESENT80_R1_3/k1_bar CMOS_PRESENT80_R1_1/k0_bar CMOS_PRESENT80_R1_1/x0_bar
+ CMOS_PRESENT80_R1_2/s3 CMOS_PRESENT80_R1_2/s2 CMOS_PRESENT80_R1_0/k3_bar CMOS_PRESENT80_R1_0/x3_bar
+ CMOS_PRESENT80_R1_2/s1 CMOS_PRESENT80_R1_2/k1_bar CMOS_PRESENT80_R1_2/x1_bar CMOS_PRESENT80_R1_2/s0
+ CMOS_PRESENT80_R1_3/VDD CMOS_PRESENT80_R1_0/x0_bar CMOS_PRESENT80_R1_1/k3 CMOS_PRESENT80_R1_0/k0_bar
+ CMOS_PRESENT80_R1_2/x3 CMOS_PRESENT80_R1_1/k2 CMOS_PRESENT80_R1_3/k2_bar CMOS_PRESENT80_R1_2/x2
+ CMOS_PRESENT80_R1_1/k1 CMOS_PRESENT80_R1_2/x1 CMOS_PRESENT80_R1_1/k0 CMOS_PRESENT80_R1_2/x0
+ CMOS_PRESENT80_R1_3/x2_bar CMOS_PRESENT80_R1_1/k1_bar CMOS_PRESENT80_R1_1/x1_bar
+ CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND
XCMOS_PRESENT80_R1_0 CMOS_PRESENT80_R1_0/k0 CMOS_PRESENT80_R1_0/k0_bar CMOS_PRESENT80_R1_0/x0
+ CMOS_PRESENT80_R1_0/x0_bar CMOS_PRESENT80_R1_0/x1_bar CMOS_PRESENT80_R1_0/x1 CMOS_PRESENT80_R1_0/k1_bar
+ CMOS_PRESENT80_R1_0/k1 CMOS_PRESENT80_R1_0/k2 CMOS_PRESENT80_R1_0/k2_bar CMOS_PRESENT80_R1_0/x2
+ CMOS_PRESENT80_R1_0/x2_bar CMOS_PRESENT80_R1_0/x3_bar CMOS_PRESENT80_R1_0/x3 CMOS_PRESENT80_R1_0/k3_bar
+ CMOS_PRESENT80_R1_0/k3 CMOS_PRESENT80_R1_0/s2 CMOS_PRESENT80_R1_0/s1 CMOS_PRESENT80_R1_0/s0
+ CMOS_PRESENT80_R1_0/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_2 CMOS_PRESENT80_R1_2/k0 CMOS_PRESENT80_R1_2/k0_bar CMOS_PRESENT80_R1_2/x0
+ CMOS_PRESENT80_R1_2/x0_bar CMOS_PRESENT80_R1_2/x1_bar CMOS_PRESENT80_R1_2/x1 CMOS_PRESENT80_R1_2/k1_bar
+ CMOS_PRESENT80_R1_2/k1 CMOS_PRESENT80_R1_2/k2 CMOS_PRESENT80_R1_2/k2_bar CMOS_PRESENT80_R1_2/x2
+ CMOS_PRESENT80_R1_2/x2_bar CMOS_PRESENT80_R1_2/x3_bar CMOS_PRESENT80_R1_2/x3 CMOS_PRESENT80_R1_2/k3_bar
+ CMOS_PRESENT80_R1_2/k3 CMOS_PRESENT80_R1_2/s2 CMOS_PRESENT80_R1_2/s1 CMOS_PRESENT80_R1_2/s0
+ CMOS_PRESENT80_R1_2/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_1 CMOS_PRESENT80_R1_1/k0 CMOS_PRESENT80_R1_1/k0_bar CMOS_PRESENT80_R1_1/x0
+ CMOS_PRESENT80_R1_1/x0_bar CMOS_PRESENT80_R1_1/x1_bar CMOS_PRESENT80_R1_1/x1 CMOS_PRESENT80_R1_1/k1_bar
+ CMOS_PRESENT80_R1_1/k1 CMOS_PRESENT80_R1_1/k2 CMOS_PRESENT80_R1_1/k2_bar CMOS_PRESENT80_R1_1/x2
+ CMOS_PRESENT80_R1_1/x2_bar CMOS_PRESENT80_R1_1/x3_bar CMOS_PRESENT80_R1_1/x3 CMOS_PRESENT80_R1_1/k3_bar
+ CMOS_PRESENT80_R1_1/k3 CMOS_PRESENT80_R1_1/s2 CMOS_PRESENT80_R1_1/s1 CMOS_PRESENT80_R1_1/s0
+ CMOS_PRESENT80_R1_1/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_3 CMOS_PRESENT80_R1_3/k0 CMOS_PRESENT80_R1_3/k0_bar CMOS_PRESENT80_R1_3/x0
+ CMOS_PRESENT80_R1_3/x0_bar CMOS_PRESENT80_R1_3/x1_bar CMOS_PRESENT80_R1_3/x1 CMOS_PRESENT80_R1_3/k1_bar
+ CMOS_PRESENT80_R1_3/k1 CMOS_PRESENT80_R1_3/k2 CMOS_PRESENT80_R1_3/k2_bar CMOS_PRESENT80_R1_3/x2
+ CMOS_PRESENT80_R1_3/x2_bar CMOS_PRESENT80_R1_3/x3_bar CMOS_PRESENT80_R1_3/x3 CMOS_PRESENT80_R1_3/k3_bar
+ CMOS_PRESENT80_R1_3/k3 CMOS_PRESENT80_R1_3/s2 CMOS_PRESENT80_R1_3/s1 CMOS_PRESENT80_R1_3/s0
+ CMOS_PRESENT80_R1_3/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
.ends

.subckt CMOS_PRESENT80_SB4andSB7 CMOS_PRESENT80_R1_1/s3 CMOS_PRESENT80_R1_2/k2_bar
+ CMOS_PRESENT80_R1_1/s2 CMOS_PRESENT80_R1_2/x2_bar CMOS_PRESENT80_R1_1/s1 CMOS_PRESENT80_R1_0/k1_bar
+ CMOS_PRESENT80_R1_1/s0 CMOS_PRESENT80_R1_0/x1_bar CMOS_PRESENT80_R1_3/k3 CMOS_PRESENT80_R1_0/k3
+ CMOS_PRESENT80_R1_3/k2 CMOS_PRESENT80_R1_1/x3 CMOS_PRESENT80_R1_0/k2 CMOS_PRESENT80_R1_3/k3_bar
+ CMOS_PRESENT80_R1_3/k1 CMOS_PRESENT80_R1_3/x3_bar CMOS_PRESENT80_R1_1/x2 CMOS_PRESENT80_R1_0/k1
+ CMOS_PRESENT80_R1_3/k0 CMOS_PRESENT80_R1_1/x1 CMOS_PRESENT80_R1_0/k0 CMOS_PRESENT80_R1_1/k2_bar
+ CMOS_PRESENT80_R1_1/x2_bar CMOS_PRESENT80_R1_1/x0 CMOS_PRESENT80_R1_3/k0_bar CMOS_PRESENT80_R1_3/x0_bar
+ CMOS_PRESENT80_R1_3/s3 CMOS_PRESENT80_R1_2/k3_bar CMOS_PRESENT80_R1_0/s3 CMOS_PRESENT80_R1_2/x3_bar
+ CMOS_PRESENT80_R1_3/s2 CMOS_PRESENT80_R1_0/s2 CMOS_PRESENT80_R1_3/s1 CMOS_PRESENT80_R1_0/k2_bar
+ CMOS_PRESENT80_R1_0/s1 CMOS_PRESENT80_R1_0/x2_bar CMOS_PRESENT80_R1_3/s0 CMOS_PRESENT80_R1_2/k0_bar
+ CMOS_PRESENT80_R1_0/s0 CMOS_PRESENT80_R1_2/x0_bar CMOS_PRESENT80_R1_2/k3 CMOS_PRESENT80_R1_3/x3
+ CMOS_PRESENT80_R1_2/k2 CMOS_PRESENT80_R1_0/x3 CMOS_PRESENT80_R1_3/x2 CMOS_PRESENT80_R1_2/k1
+ CMOS_PRESENT80_R1_0/x2 CMOS_PRESENT80_R1_1/k3_bar CMOS_PRESENT80_R1_3/x1 CMOS_PRESENT80_R1_1/x3_bar
+ CMOS_PRESENT80_R1_2/k0 CMOS_PRESENT80_R1_0/x1 CMOS_PRESENT80_R1_3/k1_bar CMOS_PRESENT80_R1_3/x0
+ CMOS_PRESENT80_R1_3/x1_bar CMOS_PRESENT80_R1_0/x0 CMOS_PRESENT80_R1_1/k0_bar CMOS_PRESENT80_R1_1/x0_bar
+ CMOS_PRESENT80_R1_2/s3 CMOS_PRESENT80_R1_2/s2 CMOS_PRESENT80_R1_0/k3_bar CMOS_PRESENT80_R1_0/x3_bar
+ CMOS_PRESENT80_R1_2/s1 CMOS_PRESENT80_R1_2/k1_bar CMOS_PRESENT80_R1_2/x1_bar CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1_2/s0 CMOS_PRESENT80_R1_0/k0_bar CMOS_PRESENT80_R1_0/x0_bar CMOS_PRESENT80_R1_1/k3
+ CMOS_PRESENT80_R1_2/x3 CMOS_PRESENT80_R1_1/k2 CMOS_PRESENT80_R1_2/x2 CMOS_PRESENT80_R1_1/k1
+ CMOS_PRESENT80_R1_3/k2_bar CMOS_PRESENT80_R1_3/x2_bar CMOS_PRESENT80_R1_2/x1 CMOS_PRESENT80_R1_1/k0
+ CMOS_PRESENT80_R1_2/x0 CMOS_PRESENT80_R1_1/k1_bar CMOS_PRESENT80_R1_1/x1_bar CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND
XCMOS_PRESENT80_R1_0 CMOS_PRESENT80_R1_0/k0 CMOS_PRESENT80_R1_0/k0_bar CMOS_PRESENT80_R1_0/x0
+ CMOS_PRESENT80_R1_0/x0_bar CMOS_PRESENT80_R1_0/x1_bar CMOS_PRESENT80_R1_0/x1 CMOS_PRESENT80_R1_0/k1_bar
+ CMOS_PRESENT80_R1_0/k1 CMOS_PRESENT80_R1_0/k2 CMOS_PRESENT80_R1_0/k2_bar CMOS_PRESENT80_R1_0/x2
+ CMOS_PRESENT80_R1_0/x2_bar CMOS_PRESENT80_R1_0/x3_bar CMOS_PRESENT80_R1_0/x3 CMOS_PRESENT80_R1_0/k3_bar
+ CMOS_PRESENT80_R1_0/k3 CMOS_PRESENT80_R1_0/s2 CMOS_PRESENT80_R1_0/s1 CMOS_PRESENT80_R1_0/s0
+ CMOS_PRESENT80_R1_0/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_2 CMOS_PRESENT80_R1_2/k0 CMOS_PRESENT80_R1_2/k0_bar CMOS_PRESENT80_R1_2/x0
+ CMOS_PRESENT80_R1_2/x0_bar CMOS_PRESENT80_R1_2/x1_bar CMOS_PRESENT80_R1_2/x1 CMOS_PRESENT80_R1_2/k1_bar
+ CMOS_PRESENT80_R1_2/k1 CMOS_PRESENT80_R1_2/k2 CMOS_PRESENT80_R1_2/k2_bar CMOS_PRESENT80_R1_2/x2
+ CMOS_PRESENT80_R1_2/x2_bar CMOS_PRESENT80_R1_2/x3_bar CMOS_PRESENT80_R1_2/x3 CMOS_PRESENT80_R1_2/k3_bar
+ CMOS_PRESENT80_R1_2/k3 CMOS_PRESENT80_R1_2/s2 CMOS_PRESENT80_R1_2/s1 CMOS_PRESENT80_R1_2/s0
+ CMOS_PRESENT80_R1_2/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_1 CMOS_PRESENT80_R1_1/k0 CMOS_PRESENT80_R1_1/k0_bar CMOS_PRESENT80_R1_1/x0
+ CMOS_PRESENT80_R1_1/x0_bar CMOS_PRESENT80_R1_1/x1_bar CMOS_PRESENT80_R1_1/x1 CMOS_PRESENT80_R1_1/k1_bar
+ CMOS_PRESENT80_R1_1/k1 CMOS_PRESENT80_R1_1/k2 CMOS_PRESENT80_R1_1/k2_bar CMOS_PRESENT80_R1_1/x2
+ CMOS_PRESENT80_R1_1/x2_bar CMOS_PRESENT80_R1_1/x3_bar CMOS_PRESENT80_R1_1/x3 CMOS_PRESENT80_R1_1/k3_bar
+ CMOS_PRESENT80_R1_1/k3 CMOS_PRESENT80_R1_1/s2 CMOS_PRESENT80_R1_1/s1 CMOS_PRESENT80_R1_1/s0
+ CMOS_PRESENT80_R1_1/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_3 CMOS_PRESENT80_R1_3/k0 CMOS_PRESENT80_R1_3/k0_bar CMOS_PRESENT80_R1_3/x0
+ CMOS_PRESENT80_R1_3/x0_bar CMOS_PRESENT80_R1_3/x1_bar CMOS_PRESENT80_R1_3/x1 CMOS_PRESENT80_R1_3/k1_bar
+ CMOS_PRESENT80_R1_3/k1 CMOS_PRESENT80_R1_3/k2 CMOS_PRESENT80_R1_3/k2_bar CMOS_PRESENT80_R1_3/x2
+ CMOS_PRESENT80_R1_3/x2_bar CMOS_PRESENT80_R1_3/x3_bar CMOS_PRESENT80_R1_3/x3 CMOS_PRESENT80_R1_3/k3_bar
+ CMOS_PRESENT80_R1_3/k3 CMOS_PRESENT80_R1_3/s2 CMOS_PRESENT80_R1_3/s1 CMOS_PRESENT80_R1_3/s0
+ CMOS_PRESENT80_R1_3/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
.ends

.subckt CMOS_PRESENT80_SB0andSB3 CMOS_PRESENT80_R1_1/s3 CMOS_PRESENT80_R1_2/k2_bar
+ CMOS_PRESENT80_R1_1/s2 CMOS_PRESENT80_R1_2/x2_bar CMOS_PRESENT80_R1_1/s1 CMOS_PRESENT80_R1_0/k1_bar
+ CMOS_PRESENT80_R1_3/k3 CMOS_PRESENT80_R1_0/x1_bar CMOS_PRESENT80_R1_1/s0 CMOS_PRESENT80_R1_0/k3
+ CMOS_PRESENT80_R1_3/k2 CMOS_PRESENT80_R1_3/k3_bar CMOS_PRESENT80_R1_0/k2 CMOS_PRESENT80_R1_3/k1
+ CMOS_PRESENT80_R1_1/x3 CMOS_PRESENT80_R1_3/x3_bar CMOS_PRESENT80_R1_0/k1 CMOS_PRESENT80_R1_3/k0
+ CMOS_PRESENT80_R1_1/x2 CMOS_PRESENT80_R1_1/x1 CMOS_PRESENT80_R1_1/k2_bar CMOS_PRESENT80_R1_1/x2_bar
+ CMOS_PRESENT80_R1_0/k0 CMOS_PRESENT80_R1_1/x0 CMOS_PRESENT80_R1_3/k0_bar CMOS_PRESENT80_R1_3/x0_bar
+ CMOS_PRESENT80_R1_2/x3_bar CMOS_PRESENT80_R1_2/k3_bar CMOS_PRESENT80_R1_3/s3 CMOS_PRESENT80_R1_0/s3
+ CMOS_PRESENT80_R1_3/s2 CMOS_PRESENT80_R1_0/s2 CMOS_PRESENT80_R1_3/s1 CMOS_PRESENT80_R1_0/k2_bar
+ CMOS_PRESENT80_R1_2/k0_bar CMOS_PRESENT80_R1_3/s0 CMOS_PRESENT80_R1_0/x2_bar CMOS_PRESENT80_R1_2/x0_bar
+ CMOS_PRESENT80_R1_0/s0 CMOS_PRESENT80_R1_2/k3 CMOS_PRESENT80_R1_3/x3 CMOS_PRESENT80_R1_2/k2
+ CMOS_PRESENT80_R1_0/x3 CMOS_PRESENT80_R1_3/x2 CMOS_PRESENT80_R1_2/k1 CMOS_PRESENT80_R1_0/x2
+ CMOS_PRESENT80_R1_0/x1 CMOS_PRESENT80_R1_2/k0 CMOS_PRESENT80_R1_1/k3_bar CMOS_PRESENT80_R1_1/x3_bar
+ CMOS_PRESENT80_R1_3/x1 CMOS_PRESENT80_R1_0/x0 CMOS_PRESENT80_R1_3/k1_bar CMOS_PRESENT80_R1_3/x1_bar
+ CMOS_PRESENT80_R1_3/x0 CMOS_PRESENT80_R1_1/k0_bar CMOS_PRESENT80_R1_1/x0_bar CMOS_PRESENT80_R1_2/s3
+ CMOS_PRESENT80_R1_3/VDD CMOS_PRESENT80_R1_2/s2 CMOS_PRESENT80_R1_0/k3_bar CMOS_PRESENT80_R1_2/s1
+ CMOS_PRESENT80_R1_0/x3_bar CMOS_PRESENT80_R1_2/k1_bar CMOS_PRESENT80_R1_2/s0 CMOS_PRESENT80_R1_2/x1_bar
+ CMOS_PRESENT80_R1_1/k3 CMOS_PRESENT80_R1_0/x0_bar CMOS_PRESENT80_R1_0/k0_bar CMOS_PRESENT80_R1_2/x3
+ CMOS_PRESENT80_R1_1/k2 CMOS_PRESENT80_R1_2/x2 CMOS_PRESENT80_R1_1/k1 CMOS_PRESENT80_R1_3/k2_bar
+ CMOS_PRESENT80_R1_1/k0 CMOS_PRESENT80_R1_2/x1 CMOS_PRESENT80_R1_2/x0 CMOS_PRESENT80_R1_0/s1
+ CMOS_PRESENT80_R1_3/x2_bar CMOS_PRESENT80_R1_1/k1_bar CMOS_PRESENT80_R1_1/x1_bar
+ CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND
XCMOS_PRESENT80_R1_0 CMOS_PRESENT80_R1_0/k0 CMOS_PRESENT80_R1_0/k0_bar CMOS_PRESENT80_R1_0/x0
+ CMOS_PRESENT80_R1_0/x0_bar CMOS_PRESENT80_R1_0/x1_bar CMOS_PRESENT80_R1_0/x1 CMOS_PRESENT80_R1_0/k1_bar
+ CMOS_PRESENT80_R1_0/k1 CMOS_PRESENT80_R1_0/k2 CMOS_PRESENT80_R1_0/k2_bar CMOS_PRESENT80_R1_0/x2
+ CMOS_PRESENT80_R1_0/x2_bar CMOS_PRESENT80_R1_0/x3_bar CMOS_PRESENT80_R1_0/x3 CMOS_PRESENT80_R1_0/k3_bar
+ CMOS_PRESENT80_R1_0/k3 CMOS_PRESENT80_R1_0/s2 CMOS_PRESENT80_R1_0/s1 CMOS_PRESENT80_R1_0/s0
+ CMOS_PRESENT80_R1_0/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_2 CMOS_PRESENT80_R1_2/k0 CMOS_PRESENT80_R1_2/k0_bar CMOS_PRESENT80_R1_2/x0
+ CMOS_PRESENT80_R1_2/x0_bar CMOS_PRESENT80_R1_2/x1_bar CMOS_PRESENT80_R1_2/x1 CMOS_PRESENT80_R1_2/k1_bar
+ CMOS_PRESENT80_R1_2/k1 CMOS_PRESENT80_R1_2/k2 CMOS_PRESENT80_R1_2/k2_bar CMOS_PRESENT80_R1_2/x2
+ CMOS_PRESENT80_R1_2/x2_bar CMOS_PRESENT80_R1_2/x3_bar CMOS_PRESENT80_R1_2/x3 CMOS_PRESENT80_R1_2/k3_bar
+ CMOS_PRESENT80_R1_2/k3 CMOS_PRESENT80_R1_2/s2 CMOS_PRESENT80_R1_2/s1 CMOS_PRESENT80_R1_2/s0
+ CMOS_PRESENT80_R1_2/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_1 CMOS_PRESENT80_R1_1/k0 CMOS_PRESENT80_R1_1/k0_bar CMOS_PRESENT80_R1_1/x0
+ CMOS_PRESENT80_R1_1/x0_bar CMOS_PRESENT80_R1_1/x1_bar CMOS_PRESENT80_R1_1/x1 CMOS_PRESENT80_R1_1/k1_bar
+ CMOS_PRESENT80_R1_1/k1 CMOS_PRESENT80_R1_1/k2 CMOS_PRESENT80_R1_1/k2_bar CMOS_PRESENT80_R1_1/x2
+ CMOS_PRESENT80_R1_1/x2_bar CMOS_PRESENT80_R1_1/x3_bar CMOS_PRESENT80_R1_1/x3 CMOS_PRESENT80_R1_1/k3_bar
+ CMOS_PRESENT80_R1_1/k3 CMOS_PRESENT80_R1_1/s2 CMOS_PRESENT80_R1_1/s1 CMOS_PRESENT80_R1_1/s0
+ CMOS_PRESENT80_R1_1/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
XCMOS_PRESENT80_R1_3 CMOS_PRESENT80_R1_3/k0 CMOS_PRESENT80_R1_3/k0_bar CMOS_PRESENT80_R1_3/x0
+ CMOS_PRESENT80_R1_3/x0_bar CMOS_PRESENT80_R1_3/x1_bar CMOS_PRESENT80_R1_3/x1 CMOS_PRESENT80_R1_3/k1_bar
+ CMOS_PRESENT80_R1_3/k1 CMOS_PRESENT80_R1_3/k2 CMOS_PRESENT80_R1_3/k2_bar CMOS_PRESENT80_R1_3/x2
+ CMOS_PRESENT80_R1_3/x2_bar CMOS_PRESENT80_R1_3/x3_bar CMOS_PRESENT80_R1_3/x3 CMOS_PRESENT80_R1_3/k3_bar
+ CMOS_PRESENT80_R1_3/k3 CMOS_PRESENT80_R1_3/s2 CMOS_PRESENT80_R1_3/s1 CMOS_PRESENT80_R1_3/s0
+ CMOS_PRESENT80_R1_3/s3 CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_R1_3/VDD
+ CMOS_PRESENT80_R1
.ends

.subckt CMOS_PRESENT80_SB x0 x0_bar x1 x2 x3 x4 x5 x6 x7 x1_bar x2_bar x3_bar x4_bar
+ x5_bar x6_bar x7_bar k0 k2 k3 k4 k5 k6 k7 k0_bar k1_bar k2_bar k3_bar k4_bar k5_bar
+ k6_bar k7_bar k15_bar x15_bar x14_bar x13_bar x12_bar x11_bar x10_bar x9_bar x8_bar
+ x15 x8 x9 x10 x11 x12 x14 x13 k8 k9 k10 k11 k12 k13 k14 k15 k14_bar k13_bar k12_bar
+ k11_bar k10_bar k9_bar k8_bar x23_bar x22_bar x21_bar x20_bar x19_bar x18_bar x17_bar
+ x16_bar k23_bar k22_bar k21_bar k20_bar k19_bar x23 x22 x21 x20 x19 x18 x17 x16
+ k18_bar k17_bar k16_bar k17 k16 k23 k22 k21 k20 k19 k18 x29_bar x31_bar x31 x30
+ x29 x28 x27 x26 x25 x24 x28_bar x27_bar x26_bar x25_bar k24 k25 k31_bar k30_bar
+ k26 k27 k28 k29 k30 k31 k29_bar k28_bar k27_bar k26_bar k25_bar x24_bar x30_bar
+ k24_bar k1 x32 x33 x34 x35 x36 x37 x38 x39 k32 k33 k34 k35 k36 k37 k38 k39 x32_bar
+ x33_bar x34_bar x35_bar x36_bar x37_bar x38_bar x39_bar k32_bar k33_bar k34_bar
+ k35_bar k36_bar k37_bar k38_bar k39_bar x47_bar x46_bar x45_bar x44_bar x43_bar
+ x42_bar x41_bar x40_bar x40 x41 x42 x43 x44 x45 x46 x47 k47_bar k46_bar k45_bar
+ k44_bar k43_bar k42_bar k41_bar k40_bar k40 k41 k42 k43 k44 k45 k46 k47 x55_bar
+ x54_bar x53_bar x52_bar x51_bar x50_bar x49_bar x48_bar x55 x54 x53 x52 x51 x50
+ x49 x48 k50 k49 k48 k55_bar k54_bar k53_bar k52_bar k51_bar k50_bar k49_bar k48_bar
+ k55 k54 k53 k52 k51 x61 x60 k63_bar k62_bar k61_bar k60_bar k59_bar x56 x57 x58
+ x59 x63 k58_bar k57_bar k56_bar x63_bar x62_bar x61_bar x60_bar x56_bar x57_bar
+ x58_bar x59_bar k63 k62 k61 k60 k59 k58 k56 k57 x62 s0 s1 s2 s3 s4 s5 s6 s7 s8 s9
+ s10 s11 s12 s13 s14 s15 s16 s17 s18 s19 s20 s21 s22 s23 s24 s25 s26 s27 s28 s29
+ s30 s31 s32 s33 s34 s35 s36 s37 s38 s39 s40 s41 s42 s43 s44 s45 s46 s47 s48 s49
+ s50 s51 s52 s53 s54 s55 s56 s57 s58 s59 s60 s61 s62 s63
XCMOS_PRESENT80_SB8andSB11_0 s39 k42_bar s38 x42_bar s37 k45_bar s36 x45_bar k35 k47
+ k34 x39 k46 k35_bar k33 x35_bar x38 k45 k32 x37 k44 k38_bar x38_bar x36 k32_bar
+ x32_bar s35 k43_bar s47 x43_bar s34 s46 s33 k46_bar x46_bar s45 s32 k40_bar x40_bar
+ s44 k43 x35 k42 x47 x34 k41 x46 k39_bar x33 x39_bar k40 x45 k33_bar x32 x33_bar
+ x44 k36_bar x36_bar s43 s42 k47_bar x47_bar s41 k41_bar x41_bar CMOS_PRESENT80_SB4andSB7_0/CMOS_PRESENT80_R1_3/VDD
+ s40 k44_bar x44_bar k39 x43 k38 x42 k37 k34_bar x41 x34_bar k36 x40 k37_bar x37_bar
+ CMOS_PRESENT80_SB4andSB7_0/CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_SB8andSB11
XCMOS_PRESENT80_SB12andSB15_0 s55 x58_bar s54 k58_bar s53 k61_bar x61_bar s52 k51
+ k63 k50 k51_bar x55 k62 k49 x51_bar x54 k61 k48 x53 k54_bar x54_bar k60 x52 k48_bar
+ x48_bar s63 s51 s50 k59_bar x59_bar s49 s62 k56_bar k62_bar s48 s61 x62_bar k59
+ s60 x56_bar k58 x51 k57 x63 x62 x50 k55_bar x49 k56 x61 x55_bar x48 x49_bar x60
+ k49_bar k52_bar x52_bar s59 s58 k63_bar x63_bar s57 k57_bar x57_bar s56 CMOS_PRESENT80_SB4andSB7_0/CMOS_PRESENT80_R1_3/VDD
+ x60_bar k55 k60_bar x59 k54 k50_bar x58 k53 x57 k52 x56 x50_bar k53_bar x53_bar
+ CMOS_PRESENT80_SB4andSB7_0/CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_SB12andSB15
XCMOS_PRESENT80_SB4andSB7_0 s23 k26_bar s22 x26_bar s21 k29_bar s20 x29_bar k19 k31
+ k18 x23 k30 k19_bar k17 x19_bar x22 k29 k16 x21 k28 k22_bar x22_bar x20 k16_bar
+ x16_bar s19 k27_bar s31 x27_bar s18 s30 s17 k30_bar s29 x30_bar s16 k24_bar s28
+ x24_bar k27 x19 k26 x31 x18 k25 x30 k23_bar x17 x23_bar k24 x29 k17_bar x16 x17_bar
+ x28 k20_bar x20_bar s27 s26 k31_bar x31_bar s25 k25_bar x25_bar CMOS_PRESENT80_SB4andSB7_0/CMOS_PRESENT80_R1_3/VDD
+ s24 k28_bar x28_bar k23 x27 k22 x26 k21 k18_bar x18_bar x25 k20 x24 k21_bar x21_bar
+ CMOS_PRESENT80_SB4andSB7_0/CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND CMOS_PRESENT80_SB4andSB7
XCMOS_PRESENT80_SB0andSB3_0 s7 k10_bar s6 x10_bar s5 k13_bar k3 x13_bar s4 k15 k2
+ k3_bar k14 k1 x7 x3_bar k13 k0 x6 x5 k6_bar x6_bar k12 x4 k0_bar x0_bar x11_bar
+ k11_bar s3 s15 s2 s14 s1 k14_bar k8_bar s0 x14_bar x8_bar s12 k11 x3 k10 x15 x2
+ k9 x14 x13 k8 k7_bar x7_bar x1 x12 k1_bar x1_bar x0 k4_bar x4_bar s11 CMOS_PRESENT80_SB4andSB7_0/CMOS_PRESENT80_R1_3/VDD
+ s10 k15_bar s9 x15_bar k9_bar s8 x9_bar k7 x12_bar k12_bar x11 k6 x10 k5 k2_bar
+ k4 x9 x8 s13 x2_bar k5_bar x5_bar CMOS_PRESENT80_SB4andSB7_0/CMOS_PRESENT80_R1_3/CMOS_4in_XOR_0/CMOS_XOR_3/GND
+ CMOS_PRESENT80_SB0andSB3
.ends

