magic
tech sky130A
timestamp 1666730241
<< nwell >>
rect -940 795 -195 890
rect -770 600 -360 795
<< nmos >>
rect -850 270 -835 420
rect -685 270 -670 420
rect -610 270 -595 420
rect -535 270 -520 420
rect -460 270 -445 420
rect -295 270 -280 420
<< pmos >>
rect -685 625 -670 775
rect -610 625 -595 775
rect -535 625 -520 775
rect -460 625 -445 775
<< ndiff >>
rect -910 385 -850 420
rect -910 365 -890 385
rect -870 365 -850 385
rect -910 345 -850 365
rect -910 325 -890 345
rect -870 325 -850 345
rect -910 305 -850 325
rect -910 285 -890 305
rect -870 285 -850 305
rect -910 270 -850 285
rect -835 385 -775 420
rect -835 365 -815 385
rect -795 365 -775 385
rect -835 345 -775 365
rect -835 325 -815 345
rect -795 325 -775 345
rect -835 305 -775 325
rect -835 285 -815 305
rect -795 285 -775 305
rect -835 270 -775 285
rect -745 385 -685 420
rect -745 365 -725 385
rect -705 365 -685 385
rect -745 345 -685 365
rect -745 325 -725 345
rect -705 325 -685 345
rect -745 305 -685 325
rect -745 285 -725 305
rect -705 285 -685 305
rect -745 270 -685 285
rect -670 385 -610 420
rect -670 365 -650 385
rect -630 365 -610 385
rect -670 345 -610 365
rect -670 325 -650 345
rect -630 325 -610 345
rect -670 305 -610 325
rect -670 285 -650 305
rect -630 285 -610 305
rect -670 270 -610 285
rect -595 385 -535 420
rect -595 365 -575 385
rect -555 365 -535 385
rect -595 345 -535 365
rect -595 325 -575 345
rect -555 325 -535 345
rect -595 305 -535 325
rect -595 285 -575 305
rect -555 285 -535 305
rect -595 270 -535 285
rect -520 385 -460 420
rect -520 365 -500 385
rect -480 365 -460 385
rect -520 345 -460 365
rect -520 325 -500 345
rect -480 325 -460 345
rect -520 305 -460 325
rect -520 285 -500 305
rect -480 285 -460 305
rect -520 270 -460 285
rect -445 385 -385 420
rect -445 365 -425 385
rect -405 365 -385 385
rect -445 345 -385 365
rect -445 325 -425 345
rect -405 325 -385 345
rect -445 305 -385 325
rect -445 285 -425 305
rect -405 285 -385 305
rect -445 270 -385 285
rect -355 385 -295 420
rect -355 365 -335 385
rect -315 365 -295 385
rect -355 345 -295 365
rect -355 325 -335 345
rect -315 325 -295 345
rect -355 305 -295 325
rect -355 285 -335 305
rect -315 285 -295 305
rect -355 270 -295 285
rect -280 385 -220 420
rect -280 365 -260 385
rect -240 365 -220 385
rect -280 345 -220 365
rect -280 325 -260 345
rect -240 325 -220 345
rect -280 305 -220 325
rect -280 285 -260 305
rect -240 285 -220 305
rect -280 270 -220 285
<< pdiff >>
rect -745 740 -685 775
rect -745 720 -725 740
rect -705 720 -685 740
rect -745 700 -685 720
rect -745 680 -725 700
rect -705 680 -685 700
rect -745 660 -685 680
rect -745 640 -725 660
rect -705 640 -685 660
rect -745 625 -685 640
rect -670 740 -610 775
rect -670 720 -650 740
rect -630 720 -610 740
rect -670 700 -610 720
rect -670 680 -650 700
rect -630 680 -610 700
rect -670 660 -610 680
rect -670 640 -650 660
rect -630 640 -610 660
rect -670 625 -610 640
rect -595 740 -535 775
rect -595 720 -575 740
rect -555 720 -535 740
rect -595 700 -535 720
rect -595 680 -575 700
rect -555 680 -535 700
rect -595 660 -535 680
rect -595 640 -575 660
rect -555 640 -535 660
rect -595 625 -535 640
rect -520 740 -460 775
rect -520 720 -500 740
rect -480 720 -460 740
rect -520 700 -460 720
rect -520 680 -500 700
rect -480 680 -460 700
rect -520 660 -460 680
rect -520 640 -500 660
rect -480 640 -460 660
rect -520 625 -460 640
rect -445 740 -385 775
rect -445 720 -425 740
rect -405 720 -385 740
rect -445 700 -385 720
rect -445 680 -425 700
rect -405 680 -385 700
rect -445 660 -385 680
rect -445 640 -425 660
rect -405 640 -385 660
rect -445 625 -385 640
<< ndiffc >>
rect -890 365 -870 385
rect -890 325 -870 345
rect -890 285 -870 305
rect -815 365 -795 385
rect -815 325 -795 345
rect -815 285 -795 305
rect -725 365 -705 385
rect -725 325 -705 345
rect -725 285 -705 305
rect -650 365 -630 385
rect -650 325 -630 345
rect -650 285 -630 305
rect -575 365 -555 385
rect -575 325 -555 345
rect -575 285 -555 305
rect -500 365 -480 385
rect -500 325 -480 345
rect -500 285 -480 305
rect -425 365 -405 385
rect -425 325 -405 345
rect -425 285 -405 305
rect -335 365 -315 385
rect -335 325 -315 345
rect -335 285 -315 305
rect -260 365 -240 385
rect -260 325 -240 345
rect -260 285 -240 305
<< pdiffc >>
rect -725 720 -705 740
rect -725 680 -705 700
rect -725 640 -705 660
rect -650 720 -630 740
rect -650 680 -630 700
rect -650 640 -630 660
rect -575 720 -555 740
rect -575 680 -555 700
rect -575 640 -555 660
rect -500 720 -480 740
rect -500 680 -480 700
rect -500 640 -480 660
rect -425 720 -405 740
rect -425 680 -405 700
rect -425 640 -405 660
<< psubdiff >>
rect -910 185 -220 200
rect -910 165 -895 185
rect -875 165 -855 185
rect -835 165 -815 185
rect -795 165 -775 185
rect -755 165 -735 185
rect -715 165 -695 185
rect -675 165 -655 185
rect -635 165 -615 185
rect -595 165 -575 185
rect -555 165 -535 185
rect -515 165 -495 185
rect -475 165 -455 185
rect -435 165 -415 185
rect -395 165 -375 185
rect -355 165 -335 185
rect -315 165 -295 185
rect -275 165 -255 185
rect -235 165 -220 185
rect -910 150 -220 165
<< nsubdiff >>
rect -910 850 -220 865
rect -910 830 -895 850
rect -875 830 -855 850
rect -835 830 -815 850
rect -795 830 -775 850
rect -755 830 -735 850
rect -715 830 -695 850
rect -675 830 -655 850
rect -635 830 -615 850
rect -595 830 -575 850
rect -555 830 -535 850
rect -515 830 -495 850
rect -475 830 -455 850
rect -435 830 -415 850
rect -395 830 -375 850
rect -355 830 -335 850
rect -315 830 -295 850
rect -275 830 -255 850
rect -235 830 -220 850
rect -910 815 -220 830
<< psubdiffcont >>
rect -895 165 -875 185
rect -855 165 -835 185
rect -815 165 -795 185
rect -775 165 -755 185
rect -735 165 -715 185
rect -695 165 -675 185
rect -655 165 -635 185
rect -615 165 -595 185
rect -575 165 -555 185
rect -535 165 -515 185
rect -495 165 -475 185
rect -455 165 -435 185
rect -415 165 -395 185
rect -375 165 -355 185
rect -335 165 -315 185
rect -295 165 -275 185
rect -255 165 -235 185
<< nsubdiffcont >>
rect -895 830 -875 850
rect -855 830 -835 850
rect -815 830 -795 850
rect -775 830 -755 850
rect -735 830 -715 850
rect -695 830 -675 850
rect -655 830 -635 850
rect -615 830 -595 850
rect -575 830 -555 850
rect -535 830 -515 850
rect -495 830 -475 850
rect -455 830 -435 850
rect -415 830 -395 850
rect -375 830 -355 850
rect -335 830 -315 850
rect -295 830 -275 850
rect -255 830 -235 850
<< poly >>
rect -685 790 -595 805
rect -685 775 -670 790
rect -610 775 -595 790
rect -535 790 -445 805
rect -535 775 -520 790
rect -460 775 -445 790
rect -685 610 -670 625
rect -610 550 -595 625
rect -535 610 -520 625
rect -460 610 -445 625
rect -560 600 -520 610
rect -560 580 -550 600
rect -530 580 -520 600
rect -560 570 -520 580
rect -610 540 -570 550
rect -610 520 -600 540
rect -580 520 -570 540
rect -610 510 -570 520
rect -875 465 -835 475
rect -875 445 -865 465
rect -845 445 -835 465
rect -875 435 -835 445
rect -850 420 -835 435
rect -685 420 -670 435
rect -610 420 -595 510
rect -535 420 -520 570
rect -295 490 -255 500
rect -295 470 -285 490
rect -265 470 -255 490
rect -295 460 -255 470
rect -460 420 -445 435
rect -295 420 -280 460
rect -850 255 -835 270
rect -685 255 -670 270
rect -610 255 -595 270
rect -535 255 -520 270
rect -460 255 -445 270
rect -295 255 -280 270
rect -685 245 -645 255
rect -685 225 -675 245
rect -655 225 -645 245
rect -685 215 -645 225
rect -485 245 -445 255
rect -485 225 -475 245
rect -455 225 -445 245
rect -485 215 -445 225
<< polycont >>
rect -550 580 -530 600
rect -600 520 -580 540
rect -865 445 -845 465
rect -285 470 -265 490
rect -675 225 -655 245
rect -475 225 -455 245
<< locali >>
rect -910 850 -220 860
rect -910 830 -895 850
rect -875 830 -855 850
rect -835 830 -815 850
rect -795 830 -775 850
rect -755 830 -735 850
rect -715 830 -695 850
rect -675 830 -655 850
rect -635 830 -615 850
rect -595 830 -575 850
rect -555 830 -535 850
rect -515 830 -495 850
rect -475 830 -455 850
rect -435 830 -415 850
rect -395 830 -375 850
rect -355 830 -335 850
rect -315 830 -295 850
rect -275 830 -255 850
rect -235 830 -220 850
rect -910 820 -220 830
rect -735 740 -695 755
rect -735 720 -725 740
rect -705 720 -695 740
rect -735 700 -695 720
rect -735 680 -725 700
rect -705 680 -695 700
rect -735 660 -695 680
rect -735 640 -725 660
rect -705 640 -695 660
rect -735 630 -695 640
rect -660 740 -620 755
rect -660 720 -650 740
rect -630 720 -620 740
rect -660 700 -620 720
rect -660 680 -650 700
rect -630 680 -620 700
rect -660 660 -620 680
rect -660 640 -650 660
rect -630 640 -620 660
rect -660 625 -620 640
rect -585 740 -545 755
rect -585 720 -575 740
rect -555 720 -545 740
rect -585 700 -545 720
rect -585 680 -575 700
rect -555 680 -545 700
rect -585 660 -545 680
rect -585 640 -575 660
rect -555 640 -545 660
rect -585 630 -545 640
rect -510 740 -470 755
rect -510 720 -500 740
rect -480 720 -470 740
rect -510 700 -470 720
rect -510 680 -500 700
rect -480 680 -470 700
rect -510 660 -470 680
rect -510 640 -500 660
rect -480 640 -470 660
rect -510 625 -470 640
rect -435 740 -395 755
rect -435 720 -425 740
rect -405 720 -395 740
rect -435 700 -395 720
rect -435 680 -425 700
rect -405 680 -395 700
rect -435 660 -395 680
rect -435 640 -425 660
rect -405 640 -395 660
rect -435 630 -395 640
rect -650 600 -630 625
rect -560 600 -520 610
rect -910 580 -780 600
rect -910 530 -845 550
rect -865 475 -845 530
rect -800 500 -780 580
rect -650 580 -550 600
rect -530 580 -520 600
rect -810 490 -770 500
rect -875 465 -835 475
rect -875 445 -865 465
rect -845 445 -835 465
rect -810 470 -800 490
rect -780 470 -770 490
rect -810 460 -770 470
rect -875 435 -835 445
rect -650 440 -630 580
rect -560 570 -520 580
rect -610 540 -570 550
rect -500 540 -480 625
rect -360 600 -320 610
rect -360 580 -350 600
rect -330 580 -220 600
rect -360 570 -320 580
rect -610 520 -600 540
rect -580 520 -220 540
rect -610 510 -570 520
rect -500 440 -480 520
rect -360 490 -320 500
rect -295 490 -255 500
rect -360 470 -350 490
rect -330 470 -285 490
rect -265 470 -255 490
rect -360 460 -320 470
rect -295 460 -255 470
rect -815 420 -620 440
rect -815 400 -795 420
rect -900 385 -860 400
rect -900 365 -890 385
rect -870 365 -860 385
rect -900 345 -860 365
rect -900 325 -890 345
rect -870 325 -860 345
rect -900 305 -860 325
rect -900 285 -890 305
rect -870 285 -860 305
rect -900 275 -860 285
rect -825 385 -785 400
rect -825 365 -815 385
rect -795 365 -785 385
rect -825 345 -785 365
rect -825 325 -815 345
rect -795 325 -785 345
rect -825 305 -785 325
rect -825 285 -815 305
rect -795 285 -785 305
rect -825 275 -785 285
rect -735 385 -695 400
rect -735 365 -725 385
rect -705 365 -695 385
rect -735 345 -695 365
rect -735 325 -725 345
rect -705 325 -695 345
rect -735 305 -695 325
rect -735 285 -725 305
rect -705 285 -695 305
rect -735 275 -695 285
rect -660 385 -620 420
rect -510 420 -315 440
rect -660 365 -650 385
rect -630 365 -620 385
rect -660 345 -620 365
rect -660 325 -650 345
rect -630 325 -620 345
rect -660 305 -620 325
rect -660 285 -650 305
rect -630 285 -620 305
rect -660 275 -620 285
rect -585 385 -545 400
rect -585 365 -575 385
rect -555 365 -545 385
rect -585 345 -545 365
rect -585 325 -575 345
rect -555 325 -545 345
rect -585 305 -545 325
rect -585 285 -575 305
rect -555 285 -545 305
rect -585 275 -545 285
rect -510 385 -470 420
rect -335 400 -315 420
rect -510 365 -500 385
rect -480 365 -470 385
rect -510 345 -470 365
rect -510 325 -500 345
rect -480 325 -470 345
rect -510 305 -470 325
rect -510 285 -500 305
rect -480 285 -470 305
rect -510 275 -470 285
rect -435 385 -395 400
rect -435 365 -425 385
rect -405 365 -395 385
rect -435 345 -395 365
rect -435 325 -425 345
rect -405 325 -395 345
rect -435 305 -395 325
rect -435 285 -425 305
rect -405 285 -395 305
rect -435 275 -395 285
rect -345 385 -305 400
rect -345 365 -335 385
rect -315 365 -305 385
rect -345 345 -305 365
rect -345 325 -335 345
rect -315 325 -305 345
rect -345 305 -305 325
rect -345 285 -335 305
rect -315 285 -305 305
rect -345 275 -305 285
rect -270 385 -230 400
rect -270 365 -260 385
rect -240 365 -230 385
rect -270 345 -230 365
rect -270 325 -260 345
rect -240 325 -230 345
rect -270 305 -230 325
rect -270 285 -260 305
rect -240 285 -230 305
rect -270 275 -230 285
rect -685 245 -645 255
rect -485 245 -445 255
rect -910 225 -675 245
rect -655 225 -475 245
rect -455 225 -445 245
rect -685 215 -645 225
rect -485 215 -445 225
rect -910 185 -220 195
rect -910 165 -895 185
rect -875 165 -855 185
rect -835 165 -815 185
rect -795 165 -775 185
rect -755 165 -735 185
rect -715 165 -695 185
rect -675 165 -655 185
rect -635 165 -615 185
rect -595 165 -575 185
rect -555 165 -535 185
rect -515 165 -495 185
rect -475 165 -455 185
rect -435 165 -415 185
rect -395 165 -375 185
rect -355 165 -335 185
rect -315 165 -295 185
rect -275 165 -255 185
rect -235 165 -220 185
rect -910 155 -220 165
<< viali >>
rect -895 830 -875 850
rect -855 830 -835 850
rect -815 830 -795 850
rect -775 830 -755 850
rect -735 830 -715 850
rect -695 830 -675 850
rect -655 830 -635 850
rect -615 830 -595 850
rect -575 830 -555 850
rect -535 830 -515 850
rect -495 830 -475 850
rect -455 830 -435 850
rect -415 830 -395 850
rect -375 830 -355 850
rect -335 830 -315 850
rect -295 830 -275 850
rect -255 830 -235 850
rect -725 720 -705 740
rect -725 680 -705 700
rect -725 640 -705 660
rect -575 720 -555 740
rect -575 680 -555 700
rect -575 640 -555 660
rect -425 720 -405 740
rect -425 680 -405 700
rect -425 640 -405 660
rect -550 580 -530 600
rect -800 470 -780 490
rect -350 580 -330 600
rect -350 470 -330 490
rect -890 365 -870 385
rect -890 325 -870 345
rect -890 285 -870 305
rect -725 365 -705 385
rect -725 325 -705 345
rect -725 285 -705 305
rect -575 365 -555 385
rect -575 325 -555 345
rect -575 285 -555 305
rect -425 365 -405 385
rect -425 325 -405 345
rect -425 285 -405 305
rect -260 365 -240 385
rect -260 325 -240 345
rect -260 285 -240 305
rect -895 165 -875 185
rect -855 165 -835 185
rect -815 165 -795 185
rect -775 165 -755 185
rect -735 165 -715 185
rect -695 165 -675 185
rect -655 165 -635 185
rect -615 165 -595 185
rect -575 165 -555 185
rect -535 165 -515 185
rect -495 165 -475 185
rect -455 165 -435 185
rect -415 165 -395 185
rect -375 165 -355 185
rect -335 165 -315 185
rect -295 165 -275 185
rect -255 165 -235 185
<< metal1 >>
rect -910 850 -220 865
rect -910 830 -895 850
rect -875 830 -855 850
rect -835 830 -815 850
rect -795 830 -775 850
rect -755 830 -735 850
rect -715 830 -695 850
rect -675 830 -655 850
rect -635 830 -615 850
rect -595 830 -575 850
rect -555 830 -535 850
rect -515 830 -495 850
rect -475 830 -455 850
rect -435 830 -415 850
rect -395 830 -375 850
rect -355 830 -335 850
rect -315 830 -295 850
rect -275 830 -255 850
rect -235 830 -220 850
rect -910 815 -220 830
rect -900 385 -860 815
rect -735 740 -695 815
rect -735 720 -725 740
rect -705 720 -695 740
rect -735 700 -695 720
rect -735 680 -725 700
rect -705 680 -695 700
rect -735 660 -695 680
rect -735 640 -725 660
rect -705 640 -695 660
rect -735 630 -695 640
rect -585 740 -545 815
rect -585 720 -575 740
rect -555 720 -545 740
rect -585 700 -545 720
rect -585 680 -575 700
rect -555 680 -545 700
rect -585 660 -545 680
rect -585 640 -575 660
rect -555 640 -545 660
rect -585 630 -545 640
rect -435 740 -395 815
rect -435 720 -425 740
rect -405 720 -395 740
rect -435 700 -395 720
rect -435 680 -425 700
rect -405 680 -395 700
rect -435 660 -395 680
rect -435 640 -425 660
rect -405 640 -395 660
rect -435 630 -395 640
rect -560 600 -520 610
rect -360 600 -320 610
rect -560 580 -550 600
rect -530 580 -350 600
rect -330 580 -320 600
rect -560 570 -520 580
rect -360 570 -320 580
rect -810 490 -770 500
rect -360 490 -320 500
rect -810 470 -800 490
rect -780 470 -350 490
rect -330 470 -320 490
rect -810 460 -770 470
rect -360 460 -320 470
rect -900 365 -890 385
rect -870 365 -860 385
rect -900 345 -860 365
rect -900 325 -890 345
rect -870 325 -860 345
rect -900 305 -860 325
rect -900 285 -890 305
rect -870 285 -860 305
rect -900 275 -860 285
rect -735 385 -695 400
rect -735 365 -725 385
rect -705 365 -695 385
rect -735 345 -695 365
rect -735 325 -725 345
rect -705 325 -695 345
rect -735 305 -695 325
rect -735 285 -725 305
rect -705 285 -695 305
rect -735 275 -695 285
rect -585 385 -545 400
rect -585 365 -575 385
rect -555 365 -545 385
rect -585 345 -545 365
rect -585 325 -575 345
rect -555 325 -545 345
rect -585 305 -545 325
rect -585 285 -575 305
rect -555 285 -545 305
rect -585 275 -545 285
rect -435 385 -395 400
rect -435 365 -425 385
rect -405 365 -395 385
rect -435 345 -395 365
rect -435 325 -425 345
rect -405 325 -395 345
rect -435 305 -395 325
rect -435 285 -425 305
rect -405 285 -395 305
rect -435 275 -395 285
rect -270 385 -230 815
rect -270 365 -260 385
rect -240 365 -230 385
rect -270 345 -230 365
rect -270 325 -260 345
rect -240 325 -230 345
rect -270 305 -230 325
rect -270 285 -260 305
rect -240 285 -230 305
rect -270 275 -230 285
rect -725 200 -705 275
rect -575 200 -555 275
rect -425 200 -405 275
rect -910 185 -220 200
rect -910 165 -895 185
rect -875 165 -855 185
rect -835 165 -815 185
rect -795 165 -775 185
rect -755 165 -735 185
rect -715 165 -695 185
rect -675 165 -655 185
rect -635 165 -615 185
rect -595 165 -575 185
rect -555 165 -535 185
rect -515 165 -495 185
rect -475 165 -455 185
rect -435 165 -415 185
rect -395 165 -375 185
rect -355 165 -335 185
rect -315 165 -295 185
rect -275 165 -255 185
rect -235 165 -220 185
rect -910 150 -220 165
<< labels >>
rlabel locali -675 225 -655 245 7 Dis
port 5 w
rlabel metal1 -575 830 -555 850 7 CLK
port 7 w
rlabel locali -285 470 -265 490 7 A
port 1 w
rlabel locali -865 445 -845 465 7 A_bar
port 2 w
rlabel metal1 -575 165 -555 185 7 GND
port 6 w
rlabel viali -550 580 -530 600 7 OUT
port 3 w
rlabel locali -600 520 -580 540 7 OUT_bar
port 4 w
<< end >>
