magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -18949 1682 19176 23236
<< l67d20 >>
rect -1529 3192 -1489 3463
rect -1425 3985 -1392 4641
rect 1378 3985 1411 4641
rect 2144 3406 2184 3463
rect 2144 3192 2184 3406
rect 669 3377 799 3423
rect -144 3377 -14 3423
rect -781 3933 -764 4355
rect -781 4355 -645 4372
rect -159 4553 -142 4641
rect 2022 3933 2039 4364
rect 2022 4364 2128 4381
rect 2615 4553 2632 4641
rect -1086 3933 -1006 4067
rect 1707 3933 1787 4066
rect -971 4641 1199 4681
rect -971 4641 1199 4681
rect -971 8570 1199 8610
rect -1668 3152 516 3192
rect -1668 3152 516 3192
rect 1872 4641 4055 4681
rect 14833 4641 17016 4681
rect 12673 4641 14856 4681
rect 16993 4641 19176 4681
rect 15939 2382 18122 2422
rect 13779 2382 15962 2422
rect 11618 2382 13801 2422
rect 9458 2382 11641 2422
rect 7298 2382 9481 2422
rect 5138 2382 7321 2422
rect 2978 2382 5161 2422
rect 818 2382 3001 2422
rect 10513 4641 12696 4681
rect 10513 4641 12696 4681
rect 8353 4641 10536 4681
rect 6192 4641 8375 4681
rect 4032 4641 6215 4681
rect 1872 4641 4055 4681
rect 14833 4641 17016 4681
rect 12673 4641 14856 4681
rect 16993 4641 19176 4681
rect 8353 4641 10536 4681
rect 10513 8570 12696 8610
rect 8353 8570 10536 8610
rect 6192 8570 8375 8610
rect 4032 8570 6215 8610
rect 1872 8570 4055 8610
rect 14833 8570 17016 8610
rect 12673 8570 14856 8610
rect 16993 8570 19176 8610
rect 1697 4066 1797 4166
rect 13454 3152 15637 3192
rect 11294 3152 13477 3192
rect 9133 3152 11316 3192
rect 6973 3152 9156 3192
rect 4813 3152 6996 3192
rect 2653 3152 4836 3192
rect 493 3152 2676 3192
rect 6192 4641 8375 4681
rect 13454 3152 15637 3192
rect 11294 3152 13477 3192
rect 9133 3152 11316 3192
rect 6973 3152 9156 3192
rect 4813 3152 6996 3192
rect 2653 3152 4836 3192
rect 493 3152 2676 3192
rect 4032 4641 6215 4681
rect 13454 3152 15637 3192
rect 11294 3152 13477 3192
rect 9133 3152 11316 3192
rect 13454 3152 15637 3192
rect 11294 3152 13477 3192
rect 9133 3152 11316 3192
rect 15614 3152 17797 3192
rect 15614 3152 17797 3192
rect 15614 3152 17797 3192
rect 669 3247 799 3377
rect 15614 3152 17797 3192
rect 671 2816 801 2946
rect -2355 2382 -172 2422
rect -18949 4641 -16766 4681
rect -3828 4641 -1645 4681
rect -5988 4641 -3805 4681
rect -1094 4066 -994 4166
rect -3828 3152 -1645 3192
rect -5988 3152 -3805 3192
rect -8148 3152 -5965 3192
rect -10308 3152 -8125 3192
rect -12468 3152 -10285 3192
rect -14629 3152 -12446 3192
rect -16789 3152 -14606 3192
rect -18949 3152 -16766 3192
rect -3828 3152 -1645 3192
rect -5988 3152 -3805 3192
rect -8148 3152 -5965 3192
rect -10308 3152 -8125 3192
rect -12468 3152 -10285 3192
rect -14629 3152 -12446 3192
rect -16789 3152 -14606 3192
rect -18949 3152 -16766 3192
rect -8149 4641 -5966 4681
rect -10309 4641 -8126 4681
rect -12469 4641 -10286 4681
rect -14629 4641 -12446 4681
rect -16789 4641 -14606 4681
rect -18949 4641 -16766 4681
rect -4515 2382 -2332 2422
rect -6675 2382 -4492 2422
rect -8835 2382 -6652 2422
rect -10995 2382 -8812 2422
rect -13156 2382 -10973 2422
rect -15316 2382 -13133 2422
rect -17476 2382 -15293 2422
rect -3828 4641 -1645 4681
rect -5988 4641 -3805 4681
rect -3828 8570 -1645 8610
rect -5988 8570 -3805 8610
rect -8149 8570 -5966 8610
rect -10309 8570 -8126 8610
rect -12469 8570 -10286 8610
rect -14629 8570 -12446 8610
rect -16789 8570 -14606 8610
rect -18949 8570 -16766 8610
rect -8149 4641 -5966 4681
rect -144 3247 -14 3377
rect -10309 4641 -8126 4681
rect -12469 4641 -10286 4681
rect -14629 4641 -12446 4681
rect -143 2816 -13 2946
rect -16789 4641 -14606 4681
rect -1930 3294 -1800 3424
rect -1930 3913 -1800 4043
<< l66d20 >>
rect -669 3392 -654 3412
rect -669 3374 -654 3392
rect 634 3928 649 3969
rect 1384 3943 1411 3955
rect -1419 3943 -1392 3955
rect -1425 3952 -1392 3985
rect 1378 3952 1411 3985
rect -678 3344 -645 3377
rect 625 3959 658 3992
<< l66d44 >>
rect 18616 8582 18633 8599
rect 18616 8582 18633 8599
rect 18976 8582 18993 8599
rect 18936 8582 18953 8599
rect 18896 8582 18913 8599
rect 18856 8582 18873 8599
rect 18816 8582 18833 8599
rect 18776 8582 18793 8599
rect 18736 8582 18753 8599
rect 19136 8582 19153 8599
rect 19096 8582 19113 8599
rect 19056 8582 19073 8599
rect 19016 8582 19033 8599
rect 18976 8582 18993 8599
rect 18936 8582 18953 8599
rect 18896 8582 18913 8599
rect 18856 8582 18873 8599
rect 18816 8582 18833 8599
rect 18776 8582 18793 8599
rect 18736 8582 18753 8599
rect 19136 8582 19153 8599
rect 19096 8582 19113 8599
rect 19056 8582 19073 8599
rect 19016 8582 19033 8599
rect 18696 8582 18713 8599
rect 18656 8582 18673 8599
rect 18696 8582 18713 8599
rect 18656 8582 18673 8599
rect 18296 8582 18313 8599
rect 18336 8582 18353 8599
rect 18576 8582 18593 8599
rect 18536 8582 18553 8599
rect 18256 8582 18273 8599
rect 18496 8582 18513 8599
rect 18216 8582 18233 8599
rect 18176 8582 18193 8599
rect 18136 8582 18153 8599
rect 18096 8582 18113 8599
rect 18456 8582 18473 8599
rect 18416 8582 18433 8599
rect 18376 8582 18393 8599
rect 18576 8582 18593 8599
rect 18536 8582 18553 8599
rect 18496 8582 18513 8599
rect 18456 8582 18473 8599
rect 18416 8582 18433 8599
rect 18376 8582 18393 8599
rect 18336 8582 18353 8599
rect 18296 8582 18313 8599
rect 18256 8582 18273 8599
rect 18216 8582 18233 8599
rect 18176 8582 18193 8599
rect 18136 8582 18153 8599
rect 18096 8582 18113 8599
rect 17976 8582 17993 8599
rect 18016 8582 18033 8599
rect 18056 8582 18073 8599
rect 18016 8582 18033 8599
rect 18056 8582 18073 8599
rect 17976 8582 17993 8599
rect 16936 8582 16953 8599
rect 16896 8582 16913 8599
rect 16856 8582 16873 8599
rect 16976 8582 16993 8599
rect 16816 8582 16833 8599
rect 16936 8582 16953 8599
rect 17176 8582 17193 8599
rect 17176 8582 17193 8599
rect 17056 8582 17073 8599
rect 17136 8582 17153 8599
rect 17216 8582 17233 8599
rect 17096 8582 17113 8599
rect 17016 8582 17033 8599
rect 17056 8582 17073 8599
rect 17936 8582 17953 8599
rect 17416 8582 17433 8599
rect 16896 8582 16913 8599
rect 17376 8582 17393 8599
rect 17656 8582 17673 8599
rect 17336 8582 17353 8599
rect 17896 8582 17913 8599
rect 17296 8582 17313 8599
rect 17856 8582 17873 8599
rect 17136 8582 17153 8599
rect 17616 8582 17633 8599
rect 17856 8582 17873 8599
rect 16776 8582 16793 8599
rect 17576 8582 17593 8599
rect 17816 8582 17833 8599
rect 17816 8582 17833 8599
rect 17776 8582 17793 8599
rect 17096 8582 17113 8599
rect 17736 8582 17753 8599
rect 16856 8582 16873 8599
rect 17696 8582 17713 8599
rect 17656 8582 17673 8599
rect 17936 8582 17953 8599
rect 17616 8582 17633 8599
rect 17576 8582 17593 8599
rect 17216 8582 17233 8599
rect 17256 8582 17273 8599
rect 17256 8582 17273 8599
rect 17016 8582 17033 8599
rect 17776 8582 17793 8599
rect 17536 8582 17553 8599
rect 17496 8582 17513 8599
rect 17536 8582 17553 8599
rect 17456 8582 17473 8599
rect 17416 8582 17433 8599
rect 17496 8582 17513 8599
rect 17376 8582 17393 8599
rect 17336 8582 17353 8599
rect 17456 8582 17473 8599
rect 17296 8582 17313 8599
rect 16816 8582 16833 8599
rect 16776 8582 16793 8599
rect 17736 8582 17753 8599
rect 16976 8582 16993 8599
rect 17896 8582 17913 8599
rect 17696 8582 17713 8599
rect 15576 8582 15593 8599
rect 15576 8582 15593 8599
rect 16696 8582 16713 8599
rect 16256 8582 16273 8599
rect 16656 8582 16673 8599
rect 16616 8582 16633 8599
rect 16616 8582 16633 8599
rect 16216 8582 16233 8599
rect 16576 8582 16593 8599
rect 16456 8582 16473 8599
rect 16536 8582 16553 8599
rect 16656 8582 16673 8599
rect 16496 8582 16513 8599
rect 16176 8582 16193 8599
rect 16456 8582 16473 8599
rect 16696 8582 16713 8599
rect 16416 8582 16433 8599
rect 16136 8582 16153 8599
rect 15696 8582 15713 8599
rect 15816 8582 15833 8599
rect 15896 8582 15913 8599
rect 15776 8582 15793 8599
rect 15736 8582 15753 8599
rect 15656 8582 15673 8599
rect 15696 8582 15713 8599
rect 15816 8582 15833 8599
rect 15656 8582 15673 8599
rect 15856 8582 15873 8599
rect 15856 8582 15873 8599
rect 15736 8582 15753 8599
rect 15896 8582 15913 8599
rect 15776 8582 15793 8599
rect 16016 8582 16033 8599
rect 15976 8582 15993 8599
rect 15616 8582 15633 8599
rect 15936 8582 15953 8599
rect 16056 8582 16073 8599
rect 16016 8582 16033 8599
rect 15976 8582 15993 8599
rect 15936 8582 15953 8599
rect 16056 8582 16073 8599
rect 15616 8582 15633 8599
rect 16096 8582 16113 8599
rect 16096 8582 16113 8599
rect 16376 8582 16393 8599
rect 16336 8582 16353 8599
rect 16256 8582 16273 8599
rect 16536 8582 16553 8599
rect 16216 8582 16233 8599
rect 16336 8582 16353 8599
rect 16296 8582 16313 8599
rect 16176 8582 16193 8599
rect 16416 8582 16433 8599
rect 16576 8582 16593 8599
rect 16136 8582 16153 8599
rect 16296 8582 16313 8599
rect 16736 8582 16753 8599
rect 16496 8582 16513 8599
rect 16376 8582 16393 8599
rect 16736 8582 16753 8599
rect 15216 8582 15233 8599
rect 14416 8582 14433 8599
rect 15496 8582 15513 8599
rect 15056 8582 15073 8599
rect 14856 8582 14873 8599
rect 14816 8582 14833 8599
rect 15496 8582 15513 8599
rect 15176 8582 15193 8599
rect 15536 8582 15553 8599
rect 14776 8582 14793 8599
rect 15456 8582 15473 8599
rect 15016 8582 15033 8599
rect 15016 8582 15033 8599
rect 14736 8582 14753 8599
rect 15136 8582 15153 8599
rect 15336 8582 15353 8599
rect 15176 8582 15193 8599
rect 14696 8582 14713 8599
rect 15416 8582 15433 8599
rect 15256 8582 15273 8599
rect 15416 8582 15433 8599
rect 14656 8582 14673 8599
rect 14976 8582 14993 8599
rect 15456 8582 15473 8599
rect 15136 8582 15153 8599
rect 14616 8582 14633 8599
rect 14976 8582 14993 8599
rect 14656 8582 14673 8599
rect 15376 8582 15393 8599
rect 14576 8582 14593 8599
rect 15096 8582 15113 8599
rect 15536 8582 15553 8599
rect 14896 8582 14913 8599
rect 14536 8582 14553 8599
rect 14896 8582 14913 8599
rect 15336 8582 15353 8599
rect 14496 8582 14513 8599
rect 14616 8582 14633 8599
rect 14456 8582 14473 8599
rect 14936 8582 14953 8599
rect 14416 8582 14433 8599
rect 15056 8582 15073 8599
rect 14816 8582 14833 8599
rect 14576 8582 14593 8599
rect 14776 8582 14793 8599
rect 15376 8582 15393 8599
rect 14736 8582 14753 8599
rect 14856 8582 14873 8599
rect 14696 8582 14713 8599
rect 14536 8582 14553 8599
rect 15296 8582 15313 8599
rect 15216 8582 15233 8599
rect 15256 8582 15273 8599
rect 14496 8582 14513 8599
rect 15096 8582 15113 8599
rect 15296 8582 15313 8599
rect 14936 8582 14953 8599
rect 14456 8582 14473 8599
rect 13496 8582 13513 8599
rect 14336 8582 14353 8599
rect 13496 8582 13513 8599
rect 13976 8582 13993 8599
rect 13456 8582 13473 8599
rect 14016 8582 14033 8599
rect 13416 8582 13433 8599
rect 14256 8582 14273 8599
rect 13736 8582 13753 8599
rect 14216 8582 14233 8599
rect 13376 8582 13393 8599
rect 13936 8582 13953 8599
rect 13336 8582 13353 8599
rect 14176 8582 14193 8599
rect 13616 8582 13633 8599
rect 13896 8582 13913 8599
rect 13296 8582 13313 8599
rect 13856 8582 13873 8599
rect 13256 8582 13273 8599
rect 13816 8582 13833 8599
rect 13456 8582 13473 8599
rect 13776 8582 13793 8599
rect 13216 8582 13233 8599
rect 14136 8582 14153 8599
rect 13216 8582 13233 8599
rect 13696 8582 13713 8599
rect 14096 8582 14113 8599
rect 13736 8582 13753 8599
rect 13416 8582 13433 8599
rect 14056 8582 14073 8599
rect 13656 8582 13673 8599
rect 13576 8582 13593 8599
rect 14256 8582 14273 8599
rect 13376 8582 13393 8599
rect 14216 8582 14233 8599
rect 14176 8582 14193 8599
rect 14136 8582 14153 8599
rect 14096 8582 14113 8599
rect 14056 8582 14073 8599
rect 14016 8582 14033 8599
rect 13976 8582 13993 8599
rect 13936 8582 13953 8599
rect 13896 8582 13913 8599
rect 13856 8582 13873 8599
rect 13816 8582 13833 8599
rect 13776 8582 13793 8599
rect 13656 8582 13673 8599
rect 13336 8582 13353 8599
rect 13576 8582 13593 8599
rect 13616 8582 13633 8599
rect 13536 8582 13553 8599
rect 14296 8582 14313 8599
rect 13296 8582 13313 8599
rect 14296 8582 14313 8599
rect 13536 8582 13553 8599
rect 14376 8582 14393 8599
rect 13696 8582 13713 8599
rect 14336 8582 14353 8599
rect 13256 8582 13273 8599
rect 14376 8582 14393 8599
rect 13176 8582 13193 8599
rect 12096 8582 12113 8599
rect 12456 8582 12473 8599
rect 12496 8582 12513 8599
rect 12256 8582 12273 8599
rect 12296 8582 12313 8599
rect 13056 8582 13073 8599
rect 12536 8582 12553 8599
rect 12176 8582 12193 8599
rect 12056 8582 12073 8599
rect 12576 8582 12593 8599
rect 12096 8582 12113 8599
rect 13016 8582 13033 8599
rect 13056 8582 13073 8599
rect 13096 8582 13113 8599
rect 12536 8582 12553 8599
rect 12256 8582 12273 8599
rect 13016 8582 13033 8599
rect 13136 8582 13153 8599
rect 12496 8582 12513 8599
rect 12976 8582 12993 8599
rect 12696 8582 12713 8599
rect 12136 8582 12153 8599
rect 12856 8582 12873 8599
rect 12976 8582 12993 8599
rect 12816 8582 12833 8599
rect 12056 8582 12073 8599
rect 13136 8582 13153 8599
rect 12216 8582 12233 8599
rect 12856 8582 12873 8599
rect 12216 8582 12233 8599
rect 12736 8582 12753 8599
rect 12176 8582 12193 8599
rect 12016 8582 12033 8599
rect 12656 8582 12673 8599
rect 12816 8582 12833 8599
rect 12416 8582 12433 8599
rect 12336 8582 12353 8599
rect 13096 8582 13113 8599
rect 12896 8582 12913 8599
rect 12376 8582 12393 8599
rect 12776 8582 12793 8599
rect 12936 8582 12953 8599
rect 12776 8582 12793 8599
rect 12656 8582 12673 8599
rect 12456 8582 12473 8599
rect 12336 8582 12353 8599
rect 12136 8582 12153 8599
rect 13176 8582 13193 8599
rect 12376 8582 12393 8599
rect 12616 8582 12633 8599
rect 12696 8582 12713 8599
rect 12616 8582 12633 8599
rect 12416 8582 12433 8599
rect 12016 8582 12033 8599
rect 12736 8582 12753 8599
rect 12576 8582 12593 8599
rect 12896 8582 12913 8599
rect 12296 8582 12313 8599
rect 12936 8582 12953 8599
rect 10816 8582 10833 8599
rect 10816 8582 10833 8599
rect 11296 8582 11313 8599
rect 11136 8582 11153 8599
rect 11616 8582 11633 8599
rect 11496 8582 11513 8599
rect 11856 8582 11873 8599
rect 11456 8582 11473 8599
rect 10896 8582 10913 8599
rect 11376 8582 11393 8599
rect 11136 8582 11153 8599
rect 11776 8582 11793 8599
rect 10976 8582 10993 8599
rect 11576 8582 11593 8599
rect 11816 8582 11833 8599
rect 11976 8582 11993 8599
rect 11816 8582 11833 8599
rect 11736 8582 11753 8599
rect 11856 8582 11873 8599
rect 10896 8582 10913 8599
rect 11656 8582 11673 8599
rect 10936 8582 10953 8599
rect 10856 8582 10873 8599
rect 11176 8582 11193 8599
rect 11336 8582 11353 8599
rect 11376 8582 11393 8599
rect 10936 8582 10953 8599
rect 11296 8582 11313 8599
rect 11056 8582 11073 8599
rect 11456 8582 11473 8599
rect 11216 8582 11233 8599
rect 11016 8582 11033 8599
rect 11256 8582 11273 8599
rect 11936 8582 11953 8599
rect 10856 8582 10873 8599
rect 11896 8582 11913 8599
rect 11416 8582 11433 8599
rect 11336 8582 11353 8599
rect 11096 8582 11113 8599
rect 11576 8582 11593 8599
rect 11016 8582 11033 8599
rect 11216 8582 11233 8599
rect 11976 8582 11993 8599
rect 11616 8582 11633 8599
rect 11056 8582 11073 8599
rect 11096 8582 11113 8599
rect 11776 8582 11793 8599
rect 11656 8582 11673 8599
rect 10976 8582 10993 8599
rect 11256 8582 11273 8599
rect 11536 8582 11553 8599
rect 11696 8582 11713 8599
rect 11936 8582 11953 8599
rect 11536 8582 11553 8599
rect 11696 8582 11713 8599
rect 11176 8582 11193 8599
rect 11736 8582 11753 8599
rect 11896 8582 11913 8599
rect 11496 8582 11513 8599
rect 11416 8582 11433 8599
rect 9696 8582 9713 8599
rect 9856 8582 9873 8599
rect 10576 8582 10593 8599
rect 9696 8582 9713 8599
rect 9856 8582 9873 8599
rect 10496 8582 10513 8599
rect 10256 8582 10273 8599
rect 10656 8582 10673 8599
rect 10216 8582 10233 8599
rect 9656 8582 9673 8599
rect 9896 8582 9913 8599
rect 10616 8582 10633 8599
rect 10256 8582 10273 8599
rect 10456 8582 10473 8599
rect 10056 8582 10073 8599
rect 10416 8582 10433 8599
rect 10456 8582 10473 8599
rect 10096 8582 10113 8599
rect 10296 8582 10313 8599
rect 10416 8582 10433 8599
rect 9816 8582 9833 8599
rect 10376 8582 10393 8599
rect 9656 8582 9673 8599
rect 10536 8582 10553 8599
rect 10136 8582 10153 8599
rect 10776 8582 10793 8599
rect 10336 8582 10353 8599
rect 10376 8582 10393 8599
rect 10696 8582 10713 8599
rect 9936 8582 9953 8599
rect 9896 8582 9913 8599
rect 10336 8582 10353 8599
rect 10176 8582 10193 8599
rect 10656 8582 10673 8599
rect 9776 8582 9793 8599
rect 9976 8582 9993 8599
rect 10216 8582 10233 8599
rect 10776 8582 10793 8599
rect 10576 8582 10593 8599
rect 10296 8582 10313 8599
rect 10736 8582 10753 8599
rect 10136 8582 10153 8599
rect 10736 8582 10753 8599
rect 10616 8582 10633 8599
rect 10096 8582 10113 8599
rect 9816 8582 9833 8599
rect 10016 8582 10033 8599
rect 10536 8582 10553 8599
rect 9736 8582 9753 8599
rect 10056 8582 10073 8599
rect 9976 8582 9993 8599
rect 10496 8582 10513 8599
rect 9736 8582 9753 8599
rect 10176 8582 10193 8599
rect 9936 8582 9953 8599
rect 10016 8582 10033 8599
rect 10696 8582 10713 8599
rect 9776 8582 9793 8599
rect 9336 8582 9353 8599
rect 9496 8582 9513 8599
rect 9256 8582 9273 8599
rect 9456 8582 9473 8599
rect 8616 8582 8633 8599
rect 8536 8582 8553 8599
rect 9056 8582 9073 8599
rect 8536 8582 8553 8599
rect 9296 8582 9313 8599
rect 8496 8582 8513 8599
rect 8576 8582 8593 8599
rect 8776 8582 8793 8599
rect 8456 8582 8473 8599
rect 8616 8582 8633 8599
rect 9336 8582 9353 8599
rect 8736 8582 8753 8599
rect 9016 8582 9033 8599
rect 9136 8582 9153 8599
rect 8696 8582 8713 8599
rect 9256 8582 9273 8599
rect 8656 8582 8673 8599
rect 8896 8582 8913 8599
rect 9216 8582 9233 8599
rect 8976 8582 8993 8599
rect 9216 8582 9233 8599
rect 8856 8582 8873 8599
rect 8576 8582 8593 8599
rect 9376 8582 9393 8599
rect 8936 8582 8953 8599
rect 8896 8582 8913 8599
rect 9176 8582 9193 8599
rect 9176 8582 9193 8599
rect 8816 8582 8833 8599
rect 9136 8582 9153 8599
rect 9096 8582 9113 8599
rect 8776 8582 8793 8599
rect 8496 8582 8513 8599
rect 8856 8582 8873 8599
rect 9416 8582 9433 8599
rect 9056 8582 9073 8599
rect 8736 8582 8753 8599
rect 9016 8582 9033 8599
rect 8696 8582 8713 8599
rect 9296 8582 9313 8599
rect 8976 8582 8993 8599
rect 8816 8582 8833 8599
rect 8936 8582 8953 8599
rect 8656 8582 8673 8599
rect 9616 8582 9633 8599
rect 9576 8582 9593 8599
rect 9376 8582 9393 8599
rect 9536 8582 9553 8599
rect 9416 8582 9433 8599
rect 9496 8582 9513 8599
rect 9456 8582 9473 8599
rect 9096 8582 9113 8599
rect 9616 8582 9633 8599
rect 8456 8582 8473 8599
rect 9576 8582 9593 8599
rect 9536 8582 9553 8599
rect 7615 8582 7632 8599
rect 8335 8582 8352 8599
rect 7655 8582 7672 8599
rect 8095 8582 8112 8599
rect 7815 8582 7832 8599
rect 7695 8582 7712 8599
rect 7575 8582 7592 8599
rect 7975 8582 7992 8599
rect 7655 8582 7672 8599
rect 8055 8582 8072 8599
rect 7975 8582 7992 8599
rect 7535 8582 7552 8599
rect 8015 8582 8032 8599
rect 8135 8582 8152 8599
rect 7255 8582 7272 8599
rect 8295 8582 8312 8599
rect 7775 8582 7792 8599
rect 8416 8582 8433 8599
rect 7495 8582 7512 8599
rect 7935 8582 7952 8599
rect 7935 8582 7952 8599
rect 8055 8582 8072 8599
rect 7575 8582 7592 8599
rect 8095 8582 8112 8599
rect 7495 8582 7512 8599
rect 8255 8582 8272 8599
rect 8215 8582 8232 8599
rect 7735 8582 7752 8599
rect 8175 8582 8192 8599
rect 8416 8582 8433 8599
rect 8135 8582 8152 8599
rect 8015 8582 8032 8599
rect 8335 8582 8352 8599
rect 7375 8582 7392 8599
rect 7455 8582 7472 8599
rect 7255 8582 7272 8599
rect 7775 8582 7792 8599
rect 7735 8582 7752 8599
rect 7335 8582 7352 8599
rect 7895 8582 7912 8599
rect 7615 8582 7632 8599
rect 8295 8582 8312 8599
rect 7295 8582 7312 8599
rect 7815 8582 7832 8599
rect 8175 8582 8192 8599
rect 7455 8582 7472 8599
rect 7415 8582 7432 8599
rect 7855 8582 7872 8599
rect 7855 8582 7872 8599
rect 7375 8582 7392 8599
rect 8255 8582 8272 8599
rect 8376 8582 8393 8599
rect 7895 8582 7912 8599
rect 7335 8582 7352 8599
rect 8215 8582 8232 8599
rect 7295 8582 7312 8599
rect 8376 8582 8393 8599
rect 7535 8582 7552 8599
rect 7415 8582 7432 8599
rect 7695 8582 7712 8599
rect 6055 8582 6072 8599
rect 6055 8582 6072 8599
rect 6255 8582 6272 8599
rect 7055 8582 7072 8599
rect 7175 8582 7192 8599
rect 7095 8582 7112 8599
rect 6215 8582 6232 8599
rect 6495 8582 6512 8599
rect 6375 8582 6392 8599
rect 6175 8582 6192 8599
rect 6735 8582 6752 8599
rect 6415 8582 6432 8599
rect 6935 8582 6952 8599
rect 6775 8582 6792 8599
rect 6655 8582 6672 8599
rect 6255 8582 6272 8599
rect 6215 8582 6232 8599
rect 6935 8582 6952 8599
rect 6655 8582 6672 8599
rect 6815 8582 6832 8599
rect 6135 8582 6152 8599
rect 6455 8582 6472 8599
rect 6855 8582 6872 8599
rect 6455 8582 6472 8599
rect 7135 8582 7152 8599
rect 6135 8582 6152 8599
rect 6415 8582 6432 8599
rect 7015 8582 7032 8599
rect 6575 8582 6592 8599
rect 6095 8582 6112 8599
rect 6895 8582 6912 8599
rect 6535 8582 6552 8599
rect 7055 8582 7072 8599
rect 6095 8582 6112 8599
rect 6295 8582 6312 8599
rect 6535 8582 6552 8599
rect 6735 8582 6752 8599
rect 6575 8582 6592 8599
rect 6335 8582 6352 8599
rect 6975 8582 6992 8599
rect 6695 8582 6712 8599
rect 7175 8582 7192 8599
rect 6375 8582 6392 8599
rect 6615 8582 6632 8599
rect 7215 8582 7232 8599
rect 6295 8582 6312 8599
rect 6975 8582 6992 8599
rect 6815 8582 6832 8599
rect 6335 8582 6352 8599
rect 7135 8582 7152 8599
rect 6615 8582 6632 8599
rect 6695 8582 6712 8599
rect 6175 8582 6192 8599
rect 7095 8582 7112 8599
rect 7015 8582 7032 8599
rect 6495 8582 6512 8599
rect 6855 8582 6872 8599
rect 7215 8582 7232 8599
rect 6775 8582 6792 8599
rect 6895 8582 6912 8599
rect 5575 8582 5592 8599
rect 5695 8582 5712 8599
rect 5095 8582 5112 8599
rect 5295 8582 5312 8599
rect 5655 8582 5672 8599
rect 5415 8582 5432 8599
rect 5615 8582 5632 8599
rect 4935 8582 4952 8599
rect 5975 8582 5992 8599
rect 4895 8582 4912 8599
rect 5895 8582 5912 8599
rect 5735 8582 5752 8599
rect 5175 8582 5192 8599
rect 5935 8582 5952 8599
rect 5615 8582 5632 8599
rect 5575 8582 5592 8599
rect 5535 8582 5552 8599
rect 5855 8582 5872 8599
rect 5775 8582 5792 8599
rect 5055 8582 5072 8599
rect 5495 8582 5512 8599
rect 5455 8582 5472 8599
rect 5415 8582 5432 8599
rect 5935 8582 5952 8599
rect 4895 8582 4912 8599
rect 5775 8582 5792 8599
rect 5135 8582 5152 8599
rect 5255 8582 5272 8599
rect 5135 8582 5152 8599
rect 6015 8582 6032 8599
rect 5215 8582 5232 8599
rect 5335 8582 5352 8599
rect 5055 8582 5072 8599
rect 5455 8582 5472 8599
rect 5015 8582 5032 8599
rect 4975 8582 4992 8599
rect 4935 8582 4952 8599
rect 5535 8582 5552 8599
rect 5175 8582 5192 8599
rect 5255 8582 5272 8599
rect 5295 8582 5312 8599
rect 5495 8582 5512 8599
rect 5015 8582 5032 8599
rect 5815 8582 5832 8599
rect 6015 8582 6032 8599
rect 5815 8582 5832 8599
rect 5335 8582 5352 8599
rect 5975 8582 5992 8599
rect 5695 8582 5712 8599
rect 5375 8582 5392 8599
rect 5895 8582 5912 8599
rect 5855 8582 5872 8599
rect 5375 8582 5392 8599
rect 5095 8582 5112 8599
rect 5655 8582 5672 8599
rect 5735 8582 5752 8599
rect 5215 8582 5232 8599
rect 4975 8582 4992 8599
rect 3895 8582 3912 8599
rect 4735 8582 4752 8599
rect 4575 8582 4592 8599
rect 4695 8582 4712 8599
rect 4095 8582 4112 8599
rect 4655 8582 4672 8599
rect 4495 8582 4512 8599
rect 4815 8582 4832 8599
rect 3695 8582 3712 8599
rect 4815 8582 4832 8599
rect 3935 8582 3952 8599
rect 4295 8582 4312 8599
rect 4535 8582 4552 8599
rect 4855 8582 4872 8599
rect 3975 8582 3992 8599
rect 4615 8582 4632 8599
rect 4055 8582 4072 8599
rect 4175 8582 4192 8599
rect 4255 8582 4272 8599
rect 3855 8582 3872 8599
rect 4375 8582 4392 8599
rect 4735 8582 4752 8599
rect 3975 8582 3992 8599
rect 4775 8582 4792 8599
rect 3815 8582 3832 8599
rect 4335 8582 4352 8599
rect 4215 8582 4232 8599
rect 4455 8582 4472 8599
rect 4175 8582 4192 8599
rect 4215 8582 4232 8599
rect 3895 8582 3912 8599
rect 4335 8582 4352 8599
rect 4135 8582 4152 8599
rect 4295 8582 4312 8599
rect 4615 8582 4632 8599
rect 3735 8582 3752 8599
rect 3815 8582 3832 8599
rect 3775 8582 3792 8599
rect 4415 8582 4432 8599
rect 3775 8582 3792 8599
rect 4535 8582 4552 8599
rect 4855 8582 4872 8599
rect 3935 8582 3952 8599
rect 3735 8582 3752 8599
rect 4775 8582 4792 8599
rect 4455 8582 4472 8599
rect 4495 8582 4512 8599
rect 4375 8582 4392 8599
rect 4255 8582 4272 8599
rect 4135 8582 4152 8599
rect 4415 8582 4432 8599
rect 4015 8582 4032 8599
rect 3855 8582 3872 8599
rect 4095 8582 4112 8599
rect 4055 8582 4072 8599
rect 4695 8582 4712 8599
rect 4015 8582 4032 8599
rect 4575 8582 4592 8599
rect 3695 8582 3712 8599
rect 4655 8582 4672 8599
rect 3015 8582 3032 8599
rect 2655 8582 2672 8599
rect 3615 8582 3632 8599
rect 2735 8582 2752 8599
rect 2615 8582 2632 8599
rect 2975 8582 2992 8599
rect 2935 8582 2952 8599
rect 3175 8582 3192 8599
rect 3335 8582 3352 8599
rect 3215 8582 3232 8599
rect 3335 8582 3352 8599
rect 3455 8582 3472 8599
rect 2815 8582 2832 8599
rect 3375 8582 3392 8599
rect 3295 8582 3312 8599
rect 2775 8582 2792 8599
rect 2975 8582 2992 8599
rect 2535 8582 2552 8599
rect 3535 8582 3552 8599
rect 3135 8582 3152 8599
rect 2935 8582 2952 8599
rect 3175 8582 3192 8599
rect 2495 8582 2512 8599
rect 3615 8582 3632 8599
rect 3215 8582 3232 8599
rect 2855 8582 2872 8599
rect 3575 8582 3592 8599
rect 2855 8582 2872 8599
rect 3015 8582 3032 8599
rect 2895 8582 2912 8599
rect 3095 8582 3112 8599
rect 2895 8582 2912 8599
rect 2735 8582 2752 8599
rect 2655 8582 2672 8599
rect 3575 8582 3592 8599
rect 2575 8582 2592 8599
rect 2575 8582 2592 8599
rect 3655 8582 3672 8599
rect 2695 8582 2712 8599
rect 2495 8582 2512 8599
rect 2615 8582 2632 8599
rect 3495 8582 3512 8599
rect 3495 8582 3512 8599
rect 3455 8582 3472 8599
rect 3255 8582 3272 8599
rect 2535 8582 2552 8599
rect 2775 8582 2792 8599
rect 3535 8582 3552 8599
rect 3655 8582 3672 8599
rect 2815 8582 2832 8599
rect 3295 8582 3312 8599
rect 3415 8582 3432 8599
rect 3055 8582 3072 8599
rect 2695 8582 2712 8599
rect 3055 8582 3072 8599
rect 3095 8582 3112 8599
rect 3415 8582 3432 8599
rect 3135 8582 3152 8599
rect 3375 8582 3392 8599
rect 3255 8582 3272 8599
rect 1895 8582 1912 8599
rect 2215 8582 2232 8599
rect 2415 8582 2432 8599
rect 2095 8582 2112 8599
rect 2415 8582 2432 8599
rect 2015 8582 2032 8599
rect 2135 8582 2152 8599
rect 1935 8582 1952 8599
rect 2255 8582 2272 8599
rect 2215 8582 2232 8599
rect 316 8582 333 8599
rect 2175 8582 2192 8599
rect 2375 8582 2392 8599
rect 596 8582 613 8599
rect 476 8582 493 8599
rect 196 8582 213 8599
rect 956 8582 973 8599
rect 1036 8582 1053 8599
rect 2055 8582 2072 8599
rect 836 8582 853 8599
rect 2295 8582 2312 8599
rect 996 8582 1013 8599
rect 556 8582 573 8599
rect 1076 8582 1093 8599
rect 236 8582 253 8599
rect 2255 8582 2272 8599
rect 636 8582 653 8599
rect 276 8582 293 8599
rect 2335 8582 2352 8599
rect 676 8582 693 8599
rect 916 8582 933 8599
rect 1116 8582 1133 8599
rect 356 8582 373 8599
rect 1975 8582 1992 8599
rect 716 8582 733 8599
rect 1935 8582 1952 8599
rect 1895 8582 1912 8599
rect 2015 8582 2032 8599
rect 2135 8582 2152 8599
rect 756 8582 773 8599
rect 436 8582 453 8599
rect 1975 8582 1992 8599
rect 796 8582 813 8599
rect 2095 8582 2112 8599
rect 156 8582 173 8599
rect 2455 8582 2472 8599
rect 1156 8582 1173 8599
rect 2175 8582 2192 8599
rect 116 8582 133 8599
rect 2055 8582 2072 8599
rect 2455 8582 2472 8599
rect 396 8582 413 8599
rect 516 8582 533 8599
rect 2295 8582 2312 8599
rect 876 8582 893 8599
rect 2335 8582 2352 8599
rect 2375 8582 2392 8599
rect 6055 4652 6072 4669
rect 6055 4652 6072 4669
rect 6055 4652 6072 4669
rect 6055 4652 6072 4669
rect 6655 4652 6672 4669
rect 6655 4652 6672 4669
rect 6655 4652 6672 4669
rect 6655 4652 6672 4669
rect 7015 4652 7032 4669
rect 6735 4652 6752 4669
rect 6895 4652 6912 4669
rect 6975 4652 6992 4669
rect 6815 4652 6832 4669
rect 7055 4652 7072 4669
rect 6975 4652 6992 4669
rect 6975 4652 6992 4669
rect 7015 4652 7032 4669
rect 6735 4652 6752 4669
rect 7175 4652 7192 4669
rect 6775 4652 6792 4669
rect 6935 4652 6952 4669
rect 7215 4652 7232 4669
rect 6855 4652 6872 4669
rect 7055 4652 7072 4669
rect 7095 4652 7112 4669
rect 6855 4652 6872 4669
rect 7175 4652 7192 4669
rect 7215 4652 7232 4669
rect 6895 4652 6912 4669
rect 6695 4652 6712 4669
rect 6855 4652 6872 4669
rect 7055 4652 7072 4669
rect 6815 4652 6832 4669
rect 7215 4652 7232 4669
rect 6735 4652 6752 4669
rect 6935 4652 6952 4669
rect 7095 4652 7112 4669
rect 7175 4652 7192 4669
rect 6935 4652 6952 4669
rect 6775 4652 6792 4669
rect 6855 4652 6872 4669
rect 7135 4652 7152 4669
rect 6815 4652 6832 4669
rect 6775 4652 6792 4669
rect 6895 4652 6912 4669
rect 7015 4652 7032 4669
rect 6895 4652 6912 4669
rect 7135 4652 7152 4669
rect 7055 4652 7072 4669
rect 6695 4652 6712 4669
rect 6735 4652 6752 4669
rect 7015 4652 7032 4669
rect 6975 4652 6992 4669
rect 6815 4652 6832 4669
rect 7135 4652 7152 4669
rect 6695 4652 6712 4669
rect 7095 4652 7112 4669
rect 6935 4652 6952 4669
rect 7215 4652 7232 4669
rect 6775 4652 6792 4669
rect 7095 4652 7112 4669
rect 6695 4652 6712 4669
rect 7175 4652 7192 4669
rect 7135 4652 7152 4669
rect 6295 4652 6312 4669
rect 6375 4652 6392 4669
rect 6535 4652 6552 4669
rect 6495 4652 6512 4669
rect 6255 4652 6272 4669
rect 6415 4652 6432 4669
rect 6175 4652 6192 4669
rect 6135 4652 6152 4669
rect 6095 4652 6112 4669
rect 6255 4652 6272 4669
rect 6615 4652 6632 4669
rect 6175 4652 6192 4669
rect 6455 4652 6472 4669
rect 6135 4652 6152 4669
rect 6095 4652 6112 4669
rect 6295 4652 6312 4669
rect 6495 4652 6512 4669
rect 6215 4652 6232 4669
rect 6575 4652 6592 4669
rect 6535 4652 6552 4669
rect 6335 4652 6352 4669
rect 6575 4652 6592 4669
rect 6335 4652 6352 4669
rect 6455 4652 6472 4669
rect 6215 4652 6232 4669
rect 6415 4652 6432 4669
rect 6615 4652 6632 4669
rect 6255 4652 6272 4669
rect 6415 4652 6432 4669
rect 6455 4652 6472 4669
rect 6175 4652 6192 4669
rect 6455 4652 6472 4669
rect 6135 4652 6152 4669
rect 6095 4652 6112 4669
rect 6295 4652 6312 4669
rect 6335 4652 6352 4669
rect 6335 4652 6352 4669
rect 6175 4652 6192 4669
rect 6495 4652 6512 4669
rect 6375 4652 6392 4669
rect 6375 4652 6392 4669
rect 6215 4652 6232 4669
rect 6615 4652 6632 4669
rect 6135 4652 6152 4669
rect 6415 4652 6432 4669
rect 6575 4652 6592 4669
rect 6535 4652 6552 4669
rect 6095 4652 6112 4669
rect 6535 4652 6552 4669
rect 6575 4652 6592 4669
rect 6375 4652 6392 4669
rect 6615 4652 6632 4669
rect 6295 4652 6312 4669
rect 6495 4652 6512 4669
rect 6255 4652 6272 4669
rect 6215 4652 6232 4669
rect 5455 4652 5472 4669
rect 5455 4652 5472 4669
rect 5455 4652 5472 4669
rect 5455 4652 5472 4669
rect 5655 4652 5672 4669
rect 5655 4652 5672 4669
rect 5815 4652 5832 4669
rect 5975 4652 5992 4669
rect 5735 4652 5752 4669
rect 5975 4652 5992 4669
rect 5535 4652 5552 4669
rect 5775 4652 5792 4669
rect 6015 4652 6032 4669
rect 5815 4652 5832 4669
rect 5855 4652 5872 4669
rect 5695 4652 5712 4669
rect 5735 4652 5752 4669
rect 5895 4652 5912 4669
rect 5615 4652 5632 4669
rect 5775 4652 5792 4669
rect 5615 4652 5632 4669
rect 5495 4652 5512 4669
rect 5615 4652 5632 4669
rect 6015 4652 6032 4669
rect 5535 4652 5552 4669
rect 5495 4652 5512 4669
rect 5815 4652 5832 4669
rect 5935 4652 5952 4669
rect 5655 4652 5672 4669
rect 5575 4652 5592 4669
rect 5895 4652 5912 4669
rect 5655 4652 5672 4669
rect 5615 4652 5632 4669
rect 5575 4652 5592 4669
rect 5575 4652 5592 4669
rect 5735 4652 5752 4669
rect 5935 4652 5952 4669
rect 5575 4652 5592 4669
rect 5855 4652 5872 4669
rect 5895 4652 5912 4669
rect 5695 4652 5712 4669
rect 5935 4652 5952 4669
rect 5775 4652 5792 4669
rect 5855 4652 5872 4669
rect 6015 4652 6032 4669
rect 5975 4652 5992 4669
rect 5815 4652 5832 4669
rect 5855 4652 5872 4669
rect 5535 4652 5552 4669
rect 5775 4652 5792 4669
rect 5695 4652 5712 4669
rect 5495 4652 5512 4669
rect 6015 4652 6032 4669
rect 5975 4652 5992 4669
rect 5695 4652 5712 4669
rect 5895 4652 5912 4669
rect 5935 4652 5952 4669
rect 5495 4652 5512 4669
rect 5735 4652 5752 4669
rect 5535 4652 5552 4669
rect 5415 4652 5432 4669
rect 5375 4652 5392 4669
rect 4935 4652 4952 4669
rect 5415 4652 5432 4669
rect 5335 4652 5352 4669
rect 4895 4652 4912 4669
rect 5295 4652 5312 4669
rect 5255 4652 5272 4669
rect 4895 4652 4912 4669
rect 5215 4652 5232 4669
rect 5175 4652 5192 4669
rect 5295 4652 5312 4669
rect 5135 4652 5152 4669
rect 5255 4652 5272 4669
rect 5215 4652 5232 4669
rect 5375 4652 5392 4669
rect 5175 4652 5192 4669
rect 5135 4652 5152 4669
rect 5055 4652 5072 4669
rect 5055 4652 5072 4669
rect 5335 4652 5352 4669
rect 5095 4652 5112 4669
rect 5015 4652 5032 4669
rect 5095 4652 5112 4669
rect 4935 4652 4952 4669
rect 4975 4652 4992 4669
rect 5215 4652 5232 4669
rect 5255 4652 5272 4669
rect 5175 4652 5192 4669
rect 5335 4652 5352 4669
rect 5295 4652 5312 4669
rect 5135 4652 5152 4669
rect 4975 4652 4992 4669
rect 5415 4652 5432 4669
rect 5415 4652 5432 4669
rect 4895 4652 4912 4669
rect 5135 4652 5152 4669
rect 5015 4652 5032 4669
rect 5375 4652 5392 4669
rect 5095 4652 5112 4669
rect 4935 4652 4952 4669
rect 4895 4652 4912 4669
rect 5055 4652 5072 4669
rect 4975 4652 4992 4669
rect 5255 4652 5272 4669
rect 5215 4652 5232 4669
rect 5055 4652 5072 4669
rect 5015 4652 5032 4669
rect 4935 4652 4952 4669
rect 5175 4652 5192 4669
rect 5295 4652 5312 4669
rect 5015 4652 5032 4669
rect 5335 4652 5352 4669
rect 5375 4652 5392 4669
rect 5095 4652 5112 4669
rect 4975 4652 4992 4669
rect 9216 4652 9233 4669
rect 9056 4652 9073 4669
rect 9136 4652 9153 4669
rect 9376 4652 9393 4669
rect 9296 4652 9313 4669
rect 9176 4652 9193 4669
rect 9176 4652 9193 4669
rect 9136 4652 9153 4669
rect 9096 4652 9113 4669
rect 9376 4652 9393 4669
rect 9416 4652 9433 4669
rect 9056 4652 9073 4669
rect 9336 4652 9353 4669
rect 9376 4652 9393 4669
rect 9416 4652 9433 4669
rect 9096 4652 9113 4669
rect 9336 4652 9353 4669
rect 9256 4652 9273 4669
rect 9056 4652 9073 4669
rect 9296 4652 9313 4669
rect 9296 4652 9313 4669
rect 9336 4652 9353 4669
rect 9416 4652 9433 4669
rect 9096 4652 9113 4669
rect 9616 4652 9633 4669
rect 9256 4652 9273 4669
rect 9576 4652 9593 4669
rect 9216 4652 9233 4669
rect 9536 4652 9553 4669
rect 9216 4652 9233 4669
rect 9376 4652 9393 4669
rect 9496 4652 9513 4669
rect 9176 4652 9193 4669
rect 9176 4652 9193 4669
rect 9136 4652 9153 4669
rect 9096 4652 9113 4669
rect 9416 4652 9433 4669
rect 9056 4652 9073 4669
rect 9456 4652 9473 4669
rect 9296 4652 9313 4669
rect 9616 4652 9633 4669
rect 9576 4652 9593 4669
rect 9616 4652 9633 4669
rect 9576 4652 9593 4669
rect 9536 4652 9553 4669
rect 9496 4652 9513 4669
rect 9456 4652 9473 4669
rect 9616 4652 9633 4669
rect 9576 4652 9593 4669
rect 9536 4652 9553 4669
rect 9496 4652 9513 4669
rect 9456 4652 9473 4669
rect 9536 4652 9553 4669
rect 9496 4652 9513 4669
rect 9456 4652 9473 4669
rect 9136 4652 9153 4669
rect 9256 4652 9273 4669
rect 9336 4652 9353 4669
rect 9216 4652 9233 4669
rect 9256 4652 9273 4669
rect 8616 4652 8633 4669
rect 8616 4652 8633 4669
rect 8896 4652 8913 4669
rect 8856 4652 8873 4669
rect 8896 4652 8913 4669
rect 8816 4652 8833 4669
rect 8776 4652 8793 4669
rect 8856 4652 8873 4669
rect 8736 4652 8753 4669
rect 8696 4652 8713 4669
rect 8816 4652 8833 4669
rect 8656 4652 8673 4669
rect 8456 4652 8473 4669
rect 8776 4652 8793 4669
rect 8736 4652 8753 4669
rect 9016 4652 9033 4669
rect 8696 4652 8713 4669
rect 8656 4652 8673 4669
rect 8976 4652 8993 4669
rect 8576 4652 8593 4669
rect 8936 4652 8953 4669
rect 8496 4652 8513 4669
rect 9016 4652 9033 4669
rect 8976 4652 8993 4669
rect 8936 4652 8953 4669
rect 8536 4652 8553 4669
rect 8536 4652 8553 4669
rect 8496 4652 8513 4669
rect 8576 4652 8593 4669
rect 8456 4652 8473 4669
rect 8616 4652 8633 4669
rect 8616 4652 8633 4669
rect 8896 4652 8913 4669
rect 8856 4652 8873 4669
rect 8896 4652 8913 4669
rect 8816 4652 8833 4669
rect 8776 4652 8793 4669
rect 8856 4652 8873 4669
rect 8736 4652 8753 4669
rect 8696 4652 8713 4669
rect 8816 4652 8833 4669
rect 8656 4652 8673 4669
rect 8776 4652 8793 4669
rect 8736 4652 8753 4669
rect 9016 4652 9033 4669
rect 8696 4652 8713 4669
rect 8656 4652 8673 4669
rect 8976 4652 8993 4669
rect 8936 4652 8953 4669
rect 9016 4652 9033 4669
rect 8976 4652 8993 4669
rect 8936 4652 8953 4669
rect 8536 4652 8553 4669
rect 8536 4652 8553 4669
rect 8496 4652 8513 4669
rect 8576 4652 8593 4669
rect 8456 4652 8473 4669
rect 8496 4652 8513 4669
rect 8456 4652 8473 4669
rect 8576 4652 8593 4669
rect 7935 4652 7952 4669
rect 7975 4652 7992 4669
rect 8055 4652 8072 4669
rect 8255 4652 8272 4669
rect 7895 4652 7912 4669
rect 8416 4652 8433 4669
rect 8015 4652 8032 4669
rect 8135 4652 8152 4669
rect 7975 4652 7992 4669
rect 8015 4652 8032 4669
rect 8295 4652 8312 4669
rect 7935 4652 7952 4669
rect 8215 4652 8232 4669
rect 7935 4652 7952 4669
rect 7855 4652 7872 4669
rect 8095 4652 8112 4669
rect 8376 4652 8393 4669
rect 8255 4652 8272 4669
rect 8175 4652 8192 4669
rect 8416 4652 8433 4669
rect 8015 4652 8032 4669
rect 8335 4652 8352 4669
rect 8416 4652 8433 4669
rect 8055 4652 8072 4669
rect 8135 4652 8152 4669
rect 8215 4652 8232 4669
rect 7895 4652 7912 4669
rect 8335 4652 8352 4669
rect 8335 4652 8352 4669
rect 7895 4652 7912 4669
rect 8055 4652 8072 4669
rect 8175 4652 8192 4669
rect 8295 4652 8312 4669
rect 8295 4652 8312 4669
rect 8255 4652 8272 4669
rect 8376 4652 8393 4669
rect 8135 4652 8152 4669
rect 8255 4652 8272 4669
rect 8215 4652 8232 4669
rect 8175 4652 8192 4669
rect 7895 4652 7912 4669
rect 7855 4652 7872 4669
rect 8175 4652 8192 4669
rect 7855 4652 7872 4669
rect 8376 4652 8393 4669
rect 8135 4652 8152 4669
rect 8095 4652 8112 4669
rect 8095 4652 8112 4669
rect 8416 4652 8433 4669
rect 8376 4652 8393 4669
rect 7855 4652 7872 4669
rect 8055 4652 8072 4669
rect 8015 4652 8032 4669
rect 8215 4652 8232 4669
rect 7975 4652 7992 4669
rect 8095 4652 8112 4669
rect 7975 4652 7992 4669
rect 8295 4652 8312 4669
rect 8335 4652 8352 4669
rect 7935 4652 7952 4669
rect 7815 4652 7832 4669
rect 7815 4652 7832 4669
rect 7655 4652 7672 4669
rect 7695 4652 7712 4669
rect 7575 4652 7592 4669
rect 7255 4652 7272 4669
rect 7735 4652 7752 4669
rect 7255 4652 7272 4669
rect 7815 4652 7832 4669
rect 7615 4652 7632 4669
rect 7655 4652 7672 4669
rect 7695 4652 7712 4669
rect 7535 4652 7552 4669
rect 7255 4652 7272 4669
rect 7775 4652 7792 4669
rect 7495 4652 7512 4669
rect 7575 4652 7592 4669
rect 7495 4652 7512 4669
rect 7735 4652 7752 4669
rect 7375 4652 7392 4669
rect 7255 4652 7272 4669
rect 7775 4652 7792 4669
rect 7335 4652 7352 4669
rect 7615 4652 7632 4669
rect 7295 4652 7312 4669
rect 7415 4652 7432 4669
rect 7375 4652 7392 4669
rect 7535 4652 7552 4669
rect 7335 4652 7352 4669
rect 7775 4652 7792 4669
rect 7495 4652 7512 4669
rect 7295 4652 7312 4669
rect 7495 4652 7512 4669
rect 7735 4652 7752 4669
rect 7375 4652 7392 4669
rect 7535 4652 7552 4669
rect 7335 4652 7352 4669
rect 7415 4652 7432 4669
rect 7295 4652 7312 4669
rect 7415 4652 7432 4669
rect 7375 4652 7392 4669
rect 7335 4652 7352 4669
rect 7295 4652 7312 4669
rect 7535 4652 7552 4669
rect 7415 4652 7432 4669
rect 7455 4652 7472 4669
rect 7455 4652 7472 4669
rect 7815 4652 7832 4669
rect 7695 4652 7712 4669
rect 7455 4652 7472 4669
rect 7775 4652 7792 4669
rect 7735 4652 7752 4669
rect 7655 4652 7672 4669
rect 7695 4652 7712 4669
rect 7655 4652 7672 4669
rect 7615 4652 7632 4669
rect 7615 4652 7632 4669
rect 7455 4652 7472 4669
rect 7575 4652 7592 4669
rect 7575 4652 7592 4669
rect 1895 4652 1912 4669
rect 2135 4652 2152 4669
rect 2095 4652 2112 4669
rect 2175 4652 2192 4669
rect 2055 4652 2072 4669
rect 2215 4652 2232 4669
rect 2015 4652 2032 4669
rect 2095 4652 2112 4669
rect 2215 4652 2232 4669
rect 2055 4652 2072 4669
rect 1975 4652 1992 4669
rect 2295 4652 2312 4669
rect 1935 4652 1952 4669
rect 2015 4652 2032 4669
rect 1895 4652 1912 4669
rect 2255 4652 2272 4669
rect 2455 4652 2472 4669
rect 2455 4652 2472 4669
rect 2415 4652 2432 4669
rect 2135 4652 2152 4669
rect 2375 4652 2392 4669
rect 2175 4652 2192 4669
rect 2415 4652 2432 4669
rect 1975 4652 1992 4669
rect 2335 4652 2352 4669
rect 2335 4652 2352 4669
rect 2295 4652 2312 4669
rect 2375 4652 2392 4669
rect 1935 4652 1952 4669
rect 2255 4652 2272 4669
rect 1895 4652 1912 4669
rect 2455 4652 2472 4669
rect 2335 4652 2352 4669
rect 2415 4652 2432 4669
rect 2335 4652 2352 4669
rect 1895 4652 1912 4669
rect 2295 4652 2312 4669
rect 1975 4652 1992 4669
rect 2135 4652 2152 4669
rect 2255 4652 2272 4669
rect 2055 4652 2072 4669
rect 1975 4652 1992 4669
rect 2415 4652 2432 4669
rect 2215 4652 2232 4669
rect 2015 4652 2032 4669
rect 2135 4652 2152 4669
rect 2095 4652 2112 4669
rect 2295 4652 2312 4669
rect 2255 4652 2272 4669
rect 2055 4652 2072 4669
rect 2015 4652 2032 4669
rect 2175 4652 2192 4669
rect 2455 4652 2472 4669
rect 2175 4652 2192 4669
rect 1935 4652 1952 4669
rect 2095 4652 2112 4669
rect 1935 4652 1952 4669
rect 2215 4652 2232 4669
rect 2375 4652 2392 4669
rect 2375 4652 2392 4669
rect 236 4652 253 4669
rect 316 4652 333 4669
rect 956 4652 973 4669
rect 556 4652 573 4669
rect 276 4652 293 4669
rect 716 4652 733 4669
rect 436 4652 453 4669
rect 1156 4652 1173 4669
rect 516 4652 533 4669
rect 356 4652 373 4669
rect 1116 4652 1133 4669
rect 876 4652 893 4669
rect 996 4652 1013 4669
rect 316 4652 333 4669
rect 356 4652 373 4669
rect 476 4652 493 4669
rect 396 4652 413 4669
rect 116 4652 133 4669
rect 396 4652 413 4669
rect 436 4652 453 4669
rect 476 4652 493 4669
rect 516 4652 533 4669
rect 196 4652 213 4669
rect 556 4652 573 4669
rect 596 4652 613 4669
rect 596 4652 613 4669
rect 636 4652 653 4669
rect 676 4652 693 4669
rect 796 4652 813 4669
rect 1036 4652 1053 4669
rect 156 4652 173 4669
rect 716 4652 733 4669
rect 916 4652 933 4669
rect 756 4652 773 4669
rect 796 4652 813 4669
rect 836 4652 853 4669
rect 876 4652 893 4669
rect 276 4652 293 4669
rect 916 4652 933 4669
rect 956 4652 973 4669
rect 236 4652 253 4669
rect 996 4652 1013 4669
rect 1076 4652 1093 4669
rect 1036 4652 1053 4669
rect 1076 4652 1093 4669
rect 676 4652 693 4669
rect 1116 4652 1133 4669
rect 836 4652 853 4669
rect 1156 4652 1173 4669
rect 116 4652 133 4669
rect 156 4652 173 4669
rect 636 4652 653 4669
rect 756 4652 773 4669
rect 196 4652 213 4669
rect 4455 4652 4472 4669
rect 4575 4652 4592 4669
rect 4615 4652 4632 4669
rect 4535 4652 4552 4669
rect 4655 4652 4672 4669
rect 4815 4652 4832 4669
rect 4455 4652 4472 4669
rect 4855 4652 4872 4669
rect 4335 4652 4352 4669
rect 4535 4652 4552 4669
rect 4415 4652 4432 4669
rect 4855 4652 4872 4669
rect 4375 4652 4392 4669
rect 4335 4652 4352 4669
rect 4295 4652 4312 4669
rect 4295 4652 4312 4669
rect 4455 4652 4472 4669
rect 4375 4652 4392 4669
rect 4855 4652 4872 4669
rect 4415 4652 4432 4669
rect 4735 4652 4752 4669
rect 4695 4652 4712 4669
rect 4495 4652 4512 4669
rect 4695 4652 4712 4669
rect 4695 4652 4712 4669
rect 4735 4652 4752 4669
rect 4775 4652 4792 4669
rect 4855 4652 4872 4669
rect 4415 4652 4432 4669
rect 4655 4652 4672 4669
rect 4495 4652 4512 4669
rect 4535 4652 4552 4669
rect 4375 4652 4392 4669
rect 4615 4652 4632 4669
rect 4335 4652 4352 4669
rect 4815 4652 4832 4669
rect 4535 4652 4552 4669
rect 4775 4652 4792 4669
rect 4415 4652 4432 4669
rect 4775 4652 4792 4669
rect 4735 4652 4752 4669
rect 4655 4652 4672 4669
rect 4295 4652 4312 4669
rect 4615 4652 4632 4669
rect 4815 4652 4832 4669
rect 4575 4652 4592 4669
rect 4815 4652 4832 4669
rect 4495 4652 4512 4669
rect 4655 4652 4672 4669
rect 4695 4652 4712 4669
rect 4495 4652 4512 4669
rect 4575 4652 4592 4669
rect 4775 4652 4792 4669
rect 4455 4652 4472 4669
rect 4615 4652 4632 4669
rect 4375 4652 4392 4669
rect 4335 4652 4352 4669
rect 4295 4652 4312 4669
rect 4575 4652 4592 4669
rect 4735 4652 4752 4669
rect 3815 4652 3832 4669
rect 3775 4652 3792 4669
rect 3735 4652 3752 4669
rect 3695 4652 3712 4669
rect 4015 4652 4032 4669
rect 3975 4652 3992 4669
rect 3935 4652 3952 4669
rect 3895 4652 3912 4669
rect 3855 4652 3872 4669
rect 3815 4652 3832 4669
rect 4055 4652 4072 4669
rect 4255 4652 4272 4669
rect 4215 4652 4232 4669
rect 4175 4652 4192 4669
rect 4095 4652 4112 4669
rect 4135 4652 4152 4669
rect 3775 4652 3792 4669
rect 4095 4652 4112 4669
rect 4055 4652 4072 4669
rect 4255 4652 4272 4669
rect 4215 4652 4232 4669
rect 4015 4652 4032 4669
rect 4175 4652 4192 4669
rect 4095 4652 4112 4669
rect 3975 4652 3992 4669
rect 4135 4652 4152 4669
rect 3775 4652 3792 4669
rect 3935 4652 3952 4669
rect 4095 4652 4112 4669
rect 3735 4652 3752 4669
rect 4055 4652 4072 4669
rect 3895 4652 3912 4669
rect 3695 4652 3712 4669
rect 3815 4652 3832 4669
rect 4255 4652 4272 4669
rect 4015 4652 4032 4669
rect 3975 4652 3992 4669
rect 3855 4652 3872 4669
rect 4215 4652 4232 4669
rect 3935 4652 3952 4669
rect 4175 4652 4192 4669
rect 3895 4652 3912 4669
rect 3775 4652 3792 4669
rect 4135 4652 4152 4669
rect 3855 4652 3872 4669
rect 3815 4652 3832 4669
rect 3735 4652 3752 4669
rect 3695 4652 3712 4669
rect 3975 4652 3992 4669
rect 4215 4652 4232 4669
rect 3935 4652 3952 4669
rect 4175 4652 4192 4669
rect 3895 4652 3912 4669
rect 4135 4652 4152 4669
rect 3855 4652 3872 4669
rect 3735 4652 3752 4669
rect 4055 4652 4072 4669
rect 3695 4652 3712 4669
rect 4255 4652 4272 4669
rect 4015 4652 4032 4669
rect 3215 4652 3232 4669
rect 3255 4652 3272 4669
rect 3335 4652 3352 4669
rect 3535 4652 3552 4669
rect 3415 4652 3432 4669
rect 3255 4652 3272 4669
rect 3455 4652 3472 4669
rect 3095 4652 3112 4669
rect 3335 4652 3352 4669
rect 3255 4652 3272 4669
rect 3615 4652 3632 4669
rect 3655 4652 3672 4669
rect 3255 4652 3272 4669
rect 3215 4652 3232 4669
rect 3575 4652 3592 4669
rect 3295 4652 3312 4669
rect 3375 4652 3392 4669
rect 3655 4652 3672 4669
rect 3495 4652 3512 4669
rect 3415 4652 3432 4669
rect 3495 4652 3512 4669
rect 3135 4652 3152 4669
rect 3535 4652 3552 4669
rect 3215 4652 3232 4669
rect 3575 4652 3592 4669
rect 3415 4652 3432 4669
rect 3095 4652 3112 4669
rect 3135 4652 3152 4669
rect 3335 4652 3352 4669
rect 3215 4652 3232 4669
rect 3135 4652 3152 4669
rect 3095 4652 3112 4669
rect 3495 4652 3512 4669
rect 3615 4652 3632 4669
rect 3415 4652 3432 4669
rect 3175 4652 3192 4669
rect 3455 4652 3472 4669
rect 3175 4652 3192 4669
rect 3375 4652 3392 4669
rect 3175 4652 3192 4669
rect 3535 4652 3552 4669
rect 3615 4652 3632 4669
rect 3495 4652 3512 4669
rect 3335 4652 3352 4669
rect 3375 4652 3392 4669
rect 3175 4652 3192 4669
rect 3295 4652 3312 4669
rect 3295 4652 3312 4669
rect 3655 4652 3672 4669
rect 3375 4652 3392 4669
rect 3135 4652 3152 4669
rect 3295 4652 3312 4669
rect 3575 4652 3592 4669
rect 3615 4652 3632 4669
rect 3455 4652 3472 4669
rect 3655 4652 3672 4669
rect 3535 4652 3552 4669
rect 3575 4652 3592 4669
rect 3095 4652 3112 4669
rect 3455 4652 3472 4669
rect 2815 4652 2832 4669
rect 2975 4652 2992 4669
rect 2895 4652 2912 4669
rect 2775 4652 2792 4669
rect 2735 4652 2752 4669
rect 3015 4652 3032 4669
rect 3055 4652 3072 4669
rect 2535 4652 2552 4669
rect 2615 4652 2632 4669
rect 2735 4652 2752 4669
rect 2495 4652 2512 4669
rect 2855 4652 2872 4669
rect 2575 4652 2592 4669
rect 2815 4652 2832 4669
rect 2975 4652 2992 4669
rect 2695 4652 2712 4669
rect 2815 4652 2832 4669
rect 2655 4652 2672 4669
rect 2775 4652 2792 4669
rect 2935 4652 2952 4669
rect 2855 4652 2872 4669
rect 2655 4652 2672 4669
rect 2495 4652 2512 4669
rect 2535 4652 2552 4669
rect 3055 4652 3072 4669
rect 2695 4652 2712 4669
rect 2615 4652 2632 4669
rect 2895 4652 2912 4669
rect 2575 4652 2592 4669
rect 3015 4652 3032 4669
rect 2935 4652 2952 4669
rect 3055 4652 3072 4669
rect 2775 4652 2792 4669
rect 2495 4652 2512 4669
rect 2735 4652 2752 4669
rect 2895 4652 2912 4669
rect 2855 4652 2872 4669
rect 3015 4652 3032 4669
rect 2575 4652 2592 4669
rect 2655 4652 2672 4669
rect 2735 4652 2752 4669
rect 2975 4652 2992 4669
rect 2815 4652 2832 4669
rect 2695 4652 2712 4669
rect 2615 4652 2632 4669
rect 2695 4652 2712 4669
rect 2935 4652 2952 4669
rect 2775 4652 2792 4669
rect 2655 4652 2672 4669
rect 2535 4652 2552 4669
rect 3055 4652 3072 4669
rect 2615 4652 2632 4669
rect 2895 4652 2912 4669
rect 3015 4652 3032 4669
rect 2935 4652 2952 4669
rect 2855 4652 2872 4669
rect 2975 4652 2992 4669
rect 2575 4652 2592 4669
rect 2535 4652 2552 4669
rect 2495 4652 2512 4669
rect 2481 2394 2498 2411
rect 2481 2394 2498 2411
rect 4836 3163 4853 3180
rect 4836 3163 4853 3180
rect 4836 3163 4853 3180
rect 4836 3163 4853 3180
rect 4276 3163 4293 3180
rect 4276 3163 4293 3180
rect 4276 3163 4293 3180
rect 4276 3163 4293 3180
rect 4796 3163 4813 3180
rect 4796 3163 4813 3180
rect 4636 3163 4653 3180
rect 4756 3163 4773 3180
rect 4636 3163 4653 3180
rect 4716 3163 4733 3180
rect 4716 3163 4733 3180
rect 4596 3163 4613 3180
rect 4436 3163 4453 3180
rect 4356 3163 4373 3180
rect 4676 3163 4693 3180
rect 4756 3163 4773 3180
rect 4676 3163 4693 3180
rect 4316 3163 4333 3180
rect 4516 3163 4533 3180
rect 4556 3163 4573 3180
rect 4356 3163 4373 3180
rect 4756 3163 4773 3180
rect 4556 3163 4573 3180
rect 4476 3163 4493 3180
rect 4636 3163 4653 3180
rect 4356 3163 4373 3180
rect 4756 3163 4773 3180
rect 4516 3163 4533 3180
rect 4716 3163 4733 3180
rect 4316 3163 4333 3180
rect 4516 3163 4533 3180
rect 4316 3163 4333 3180
rect 4476 3163 4493 3180
rect 4596 3163 4613 3180
rect 4676 3163 4693 3180
rect 4556 3163 4573 3180
rect 4596 3163 4613 3180
rect 4396 3163 4413 3180
rect 4796 3163 4813 3180
rect 4796 3163 4813 3180
rect 4516 3163 4533 3180
rect 4476 3163 4493 3180
rect 4556 3163 4573 3180
rect 4436 3163 4453 3180
rect 4476 3163 4493 3180
rect 4676 3163 4693 3180
rect 4436 3163 4453 3180
rect 4316 3163 4333 3180
rect 4396 3163 4413 3180
rect 4436 3163 4453 3180
rect 4636 3163 4653 3180
rect 4716 3163 4733 3180
rect 4596 3163 4613 3180
rect 4356 3163 4373 3180
rect 4396 3163 4413 3180
rect 4396 3163 4413 3180
rect 3836 3163 3853 3180
rect 3876 3163 3893 3180
rect 3796 3163 3813 3180
rect 4036 3163 4053 3180
rect 4236 3163 4253 3180
rect 3916 3163 3933 3180
rect 3956 3163 3973 3180
rect 4116 3163 4133 3180
rect 3956 3163 3973 3180
rect 3836 3163 3853 3180
rect 3756 3163 3773 3180
rect 4116 3163 4133 3180
rect 4196 3163 4213 3180
rect 3796 3163 3813 3180
rect 3796 3163 3813 3180
rect 3756 3163 3773 3180
rect 4076 3163 4093 3180
rect 3836 3163 3853 3180
rect 4236 3163 4253 3180
rect 4076 3163 4093 3180
rect 4196 3163 4213 3180
rect 4196 3163 4213 3180
rect 3916 3163 3933 3180
rect 4156 3163 4173 3180
rect 3756 3163 3773 3180
rect 4156 3163 4173 3180
rect 4156 3163 4173 3180
rect 4036 3163 4053 3180
rect 4236 3163 4253 3180
rect 4156 3163 4173 3180
rect 4076 3163 4093 3180
rect 4036 3163 4053 3180
rect 3956 3163 3973 3180
rect 3876 3163 3893 3180
rect 4196 3163 4213 3180
rect 3876 3163 3893 3180
rect 3756 3163 3773 3180
rect 4116 3163 4133 3180
rect 3876 3163 3893 3180
rect 4076 3163 4093 3180
rect 3796 3163 3813 3180
rect 4036 3163 4053 3180
rect 3916 3163 3933 3180
rect 3996 3163 4013 3180
rect 4116 3163 4133 3180
rect 3836 3163 3853 3180
rect 3996 3163 4013 3180
rect 3996 3163 4013 3180
rect 3996 3163 4013 3180
rect 3956 3163 3973 3180
rect 4236 3163 4253 3180
rect 3916 3163 3933 3180
rect 3196 3163 3213 3180
rect 3196 3163 3213 3180
rect 3196 3163 3213 3180
rect 3196 3163 3213 3180
rect 3356 3163 3373 3180
rect 3636 3163 3653 3180
rect 3396 3163 3413 3180
rect 3596 3163 3613 3180
rect 3276 3163 3293 3180
rect 3676 3163 3693 3180
rect 3396 3163 3413 3180
rect 3316 3163 3333 3180
rect 3476 3163 3493 3180
rect 3396 3163 3413 3180
rect 3636 3163 3653 3180
rect 3716 3163 3733 3180
rect 3636 3163 3653 3180
rect 3316 3163 3333 3180
rect 3556 3163 3573 3180
rect 3596 3163 3613 3180
rect 3636 3163 3653 3180
rect 3596 3163 3613 3180
rect 3556 3163 3573 3180
rect 3236 3163 3253 3180
rect 3436 3163 3453 3180
rect 3716 3163 3733 3180
rect 3516 3163 3533 3180
rect 3716 3163 3733 3180
rect 3556 3163 3573 3180
rect 3436 3163 3453 3180
rect 3676 3163 3693 3180
rect 3556 3163 3573 3180
rect 3316 3163 3333 3180
rect 3516 3163 3533 3180
rect 3276 3163 3293 3180
rect 3356 3163 3373 3180
rect 3596 3163 3613 3180
rect 3396 3163 3413 3180
rect 3476 3163 3493 3180
rect 3236 3163 3253 3180
rect 3316 3163 3333 3180
rect 3476 3163 3493 3180
rect 3716 3163 3733 3180
rect 3436 3163 3453 3180
rect 3276 3163 3293 3180
rect 3236 3163 3253 3180
rect 3476 3163 3493 3180
rect 3236 3163 3253 3180
rect 3276 3163 3293 3180
rect 3356 3163 3373 3180
rect 3516 3163 3533 3180
rect 3516 3163 3533 3180
rect 3676 3163 3693 3180
rect 3436 3163 3453 3180
rect 3676 3163 3693 3180
rect 3356 3163 3373 3180
rect 3076 3163 3093 3180
rect 3116 3163 3133 3180
rect 2876 3163 2893 3180
rect 2996 3163 3013 3180
rect 3036 3163 3053 3180
rect 3076 3163 3093 3180
rect 3116 3163 3133 3180
rect 3116 3163 3133 3180
rect 2796 3163 2813 3180
rect 2996 3163 3013 3180
rect 2796 3163 2813 3180
rect 2676 3163 2693 3180
rect 2876 3163 2893 3180
rect 3116 3163 3133 3180
rect 2836 3163 2853 3180
rect 2916 3163 2933 3180
rect 3036 3163 3053 3180
rect 3076 3163 3093 3180
rect 2916 3163 2933 3180
rect 2796 3163 2813 3180
rect 2756 3163 2773 3180
rect 2716 3163 2733 3180
rect 3076 3163 3093 3180
rect 2836 3163 2853 3180
rect 3036 3163 3053 3180
rect 2836 3163 2853 3180
rect 2676 3163 2693 3180
rect 2836 3163 2853 3180
rect 2796 3163 2813 3180
rect 2956 3163 2973 3180
rect 2676 3163 2693 3180
rect 2876 3163 2893 3180
rect 2716 3163 2733 3180
rect 2956 3163 2973 3180
rect 2916 3163 2933 3180
rect 2716 3163 2733 3180
rect 2956 3163 2973 3180
rect 2956 3163 2973 3180
rect 3036 3163 3053 3180
rect 3156 3163 3173 3180
rect 2676 3163 2693 3180
rect 2876 3163 2893 3180
rect 2756 3163 2773 3180
rect 2996 3163 3013 3180
rect 2716 3163 2733 3180
rect 2996 3163 3013 3180
rect 3156 3163 3173 3180
rect 3156 3163 3173 3180
rect 2756 3163 2773 3180
rect 2916 3163 2933 3180
rect 3156 3163 3173 3180
rect 2756 3163 2773 3180
rect 2116 3163 2133 3180
rect 2116 3163 2133 3180
rect 2116 3163 2133 3180
rect 2116 3163 2133 3180
rect 2236 3163 2253 3180
rect 2196 3163 2213 3180
rect 2556 3163 2573 3180
rect 2636 3163 2653 3180
rect 2596 3163 2613 3180
rect 2276 3163 2293 3180
rect 2276 3163 2293 3180
rect 2516 3163 2533 3180
rect 2436 3163 2453 3180
rect 2316 3163 2333 3180
rect 2596 3163 2613 3180
rect 2596 3163 2613 3180
rect 2156 3163 2173 3180
rect 2596 3163 2613 3180
rect 2636 3163 2653 3180
rect 2636 3163 2653 3180
rect 2516 3163 2533 3180
rect 2476 3163 2493 3180
rect 2396 3163 2413 3180
rect 2396 3163 2413 3180
rect 2436 3163 2453 3180
rect 2396 3163 2413 3180
rect 2436 3163 2453 3180
rect 2196 3163 2213 3180
rect 2396 3163 2413 3180
rect 2516 3163 2533 3180
rect 2436 3163 2453 3180
rect 2356 3163 2373 3180
rect 2236 3163 2253 3180
rect 2556 3163 2573 3180
rect 2476 3163 2493 3180
rect 2356 3163 2373 3180
rect 2316 3163 2333 3180
rect 2516 3163 2533 3180
rect 2156 3163 2173 3180
rect 2276 3163 2293 3180
rect 2356 3163 2373 3180
rect 2476 3163 2493 3180
rect 2236 3163 2253 3180
rect 2156 3163 2173 3180
rect 2476 3163 2493 3180
rect 2556 3163 2573 3180
rect 2636 3163 2653 3180
rect 2156 3163 2173 3180
rect 2316 3163 2333 3180
rect 2316 3163 2333 3180
rect 2356 3163 2373 3180
rect 2276 3163 2293 3180
rect 2556 3163 2573 3180
rect 2196 3163 2213 3180
rect 2236 3163 2253 3180
rect 2196 3163 2213 3180
rect 1676 3163 1693 3180
rect 1876 3163 1893 3180
rect 1796 3163 1813 3180
rect 2076 3163 2093 3180
rect 1636 3163 1653 3180
rect 1676 3163 1693 3180
rect 1916 3163 1933 3180
rect 1876 3163 1893 3180
rect 1956 3163 1973 3180
rect 1996 3163 2013 3180
rect 1756 3163 1773 3180
rect 1836 3163 1853 3180
rect 1636 3163 1653 3180
rect 1876 3163 1893 3180
rect 2076 3163 2093 3180
rect 1716 3163 1733 3180
rect 1836 3163 1853 3180
rect 1996 3163 2013 3180
rect 1876 3163 1893 3180
rect 1596 3163 1613 3180
rect 1596 3163 1613 3180
rect 1956 3163 1973 3180
rect 1796 3163 1813 3180
rect 2076 3163 2093 3180
rect 1636 3163 1653 3180
rect 1716 3163 1733 3180
rect 1596 3163 1613 3180
rect 1636 3163 1653 3180
rect 1916 3163 1933 3180
rect 2036 3163 2053 3180
rect 1756 3163 1773 3180
rect 2076 3163 2093 3180
rect 2036 3163 2053 3180
rect 1956 3163 1973 3180
rect 1996 3163 2013 3180
rect 1596 3163 1613 3180
rect 1756 3163 1773 3180
rect 1676 3163 1693 3180
rect 1836 3163 1853 3180
rect 1796 3163 1813 3180
rect 1916 3163 1933 3180
rect 2036 3163 2053 3180
rect 1716 3163 1733 3180
rect 1836 3163 1853 3180
rect 1676 3163 1693 3180
rect 1956 3163 1973 3180
rect 1996 3163 2013 3180
rect 1796 3163 1813 3180
rect 2036 3163 2053 3180
rect 1916 3163 1933 3180
rect 1716 3163 1733 3180
rect 1756 3163 1773 3180
rect 1036 3163 1053 3180
rect 1036 3163 1053 3180
rect 1036 3163 1053 3180
rect 1036 3163 1053 3180
rect 1276 3163 1293 3180
rect 1476 3163 1493 3180
rect 1436 3163 1453 3180
rect 1476 3163 1493 3180
rect 1076 3163 1093 3180
rect 1116 3163 1133 3180
rect 1076 3163 1093 3180
rect 1156 3163 1173 3180
rect 1516 3163 1533 3180
rect 1156 3163 1173 3180
rect 1396 3163 1413 3180
rect 1556 3163 1573 3180
rect 1436 3163 1453 3180
rect 1276 3163 1293 3180
rect 1316 3163 1333 3180
rect 1196 3163 1213 3180
rect 1316 3163 1333 3180
rect 1356 3163 1373 3180
rect 1196 3163 1213 3180
rect 1236 3163 1253 3180
rect 1516 3163 1533 3180
rect 1236 3163 1253 3180
rect 1396 3163 1413 3180
rect 1556 3163 1573 3180
rect 1276 3163 1293 3180
rect 1116 3163 1133 3180
rect 1476 3163 1493 3180
rect 1516 3163 1533 3180
rect 1076 3163 1093 3180
rect 1396 3163 1413 3180
rect 1316 3163 1333 3180
rect 1276 3163 1293 3180
rect 1436 3163 1453 3180
rect 1556 3163 1573 3180
rect 1156 3163 1173 3180
rect 1236 3163 1253 3180
rect 1196 3163 1213 3180
rect 1316 3163 1333 3180
rect 1356 3163 1373 3180
rect 1356 3163 1373 3180
rect 1396 3163 1413 3180
rect 1356 3163 1373 3180
rect 1116 3163 1133 3180
rect 1196 3163 1213 3180
rect 1476 3163 1493 3180
rect 1116 3163 1133 3180
rect 1436 3163 1453 3180
rect 1556 3163 1573 3180
rect 1516 3163 1533 3180
rect 1076 3163 1093 3180
rect 1236 3163 1253 3180
rect 1156 3163 1173 3180
rect 516 3163 533 3180
rect 836 3163 853 3180
rect 556 3163 573 3180
rect 836 3163 853 3180
rect 676 3163 693 3180
rect 596 3163 613 3180
rect 836 3163 853 3180
rect 716 3163 733 3180
rect 596 3163 613 3180
rect 556 3163 573 3180
rect 516 3163 533 3180
rect 916 3163 933 3180
rect 716 3163 733 3180
rect 916 3163 933 3180
rect 756 3163 773 3180
rect 756 3163 773 3180
rect 676 3163 693 3180
rect 516 3163 533 3180
rect 796 3163 813 3180
rect 756 3163 773 3180
rect 996 3163 1013 3180
rect 676 3163 693 3180
rect 636 3163 653 3180
rect 796 3163 813 3180
rect 876 3163 893 3180
rect 916 3163 933 3180
rect 876 3163 893 3180
rect 636 3163 653 3180
rect 756 3163 773 3180
rect 796 3163 813 3180
rect 716 3163 733 3180
rect 836 3163 853 3180
rect 996 3163 1013 3180
rect 716 3163 733 3180
rect 596 3163 613 3180
rect 676 3163 693 3180
rect 556 3163 573 3180
rect 516 3163 533 3180
rect 796 3163 813 3180
rect 956 3163 973 3180
rect 996 3163 1013 3180
rect 636 3163 653 3180
rect 916 3163 933 3180
rect 956 3163 973 3180
rect 996 3163 1013 3180
rect 596 3163 613 3180
rect 956 3163 973 3180
rect 876 3163 893 3180
rect 636 3163 653 3180
rect 876 3163 893 3180
rect 956 3163 973 3180
rect 556 3163 573 3180
rect 276 3163 293 3180
rect 476 3163 493 3180
rect 356 3163 373 3180
rect 396 3163 413 3180
rect 276 3163 293 3180
rect 356 3163 373 3180
rect 156 3163 173 3180
rect 236 3163 253 3180
rect 236 3163 253 3180
rect 276 3163 293 3180
rect 156 3163 173 3180
rect 116 3163 133 3180
rect 236 3163 253 3180
rect 396 3163 413 3180
rect 316 3163 333 3180
rect 476 3163 493 3180
rect 116 3163 133 3180
rect 436 3163 453 3180
rect 436 3163 453 3180
rect 236 3163 253 3180
rect 276 3163 293 3180
rect 156 3163 173 3180
rect 356 3163 373 3180
rect 396 3163 413 3180
rect 476 3163 493 3180
rect 436 3163 453 3180
rect 316 3163 333 3180
rect 116 3163 133 3180
rect 476 3163 493 3180
rect 396 3163 413 3180
rect 356 3163 373 3180
rect 156 3163 173 3180
rect 196 3163 213 3180
rect 196 3163 213 3180
rect 196 3163 213 3180
rect 196 3163 213 3180
rect 316 3163 333 3180
rect 436 3163 453 3180
rect 316 3163 333 3180
rect 116 3163 133 3180
rect 1641 2394 1658 2411
rect 1161 2394 1178 2411
rect 1201 2394 1218 2411
rect 841 2394 858 2411
rect 1841 2394 1858 2411
rect 1481 2394 1498 2411
rect 1001 2394 1018 2411
rect 1001 2394 1018 2411
rect 1201 2394 1218 2411
rect 1361 2394 1378 2411
rect 1801 2394 1818 2411
rect 1121 2394 1138 2411
rect 1321 2394 1338 2411
rect 1721 2394 1738 2411
rect 1601 2394 1618 2411
rect 1241 2394 1258 2411
rect 2441 2394 2458 2411
rect 2001 2394 2018 2411
rect 2241 2394 2258 2411
rect 2201 2394 2218 2411
rect 2361 2394 2378 2411
rect 2001 2394 2018 2411
rect 2121 2394 2138 2411
rect 1921 2394 1938 2411
rect 1961 2394 1978 2411
rect 2161 2394 2178 2411
rect 2041 2394 2058 2411
rect 2401 2394 2418 2411
rect 2161 2394 2178 2411
rect 1921 2394 1938 2411
rect 2201 2394 2218 2411
rect 2281 2394 2298 2411
rect 2121 2394 2138 2411
rect 2321 2394 2338 2411
rect 2041 2394 2058 2411
rect 2081 2394 2098 2411
rect 2441 2394 2458 2411
rect 2361 2394 2378 2411
rect 2081 2394 2098 2411
rect 2281 2394 2298 2411
rect 1961 2394 1978 2411
rect 2401 2394 2418 2411
rect 2321 2394 2338 2411
rect 2241 2394 2258 2411
rect 961 2394 978 2411
rect 1681 2394 1698 2411
rect 881 2394 898 2411
rect 1881 2394 1898 2411
rect 1521 2394 1538 2411
rect 1041 2394 1058 2411
rect 1441 2394 1458 2411
rect 1121 2394 1138 2411
rect 1401 2394 1418 2411
rect 1681 2394 1698 2411
rect 1361 2394 1378 2411
rect 1081 2394 1098 2411
rect 841 2394 858 2411
rect 1081 2394 1098 2411
rect 1481 2394 1498 2411
rect 1521 2394 1538 2411
rect 1801 2394 1818 2411
rect 1881 2394 1898 2411
rect 1321 2394 1338 2411
rect 1721 2394 1738 2411
rect 921 2394 938 2411
rect 1441 2394 1458 2411
rect 1841 2394 1858 2411
rect 1761 2394 1778 2411
rect 1281 2394 1298 2411
rect 1641 2394 1658 2411
rect 1161 2394 1178 2411
rect 1561 2394 1578 2411
rect 1241 2394 1258 2411
rect 1601 2394 1618 2411
rect 1761 2394 1778 2411
rect 1401 2394 1418 2411
rect 921 2394 938 2411
rect 961 2394 978 2411
rect 1041 2394 1058 2411
rect 1561 2394 1578 2411
rect 881 2394 898 2411
rect 1281 2394 1298 2411
rect 3681 2394 3698 2411
rect 3681 2394 3698 2411
rect 2721 2394 2738 2411
rect 2921 2394 2938 2411
rect 2801 2394 2818 2411
rect 2761 2394 2778 2411
rect 2521 2394 2538 2411
rect 2601 2394 2618 2411
rect 2561 2394 2578 2411
rect 2641 2394 2658 2411
rect 2881 2394 2898 2411
rect 2961 2394 2978 2411
rect 2681 2394 2698 2411
rect 2601 2394 2618 2411
rect 2961 2394 2978 2411
rect 2681 2394 2698 2411
rect 2921 2394 2938 2411
rect 2521 2394 2538 2411
rect 2841 2394 2858 2411
rect 3561 2394 3578 2411
rect 3041 2394 3058 2411
rect 3121 2394 3138 2411
rect 3361 2394 3378 2411
rect 3081 2394 3098 2411
rect 3241 2394 3258 2411
rect 3561 2394 3578 2411
rect 3441 2394 3458 2411
rect 3481 2394 3498 2411
rect 3001 2394 3018 2411
rect 3641 2394 3658 2411
rect 3481 2394 3498 2411
rect 3401 2394 3418 2411
rect 3161 2394 3178 2411
rect 3321 2394 3338 2411
rect 3521 2394 3538 2411
rect 3081 2394 3098 2411
rect 3641 2394 3658 2411
rect 3521 2394 3538 2411
rect 3601 2394 3618 2411
rect 3201 2394 3218 2411
rect 3441 2394 3458 2411
rect 3001 2394 3018 2411
rect 3121 2394 3138 2411
rect 3601 2394 3618 2411
rect 3281 2394 3298 2411
rect 2641 2394 2658 2411
rect 3201 2394 3218 2411
rect 3401 2394 3418 2411
rect 3281 2394 3298 2411
rect 3041 2394 3058 2411
rect 2801 2394 2818 2411
rect 3241 2394 3258 2411
rect 3321 2394 3338 2411
rect 3361 2394 3378 2411
rect 3161 2394 3178 2411
rect 2721 2394 2738 2411
rect 2761 2394 2778 2411
rect 2561 2394 2578 2411
rect 2881 2394 2898 2411
rect 2841 2394 2858 2411
rect 4001 2394 4018 2411
rect 4521 2394 4538 2411
rect 4041 2394 4058 2411
rect 4601 2394 4618 2411
rect 4201 2394 4218 2411
rect 4481 2394 4498 2411
rect 3801 2394 3818 2411
rect 4601 2394 4618 2411
rect 4281 2394 4298 2411
rect 4721 2394 4738 2411
rect 4401 2394 4418 2411
rect 4081 2394 4098 2411
rect 4801 2394 4818 2411
rect 4161 2394 4178 2411
rect 3961 2394 3978 2411
rect 4241 2394 4258 2411
rect 4321 2394 4338 2411
rect 3921 2394 3938 2411
rect 4161 2394 4178 2411
rect 4121 2394 4138 2411
rect 3881 2394 3898 2411
rect 4201 2394 4218 2411
rect 4281 2394 4298 2411
rect 4361 2394 4378 2411
rect 4401 2394 4418 2411
rect 3761 2394 3778 2411
rect 3921 2394 3938 2411
rect 4561 2394 4578 2411
rect 4841 2394 4858 2411
rect 3761 2394 3778 2411
rect 4721 2394 4738 2411
rect 4481 2394 4498 2411
rect 3841 2394 3858 2411
rect 3721 2394 3738 2411
rect 4841 2394 4858 2411
rect 3841 2394 3858 2411
rect 3881 2394 3898 2411
rect 3721 2394 3738 2411
rect 4001 2394 4018 2411
rect 4041 2394 4058 2411
rect 4681 2394 4698 2411
rect 4641 2394 4658 2411
rect 3801 2394 3818 2411
rect 4521 2394 4538 2411
rect 4761 2394 4778 2411
rect 4361 2394 4378 2411
rect 4441 2394 4458 2411
rect 4641 2394 4658 2411
rect 4081 2394 4098 2411
rect 4801 2394 4818 2411
rect 4441 2394 4458 2411
rect 4681 2394 4698 2411
rect 4321 2394 4338 2411
rect 4121 2394 4138 2411
rect 4761 2394 4778 2411
rect 4241 2394 4258 2411
rect 4561 2394 4578 2411
rect 3961 2394 3978 2411
rect 7436 3163 7453 3180
rect 7276 3163 7293 3180
rect 7316 3163 7333 3180
rect 7276 3163 7293 3180
rect 7316 3163 7333 3180
rect 7356 3163 7373 3180
rect 7116 3163 7133 3180
rect 7236 3163 7253 3180
rect 7036 3163 7053 3180
rect 6996 3163 7013 3180
rect 7236 3163 7253 3180
rect 7476 3163 7493 3180
rect 7196 3163 7213 3180
rect 7196 3163 7213 3180
rect 7076 3163 7093 3180
rect 7116 3163 7133 3180
rect 6996 3163 7013 3180
rect 7076 3163 7093 3180
rect 7356 3163 7373 3180
rect 7276 3163 7293 3180
rect 7356 3163 7373 3180
rect 7156 3163 7173 3180
rect 7236 3163 7253 3180
rect 7476 3163 7493 3180
rect 7036 3163 7053 3180
rect 7036 3163 7053 3180
rect 6436 3163 6453 3180
rect 6436 3163 6453 3180
rect 6436 3163 6453 3180
rect 6436 3163 6453 3180
rect 6476 3163 6493 3180
rect 6516 3163 6533 3180
rect 6516 3163 6533 3180
rect 6636 3163 6653 3180
rect 6476 3163 6493 3180
rect 6596 3163 6613 3180
rect 6556 3163 6573 3180
rect 6636 3163 6653 3180
rect 6556 3163 6573 3180
rect 6596 3163 6613 3180
rect 6476 3163 6493 3180
rect 6636 3163 6653 3180
rect 6596 3163 6613 3180
rect 6556 3163 6573 3180
rect 6516 3163 6533 3180
rect 6476 3163 6493 3180
rect 6676 3163 6693 3180
rect 6676 3163 6693 3180
rect 6676 3163 6693 3180
rect 6676 3163 6693 3180
rect 6796 3163 6813 3180
rect 6756 3163 6773 3180
rect 6716 3163 6733 3180
rect 6956 3163 6973 3180
rect 6916 3163 6933 3180
rect 6876 3163 6893 3180
rect 6836 3163 6853 3180
rect 6796 3163 6813 3180
rect 6756 3163 6773 3180
rect 6716 3163 6733 3180
rect 6956 3163 6973 3180
rect 6916 3163 6933 3180
rect 6876 3163 6893 3180
rect 6836 3163 6853 3180
rect 6716 3163 6733 3180
rect 6956 3163 6973 3180
rect 6916 3163 6933 3180
rect 6876 3163 6893 3180
rect 6836 3163 6853 3180
rect 6796 3163 6813 3180
rect 6756 3163 6773 3180
rect 6716 3163 6733 3180
rect 6916 3163 6933 3180
rect 6956 3163 6973 3180
rect 6836 3163 6853 3180
rect 6636 3163 6653 3180
rect 6796 3163 6813 3180
rect 6756 3163 6773 3180
rect 6596 3163 6613 3180
rect 6556 3163 6573 3180
rect 6876 3163 6893 3180
rect 6516 3163 6533 3180
rect 6236 3163 6253 3180
rect 6236 3163 6253 3180
rect 5956 3163 5973 3180
rect 5916 3163 5933 3180
rect 5956 3163 5973 3180
rect 6036 3163 6053 3180
rect 6156 3163 6173 3180
rect 6356 3163 6373 3180
rect 6396 3163 6413 3180
rect 6276 3163 6293 3180
rect 6156 3163 6173 3180
rect 5916 3163 5933 3180
rect 6036 3163 6053 3180
rect 6156 3163 6173 3180
rect 5996 3163 6013 3180
rect 6316 3163 6333 3180
rect 6196 3163 6213 3180
rect 6396 3163 6413 3180
rect 6396 3163 6413 3180
rect 6356 3163 6373 3180
rect 6116 3163 6133 3180
rect 6316 3163 6333 3180
rect 6356 3163 6373 3180
rect 6356 3163 6373 3180
rect 6076 3163 6093 3180
rect 6036 3163 6053 3180
rect 6076 3163 6093 3180
rect 6196 3163 6213 3180
rect 5956 3163 5973 3180
rect 5996 3163 6013 3180
rect 6316 3163 6333 3180
rect 6076 3163 6093 3180
rect 5996 3163 6013 3180
rect 6076 3163 6093 3180
rect 5956 3163 5973 3180
rect 6196 3163 6213 3180
rect 6276 3163 6293 3180
rect 5916 3163 5933 3180
rect 6316 3163 6333 3180
rect 6116 3163 6133 3180
rect 6236 3163 6253 3180
rect 6156 3163 6173 3180
rect 5996 3163 6013 3180
rect 5916 3163 5933 3180
rect 6236 3163 6253 3180
rect 6116 3163 6133 3180
rect 6036 3163 6053 3180
rect 6276 3163 6293 3180
rect 6276 3163 6293 3180
rect 6396 3163 6413 3180
rect 6196 3163 6213 3180
rect 6116 3163 6133 3180
rect 5356 3163 5373 3180
rect 5356 3163 5373 3180
rect 5356 3163 5373 3180
rect 5356 3163 5373 3180
rect 5396 3163 5413 3180
rect 5756 3163 5773 3180
rect 5796 3163 5813 3180
rect 5436 3163 5453 3180
rect 5796 3163 5813 3180
rect 5476 3163 5493 3180
rect 5756 3163 5773 3180
rect 5516 3163 5533 3180
rect 5636 3163 5653 3180
rect 5436 3163 5453 3180
rect 5756 3163 5773 3180
rect 5596 3163 5613 3180
rect 5716 3163 5733 3180
rect 5556 3163 5573 3180
rect 5876 3163 5893 3180
rect 5396 3163 5413 3180
rect 5476 3163 5493 3180
rect 5436 3163 5453 3180
rect 5556 3163 5573 3180
rect 5716 3163 5733 3180
rect 5796 3163 5813 3180
rect 5876 3163 5893 3180
rect 5396 3163 5413 3180
rect 5716 3163 5733 3180
rect 5836 3163 5853 3180
rect 5676 3163 5693 3180
rect 5796 3163 5813 3180
rect 5676 3163 5693 3180
rect 5676 3163 5693 3180
rect 5716 3163 5733 3180
rect 5636 3163 5653 3180
rect 5556 3163 5573 3180
rect 5876 3163 5893 3180
rect 5596 3163 5613 3180
rect 5516 3163 5533 3180
rect 5396 3163 5413 3180
rect 5516 3163 5533 3180
rect 5756 3163 5773 3180
rect 5636 3163 5653 3180
rect 5676 3163 5693 3180
rect 5596 3163 5613 3180
rect 5596 3163 5613 3180
rect 5836 3163 5853 3180
rect 5836 3163 5853 3180
rect 5476 3163 5493 3180
rect 5556 3163 5573 3180
rect 5636 3163 5653 3180
rect 5836 3163 5853 3180
rect 5476 3163 5493 3180
rect 5876 3163 5893 3180
rect 5436 3163 5453 3180
rect 5516 3163 5533 3180
rect 5076 3163 5093 3180
rect 5316 3163 5333 3180
rect 5236 3163 5253 3180
rect 5076 3163 5093 3180
rect 4956 3163 4973 3180
rect 4956 3163 4973 3180
rect 7241 2394 7258 2411
rect 5116 3163 5133 3180
rect 7241 2394 7258 2411
rect 5036 3163 5053 3180
rect 5196 3163 5213 3180
rect 5156 3163 5173 3180
rect 5156 3163 5173 3180
rect 4916 3163 4933 3180
rect 5196 3163 5213 3180
rect 4876 3163 4893 3180
rect 4996 3163 5013 3180
rect 5196 3163 5213 3180
rect 5316 3163 5333 3180
rect 5196 3163 5213 3180
rect 4916 3163 4933 3180
rect 5116 3163 5133 3180
rect 5036 3163 5053 3180
rect 4876 3163 4893 3180
rect 5156 3163 5173 3180
rect 4916 3163 4933 3180
rect 5316 3163 5333 3180
rect 4996 3163 5013 3180
rect 4876 3163 4893 3180
rect 4956 3163 4973 3180
rect 5316 3163 5333 3180
rect 5036 3163 5053 3180
rect 5076 3163 5093 3180
rect 5276 3163 5293 3180
rect 5276 3163 5293 3180
rect 5236 3163 5253 3180
rect 5156 3163 5173 3180
rect 4876 3163 4893 3180
rect 5236 3163 5253 3180
rect 5276 3163 5293 3180
rect 5076 3163 5093 3180
rect 5116 3163 5133 3180
rect 5036 3163 5053 3180
rect 4916 3163 4933 3180
rect 4956 3163 4973 3180
rect 4996 3163 5013 3180
rect 5116 3163 5133 3180
rect 4996 3163 5013 3180
rect 5236 3163 5253 3180
rect 5276 3163 5293 3180
rect 9236 3163 9253 3180
rect 9236 3163 9253 3180
rect 9396 3163 9413 3180
rect 9436 3163 9453 3180
rect 9156 3163 9173 3180
rect 9596 3163 9613 3180
rect 9316 3163 9333 3180
rect 9476 3163 9493 3180
rect 9516 3163 9533 3180
rect 9356 3163 9373 3180
rect 9276 3163 9293 3180
rect 9276 3163 9293 3180
rect 9396 3163 9413 3180
rect 9476 3163 9493 3180
rect 9316 3163 9333 3180
rect 9436 3163 9453 3180
rect 9596 3163 9613 3180
rect 9476 3163 9493 3180
rect 9356 3163 9373 3180
rect 9556 3163 9573 3180
rect 9156 3163 9173 3180
rect 9156 3163 9173 3180
rect 9316 3163 9333 3180
rect 9276 3163 9293 3180
rect 9556 3163 9573 3180
rect 9596 3163 9613 3180
rect 9356 3163 9373 3180
rect 9436 3163 9453 3180
rect 9356 3163 9373 3180
rect 9196 3163 9213 3180
rect 9276 3163 9293 3180
rect 9396 3163 9413 3180
rect 9156 3163 9173 3180
rect 9436 3163 9453 3180
rect 9476 3163 9493 3180
rect 9396 3163 9413 3180
rect 9516 3163 9533 3180
rect 9236 3163 9253 3180
rect 9236 3163 9253 3180
rect 9556 3163 9573 3180
rect 9316 3163 9333 3180
rect 9596 3163 9613 3180
rect 9516 3163 9533 3180
rect 9196 3163 9213 3180
rect 9196 3163 9213 3180
rect 9196 3163 9213 3180
rect 9516 3163 9533 3180
rect 9556 3163 9573 3180
rect 8596 3163 8613 3180
rect 8596 3163 8613 3180
rect 8596 3163 8613 3180
rect 8596 3163 8613 3180
rect 8956 3163 8973 3180
rect 8956 3163 8973 3180
rect 8876 3163 8893 3180
rect 8716 3163 8733 3180
rect 8756 3163 8773 3180
rect 8916 3163 8933 3180
rect 8796 3163 8813 3180
rect 8956 3163 8973 3180
rect 8876 3163 8893 3180
rect 9116 3163 9133 3180
rect 8756 3163 8773 3180
rect 9076 3163 9093 3180
rect 9036 3163 9053 3180
rect 8956 3163 8973 3180
rect 8676 3163 8693 3180
rect 9076 3163 9093 3180
rect 8756 3163 8773 3180
rect 8796 3163 8813 3180
rect 8836 3163 8853 3180
rect 8636 3163 8653 3180
rect 8716 3163 8733 3180
rect 8716 3163 8733 3180
rect 8876 3163 8893 3180
rect 8836 3163 8853 3180
rect 8636 3163 8653 3180
rect 8916 3163 8933 3180
rect 9036 3163 9053 3180
rect 9036 3163 9053 3180
rect 8676 3163 8693 3180
rect 9116 3163 9133 3180
rect 8836 3163 8853 3180
rect 8996 3163 9013 3180
rect 8796 3163 8813 3180
rect 9036 3163 9053 3180
rect 9116 3163 9133 3180
rect 8636 3163 8653 3180
rect 8716 3163 8733 3180
rect 8916 3163 8933 3180
rect 8836 3163 8853 3180
rect 8996 3163 9013 3180
rect 9116 3163 9133 3180
rect 8676 3163 8693 3180
rect 9076 3163 9093 3180
rect 8996 3163 9013 3180
rect 8676 3163 8693 3180
rect 8916 3163 8933 3180
rect 8756 3163 8773 3180
rect 8796 3163 8813 3180
rect 8636 3163 8653 3180
rect 8996 3163 9013 3180
rect 9076 3163 9093 3180
rect 8876 3163 8893 3180
rect 8316 3163 8333 3180
rect 8196 3163 8213 3180
rect 8116 3163 8133 3180
rect 8196 3163 8213 3180
rect 8076 3163 8093 3180
rect 8396 3163 8413 3180
rect 8156 3163 8173 3180
rect 8276 3163 8293 3180
rect 8196 3163 8213 3180
rect 8556 3163 8573 3180
rect 8316 3163 8333 3180
rect 8316 3163 8333 3180
rect 8276 3163 8293 3180
rect 8516 3163 8533 3180
rect 8356 3163 8373 3180
rect 8476 3163 8493 3180
rect 8236 3163 8253 3180
rect 8396 3163 8413 3180
rect 8436 3163 8453 3180
rect 8076 3163 8093 3180
rect 8156 3163 8173 3180
rect 8116 3163 8133 3180
rect 8116 3163 8133 3180
rect 8076 3163 8093 3180
rect 8396 3163 8413 3180
rect 8236 3163 8253 3180
rect 8516 3163 8533 3180
rect 8556 3163 8573 3180
rect 8556 3163 8573 3180
rect 8276 3163 8293 3180
rect 8276 3163 8293 3180
rect 8476 3163 8493 3180
rect 8556 3163 8573 3180
rect 8156 3163 8173 3180
rect 8396 3163 8413 3180
rect 8316 3163 8333 3180
rect 8116 3163 8133 3180
rect 8236 3163 8253 3180
rect 8236 3163 8253 3180
rect 8516 3163 8533 3180
rect 8476 3163 8493 3180
rect 8436 3163 8453 3180
rect 8476 3163 8493 3180
rect 8156 3163 8173 3180
rect 8356 3163 8373 3180
rect 8436 3163 8453 3180
rect 8196 3163 8213 3180
rect 8436 3163 8453 3180
rect 8516 3163 8533 3180
rect 8356 3163 8373 3180
rect 8076 3163 8093 3180
rect 8356 3163 8373 3180
rect 7516 3163 7533 3180
rect 7516 3163 7533 3180
rect 7516 3163 7533 3180
rect 7516 3163 7533 3180
rect 7636 3163 7653 3180
rect 7916 3163 7933 3180
rect 7676 3163 7693 3180
rect 7716 3163 7733 3180
rect 7956 3163 7973 3180
rect 7596 3163 7613 3180
rect 7876 3163 7893 3180
rect 7596 3163 7613 3180
rect 7876 3163 7893 3180
rect 7756 3163 7773 3180
rect 8036 3163 8053 3180
rect 8036 3163 8053 3180
rect 7916 3163 7933 3180
rect 7956 3163 7973 3180
rect 7956 3163 7973 3180
rect 8036 3163 8053 3180
rect 7836 3163 7853 3180
rect 7716 3163 7733 3180
rect 7996 3163 8013 3180
rect 7836 3163 7853 3180
rect 7716 3163 7733 3180
rect 7756 3163 7773 3180
rect 7876 3163 7893 3180
rect 7596 3163 7613 3180
rect 7556 3163 7573 3180
rect 7716 3163 7733 3180
rect 7796 3163 7813 3180
rect 7556 3163 7573 3180
rect 7676 3163 7693 3180
rect 7556 3163 7573 3180
rect 7796 3163 7813 3180
rect 7796 3163 7813 3180
rect 7876 3163 7893 3180
rect 7996 3163 8013 3180
rect 7836 3163 7853 3180
rect 7756 3163 7773 3180
rect 7916 3163 7933 3180
rect 8036 3163 8053 3180
rect 7956 3163 7973 3180
rect 7676 3163 7693 3180
rect 7636 3163 7653 3180
rect 7676 3163 7693 3180
rect 7796 3163 7813 3180
rect 7996 3163 8013 3180
rect 7836 3163 7853 3180
rect 7636 3163 7653 3180
rect 7556 3163 7573 3180
rect 7996 3163 8013 3180
rect 7916 3163 7933 3180
rect 7596 3163 7613 3180
rect 7636 3163 7653 3180
rect 7756 3163 7773 3180
rect 7396 3163 7413 3180
rect 7156 3163 7173 3180
rect 6996 3163 7013 3180
rect 7076 3163 7093 3180
rect 7356 3163 7373 3180
rect 7196 3163 7213 3180
rect 7236 3163 7253 3180
rect 7076 3163 7093 3180
rect 7396 3163 7413 3180
rect 7436 3163 7453 3180
rect 7276 3163 7293 3180
rect 7316 3163 7333 3180
rect 7316 3163 7333 3180
rect 7116 3163 7133 3180
rect 7116 3163 7133 3180
rect 7156 3163 7173 3180
rect 7396 3163 7413 3180
rect 7156 3163 7173 3180
rect 7436 3163 7453 3180
rect 7476 3163 7493 3180
rect 6996 3163 7013 3180
rect 7036 3163 7053 3180
rect 7396 3163 7413 3180
rect 7436 3163 7453 3180
rect 7196 3163 7213 3180
rect 7476 3163 7493 3180
rect 9276 3163 9293 3180
rect 9556 3163 9573 3180
rect 9356 3163 9373 3180
rect 9476 3163 9493 3180
rect 9316 3163 9333 3180
rect 9596 3163 9613 3180
rect 9196 3163 9213 3180
rect 8996 3163 9013 3180
rect 9516 3163 9533 3180
rect 9516 3163 9533 3180
rect 8996 3163 9013 3180
rect 9196 3163 9213 3180
rect 9076 3163 9093 3180
rect 9276 3163 9293 3180
rect 9236 3163 9253 3180
rect 9196 3163 9213 3180
rect 9556 3163 9573 3180
rect 9156 3163 9173 3180
rect 9036 3163 9053 3180
rect 9196 3163 9213 3180
rect 9396 3163 9413 3180
rect 9356 3163 9373 3180
rect 9396 3163 9413 3180
rect 9116 3163 9133 3180
rect 9156 3163 9173 3180
rect 9556 3163 9573 3180
rect 9516 3163 9533 3180
rect 9276 3163 9293 3180
rect 9596 3163 9613 3180
rect 9556 3163 9573 3180
rect 9436 3163 9453 3180
rect 9436 3163 9453 3180
rect 9276 3163 9293 3180
rect 9036 3163 9053 3180
rect 9156 3163 9173 3180
rect 9476 3163 9493 3180
rect 9316 3163 9333 3180
rect 9396 3163 9413 3180
rect 9156 3163 9173 3180
rect 8956 3163 8973 3180
rect 9036 3163 9053 3180
rect 8956 3163 8973 3180
rect 9476 3163 9493 3180
rect 9356 3163 9373 3180
rect 9396 3163 9413 3180
rect 8996 3163 9013 3180
rect 9596 3163 9613 3180
rect 9316 3163 9333 3180
rect 9116 3163 9133 3180
rect 8956 3163 8973 3180
rect 9516 3163 9533 3180
rect 9436 3163 9453 3180
rect 9116 3163 9133 3180
rect 9316 3163 9333 3180
rect 9436 3163 9453 3180
rect 9236 3163 9253 3180
rect 9596 3163 9613 3180
rect 9076 3163 9093 3180
rect 9076 3163 9093 3180
rect 9036 3163 9053 3180
rect 9236 3163 9253 3180
rect 9116 3163 9133 3180
rect 8956 3163 8973 3180
rect 9476 3163 9493 3180
rect 9236 3163 9253 3180
rect 8996 3163 9013 3180
rect 9076 3163 9093 3180
rect 9356 3163 9373 3180
rect 8796 3163 8813 3180
rect 8596 3163 8613 3180
rect 8476 3163 8493 3180
rect 8876 3163 8893 3180
rect 8316 3163 8333 3180
rect 8156 3163 8173 3180
rect 8596 3163 8613 3180
rect 8916 3163 8933 3180
rect 8316 3163 8333 3180
rect 8036 3163 8053 3180
rect 8156 3163 8173 3180
rect 8596 3163 8613 3180
rect 8836 3163 8853 3180
rect 8036 3163 8053 3180
rect 7996 3163 8013 3180
rect 8276 3163 8293 3180
rect 8356 3163 8373 3180
rect 8316 3163 8333 3180
rect 8396 3163 8413 3180
rect 8516 3163 8533 3180
rect 8436 3163 8453 3180
rect 8276 3163 8293 3180
rect 8836 3163 8853 3180
rect 8196 3163 8213 3180
rect 8356 3163 8373 3180
rect 8196 3163 8213 3180
rect 8036 3163 8053 3180
rect 8876 3163 8893 3180
rect 8796 3163 8813 3180
rect 8316 3163 8333 3180
rect 8476 3163 8493 3180
rect 8716 3163 8733 3180
rect 8436 3163 8453 3180
rect 8916 3163 8933 3180
rect 8836 3163 8853 3180
rect 8236 3163 8253 3180
rect 7996 3163 8013 3180
rect 8756 3163 8773 3180
rect 8516 3163 8533 3180
rect 8116 3163 8133 3180
rect 8396 3163 8413 3180
rect 8916 3163 8933 3180
rect 8116 3163 8133 3180
rect 8356 3163 8373 3180
rect 8876 3163 8893 3180
rect 8436 3163 8453 3180
rect 8796 3163 8813 3180
rect 8676 3163 8693 3180
rect 8636 3163 8653 3180
rect 8076 3163 8093 3180
rect 8916 3163 8933 3180
rect 8076 3163 8093 3180
rect 8196 3163 8213 3180
rect 8156 3163 8173 3180
rect 8636 3163 8653 3180
rect 8876 3163 8893 3180
rect 8556 3163 8573 3180
rect 8676 3163 8693 3180
rect 8116 3163 8133 3180
rect 8356 3163 8373 3180
rect 8236 3163 8253 3180
rect 8076 3163 8093 3180
rect 8116 3163 8133 3180
rect 8476 3163 8493 3180
rect 8756 3163 8773 3180
rect 8716 3163 8733 3180
rect 8796 3163 8813 3180
rect 8076 3163 8093 3180
rect 8236 3163 8253 3180
rect 8276 3163 8293 3180
rect 8396 3163 8413 3180
rect 8836 3163 8853 3180
rect 8396 3163 8413 3180
rect 8516 3163 8533 3180
rect 8636 3163 8653 3180
rect 7996 3163 8013 3180
rect 8156 3163 8173 3180
rect 8636 3163 8653 3180
rect 8236 3163 8253 3180
rect 8476 3163 8493 3180
rect 8556 3163 8573 3180
rect 8276 3163 8293 3180
rect 7996 3163 8013 3180
rect 8676 3163 8693 3180
rect 8676 3163 8693 3180
rect 8516 3163 8533 3180
rect 8716 3163 8733 3180
rect 8196 3163 8213 3180
rect 8436 3163 8453 3180
rect 8596 3163 8613 3180
rect 8716 3163 8733 3180
rect 8756 3163 8773 3180
rect 8756 3163 8773 3180
rect 8556 3163 8573 3180
rect 8556 3163 8573 3180
rect 8036 3163 8053 3180
rect 4921 2394 4938 2411
rect 4921 2394 4938 2411
rect 4881 2394 4898 2411
rect 4881 2394 4898 2411
rect 4961 2394 4978 2411
rect 5041 2394 5058 2411
rect 5121 2394 5138 2411
rect 5121 2394 5138 2411
rect 5081 2394 5098 2411
rect 4961 2394 4978 2411
rect 5081 2394 5098 2411
rect 5001 2394 5018 2411
rect 5841 2394 5858 2411
rect 5641 2394 5658 2411
rect 5401 2394 5418 2411
rect 5241 2394 5258 2411
rect 6001 2394 6018 2411
rect 5521 2394 5538 2411
rect 5681 2394 5698 2411
rect 5921 2394 5938 2411
rect 5881 2394 5898 2411
rect 5761 2394 5778 2411
rect 5561 2394 5578 2411
rect 5601 2394 5618 2411
rect 5801 2394 5818 2411
rect 5481 2394 5498 2411
rect 5401 2394 5418 2411
rect 5361 2394 5378 2411
rect 5521 2394 5538 2411
rect 5961 2394 5978 2411
rect 5321 2394 5338 2411
rect 5761 2394 5778 2411
rect 5321 2394 5338 2411
rect 5961 2394 5978 2411
rect 5721 2394 5738 2411
rect 5201 2394 5218 2411
rect 5561 2394 5578 2411
rect 5441 2394 5458 2411
rect 5841 2394 5858 2411
rect 5641 2394 5658 2411
rect 5161 2394 5178 2411
rect 5481 2394 5498 2411
rect 6041 2394 6058 2411
rect 5441 2394 5458 2411
rect 5241 2394 5258 2411
rect 5721 2394 5738 2411
rect 5281 2394 5298 2411
rect 6041 2394 6058 2411
rect 5281 2394 5298 2411
rect 6001 2394 6018 2411
rect 5601 2394 5618 2411
rect 5681 2394 5698 2411
rect 5361 2394 5378 2411
rect 5161 2394 5178 2411
rect 5921 2394 5938 2411
rect 5881 2394 5898 2411
rect 5801 2394 5818 2411
rect 5201 2394 5218 2411
rect 5041 2394 5058 2411
rect 5001 2394 5018 2411
rect 6761 2394 6778 2411
rect 6881 2394 6898 2411
rect 6761 2394 6778 2411
rect 6961 2394 6978 2411
rect 6681 2394 6698 2411
rect 6321 2394 6338 2411
rect 6281 2394 6298 2411
rect 7041 2394 7058 2411
rect 6241 2394 6258 2411
rect 6441 2394 6458 2411
rect 6121 2394 6138 2411
rect 6401 2394 6418 2411
rect 6401 2394 6418 2411
rect 6081 2394 6098 2411
rect 6481 2394 6498 2411
rect 6161 2394 6178 2411
rect 6161 2394 6178 2411
rect 7001 2394 7018 2411
rect 6081 2394 6098 2411
rect 7161 2394 7178 2411
rect 6841 2394 6858 2411
rect 6121 2394 6138 2411
rect 6481 2394 6498 2411
rect 6721 2394 6738 2411
rect 6641 2394 6658 2411
rect 6721 2394 6738 2411
rect 7121 2394 7138 2411
rect 6361 2394 6378 2411
rect 6201 2394 6218 2411
rect 6641 2394 6658 2411
rect 7201 2394 7218 2411
rect 7081 2394 7098 2411
rect 7161 2394 7178 2411
rect 6601 2394 6618 2411
rect 6881 2394 6898 2411
rect 6201 2394 6218 2411
rect 7121 2394 7138 2411
rect 6321 2394 6338 2411
rect 6281 2394 6298 2411
rect 6521 2394 6538 2411
rect 6241 2394 6258 2411
rect 6361 2394 6378 2411
rect 6561 2394 6578 2411
rect 6801 2394 6818 2411
rect 6441 2394 6458 2411
rect 7081 2394 7098 2411
rect 7041 2394 7058 2411
rect 6601 2394 6618 2411
rect 6801 2394 6818 2411
rect 6561 2394 6578 2411
rect 6841 2394 6858 2411
rect 7001 2394 7018 2411
rect 7201 2394 7218 2411
rect 6961 2394 6978 2411
rect 6921 2394 6938 2411
rect 6681 2394 6698 2411
rect 6921 2394 6938 2411
rect 6521 2394 6538 2411
rect 8441 2394 8458 2411
rect 8441 2394 8458 2411
rect 7961 2394 7978 2411
rect 7881 2394 7898 2411
rect 8081 2394 8098 2411
rect 7401 2394 7418 2411
rect 7681 2394 7698 2411
rect 7841 2394 7858 2411
rect 7641 2394 7658 2411
rect 8241 2394 8258 2411
rect 7761 2394 7778 2411
rect 7281 2394 7298 2411
rect 7441 2394 7458 2411
rect 7441 2394 7458 2411
rect 7281 2394 7298 2411
rect 8401 2394 8418 2411
rect 8401 2394 8418 2411
rect 7361 2394 7378 2411
rect 7601 2394 7618 2411
rect 8321 2394 8338 2411
rect 7321 2394 7338 2411
rect 8361 2394 8378 2411
rect 8041 2394 8058 2411
rect 7881 2394 7898 2411
rect 8281 2394 8298 2411
rect 8201 2394 8218 2411
rect 8001 2394 8018 2411
rect 8241 2394 8258 2411
rect 7921 2394 7938 2411
rect 7721 2394 7738 2411
rect 8281 2394 8298 2411
rect 7761 2394 7778 2411
rect 7681 2394 7698 2411
rect 7961 2394 7978 2411
rect 7801 2394 7818 2411
rect 7641 2394 7658 2411
rect 8201 2394 8218 2411
rect 7601 2394 7618 2411
rect 8161 2394 8178 2411
rect 7721 2394 7738 2411
rect 7401 2394 7418 2411
rect 8121 2394 8138 2411
rect 7561 2394 7578 2411
rect 7361 2394 7378 2411
rect 8121 2394 8138 2411
rect 7921 2394 7938 2411
rect 7321 2394 7338 2411
rect 7841 2394 7858 2411
rect 8081 2394 8098 2411
rect 7521 2394 7538 2411
rect 7561 2394 7578 2411
rect 8041 2394 8058 2411
rect 8161 2394 8178 2411
rect 7521 2394 7538 2411
rect 7801 2394 7818 2411
rect 8361 2394 8378 2411
rect 7481 2394 7498 2411
rect 7481 2394 7498 2411
rect 8001 2394 8018 2411
rect 8321 2394 8338 2411
rect 9081 2394 9098 2411
rect 9041 2394 9058 2411
rect 9601 2394 9618 2411
rect 9481 2394 9498 2411
rect 8641 2394 8658 2411
rect 9441 2394 9458 2411
rect 9401 2394 9418 2411
rect 8601 2394 8618 2411
rect 9361 2394 9378 2411
rect 9321 2394 9338 2411
rect 8881 2394 8898 2411
rect 8601 2394 8618 2411
rect 9001 2394 9018 2411
rect 9281 2394 9298 2411
rect 9241 2394 9258 2411
rect 8961 2394 8978 2411
rect 9201 2394 9218 2411
rect 9161 2394 9178 2411
rect 8921 2394 8938 2411
rect 9121 2394 9138 2411
rect 9081 2394 9098 2411
rect 8881 2394 8898 2411
rect 9041 2394 9058 2411
rect 8841 2394 8858 2411
rect 8561 2394 8578 2411
rect 8521 2394 8538 2411
rect 8801 2394 8818 2411
rect 9441 2394 9458 2411
rect 8521 2394 8538 2411
rect 8841 2394 8858 2411
rect 9401 2394 9418 2411
rect 8481 2394 8498 2411
rect 8481 2394 8498 2411
rect 9481 2394 9498 2411
rect 8561 2394 8578 2411
rect 9521 2394 9538 2411
rect 8761 2394 8778 2411
rect 9561 2394 9578 2411
rect 9001 2394 9018 2411
rect 8721 2394 8738 2411
rect 8921 2394 8938 2411
rect 8961 2394 8978 2411
rect 8681 2394 8698 2411
rect 8641 2394 8658 2411
rect 9561 2394 9578 2411
rect 9361 2394 9378 2411
rect 8801 2394 8818 2411
rect 9321 2394 9338 2411
rect 9281 2394 9298 2411
rect 8761 2394 8778 2411
rect 9601 2394 9618 2411
rect 9241 2394 9258 2411
rect 9201 2394 9218 2411
rect 8721 2394 8738 2411
rect 9161 2394 9178 2411
rect 9121 2394 9138 2411
rect 9521 2394 9538 2411
rect 8681 2394 8698 2411
rect 15576 4652 15593 4669
rect 15576 4652 15593 4669
rect 15576 4652 15593 4669
rect 15576 4652 15593 4669
rect 16176 4652 16193 4669
rect 16176 4652 16193 4669
rect 16176 4652 16193 4669
rect 16176 4652 16193 4669
rect 16656 4652 16673 4669
rect 16616 4652 16633 4669
rect 16616 4652 16633 4669
rect 16216 4652 16233 4669
rect 16576 4652 16593 4669
rect 16456 4652 16473 4669
rect 16536 4652 16553 4669
rect 16656 4652 16673 4669
rect 16496 4652 16513 4669
rect 16456 4652 16473 4669
rect 16456 4652 16473 4669
rect 16696 4652 16713 4669
rect 16416 4652 16433 4669
rect 16536 4652 16553 4669
rect 16496 4652 16513 4669
rect 16376 4652 16393 4669
rect 16456 4652 16473 4669
rect 16696 4652 16713 4669
rect 16416 4652 16433 4669
rect 16656 4652 16673 4669
rect 16576 4652 16593 4669
rect 16416 4652 16433 4669
rect 16376 4652 16393 4669
rect 16336 4652 16353 4669
rect 16536 4652 16553 4669
rect 16336 4652 16353 4669
rect 16296 4652 16313 4669
rect 16496 4652 16513 4669
rect 16736 4652 16753 4669
rect 16256 4652 16273 4669
rect 16696 4652 16713 4669
rect 16656 4652 16673 4669
rect 16616 4652 16633 4669
rect 16616 4652 16633 4669
rect 16216 4652 16233 4669
rect 16576 4652 16593 4669
rect 16296 4652 16313 4669
rect 16736 4652 16753 4669
rect 16256 4652 16273 4669
rect 16216 4652 16233 4669
rect 16376 4652 16393 4669
rect 16336 4652 16353 4669
rect 16256 4652 16273 4669
rect 16536 4652 16553 4669
rect 16216 4652 16233 4669
rect 16336 4652 16353 4669
rect 16296 4652 16313 4669
rect 16696 4652 16713 4669
rect 16416 4652 16433 4669
rect 16576 4652 16593 4669
rect 16256 4652 16273 4669
rect 16296 4652 16313 4669
rect 16736 4652 16753 4669
rect 16496 4652 16513 4669
rect 16376 4652 16393 4669
rect 16736 4652 16753 4669
rect 15936 4652 15953 4669
rect 16056 4652 16073 4669
rect 16016 4652 16033 4669
rect 15976 4652 15993 4669
rect 15936 4652 15953 4669
rect 16056 4652 16073 4669
rect 16096 4652 16113 4669
rect 16096 4652 16113 4669
rect 16136 4652 16153 4669
rect 16136 4652 16153 4669
rect 15696 4652 15713 4669
rect 15816 4652 15833 4669
rect 15896 4652 15913 4669
rect 15776 4652 15793 4669
rect 15736 4652 15753 4669
rect 15656 4652 15673 4669
rect 15696 4652 15713 4669
rect 15816 4652 15833 4669
rect 15656 4652 15673 4669
rect 15856 4652 15873 4669
rect 15856 4652 15873 4669
rect 15736 4652 15753 4669
rect 15896 4652 15913 4669
rect 15776 4652 15793 4669
rect 15616 4652 15633 4669
rect 15616 4652 15633 4669
rect 16016 4652 16033 4669
rect 16136 4652 16153 4669
rect 15696 4652 15713 4669
rect 15816 4652 15833 4669
rect 15896 4652 15913 4669
rect 15776 4652 15793 4669
rect 15736 4652 15753 4669
rect 15656 4652 15673 4669
rect 15696 4652 15713 4669
rect 15816 4652 15833 4669
rect 15656 4652 15673 4669
rect 15856 4652 15873 4669
rect 15856 4652 15873 4669
rect 15736 4652 15753 4669
rect 15896 4652 15913 4669
rect 15776 4652 15793 4669
rect 16016 4652 16033 4669
rect 15976 4652 15993 4669
rect 15616 4652 15633 4669
rect 15936 4652 15953 4669
rect 16056 4652 16073 4669
rect 16016 4652 16033 4669
rect 15976 4652 15993 4669
rect 15936 4652 15953 4669
rect 16056 4652 16073 4669
rect 15616 4652 15633 4669
rect 16096 4652 16113 4669
rect 16096 4652 16113 4669
rect 15976 4652 15993 4669
rect 16136 4652 16153 4669
rect 14976 4652 14993 4669
rect 14976 4652 14993 4669
rect 14976 4652 14993 4669
rect 14976 4652 14993 4669
rect 15056 4652 15073 4669
rect 15016 4652 15033 4669
rect 15016 4652 15033 4669
rect 15056 4652 15073 4669
rect 15136 4652 15153 4669
rect 15176 4652 15193 4669
rect 15416 4652 15433 4669
rect 15376 4652 15393 4669
rect 15416 4652 15433 4669
rect 15496 4652 15513 4669
rect 15136 4652 15153 4669
rect 15096 4652 15113 4669
rect 15296 4652 15313 4669
rect 15216 4652 15233 4669
rect 15256 4652 15273 4669
rect 15376 4652 15393 4669
rect 15096 4652 15113 4669
rect 15296 4652 15313 4669
rect 15096 4652 15113 4669
rect 15496 4652 15513 4669
rect 15216 4652 15233 4669
rect 15536 4652 15553 4669
rect 15496 4652 15513 4669
rect 15056 4652 15073 4669
rect 15056 4652 15073 4669
rect 15336 4652 15353 4669
rect 15496 4652 15513 4669
rect 15176 4652 15193 4669
rect 15536 4652 15553 4669
rect 15456 4652 15473 4669
rect 15456 4652 15473 4669
rect 15016 4652 15033 4669
rect 15016 4652 15033 4669
rect 15336 4652 15353 4669
rect 15136 4652 15153 4669
rect 15336 4652 15353 4669
rect 15176 4652 15193 4669
rect 15216 4652 15233 4669
rect 15416 4652 15433 4669
rect 15256 4652 15273 4669
rect 15416 4652 15433 4669
rect 15456 4652 15473 4669
rect 15216 4652 15233 4669
rect 15456 4652 15473 4669
rect 15136 4652 15153 4669
rect 15176 4652 15193 4669
rect 15256 4652 15273 4669
rect 15536 4652 15553 4669
rect 15376 4652 15393 4669
rect 15296 4652 15313 4669
rect 15096 4652 15113 4669
rect 15536 4652 15553 4669
rect 15256 4652 15273 4669
rect 15376 4652 15393 4669
rect 15296 4652 15313 4669
rect 15336 4652 15353 4669
rect 14936 4652 14953 4669
rect 14896 4652 14913 4669
rect 14896 4652 14913 4669
rect 14856 4652 14873 4669
rect 14656 4652 14673 4669
rect 14616 4652 14633 4669
rect 14576 4652 14593 4669
rect 14536 4652 14553 4669
rect 14496 4652 14513 4669
rect 14456 4652 14473 4669
rect 14416 4652 14433 4669
rect 14816 4652 14833 4669
rect 14776 4652 14793 4669
rect 14736 4652 14753 4669
rect 14696 4652 14713 4669
rect 14656 4652 14673 4669
rect 14616 4652 14633 4669
rect 14576 4652 14593 4669
rect 14536 4652 14553 4669
rect 14496 4652 14513 4669
rect 14456 4652 14473 4669
rect 14416 4652 14433 4669
rect 14816 4652 14833 4669
rect 14776 4652 14793 4669
rect 14736 4652 14753 4669
rect 14696 4652 14713 4669
rect 14496 4652 14513 4669
rect 14616 4652 14633 4669
rect 14456 4652 14473 4669
rect 14936 4652 14953 4669
rect 14416 4652 14433 4669
rect 14816 4652 14833 4669
rect 14576 4652 14593 4669
rect 14776 4652 14793 4669
rect 14736 4652 14753 4669
rect 14856 4652 14873 4669
rect 14696 4652 14713 4669
rect 14536 4652 14553 4669
rect 14496 4652 14513 4669
rect 14936 4652 14953 4669
rect 14456 4652 14473 4669
rect 14416 4652 14433 4669
rect 14856 4652 14873 4669
rect 14816 4652 14833 4669
rect 14776 4652 14793 4669
rect 14736 4652 14753 4669
rect 14696 4652 14713 4669
rect 14656 4652 14673 4669
rect 14856 4652 14873 4669
rect 14616 4652 14633 4669
rect 14936 4652 14953 4669
rect 14656 4652 14673 4669
rect 14576 4652 14593 4669
rect 14896 4652 14913 4669
rect 14536 4652 14553 4669
rect 14896 4652 14913 4669
rect 18776 4652 18793 4669
rect 18616 4652 18633 4669
rect 18616 4652 18633 4669
rect 18976 4652 18993 4669
rect 18936 4652 18953 4669
rect 18896 4652 18913 4669
rect 18856 4652 18873 4669
rect 18816 4652 18833 4669
rect 18776 4652 18793 4669
rect 18736 4652 18753 4669
rect 19136 4652 19153 4669
rect 19096 4652 19113 4669
rect 19056 4652 19073 4669
rect 19016 4652 19033 4669
rect 18976 4652 18993 4669
rect 18936 4652 18953 4669
rect 18896 4652 18913 4669
rect 18856 4652 18873 4669
rect 18816 4652 18833 4669
rect 18776 4652 18793 4669
rect 18736 4652 18753 4669
rect 19136 4652 19153 4669
rect 19096 4652 19113 4669
rect 19056 4652 19073 4669
rect 19016 4652 19033 4669
rect 18696 4652 18713 4669
rect 18656 4652 18673 4669
rect 18696 4652 18713 4669
rect 18656 4652 18673 4669
rect 18736 4652 18753 4669
rect 19136 4652 19153 4669
rect 18576 4652 18593 4669
rect 19096 4652 19113 4669
rect 19056 4652 19073 4669
rect 19016 4652 19033 4669
rect 18976 4652 18993 4669
rect 18576 4652 18593 4669
rect 18936 4652 18953 4669
rect 18896 4652 18913 4669
rect 18856 4652 18873 4669
rect 18816 4652 18833 4669
rect 18776 4652 18793 4669
rect 18576 4652 18593 4669
rect 18736 4652 18753 4669
rect 19136 4652 19153 4669
rect 19096 4652 19113 4669
rect 19056 4652 19073 4669
rect 19016 4652 19033 4669
rect 18696 4652 18713 4669
rect 18656 4652 18673 4669
rect 18696 4652 18713 4669
rect 18656 4652 18673 4669
rect 18976 4652 18993 4669
rect 18936 4652 18953 4669
rect 18576 4652 18593 4669
rect 18896 4652 18913 4669
rect 18856 4652 18873 4669
rect 18816 4652 18833 4669
rect 18616 4652 18633 4669
rect 18616 4652 18633 4669
rect 18296 4652 18313 4669
rect 18336 4652 18353 4669
rect 18536 4652 18553 4669
rect 18256 4652 18273 4669
rect 18496 4652 18513 4669
rect 18216 4652 18233 4669
rect 18176 4652 18193 4669
rect 18136 4652 18153 4669
rect 18096 4652 18113 4669
rect 18456 4652 18473 4669
rect 18416 4652 18433 4669
rect 18376 4652 18393 4669
rect 18536 4652 18553 4669
rect 18496 4652 18513 4669
rect 18456 4652 18473 4669
rect 18416 4652 18433 4669
rect 18376 4652 18393 4669
rect 18336 4652 18353 4669
rect 18296 4652 18313 4669
rect 18256 4652 18273 4669
rect 18216 4652 18233 4669
rect 18176 4652 18193 4669
rect 18136 4652 18153 4669
rect 18096 4652 18113 4669
rect 17976 4652 17993 4669
rect 18016 4652 18033 4669
rect 18056 4652 18073 4669
rect 18016 4652 18033 4669
rect 18056 4652 18073 4669
rect 17976 4652 17993 4669
rect 18016 4652 18033 4669
rect 18056 4652 18073 4669
rect 17976 4652 17993 4669
rect 18296 4652 18313 4669
rect 18336 4652 18353 4669
rect 18536 4652 18553 4669
rect 18256 4652 18273 4669
rect 18496 4652 18513 4669
rect 18216 4652 18233 4669
rect 18176 4652 18193 4669
rect 18136 4652 18153 4669
rect 18096 4652 18113 4669
rect 18456 4652 18473 4669
rect 18416 4652 18433 4669
rect 18376 4652 18393 4669
rect 17976 4652 17993 4669
rect 18016 4652 18033 4669
rect 18056 4652 18073 4669
rect 18536 4652 18553 4669
rect 18496 4652 18513 4669
rect 18456 4652 18473 4669
rect 18416 4652 18433 4669
rect 18376 4652 18393 4669
rect 18336 4652 18353 4669
rect 18296 4652 18313 4669
rect 18256 4652 18273 4669
rect 18216 4652 18233 4669
rect 18176 4652 18193 4669
rect 18136 4652 18153 4669
rect 18096 4652 18113 4669
rect 17656 4652 17673 4669
rect 17936 4652 17953 4669
rect 17616 4652 17633 4669
rect 17576 4652 17593 4669
rect 17376 4652 17393 4669
rect 17616 4652 17633 4669
rect 17456 4652 17473 4669
rect 17776 4652 17793 4669
rect 17776 4652 17793 4669
rect 17536 4652 17553 4669
rect 17536 4652 17553 4669
rect 17936 4652 17953 4669
rect 17416 4652 17433 4669
rect 17496 4652 17513 4669
rect 17496 4652 17513 4669
rect 17376 4652 17393 4669
rect 17656 4652 17673 4669
rect 17736 4652 17753 4669
rect 17896 4652 17913 4669
rect 17936 4652 17953 4669
rect 17416 4652 17433 4669
rect 17856 4652 17873 4669
rect 17536 4652 17553 4669
rect 17616 4652 17633 4669
rect 17856 4652 17873 4669
rect 17536 4652 17553 4669
rect 17576 4652 17593 4669
rect 17816 4652 17833 4669
rect 17816 4652 17833 4669
rect 17776 4652 17793 4669
rect 17376 4652 17393 4669
rect 17736 4652 17753 4669
rect 17456 4652 17473 4669
rect 17696 4652 17713 4669
rect 17656 4652 17673 4669
rect 17656 4652 17673 4669
rect 17896 4652 17913 4669
rect 17936 4652 17953 4669
rect 17896 4652 17913 4669
rect 17416 4652 17433 4669
rect 17496 4652 17513 4669
rect 17376 4652 17393 4669
rect 17696 4652 17713 4669
rect 17456 4652 17473 4669
rect 17856 4652 17873 4669
rect 17456 4652 17473 4669
rect 17616 4652 17633 4669
rect 17736 4652 17753 4669
rect 17856 4652 17873 4669
rect 17896 4652 17913 4669
rect 17696 4652 17713 4669
rect 17416 4652 17433 4669
rect 17576 4652 17593 4669
rect 17816 4652 17833 4669
rect 17816 4652 17833 4669
rect 17776 4652 17793 4669
rect 17576 4652 17593 4669
rect 17736 4652 17753 4669
rect 17496 4652 17513 4669
rect 17696 4652 17713 4669
rect 16776 4652 16793 4669
rect 16856 4652 16873 4669
rect 16816 4652 16833 4669
rect 16776 4652 16793 4669
rect 17216 4652 17233 4669
rect 17256 4652 17273 4669
rect 17256 4652 17273 4669
rect 17016 4652 17033 4669
rect 16976 4652 16993 4669
rect 17336 4652 17353 4669
rect 17296 4652 17313 4669
rect 16936 4652 16953 4669
rect 16896 4652 16913 4669
rect 16856 4652 16873 4669
rect 16976 4652 16993 4669
rect 16816 4652 16833 4669
rect 16936 4652 16953 4669
rect 17176 4652 17193 4669
rect 17176 4652 17193 4669
rect 17056 4652 17073 4669
rect 17136 4652 17153 4669
rect 17216 4652 17233 4669
rect 17096 4652 17113 4669
rect 17016 4652 17033 4669
rect 17056 4652 17073 4669
rect 16896 4652 16913 4669
rect 17336 4652 17353 4669
rect 17296 4652 17313 4669
rect 17136 4652 17153 4669
rect 16776 4652 16793 4669
rect 17096 4652 17113 4669
rect 16856 4652 16873 4669
rect 17216 4652 17233 4669
rect 17256 4652 17273 4669
rect 17256 4652 17273 4669
rect 17016 4652 17033 4669
rect 17056 4652 17073 4669
rect 16936 4652 16953 4669
rect 17336 4652 17353 4669
rect 16896 4652 16913 4669
rect 17296 4652 17313 4669
rect 17136 4652 17153 4669
rect 17096 4652 17113 4669
rect 16856 4652 16873 4669
rect 16976 4652 16993 4669
rect 16816 4652 16833 4669
rect 17336 4652 17353 4669
rect 17296 4652 17313 4669
rect 16816 4652 16833 4669
rect 16776 4652 16793 4669
rect 16976 4652 16993 4669
rect 17176 4652 17193 4669
rect 17176 4652 17193 4669
rect 17056 4652 17073 4669
rect 16936 4652 16953 4669
rect 16896 4652 16913 4669
rect 17136 4652 17153 4669
rect 17216 4652 17233 4669
rect 17096 4652 17113 4669
rect 17016 4652 17033 4669
rect 10816 4652 10833 4669
rect 10816 4652 10833 4669
rect 10816 4652 10833 4669
rect 10816 4652 10833 4669
rect 11416 4652 11433 4669
rect 11416 4652 11433 4669
rect 11416 4652 11433 4669
rect 11416 4652 11433 4669
rect 11456 4652 11473 4669
rect 11776 4652 11793 4669
rect 11816 4652 11833 4669
rect 11656 4652 11673 4669
rect 11776 4652 11793 4669
rect 11456 4652 11473 4669
rect 11776 4652 11793 4669
rect 11576 4652 11593 4669
rect 11896 4652 11913 4669
rect 11976 4652 11993 4669
rect 11696 4652 11713 4669
rect 11456 4652 11473 4669
rect 11976 4652 11993 4669
rect 11616 4652 11633 4669
rect 11656 4652 11673 4669
rect 11656 4652 11673 4669
rect 11456 4652 11473 4669
rect 11536 4652 11553 4669
rect 11936 4652 11953 4669
rect 11536 4652 11553 4669
rect 11936 4652 11953 4669
rect 11736 4652 11753 4669
rect 11896 4652 11913 4669
rect 11616 4652 11633 4669
rect 11536 4652 11553 4669
rect 11536 4652 11553 4669
rect 11616 4652 11633 4669
rect 11856 4652 11873 4669
rect 11896 4652 11913 4669
rect 11736 4652 11753 4669
rect 11696 4652 11713 4669
rect 11856 4652 11873 4669
rect 11816 4652 11833 4669
rect 11976 4652 11993 4669
rect 11736 4652 11753 4669
rect 11496 4652 11513 4669
rect 11656 4652 11673 4669
rect 11856 4652 11873 4669
rect 11576 4652 11593 4669
rect 11616 4652 11633 4669
rect 11496 4652 11513 4669
rect 11576 4652 11593 4669
rect 11736 4652 11753 4669
rect 11976 4652 11993 4669
rect 11936 4652 11953 4669
rect 11816 4652 11833 4669
rect 11576 4652 11593 4669
rect 11776 4652 11793 4669
rect 11936 4652 11953 4669
rect 11896 4652 11913 4669
rect 11856 4652 11873 4669
rect 11816 4652 11833 4669
rect 11696 4652 11713 4669
rect 11696 4652 11713 4669
rect 11496 4652 11513 4669
rect 11496 4652 11513 4669
rect 11376 4652 11393 4669
rect 11336 4652 11353 4669
rect 11376 4652 11393 4669
rect 11296 4652 11313 4669
rect 11176 4652 11193 4669
rect 11176 4652 11193 4669
rect 11216 4652 11233 4669
rect 11136 4652 11153 4669
rect 10856 4652 10873 4669
rect 10856 4652 10873 4669
rect 11096 4652 11113 4669
rect 11096 4652 11113 4669
rect 10936 4652 10953 4669
rect 11056 4652 11073 4669
rect 11256 4652 11273 4669
rect 11256 4652 11273 4669
rect 11216 4652 11233 4669
rect 11056 4652 11073 4669
rect 11056 4652 11073 4669
rect 10976 4652 10993 4669
rect 11176 4652 11193 4669
rect 11336 4652 11353 4669
rect 11216 4652 11233 4669
rect 11136 4652 11153 4669
rect 11376 4652 11393 4669
rect 11256 4652 11273 4669
rect 10856 4652 10873 4669
rect 10976 4652 10993 4669
rect 11096 4652 11113 4669
rect 11016 4652 11033 4669
rect 11096 4652 11113 4669
rect 11256 4652 11273 4669
rect 11176 4652 11193 4669
rect 11336 4652 11353 4669
rect 11016 4652 11033 4669
rect 11296 4652 11313 4669
rect 10896 4652 10913 4669
rect 11376 4652 11393 4669
rect 11136 4652 11153 4669
rect 10976 4652 10993 4669
rect 10896 4652 10913 4669
rect 10936 4652 10953 4669
rect 10856 4652 10873 4669
rect 11336 4652 11353 4669
rect 10936 4652 10953 4669
rect 11296 4652 11313 4669
rect 11056 4652 11073 4669
rect 11216 4652 11233 4669
rect 11016 4652 11033 4669
rect 10896 4652 10913 4669
rect 11136 4652 11153 4669
rect 10896 4652 10913 4669
rect 11016 4652 11033 4669
rect 11296 4652 11313 4669
rect 10976 4652 10993 4669
rect 10936 4652 10953 4669
rect 10216 4652 10233 4669
rect 10216 4652 10233 4669
rect 10216 4652 10233 4669
rect 10216 4652 10233 4669
rect 10536 4652 10553 4669
rect 10776 4652 10793 4669
rect 10376 4652 10393 4669
rect 10776 4652 10793 4669
rect 10336 4652 10353 4669
rect 10656 4652 10673 4669
rect 10456 4652 10473 4669
rect 10776 4652 10793 4669
rect 10296 4652 10313 4669
rect 10416 4652 10433 4669
rect 10616 4652 10633 4669
rect 10376 4652 10393 4669
rect 10536 4652 10553 4669
rect 10576 4652 10593 4669
rect 10496 4652 10513 4669
rect 10576 4652 10593 4669
rect 10456 4652 10473 4669
rect 10736 4652 10753 4669
rect 10256 4652 10273 4669
rect 10616 4652 10633 4669
rect 10576 4652 10593 4669
rect 10696 4652 10713 4669
rect 10496 4652 10513 4669
rect 10736 4652 10753 4669
rect 10736 4652 10753 4669
rect 10576 4652 10593 4669
rect 10656 4652 10673 4669
rect 10336 4652 10353 4669
rect 10696 4652 10713 4669
rect 10736 4652 10753 4669
rect 10536 4652 10553 4669
rect 10696 4652 10713 4669
rect 10296 4652 10313 4669
rect 10496 4652 10513 4669
rect 10656 4652 10673 4669
rect 10256 4652 10273 4669
rect 10336 4652 10353 4669
rect 10296 4652 10313 4669
rect 10256 4652 10273 4669
rect 10656 4652 10673 4669
rect 10616 4652 10633 4669
rect 10456 4652 10473 4669
rect 10416 4652 10433 4669
rect 10696 4652 10713 4669
rect 10496 4652 10513 4669
rect 10456 4652 10473 4669
rect 10616 4652 10633 4669
rect 10416 4652 10433 4669
rect 10536 4652 10553 4669
rect 10376 4652 10393 4669
rect 10776 4652 10793 4669
rect 10336 4652 10353 4669
rect 10296 4652 10313 4669
rect 10256 4652 10273 4669
rect 10416 4652 10433 4669
rect 10376 4652 10393 4669
rect 9976 4652 9993 4669
rect 9856 4652 9873 4669
rect 9696 4652 9713 4669
rect 10136 4652 10153 4669
rect 10096 4652 10113 4669
rect 9656 4652 9673 4669
rect 9816 4652 9833 4669
rect 9936 4652 9953 4669
rect 9776 4652 9793 4669
rect 9736 4652 9753 4669
rect 9896 4652 9913 4669
rect 9936 4652 9953 4669
rect 9896 4652 9913 4669
rect 9856 4652 9873 4669
rect 9816 4652 9833 4669
rect 9776 4652 9793 4669
rect 9736 4652 9753 4669
rect 9696 4652 9713 4669
rect 9656 4652 9673 4669
rect 9856 4652 9873 4669
rect 9896 4652 9913 4669
rect 9816 4652 9833 4669
rect 10136 4652 10153 4669
rect 9776 4652 9793 4669
rect 10096 4652 10113 4669
rect 9736 4652 9753 4669
rect 9856 4652 9873 4669
rect 9696 4652 9713 4669
rect 9656 4652 9673 4669
rect 10096 4652 10113 4669
rect 9936 4652 9953 4669
rect 9976 4652 9993 4669
rect 10136 4652 10153 4669
rect 9816 4652 9833 4669
rect 10056 4652 10073 4669
rect 10176 4652 10193 4669
rect 10016 4652 10033 4669
rect 9776 4652 9793 4669
rect 10056 4652 10073 4669
rect 9736 4652 9753 4669
rect 9976 4652 9993 4669
rect 10056 4652 10073 4669
rect 10016 4652 10033 4669
rect 9936 4652 9953 4669
rect 10016 4652 10033 4669
rect 9896 4652 9913 4669
rect 9696 4652 9713 4669
rect 9656 4652 9673 4669
rect 10176 4652 10193 4669
rect 10056 4652 10073 4669
rect 10176 4652 10193 4669
rect 10136 4652 10153 4669
rect 10096 4652 10113 4669
rect 9976 4652 9993 4669
rect 10016 4652 10033 4669
rect 10176 4652 10193 4669
rect 13896 4652 13913 4669
rect 13856 4652 13873 4669
rect 13816 4652 13833 4669
rect 14176 4652 14193 4669
rect 13896 4652 13913 4669
rect 13856 4652 13873 4669
rect 13816 4652 13833 4669
rect 13936 4652 13953 4669
rect 14136 4652 14153 4669
rect 14096 4652 14113 4669
rect 14056 4652 14073 4669
rect 14256 4652 14273 4669
rect 14296 4652 14313 4669
rect 14296 4652 14313 4669
rect 14376 4652 14393 4669
rect 14336 4652 14353 4669
rect 14376 4652 14393 4669
rect 14336 4652 14353 4669
rect 13976 4652 13993 4669
rect 14016 4652 14033 4669
rect 14256 4652 14273 4669
rect 14216 4652 14233 4669
rect 14216 4652 14233 4669
rect 14296 4652 14313 4669
rect 14296 4652 14313 4669
rect 14376 4652 14393 4669
rect 14336 4652 14353 4669
rect 14376 4652 14393 4669
rect 14336 4652 14353 4669
rect 13976 4652 13993 4669
rect 14016 4652 14033 4669
rect 14256 4652 14273 4669
rect 14216 4652 14233 4669
rect 13936 4652 13953 4669
rect 14176 4652 14193 4669
rect 13896 4652 13913 4669
rect 13856 4652 13873 4669
rect 13816 4652 13833 4669
rect 14176 4652 14193 4669
rect 14136 4652 14153 4669
rect 14096 4652 14113 4669
rect 14056 4652 14073 4669
rect 14256 4652 14273 4669
rect 14216 4652 14233 4669
rect 14176 4652 14193 4669
rect 14136 4652 14153 4669
rect 14096 4652 14113 4669
rect 14056 4652 14073 4669
rect 14016 4652 14033 4669
rect 13976 4652 13993 4669
rect 13936 4652 13953 4669
rect 13896 4652 13913 4669
rect 13856 4652 13873 4669
rect 13816 4652 13833 4669
rect 14136 4652 14153 4669
rect 14096 4652 14113 4669
rect 14056 4652 14073 4669
rect 14016 4652 14033 4669
rect 13976 4652 13993 4669
rect 13936 4652 13953 4669
rect 13536 4652 13553 4669
rect 13696 4652 13713 4669
rect 13256 4652 13273 4669
rect 13496 4652 13513 4669
rect 13496 4652 13513 4669
rect 13456 4652 13473 4669
rect 13416 4652 13433 4669
rect 13736 4652 13753 4669
rect 13376 4652 13393 4669
rect 13336 4652 13353 4669
rect 13616 4652 13633 4669
rect 13296 4652 13313 4669
rect 13256 4652 13273 4669
rect 13456 4652 13473 4669
rect 13216 4652 13233 4669
rect 13216 4652 13233 4669
rect 13696 4652 13713 4669
rect 13736 4652 13753 4669
rect 13416 4652 13433 4669
rect 13656 4652 13673 4669
rect 13576 4652 13593 4669
rect 13376 4652 13393 4669
rect 13776 4652 13793 4669
rect 13776 4652 13793 4669
rect 13656 4652 13673 4669
rect 13336 4652 13353 4669
rect 13576 4652 13593 4669
rect 13536 4652 13553 4669
rect 13296 4652 13313 4669
rect 13536 4652 13553 4669
rect 13696 4652 13713 4669
rect 13256 4652 13273 4669
rect 13496 4652 13513 4669
rect 13496 4652 13513 4669
rect 13456 4652 13473 4669
rect 13416 4652 13433 4669
rect 13736 4652 13753 4669
rect 13376 4652 13393 4669
rect 13336 4652 13353 4669
rect 13616 4652 13633 4669
rect 13296 4652 13313 4669
rect 13256 4652 13273 4669
rect 13456 4652 13473 4669
rect 13216 4652 13233 4669
rect 13216 4652 13233 4669
rect 13696 4652 13713 4669
rect 13736 4652 13753 4669
rect 13416 4652 13433 4669
rect 13656 4652 13673 4669
rect 13576 4652 13593 4669
rect 13376 4652 13393 4669
rect 13616 4652 13633 4669
rect 13616 4652 13633 4669
rect 13776 4652 13793 4669
rect 13776 4652 13793 4669
rect 13656 4652 13673 4669
rect 13336 4652 13353 4669
rect 13576 4652 13593 4669
rect 13536 4652 13553 4669
rect 13296 4652 13313 4669
rect 12696 4652 12713 4669
rect 12936 4652 12953 4669
rect 12776 4652 12793 4669
rect 12616 4652 12633 4669
rect 12616 4652 12633 4669
rect 12776 4652 12793 4669
rect 12816 4652 12833 4669
rect 12656 4652 12673 4669
rect 12656 4652 12673 4669
rect 12896 4652 12913 4669
rect 12696 4652 12713 4669
rect 12936 4652 12953 4669
rect 13176 4652 13193 4669
rect 12696 4652 12713 4669
rect 13136 4652 13153 4669
rect 13056 4652 13073 4669
rect 13096 4652 13113 4669
rect 13096 4652 13113 4669
rect 13016 4652 13033 4669
rect 13176 4652 13193 4669
rect 12616 4652 12633 4669
rect 13056 4652 13073 4669
rect 13016 4652 13033 4669
rect 13136 4652 13153 4669
rect 12976 4652 12993 4669
rect 12976 4652 12993 4669
rect 12776 4652 12793 4669
rect 12736 4652 12753 4669
rect 13176 4652 13193 4669
rect 12896 4652 12913 4669
rect 12856 4652 12873 4669
rect 12816 4652 12833 4669
rect 13136 4652 13153 4669
rect 13096 4652 13113 4669
rect 13176 4652 13193 4669
rect 13096 4652 13113 4669
rect 12856 4652 12873 4669
rect 12856 4652 12873 4669
rect 13056 4652 13073 4669
rect 12736 4652 12753 4669
rect 12816 4652 12833 4669
rect 13056 4652 13073 4669
rect 12656 4652 12673 4669
rect 13016 4652 13033 4669
rect 12616 4652 12633 4669
rect 12896 4652 12913 4669
rect 12776 4652 12793 4669
rect 12696 4652 12713 4669
rect 12736 4652 12753 4669
rect 13136 4652 13153 4669
rect 12976 4652 12993 4669
rect 13016 4652 13033 4669
rect 12896 4652 12913 4669
rect 12936 4652 12953 4669
rect 12936 4652 12953 4669
rect 12856 4652 12873 4669
rect 12976 4652 12993 4669
rect 12736 4652 12753 4669
rect 12816 4652 12833 4669
rect 12656 4652 12673 4669
rect 12336 4652 12353 4669
rect 12456 4652 12473 4669
rect 12136 4652 12153 4669
rect 12376 4652 12393 4669
rect 12416 4652 12433 4669
rect 12056 4652 12073 4669
rect 12016 4652 12033 4669
rect 12536 4652 12553 4669
rect 12216 4652 12233 4669
rect 12016 4652 12033 4669
rect 12496 4652 12513 4669
rect 12056 4652 12073 4669
rect 12016 4652 12033 4669
rect 12536 4652 12553 4669
rect 12216 4652 12233 4669
rect 12416 4652 12433 4669
rect 12376 4652 12393 4669
rect 12016 4652 12033 4669
rect 12496 4652 12513 4669
rect 12336 4652 12353 4669
rect 12576 4652 12593 4669
rect 12296 4652 12313 4669
rect 12096 4652 12113 4669
rect 12456 4652 12473 4669
rect 12256 4652 12273 4669
rect 12296 4652 12313 4669
rect 12536 4652 12553 4669
rect 12176 4652 12193 4669
rect 12576 4652 12593 4669
rect 12096 4652 12113 4669
rect 12256 4652 12273 4669
rect 12496 4652 12513 4669
rect 12576 4652 12593 4669
rect 12456 4652 12473 4669
rect 12536 4652 12553 4669
rect 12496 4652 12513 4669
rect 12176 4652 12193 4669
rect 12456 4652 12473 4669
rect 12416 4652 12433 4669
rect 12136 4652 12153 4669
rect 12416 4652 12433 4669
rect 12056 4652 12073 4669
rect 12376 4652 12393 4669
rect 12336 4652 12353 4669
rect 12296 4652 12313 4669
rect 12296 4652 12313 4669
rect 12256 4652 12273 4669
rect 12136 4652 12153 4669
rect 12216 4652 12233 4669
rect 12176 4652 12193 4669
rect 12136 4652 12153 4669
rect 12376 4652 12393 4669
rect 12096 4652 12113 4669
rect 12216 4652 12233 4669
rect 12096 4652 12113 4669
rect 12256 4652 12273 4669
rect 12576 4652 12593 4669
rect 12056 4652 12073 4669
rect 12336 4652 12353 4669
rect 12176 4652 12193 4669
rect 11156 3163 11173 3180
rect 10796 3163 10813 3180
rect 11116 3163 11133 3180
rect 11076 3163 11093 3180
rect 11036 3163 11053 3180
rect 10996 3163 11013 3180
rect 10956 3163 10973 3180
rect 10916 3163 10933 3180
rect 10876 3163 10893 3180
rect 11116 3163 11133 3180
rect 11076 3163 11093 3180
rect 11036 3163 11053 3180
rect 10796 3163 10813 3180
rect 11076 3163 11093 3180
rect 10956 3163 10973 3180
rect 11276 3163 11293 3180
rect 11276 3163 11293 3180
rect 11156 3163 11173 3180
rect 11156 3163 11173 3180
rect 10916 3163 10933 3180
rect 10876 3163 10893 3180
rect 10996 3163 11013 3180
rect 11196 3163 11213 3180
rect 11116 3163 11133 3180
rect 11036 3163 11053 3180
rect 10956 3163 10973 3180
rect 10876 3163 10893 3180
rect 10996 3163 11013 3180
rect 11236 3163 11253 3180
rect 11236 3163 11253 3180
rect 10916 3163 10933 3180
rect 10916 3163 10933 3180
rect 10796 3163 10813 3180
rect 11236 3163 11253 3180
rect 10876 3163 10893 3180
rect 11156 3163 11173 3180
rect 10676 3163 10693 3180
rect 10236 3163 10253 3180
rect 10276 3163 10293 3180
rect 10476 3163 10493 3180
rect 10436 3163 10453 3180
rect 10316 3163 10333 3180
rect 10556 3163 10573 3180
rect 10396 3163 10413 3180
rect 10716 3163 10733 3180
rect 10716 3163 10733 3180
rect 10516 3163 10533 3180
rect 10716 3163 10733 3180
rect 10476 3163 10493 3180
rect 10356 3163 10373 3180
rect 10556 3163 10573 3180
rect 10316 3163 10333 3180
rect 10436 3163 10453 3180
rect 10396 3163 10413 3180
rect 10436 3163 10453 3180
rect 10356 3163 10373 3180
rect 10236 3163 10253 3180
rect 10596 3163 10613 3180
rect 10676 3163 10693 3180
rect 10396 3163 10413 3180
rect 10276 3163 10293 3180
rect 10276 3163 10293 3180
rect 10636 3163 10653 3180
rect 10396 3163 10413 3180
rect 10556 3163 10573 3180
rect 10516 3163 10533 3180
rect 10636 3163 10653 3180
rect 10676 3163 10693 3180
rect 10236 3163 10253 3180
rect 10516 3163 10533 3180
rect 10676 3163 10693 3180
rect 10716 3163 10733 3180
rect 10596 3163 10613 3180
rect 10516 3163 10533 3180
rect 10636 3163 10653 3180
rect 10276 3163 10293 3180
rect 10316 3163 10333 3180
rect 10476 3163 10493 3180
rect 10436 3163 10453 3180
rect 10636 3163 10653 3180
rect 10476 3163 10493 3180
rect 10316 3163 10333 3180
rect 10356 3163 10373 3180
rect 10596 3163 10613 3180
rect 10356 3163 10373 3180
rect 10596 3163 10613 3180
rect 10556 3163 10573 3180
rect 10236 3163 10253 3180
rect 9676 3163 9693 3180
rect 9676 3163 9693 3180
rect 9676 3163 9693 3180
rect 9676 3163 9693 3180
rect 10116 3163 10133 3180
rect 9916 3163 9933 3180
rect 9836 3163 9853 3180
rect 9876 3163 9893 3180
rect 9836 3163 9853 3180
rect 9716 3163 9733 3180
rect 9956 3163 9973 3180
rect 9796 3163 9813 3180
rect 9996 3163 10013 3180
rect 9916 3163 9933 3180
rect 9796 3163 9813 3180
rect 10076 3163 10093 3180
rect 10196 3163 10213 3180
rect 9956 3163 9973 3180
rect 10196 3163 10213 3180
rect 9956 3163 9973 3180
rect 10156 3163 10173 3180
rect 9996 3163 10013 3180
rect 9796 3163 9813 3180
rect 9916 3163 9933 3180
rect 9916 3163 9933 3180
rect 9876 3163 9893 3180
rect 10076 3163 10093 3180
rect 9756 3163 9773 3180
rect 9836 3163 9853 3180
rect 10116 3163 10133 3180
rect 9756 3163 9773 3180
rect 9796 3163 9813 3180
rect 10036 3163 10053 3180
rect 9876 3163 9893 3180
rect 10036 3163 10053 3180
rect 10196 3163 10213 3180
rect 9716 3163 9733 3180
rect 9716 3163 9733 3180
rect 9996 3163 10013 3180
rect 9876 3163 9893 3180
rect 10196 3163 10213 3180
rect 9756 3163 9773 3180
rect 9756 3163 9773 3180
rect 10156 3163 10173 3180
rect 10156 3163 10173 3180
rect 10116 3163 10133 3180
rect 10036 3163 10053 3180
rect 10036 3163 10053 3180
rect 10076 3163 10093 3180
rect 9716 3163 9733 3180
rect 9956 3163 9973 3180
rect 9836 3163 9853 3180
rect 10156 3163 10173 3180
rect 10076 3163 10093 3180
rect 9996 3163 10013 3180
rect 10116 3163 10133 3180
rect 9636 3163 9653 3180
rect 9636 3163 9653 3180
rect 9636 3163 9653 3180
rect 9636 3163 9653 3180
rect 14277 3163 14294 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 14357 3163 14374 3180
rect 13997 3163 14014 3180
rect 14277 3163 14294 3180
rect 14357 3163 14374 3180
rect 14317 3163 14334 3180
rect 14357 3163 14374 3180
rect 14277 3163 14294 3180
rect 14317 3163 14334 3180
rect 14237 3163 14254 3180
rect 14277 3163 14294 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14357 3163 14374 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14317 3163 14334 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14317 3163 14334 3180
rect 13837 3163 13854 3180
rect 13957 3163 13974 3180
rect 13917 3163 13934 3180
rect 13877 3163 13894 3180
rect 13837 3163 13854 3180
rect 13917 3163 13934 3180
rect 13917 3163 13934 3180
rect 13517 3163 13534 3180
rect 13597 3163 13614 3180
rect 13597 3163 13614 3180
rect 13877 3163 13894 3180
rect 13677 3163 13694 3180
rect 13837 3163 13854 3180
rect 13837 3163 13854 3180
rect 13557 3163 13574 3180
rect 13957 3163 13974 3180
rect 13877 3163 13894 3180
rect 13957 3163 13974 3180
rect 13637 3163 13654 3180
rect 13957 3163 13974 3180
rect 13917 3163 13934 3180
rect 13757 3163 13774 3180
rect 13877 3163 13894 3180
rect 13477 3163 13494 3180
rect 13797 3163 13814 3180
rect 13717 3163 13734 3180
rect 13797 3163 13814 3180
rect 13797 3163 13814 3180
rect 13757 3163 13774 3180
rect 13757 3163 13774 3180
rect 13717 3163 13734 3180
rect 13677 3163 13694 3180
rect 13637 3163 13654 3180
rect 13677 3163 13694 3180
rect 13597 3163 13614 3180
rect 13557 3163 13574 3180
rect 13517 3163 13534 3180
rect 13477 3163 13494 3180
rect 13557 3163 13574 3180
rect 13717 3163 13734 3180
rect 13637 3163 13654 3180
rect 13677 3163 13694 3180
rect 13597 3163 13614 3180
rect 13717 3163 13734 3180
rect 13637 3163 13654 3180
rect 13517 3163 13534 3180
rect 13557 3163 13574 3180
rect 13477 3163 13494 3180
rect 13757 3163 13774 3180
rect 13517 3163 13534 3180
rect 13797 3163 13814 3180
rect 13477 3163 13494 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 13237 3163 13254 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13397 3163 13414 3180
rect 13037 3163 13054 3180
rect 13397 3163 13414 3180
rect 13197 3163 13214 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13357 3163 13374 3180
rect 13117 3163 13134 3180
rect 13437 3163 13454 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13037 3163 13054 3180
rect 13277 3163 13294 3180
rect 12997 3163 13014 3180
rect 13277 3163 13294 3180
rect 12957 3163 12974 3180
rect 13237 3163 13254 3180
rect 13197 3163 13214 3180
rect 13277 3163 13294 3180
rect 12957 3163 12974 3180
rect 13237 3163 13254 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13437 3163 13454 3180
rect 12997 3163 13014 3180
rect 13277 3163 13294 3180
rect 12997 3163 13014 3180
rect 13437 3163 13454 3180
rect 13197 3163 13214 3180
rect 13117 3163 13134 3180
rect 13117 3163 13134 3180
rect 13037 3163 13054 3180
rect 13037 3163 13054 3180
rect 13117 3163 13134 3180
rect 12957 3163 12974 3180
rect 13197 3163 13214 3180
rect 13077 3163 13094 3180
rect 13157 3163 13174 3180
rect 12997 3163 13014 3180
rect 13397 3163 13414 3180
rect 13357 3163 13374 3180
rect 13357 3163 13374 3180
rect 13357 3163 13374 3180
rect 13237 3163 13254 3180
rect 13437 3163 13454 3180
rect 12957 3163 12974 3180
rect 13397 3163 13414 3180
rect 12637 3163 12654 3180
rect 12677 3163 12694 3180
rect 12437 3163 12454 3180
rect 12517 3163 12534 3180
rect 12757 3163 12774 3180
rect 12637 3163 12654 3180
rect 12437 3163 12454 3180
rect 12757 3163 12774 3180
rect 12637 3163 12654 3180
rect 12517 3163 12534 3180
rect 12637 3163 12654 3180
rect 12797 3163 12814 3180
rect 12597 3163 12614 3180
rect 12477 3163 12494 3180
rect 12837 3163 12854 3180
rect 12797 3163 12814 3180
rect 12397 3163 12414 3180
rect 12597 3163 12614 3180
rect 12717 3163 12734 3180
rect 12877 3163 12894 3180
rect 12597 3163 12614 3180
rect 12877 3163 12894 3180
rect 12877 3163 12894 3180
rect 12757 3163 12774 3180
rect 12717 3163 12734 3180
rect 12557 3163 12574 3180
rect 12717 3163 12734 3180
rect 12477 3163 12494 3180
rect 12837 3163 12854 3180
rect 12477 3163 12494 3180
rect 12397 3163 12414 3180
rect 12397 3163 12414 3180
rect 12717 3163 12734 3180
rect 12557 3163 12574 3180
rect 12877 3163 12894 3180
rect 12677 3163 12694 3180
rect 12837 3163 12854 3180
rect 12797 3163 12814 3180
rect 12557 3163 12574 3180
rect 12477 3163 12494 3180
rect 12837 3163 12854 3180
rect 12757 3163 12774 3180
rect 12677 3163 12694 3180
rect 12437 3163 12454 3180
rect 12557 3163 12574 3180
rect 12397 3163 12414 3180
rect 12677 3163 12694 3180
rect 12797 3163 12814 3180
rect 12597 3163 12614 3180
rect 12517 3163 12534 3180
rect 12517 3163 12534 3180
rect 12437 3163 12454 3180
rect 11837 3163 11854 3180
rect 11837 3163 11854 3180
rect 11837 3163 11854 3180
rect 11837 3163 11854 3180
rect 12197 3163 12214 3180
rect 12277 3163 12294 3180
rect 12117 3163 12134 3180
rect 12237 3163 12254 3180
rect 11917 3163 11934 3180
rect 12037 3163 12054 3180
rect 11877 3163 11894 3180
rect 12357 3163 12374 3180
rect 12157 3163 12174 3180
rect 12357 3163 12374 3180
rect 12317 3163 12334 3180
rect 11957 3163 11974 3180
rect 12237 3163 12254 3180
rect 12317 3163 12334 3180
rect 11997 3163 12014 3180
rect 12237 3163 12254 3180
rect 12277 3163 12294 3180
rect 12197 3163 12214 3180
rect 11997 3163 12014 3180
rect 12117 3163 12134 3180
rect 11877 3163 11894 3180
rect 11877 3163 11894 3180
rect 12037 3163 12054 3180
rect 12197 3163 12214 3180
rect 12157 3163 12174 3180
rect 12077 3163 12094 3180
rect 12117 3163 12134 3180
rect 12077 3163 12094 3180
rect 12037 3163 12054 3180
rect 12197 3163 12214 3180
rect 11997 3163 12014 3180
rect 11957 3163 11974 3180
rect 12357 3163 12374 3180
rect 12317 3163 12334 3180
rect 12277 3163 12294 3180
rect 12317 3163 12334 3180
rect 12237 3163 12254 3180
rect 12077 3163 12094 3180
rect 11957 3163 11974 3180
rect 12357 3163 12374 3180
rect 12157 3163 12174 3180
rect 11997 3163 12014 3180
rect 11917 3163 11934 3180
rect 12037 3163 12054 3180
rect 12157 3163 12174 3180
rect 12117 3163 12134 3180
rect 11917 3163 11934 3180
rect 11957 3163 11974 3180
rect 12277 3163 12294 3180
rect 11917 3163 11934 3180
rect 12077 3163 12094 3180
rect 11877 3163 11894 3180
rect 11317 3163 11334 3180
rect 11397 3163 11414 3180
rect 11397 3163 11414 3180
rect 11637 3163 11654 3180
rect 11397 3163 11414 3180
rect 11717 3163 11734 3180
rect 11557 3163 11574 3180
rect 11637 3163 11654 3180
rect 11597 3163 11614 3180
rect 11477 3163 11494 3180
rect 11637 3163 11654 3180
rect 11757 3163 11774 3180
rect 11797 3163 11814 3180
rect 11557 3163 11574 3180
rect 11357 3163 11374 3180
rect 11437 3163 11454 3180
rect 11677 3163 11694 3180
rect 11397 3163 11414 3180
rect 11717 3163 11734 3180
rect 11517 3163 11534 3180
rect 11637 3163 11654 3180
rect 11357 3163 11374 3180
rect 11557 3163 11574 3180
rect 11677 3163 11694 3180
rect 11317 3163 11334 3180
rect 11797 3163 11814 3180
rect 11477 3163 11494 3180
rect 11437 3163 11454 3180
rect 11517 3163 11534 3180
rect 11437 3163 11454 3180
rect 11757 3163 11774 3180
rect 11437 3163 11454 3180
rect 11797 3163 11814 3180
rect 11477 3163 11494 3180
rect 11517 3163 11534 3180
rect 11317 3163 11334 3180
rect 11677 3163 11694 3180
rect 11757 3163 11774 3180
rect 11717 3163 11734 3180
rect 11597 3163 11614 3180
rect 11317 3163 11334 3180
rect 11357 3163 11374 3180
rect 11717 3163 11734 3180
rect 11797 3163 11814 3180
rect 11357 3163 11374 3180
rect 11517 3163 11534 3180
rect 11557 3163 11574 3180
rect 11597 3163 11614 3180
rect 11477 3163 11494 3180
rect 11597 3163 11614 3180
rect 11677 3163 11694 3180
rect 11757 3163 11774 3180
rect 10756 3163 10773 3180
rect 10756 3163 10773 3180
rect 10756 3163 10773 3180
rect 10756 3163 10773 3180
rect 11196 3163 11213 3180
rect 10836 3163 10853 3180
rect 10836 3163 10853 3180
rect 11036 3163 11053 3180
rect 10796 3163 10813 3180
rect 10836 3163 10853 3180
rect 11196 3163 11213 3180
rect 10836 3163 10853 3180
rect 11116 3163 11133 3180
rect 10996 3163 11013 3180
rect 11076 3163 11093 3180
rect 10956 3163 10973 3180
rect 11276 3163 11293 3180
rect 11236 3163 11253 3180
rect 11196 3163 11213 3180
rect 11276 3163 11293 3180
rect 11797 3163 11814 3180
rect 11797 3163 11814 3180
rect 11797 3163 11814 3180
rect 11797 3163 11814 3180
rect 14357 3163 14374 3180
rect 14317 3163 14334 3180
rect 14357 3163 14374 3180
rect 14277 3163 14294 3180
rect 14317 3163 14334 3180
rect 14237 3163 14254 3180
rect 14277 3163 14294 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14357 3163 14374 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14317 3163 14334 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14317 3163 14334 3180
rect 13837 3163 13854 3180
rect 13957 3163 13974 3180
rect 13917 3163 13934 3180
rect 13877 3163 13894 3180
rect 13837 3163 13854 3180
rect 13917 3163 13934 3180
rect 13917 3163 13934 3180
rect 13877 3163 13894 3180
rect 13837 3163 13854 3180
rect 13837 3163 13854 3180
rect 13957 3163 13974 3180
rect 13877 3163 13894 3180
rect 13957 3163 13974 3180
rect 13957 3163 13974 3180
rect 13917 3163 13934 3180
rect 13757 3163 13774 3180
rect 13877 3163 13894 3180
rect 13797 3163 13814 3180
rect 13717 3163 13734 3180
rect 13797 3163 13814 3180
rect 13797 3163 13814 3180
rect 13757 3163 13774 3180
rect 13757 3163 13774 3180
rect 13717 3163 13734 3180
rect 13717 3163 13734 3180
rect 13717 3163 13734 3180
rect 13757 3163 13774 3180
rect 13797 3163 13814 3180
rect 14277 3163 14294 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 14357 3163 14374 3180
rect 13997 3163 14014 3180
rect 14277 3163 14294 3180
rect 12757 3163 12774 3180
rect 12757 3163 12774 3180
rect 12757 3163 12774 3180
rect 12757 3163 12774 3180
rect 12837 3163 12854 3180
rect 12837 3163 12854 3180
rect 12797 3163 12814 3180
rect 12797 3163 12814 3180
rect 13517 3163 13534 3180
rect 13597 3163 13614 3180
rect 13597 3163 13614 3180
rect 13677 3163 13694 3180
rect 13557 3163 13574 3180
rect 13637 3163 13654 3180
rect 12877 3163 12894 3180
rect 13477 3163 13494 3180
rect 13677 3163 13694 3180
rect 13637 3163 13654 3180
rect 13677 3163 13694 3180
rect 13597 3163 13614 3180
rect 13557 3163 13574 3180
rect 13517 3163 13534 3180
rect 13477 3163 13494 3180
rect 13557 3163 13574 3180
rect 13637 3163 13654 3180
rect 13677 3163 13694 3180
rect 13597 3163 13614 3180
rect 13637 3163 13654 3180
rect 13517 3163 13534 3180
rect 13557 3163 13574 3180
rect 13477 3163 13494 3180
rect 13517 3163 13534 3180
rect 13477 3163 13494 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 13237 3163 13254 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13397 3163 13414 3180
rect 13037 3163 13054 3180
rect 13397 3163 13414 3180
rect 13197 3163 13214 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13357 3163 13374 3180
rect 13117 3163 13134 3180
rect 13437 3163 13454 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13037 3163 13054 3180
rect 13277 3163 13294 3180
rect 12997 3163 13014 3180
rect 13277 3163 13294 3180
rect 12957 3163 12974 3180
rect 13237 3163 13254 3180
rect 13197 3163 13214 3180
rect 13277 3163 13294 3180
rect 12957 3163 12974 3180
rect 13237 3163 13254 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13437 3163 13454 3180
rect 12997 3163 13014 3180
rect 13277 3163 13294 3180
rect 12997 3163 13014 3180
rect 13437 3163 13454 3180
rect 13197 3163 13214 3180
rect 13117 3163 13134 3180
rect 13117 3163 13134 3180
rect 13037 3163 13054 3180
rect 13037 3163 13054 3180
rect 12837 3163 12854 3180
rect 13117 3163 13134 3180
rect 12957 3163 12974 3180
rect 13197 3163 13214 3180
rect 13077 3163 13094 3180
rect 13157 3163 13174 3180
rect 12997 3163 13014 3180
rect 13397 3163 13414 3180
rect 13357 3163 13374 3180
rect 12797 3163 12814 3180
rect 13357 3163 13374 3180
rect 13357 3163 13374 3180
rect 13237 3163 13254 3180
rect 13437 3163 13454 3180
rect 12877 3163 12894 3180
rect 12957 3163 12974 3180
rect 13397 3163 13414 3180
rect 12877 3163 12894 3180
rect 12877 3163 12894 3180
rect 12797 3163 12814 3180
rect 12837 3163 12854 3180
rect 12197 3163 12214 3180
rect 12557 3163 12574 3180
rect 12477 3163 12494 3180
rect 11997 3163 12014 3180
rect 12437 3163 12454 3180
rect 11997 3163 12014 3180
rect 12237 3163 12254 3180
rect 12437 3163 12454 3180
rect 11957 3163 11974 3180
rect 11957 3163 11974 3180
rect 12597 3163 12614 3180
rect 12357 3163 12374 3180
rect 11837 3163 11854 3180
rect 12277 3163 12294 3180
rect 12317 3163 12334 3180
rect 12557 3163 12574 3180
rect 12277 3163 12294 3180
rect 11837 3163 11854 3180
rect 12197 3163 12214 3180
rect 12317 3163 12334 3180
rect 12557 3163 12574 3180
rect 12237 3163 12254 3180
rect 11837 3163 11854 3180
rect 12077 3163 12094 3180
rect 12677 3163 12694 3180
rect 11957 3163 11974 3180
rect 12397 3163 12414 3180
rect 11997 3163 12014 3180
rect 12397 3163 12414 3180
rect 12317 3163 12334 3180
rect 12117 3163 12134 3180
rect 12237 3163 12254 3180
rect 12197 3163 12214 3180
rect 11877 3163 11894 3180
rect 11997 3163 12014 3180
rect 12677 3163 12694 3180
rect 11837 3163 11854 3180
rect 11877 3163 11894 3180
rect 11917 3163 11934 3180
rect 12397 3163 12414 3180
rect 12277 3163 12294 3180
rect 12037 3163 12054 3180
rect 12037 3163 12054 3180
rect 12357 3163 12374 3180
rect 12717 3163 12734 3180
rect 12677 3163 12694 3180
rect 12157 3163 12174 3180
rect 12197 3163 12214 3180
rect 12117 3163 12134 3180
rect 12397 3163 12414 3180
rect 12117 3163 12134 3180
rect 12157 3163 12174 3180
rect 12717 3163 12734 3180
rect 12597 3163 12614 3180
rect 11917 3163 11934 3180
rect 12157 3163 12174 3180
rect 12237 3163 12254 3180
rect 12077 3163 12094 3180
rect 11957 3163 11974 3180
rect 12717 3163 12734 3180
rect 12117 3163 12134 3180
rect 12517 3163 12534 3180
rect 12277 3163 12294 3180
rect 12077 3163 12094 3180
rect 11917 3163 11934 3180
rect 12637 3163 12654 3180
rect 11917 3163 11934 3180
rect 12677 3163 12694 3180
rect 12557 3163 12574 3180
rect 12437 3163 12454 3180
rect 12077 3163 12094 3180
rect 12517 3163 12534 3180
rect 12037 3163 12054 3180
rect 12717 3163 12734 3180
rect 11877 3163 11894 3180
rect 12637 3163 12654 3180
rect 12477 3163 12494 3180
rect 12437 3163 12454 3180
rect 11877 3163 11894 3180
rect 12037 3163 12054 3180
rect 12477 3163 12494 3180
rect 12637 3163 12654 3180
rect 12357 3163 12374 3180
rect 12517 3163 12534 3180
rect 12597 3163 12614 3180
rect 12637 3163 12654 3180
rect 12157 3163 12174 3180
rect 12317 3163 12334 3180
rect 12517 3163 12534 3180
rect 12597 3163 12614 3180
rect 12357 3163 12374 3180
rect 12477 3163 12494 3180
rect 10836 3163 10853 3180
rect 10836 3163 10853 3180
rect 10836 3163 10853 3180
rect 10836 3163 10853 3180
rect 11757 3163 11774 3180
rect 11717 3163 11734 3180
rect 11597 3163 11614 3180
rect 11317 3163 11334 3180
rect 11357 3163 11374 3180
rect 11717 3163 11734 3180
rect 11357 3163 11374 3180
rect 11517 3163 11534 3180
rect 11557 3163 11574 3180
rect 11597 3163 11614 3180
rect 11477 3163 11494 3180
rect 11597 3163 11614 3180
rect 11677 3163 11694 3180
rect 11757 3163 11774 3180
rect 11196 3163 11213 3180
rect 11477 3163 11494 3180
rect 11517 3163 11534 3180
rect 11036 3163 11053 3180
rect 11317 3163 11334 3180
rect 11196 3163 11213 3180
rect 11677 3163 11694 3180
rect 11116 3163 11133 3180
rect 10996 3163 11013 3180
rect 11076 3163 11093 3180
rect 10956 3163 10973 3180
rect 11276 3163 11293 3180
rect 11236 3163 11253 3180
rect 11196 3163 11213 3180
rect 11276 3163 11293 3180
rect 11156 3163 11173 3180
rect 11116 3163 11133 3180
rect 11076 3163 11093 3180
rect 11036 3163 11053 3180
rect 10996 3163 11013 3180
rect 10956 3163 10973 3180
rect 10916 3163 10933 3180
rect 10876 3163 10893 3180
rect 11116 3163 11133 3180
rect 11076 3163 11093 3180
rect 11036 3163 11053 3180
rect 11076 3163 11093 3180
rect 10956 3163 10973 3180
rect 11276 3163 11293 3180
rect 11276 3163 11293 3180
rect 11156 3163 11173 3180
rect 11156 3163 11173 3180
rect 10916 3163 10933 3180
rect 10876 3163 10893 3180
rect 11317 3163 11334 3180
rect 10996 3163 11013 3180
rect 11196 3163 11213 3180
rect 11116 3163 11133 3180
rect 11397 3163 11414 3180
rect 11036 3163 11053 3180
rect 10956 3163 10973 3180
rect 10876 3163 10893 3180
rect 11397 3163 11414 3180
rect 10996 3163 11013 3180
rect 11236 3163 11253 3180
rect 11236 3163 11253 3180
rect 11637 3163 11654 3180
rect 10916 3163 10933 3180
rect 10916 3163 10933 3180
rect 11397 3163 11414 3180
rect 11236 3163 11253 3180
rect 10876 3163 10893 3180
rect 11156 3163 11173 3180
rect 11717 3163 11734 3180
rect 11557 3163 11574 3180
rect 11637 3163 11654 3180
rect 11597 3163 11614 3180
rect 11477 3163 11494 3180
rect 11637 3163 11654 3180
rect 11757 3163 11774 3180
rect 11557 3163 11574 3180
rect 11357 3163 11374 3180
rect 11437 3163 11454 3180
rect 11677 3163 11694 3180
rect 11397 3163 11414 3180
rect 11717 3163 11734 3180
rect 11517 3163 11534 3180
rect 11637 3163 11654 3180
rect 11357 3163 11374 3180
rect 11557 3163 11574 3180
rect 11677 3163 11694 3180
rect 11317 3163 11334 3180
rect 11477 3163 11494 3180
rect 11437 3163 11454 3180
rect 11517 3163 11534 3180
rect 11437 3163 11454 3180
rect 11757 3163 11774 3180
rect 11437 3163 11454 3180
rect 10196 3163 10213 3180
rect 9916 3163 9933 3180
rect 10756 3163 10773 3180
rect 10676 3163 10693 3180
rect 10236 3163 10253 3180
rect 9956 3163 9973 3180
rect 10276 3163 10293 3180
rect 9996 3163 10013 3180
rect 10476 3163 10493 3180
rect 10436 3163 10453 3180
rect 10116 3163 10133 3180
rect 10316 3163 10333 3180
rect 9956 3163 9973 3180
rect 10556 3163 10573 3180
rect 10396 3163 10413 3180
rect 10716 3163 10733 3180
rect 10116 3163 10133 3180
rect 10716 3163 10733 3180
rect 10516 3163 10533 3180
rect 10156 3163 10173 3180
rect 10716 3163 10733 3180
rect 10756 3163 10773 3180
rect 10476 3163 10493 3180
rect 10356 3163 10373 3180
rect 10556 3163 10573 3180
rect 10756 3163 10773 3180
rect 10316 3163 10333 3180
rect 10436 3163 10453 3180
rect 10396 3163 10413 3180
rect 10196 3163 10213 3180
rect 10436 3163 10453 3180
rect 10356 3163 10373 3180
rect 9916 3163 9933 3180
rect 10236 3163 10253 3180
rect 10116 3163 10133 3180
rect 10596 3163 10613 3180
rect 10676 3163 10693 3180
rect 10396 3163 10413 3180
rect 10796 3163 10813 3180
rect 10276 3163 10293 3180
rect 10076 3163 10093 3180
rect 10276 3163 10293 3180
rect 10156 3163 10173 3180
rect 10636 3163 10653 3180
rect 9956 3163 9973 3180
rect 10396 3163 10413 3180
rect 10156 3163 10173 3180
rect 10556 3163 10573 3180
rect 10036 3163 10053 3180
rect 10516 3163 10533 3180
rect 10076 3163 10093 3180
rect 10636 3163 10653 3180
rect 10116 3163 10133 3180
rect 10676 3163 10693 3180
rect 10236 3163 10253 3180
rect 10196 3163 10213 3180
rect 10516 3163 10533 3180
rect 10796 3163 10813 3180
rect 10676 3163 10693 3180
rect 10036 3163 10053 3180
rect 10716 3163 10733 3180
rect 9916 3163 9933 3180
rect 10596 3163 10613 3180
rect 10196 3163 10213 3180
rect 10516 3163 10533 3180
rect 9916 3163 9933 3180
rect 10636 3163 10653 3180
rect 9996 3163 10013 3180
rect 10276 3163 10293 3180
rect 9996 3163 10013 3180
rect 10036 3163 10053 3180
rect 10316 3163 10333 3180
rect 10476 3163 10493 3180
rect 10076 3163 10093 3180
rect 10436 3163 10453 3180
rect 10036 3163 10053 3180
rect 9996 3163 10013 3180
rect 10636 3163 10653 3180
rect 10476 3163 10493 3180
rect 10796 3163 10813 3180
rect 10316 3163 10333 3180
rect 10156 3163 10173 3180
rect 10356 3163 10373 3180
rect 10596 3163 10613 3180
rect 10796 3163 10813 3180
rect 10356 3163 10373 3180
rect 10076 3163 10093 3180
rect 10596 3163 10613 3180
rect 10556 3163 10573 3180
rect 10756 3163 10773 3180
rect 10236 3163 10253 3180
rect 9956 3163 9973 3180
rect 12001 2394 12018 2411
rect 12001 2394 12018 2411
rect 9876 3163 9893 3180
rect 9836 3163 9853 3180
rect 9636 3163 9653 3180
rect 9836 3163 9853 3180
rect 9876 3163 9893 3180
rect 9636 3163 9653 3180
rect 9636 3163 9653 3180
rect 9676 3163 9693 3180
rect 9716 3163 9733 3180
rect 9676 3163 9693 3180
rect 9756 3163 9773 3180
rect 9836 3163 9853 3180
rect 9636 3163 9653 3180
rect 9716 3163 9733 3180
rect 9756 3163 9773 3180
rect 9756 3163 9773 3180
rect 9796 3163 9813 3180
rect 9796 3163 9813 3180
rect 9716 3163 9733 3180
rect 9756 3163 9773 3180
rect 9796 3163 9813 3180
rect 9716 3163 9733 3180
rect 9876 3163 9893 3180
rect 9836 3163 9853 3180
rect 9796 3163 9813 3180
rect 9876 3163 9893 3180
rect 9676 3163 9693 3180
rect 9676 3163 9693 3180
rect 10641 2394 10658 2411
rect 10041 2394 10058 2411
rect 10721 2394 10738 2411
rect 10601 2394 10618 2411
rect 9801 2394 9818 2411
rect 9881 2394 9898 2411
rect 10521 2394 10538 2411
rect 10721 2394 10738 2411
rect 10201 2394 10218 2411
rect 10201 2394 10218 2411
rect 9681 2394 9698 2411
rect 9641 2394 9658 2411
rect 10441 2394 10458 2411
rect 10281 2394 10298 2411
rect 10241 2394 10258 2411
rect 10561 2394 10578 2411
rect 10121 2394 10138 2411
rect 10641 2394 10658 2411
rect 9641 2394 9658 2411
rect 10001 2394 10018 2411
rect 10281 2394 10298 2411
rect 9681 2394 9698 2411
rect 9841 2394 9858 2411
rect 10681 2394 10698 2411
rect 10081 2394 10098 2411
rect 10761 2394 10778 2411
rect 10601 2394 10618 2411
rect 9841 2394 9858 2411
rect 9801 2394 9818 2411
rect 10801 2394 10818 2411
rect 10761 2394 10778 2411
rect 10161 2394 10178 2411
rect 9721 2394 9738 2411
rect 10481 2394 10498 2411
rect 10321 2394 10338 2411
rect 9761 2394 9778 2411
rect 10081 2394 10098 2411
rect 10001 2394 10018 2411
rect 10481 2394 10498 2411
rect 10441 2394 10458 2411
rect 9721 2394 9738 2411
rect 10041 2394 10058 2411
rect 9921 2394 9938 2411
rect 9961 2394 9978 2411
rect 10241 2394 10258 2411
rect 10361 2394 10378 2411
rect 9961 2394 9978 2411
rect 9761 2394 9778 2411
rect 9881 2394 9898 2411
rect 10401 2394 10418 2411
rect 10361 2394 10378 2411
rect 10121 2394 10138 2411
rect 10521 2394 10538 2411
rect 9921 2394 9938 2411
rect 10401 2394 10418 2411
rect 10801 2394 10818 2411
rect 10561 2394 10578 2411
rect 10681 2394 10698 2411
rect 10321 2394 10338 2411
rect 10161 2394 10178 2411
rect 11121 2394 11138 2411
rect 11881 2394 11898 2411
rect 11601 2394 11618 2411
rect 11961 2394 11978 2411
rect 11041 2394 11058 2411
rect 11161 2394 11178 2411
rect 11561 2394 11578 2411
rect 11081 2394 11098 2411
rect 11001 2394 11018 2411
rect 11321 2394 11338 2411
rect 11041 2394 11058 2411
rect 11881 2394 11898 2411
rect 11721 2394 11738 2411
rect 11841 2394 11858 2411
rect 11841 2394 11858 2411
rect 11921 2394 11938 2411
rect 11801 2394 11818 2411
rect 11961 2394 11978 2411
rect 11201 2394 11218 2411
rect 11761 2394 11778 2411
rect 10961 2394 10978 2411
rect 11801 2394 11818 2411
rect 11641 2394 11658 2411
rect 11641 2394 11658 2411
rect 11721 2394 11738 2411
rect 11481 2394 11498 2411
rect 11161 2394 11178 2411
rect 10921 2394 10938 2411
rect 11681 2394 11698 2411
rect 11601 2394 11618 2411
rect 11681 2394 11698 2411
rect 10961 2394 10978 2411
rect 11761 2394 11778 2411
rect 11441 2394 11458 2411
rect 11561 2394 11578 2411
rect 11281 2394 11298 2411
rect 11521 2394 11538 2411
rect 10841 2394 10858 2411
rect 11401 2394 11418 2411
rect 11481 2394 11498 2411
rect 10921 2394 10938 2411
rect 11441 2394 11458 2411
rect 11121 2394 11138 2411
rect 11001 2394 11018 2411
rect 11401 2394 11418 2411
rect 11361 2394 11378 2411
rect 10881 2394 10898 2411
rect 11361 2394 11378 2411
rect 11521 2394 11538 2411
rect 11321 2394 11338 2411
rect 11281 2394 11298 2411
rect 11241 2394 11258 2411
rect 11921 2394 11938 2411
rect 11241 2394 11258 2411
rect 10841 2394 10858 2411
rect 11201 2394 11218 2411
rect 11081 2394 11098 2411
rect 10881 2394 10898 2411
rect 13201 2394 13218 2411
rect 13201 2394 13218 2411
rect 12361 2394 12378 2411
rect 12321 2394 12338 2411
rect 12241 2394 12258 2411
rect 12201 2394 12218 2411
rect 12081 2394 12098 2411
rect 12281 2394 12298 2411
rect 12281 2394 12298 2411
rect 12041 2394 12058 2411
rect 12041 2394 12058 2411
rect 12321 2394 12338 2411
rect 12521 2394 12538 2411
rect 12561 2394 12578 2411
rect 12161 2394 12178 2411
rect 12161 2394 12178 2411
rect 12081 2394 12098 2411
rect 12121 2394 12138 2411
rect 12401 2394 12418 2411
rect 12601 2394 12618 2411
rect 13121 2394 13138 2411
rect 13081 2394 13098 2411
rect 13041 2394 13058 2411
rect 13001 2394 13018 2411
rect 12961 2394 12978 2411
rect 12921 2394 12938 2411
rect 12881 2394 12898 2411
rect 12841 2394 12858 2411
rect 12801 2394 12818 2411
rect 12761 2394 12778 2411
rect 12721 2394 12738 2411
rect 12401 2394 12418 2411
rect 13161 2394 13178 2411
rect 13121 2394 13138 2411
rect 13081 2394 13098 2411
rect 13041 2394 13058 2411
rect 13001 2394 13018 2411
rect 12961 2394 12978 2411
rect 12921 2394 12938 2411
rect 12881 2394 12898 2411
rect 12841 2394 12858 2411
rect 12801 2394 12818 2411
rect 12761 2394 12778 2411
rect 12721 2394 12738 2411
rect 12681 2394 12698 2411
rect 13161 2394 13178 2411
rect 12361 2394 12378 2411
rect 12481 2394 12498 2411
rect 12681 2394 12698 2411
rect 12641 2394 12658 2411
rect 12601 2394 12618 2411
rect 12561 2394 12578 2411
rect 12521 2394 12538 2411
rect 12481 2394 12498 2411
rect 12241 2394 12258 2411
rect 12441 2394 12458 2411
rect 12441 2394 12458 2411
rect 12121 2394 12138 2411
rect 12641 2394 12658 2411
rect 12201 2394 12218 2411
rect 13241 2394 13258 2411
rect 14242 2394 14259 2411
rect 13802 2394 13819 2411
rect 14202 2394 14219 2411
rect 14322 2394 14339 2411
rect 14002 2394 14019 2411
rect 14242 2394 14259 2411
rect 13962 2394 13979 2411
rect 13842 2394 13859 2411
rect 13761 2394 13778 2411
rect 13641 2394 13658 2411
rect 14202 2394 14219 2411
rect 13721 2394 13738 2411
rect 14162 2394 14179 2411
rect 13601 2394 13618 2411
rect 13882 2394 13899 2411
rect 13561 2394 13578 2411
rect 13521 2394 13538 2411
rect 13481 2394 13498 2411
rect 13441 2394 13458 2411
rect 14042 2394 14059 2411
rect 14082 2394 14099 2411
rect 13401 2394 13418 2411
rect 13361 2394 13378 2411
rect 13321 2394 13338 2411
rect 14362 2394 14379 2411
rect 13842 2394 13859 2411
rect 13882 2394 13899 2411
rect 14002 2394 14019 2411
rect 13802 2394 13819 2411
rect 14362 2394 14379 2411
rect 14122 2394 14139 2411
rect 14322 2394 14339 2411
rect 13922 2394 13939 2411
rect 14282 2394 14299 2411
rect 13962 2394 13979 2411
rect 14122 2394 14139 2411
rect 13922 2394 13939 2411
rect 14082 2394 14099 2411
rect 14042 2394 14059 2411
rect 13641 2394 13658 2411
rect 13601 2394 13618 2411
rect 14162 2394 14179 2411
rect 13681 2394 13698 2411
rect 13561 2394 13578 2411
rect 13521 2394 13538 2411
rect 14282 2394 14299 2411
rect 13721 2394 13738 2411
rect 13681 2394 13698 2411
rect 13281 2394 13298 2411
rect 13241 2394 13258 2411
rect 13481 2394 13498 2411
rect 13441 2394 13458 2411
rect 13401 2394 13418 2411
rect 13361 2394 13378 2411
rect 13321 2394 13338 2411
rect 13761 2394 13778 2411
rect 13281 2394 13298 2411
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 15077 3163 15094 3180
rect 15117 3163 15134 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 14717 3163 14734 3180
rect 14997 3163 15014 3180
rect 14797 3163 14814 3180
rect 14997 3163 15014 3180
rect 14677 3163 14694 3180
rect 14957 3163 14974 3180
rect 14877 3163 14894 3180
rect 14997 3163 15014 3180
rect 14917 3163 14934 3180
rect 14917 3163 14934 3180
rect 14957 3163 14974 3180
rect 14917 3163 14934 3180
rect 14877 3163 14894 3180
rect 14877 3163 14894 3180
rect 14837 3163 14854 3180
rect 14837 3163 14854 3180
rect 14837 3163 14854 3180
rect 15037 3163 15054 3180
rect 14797 3163 14814 3180
rect 14797 3163 14814 3180
rect 14917 3163 14934 3180
rect 14757 3163 14774 3180
rect 14757 3163 14774 3180
rect 14757 3163 14774 3180
rect 15037 3163 15054 3180
rect 14717 3163 14734 3180
rect 14717 3163 14734 3180
rect 14877 3163 14894 3180
rect 15037 3163 15054 3180
rect 14677 3163 14694 3180
rect 14677 3163 14694 3180
rect 15037 3163 15054 3180
rect 14957 3163 14974 3180
rect 14837 3163 14854 3180
rect 14677 3163 14694 3180
rect 14797 3163 14814 3180
rect 14717 3163 14734 3180
rect 14997 3163 15014 3180
rect 14957 3163 14974 3180
rect 14757 3163 14774 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 15077 3163 15094 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 15077 3163 15094 3180
rect 15077 3163 15094 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15077 3163 15094 3180
rect 14397 3163 14414 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 14557 3163 14574 3180
rect 14397 3163 14414 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 14477 3163 14494 3180
rect 14437 3163 14454 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 14517 3163 14534 3180
rect 14477 3163 14494 3180
rect 14437 3163 14454 3180
rect 15077 3163 15094 3180
rect 15077 3163 15094 3180
rect 15517 3163 15534 3180
rect 14517 3163 14534 3180
rect 15477 3163 15494 3180
rect 14477 3163 14494 3180
rect 14517 3163 14534 3180
rect 14477 3163 14494 3180
rect 14597 3163 14614 3180
rect 14437 3163 14454 3180
rect 14517 3163 14534 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15077 3163 15094 3180
rect 15117 3163 15134 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 14717 3163 14734 3180
rect 14637 3163 14654 3180
rect 14637 3163 14654 3180
rect 14637 3163 14654 3180
rect 14597 3163 14614 3180
rect 14557 3163 14574 3180
rect 14637 3163 14654 3180
rect 14557 3163 14574 3180
rect 14557 3163 14574 3180
rect 14597 3163 14614 3180
rect 14597 3163 14614 3180
rect 14997 3163 15014 3180
rect 14797 3163 14814 3180
rect 14437 3163 14454 3180
rect 14997 3163 15014 3180
rect 14677 3163 14694 3180
rect 14957 3163 14974 3180
rect 14877 3163 14894 3180
rect 14997 3163 15014 3180
rect 14557 3163 14574 3180
rect 14917 3163 14934 3180
rect 14917 3163 14934 3180
rect 14957 3163 14974 3180
rect 14917 3163 14934 3180
rect 14877 3163 14894 3180
rect 14397 3163 14414 3180
rect 14877 3163 14894 3180
rect 14597 3163 14614 3180
rect 14837 3163 14854 3180
rect 14837 3163 14854 3180
rect 14397 3163 14414 3180
rect 14837 3163 14854 3180
rect 14557 3163 14574 3180
rect 15037 3163 15054 3180
rect 14797 3163 14814 3180
rect 14797 3163 14814 3180
rect 14917 3163 14934 3180
rect 14757 3163 14774 3180
rect 14757 3163 14774 3180
rect 14757 3163 14774 3180
rect 14637 3163 14654 3180
rect 15037 3163 15054 3180
rect 14717 3163 14734 3180
rect 14717 3163 14734 3180
rect 14877 3163 14894 3180
rect 15037 3163 15054 3180
rect 14677 3163 14694 3180
rect 14677 3163 14694 3180
rect 15037 3163 15054 3180
rect 14637 3163 14654 3180
rect 14957 3163 14974 3180
rect 14837 3163 14854 3180
rect 14597 3163 14614 3180
rect 14557 3163 14574 3180
rect 14677 3163 14694 3180
rect 14797 3163 14814 3180
rect 14717 3163 14734 3180
rect 14637 3163 14654 3180
rect 14597 3163 14614 3180
rect 14557 3163 14574 3180
rect 14637 3163 14654 3180
rect 14997 3163 15014 3180
rect 14957 3163 14974 3180
rect 14757 3163 14774 3180
rect 14597 3163 14614 3180
rect 16762 2394 16779 2411
rect 16762 2394 16779 2411
rect 14437 3163 14454 3180
rect 14397 3163 14414 3180
rect 14397 3163 14414 3180
rect 14397 3163 14414 3180
rect 14397 3163 14414 3180
rect 14477 3163 14494 3180
rect 14437 3163 14454 3180
rect 14517 3163 14534 3180
rect 14477 3163 14494 3180
rect 14437 3163 14454 3180
rect 14517 3163 14534 3180
rect 14477 3163 14494 3180
rect 14517 3163 14534 3180
rect 14477 3163 14494 3180
rect 14437 3163 14454 3180
rect 14517 3163 14534 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17477 3163 17494 3180
rect 17717 3163 17734 3180
rect 17717 3163 17734 3180
rect 17517 3163 17534 3180
rect 17637 3163 17654 3180
rect 17477 3163 17494 3180
rect 17677 3163 17694 3180
rect 17637 3163 17654 3180
rect 17597 3163 17614 3180
rect 17597 3163 17614 3180
rect 17557 3163 17574 3180
rect 17517 3163 17534 3180
rect 17597 3163 17614 3180
rect 17557 3163 17574 3180
rect 17637 3163 17654 3180
rect 17477 3163 17494 3180
rect 17597 3163 17614 3180
rect 17517 3163 17534 3180
rect 17517 3163 17534 3180
rect 17477 3163 17494 3180
rect 17717 3163 17734 3180
rect 17677 3163 17694 3180
rect 17677 3163 17694 3180
rect 17677 3163 17694 3180
rect 17557 3163 17574 3180
rect 17557 3163 17574 3180
rect 17637 3163 17654 3180
rect 17477 3163 17494 3180
rect 17717 3163 17734 3180
rect 17717 3163 17734 3180
rect 17557 3163 17574 3180
rect 17717 3163 17734 3180
rect 17517 3163 17534 3180
rect 17637 3163 17654 3180
rect 17477 3163 17494 3180
rect 17677 3163 17694 3180
rect 17637 3163 17654 3180
rect 17597 3163 17614 3180
rect 17597 3163 17614 3180
rect 17557 3163 17574 3180
rect 17517 3163 17534 3180
rect 17597 3163 17614 3180
rect 17557 3163 17574 3180
rect 17637 3163 17654 3180
rect 17477 3163 17494 3180
rect 17597 3163 17614 3180
rect 17517 3163 17534 3180
rect 17517 3163 17534 3180
rect 17477 3163 17494 3180
rect 17717 3163 17734 3180
rect 17677 3163 17694 3180
rect 17677 3163 17694 3180
rect 17677 3163 17694 3180
rect 17557 3163 17574 3180
rect 17717 3163 17734 3180
rect 17637 3163 17654 3180
rect 17357 3163 17374 3180
rect 17237 3163 17254 3180
rect 17357 3163 17374 3180
rect 17437 3163 17454 3180
rect 17437 3163 17454 3180
rect 17357 3163 17374 3180
rect 17357 3163 17374 3180
rect 17437 3163 17454 3180
rect 17277 3163 17294 3180
rect 17437 3163 17454 3180
rect 17397 3163 17414 3180
rect 17437 3163 17454 3180
rect 17357 3163 17374 3180
rect 17397 3163 17414 3180
rect 17317 3163 17334 3180
rect 17277 3163 17294 3180
rect 17277 3163 17294 3180
rect 17317 3163 17334 3180
rect 17317 3163 17334 3180
rect 17397 3163 17414 3180
rect 17277 3163 17294 3180
rect 17237 3163 17254 3180
rect 17397 3163 17414 3180
rect 17237 3163 17254 3180
rect 17237 3163 17254 3180
rect 17317 3163 17334 3180
rect 17237 3163 17254 3180
rect 17317 3163 17334 3180
rect 17397 3163 17414 3180
rect 17437 3163 17454 3180
rect 17437 3163 17454 3180
rect 17357 3163 17374 3180
rect 17357 3163 17374 3180
rect 17437 3163 17454 3180
rect 17277 3163 17294 3180
rect 17237 3163 17254 3180
rect 17397 3163 17414 3180
rect 17277 3163 17294 3180
rect 17317 3163 17334 3180
rect 17317 3163 17334 3180
rect 17397 3163 17414 3180
rect 17237 3163 17254 3180
rect 17357 3163 17374 3180
rect 17277 3163 17294 3180
rect 17277 3163 17294 3180
rect 17237 3163 17254 3180
rect 17397 3163 17414 3180
rect 17317 3163 17334 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 17117 3163 17134 3180
rect 17037 3163 17054 3180
rect 17117 3163 17134 3180
rect 17117 3163 17134 3180
rect 16997 3163 17014 3180
rect 17037 3163 17054 3180
rect 17077 3163 17094 3180
rect 17077 3163 17094 3180
rect 16957 3163 16974 3180
rect 16997 3163 17014 3180
rect 16957 3163 16974 3180
rect 17077 3163 17094 3180
rect 17157 3163 17174 3180
rect 17077 3163 17094 3180
rect 17037 3163 17054 3180
rect 17077 3163 17094 3180
rect 17157 3163 17174 3180
rect 17157 3163 17174 3180
rect 17157 3163 17174 3180
rect 17117 3163 17134 3180
rect 17157 3163 17174 3180
rect 16997 3163 17014 3180
rect 17117 3163 17134 3180
rect 16997 3163 17014 3180
rect 17117 3163 17134 3180
rect 16957 3163 16974 3180
rect 17077 3163 17094 3180
rect 17117 3163 17134 3180
rect 17037 3163 17054 3180
rect 16957 3163 16974 3180
rect 17157 3163 17174 3180
rect 17037 3163 17054 3180
rect 16957 3163 16974 3180
rect 17037 3163 17054 3180
rect 16997 3163 17014 3180
rect 16997 3163 17014 3180
rect 16997 3163 17014 3180
rect 17157 3163 17174 3180
rect 17077 3163 17094 3180
rect 16957 3163 16974 3180
rect 17077 3163 17094 3180
rect 17037 3163 17054 3180
rect 16957 3163 16974 3180
rect 17037 3163 17054 3180
rect 16997 3163 17014 3180
rect 16957 3163 16974 3180
rect 17117 3163 17134 3180
rect 17157 3163 17174 3180
rect 16877 3163 16894 3180
rect 16677 3163 16694 3180
rect 16757 3163 16774 3180
rect 16677 3163 16694 3180
rect 16797 3163 16814 3180
rect 16837 3163 16854 3180
rect 16877 3163 16894 3180
rect 16877 3163 16894 3180
rect 16757 3163 16774 3180
rect 16877 3163 16894 3180
rect 16877 3163 16894 3180
rect 16837 3163 16854 3180
rect 16797 3163 16814 3180
rect 16837 3163 16854 3180
rect 16877 3163 16894 3180
rect 16717 3163 16734 3180
rect 16837 3163 16854 3180
rect 16837 3163 16854 3180
rect 16717 3163 16734 3180
rect 16797 3163 16814 3180
rect 16757 3163 16774 3180
rect 16757 3163 16774 3180
rect 16677 3163 16694 3180
rect 16677 3163 16694 3180
rect 16757 3163 16774 3180
rect 16797 3163 16814 3180
rect 16677 3163 16694 3180
rect 16677 3163 16694 3180
rect 16877 3163 16894 3180
rect 16757 3163 16774 3180
rect 16837 3163 16854 3180
rect 16717 3163 16734 3180
rect 16837 3163 16854 3180
rect 16877 3163 16894 3180
rect 16717 3163 16734 3180
rect 16757 3163 16774 3180
rect 16717 3163 16734 3180
rect 16677 3163 16694 3180
rect 16797 3163 16814 3180
rect 16717 3163 16734 3180
rect 16797 3163 16814 3180
rect 16837 3163 16854 3180
rect 16797 3163 16814 3180
rect 16757 3163 16774 3180
rect 16717 3163 16734 3180
rect 16677 3163 16694 3180
rect 16717 3163 16734 3180
rect 16797 3163 16814 3180
rect 16597 3163 16614 3180
rect 16437 3163 16454 3180
rect 16517 3163 16534 3180
rect 16557 3163 16574 3180
rect 16397 3163 16414 3180
rect 16557 3163 16574 3180
rect 16477 3163 16494 3180
rect 16397 3163 16414 3180
rect 16597 3163 16614 3180
rect 16397 3163 16414 3180
rect 16597 3163 16614 3180
rect 16477 3163 16494 3180
rect 16517 3163 16534 3180
rect 16517 3163 16534 3180
rect 16557 3163 16574 3180
rect 16397 3163 16414 3180
rect 16597 3163 16614 3180
rect 16437 3163 16454 3180
rect 16477 3163 16494 3180
rect 16437 3163 16454 3180
rect 16517 3163 16534 3180
rect 16437 3163 16454 3180
rect 16437 3163 16454 3180
rect 16557 3163 16574 3180
rect 16557 3163 16574 3180
rect 16517 3163 16534 3180
rect 16437 3163 16454 3180
rect 16397 3163 16414 3180
rect 16597 3163 16614 3180
rect 16557 3163 16574 3180
rect 16597 3163 16614 3180
rect 16517 3163 16534 3180
rect 16397 3163 16414 3180
rect 16597 3163 16614 3180
rect 16477 3163 16494 3180
rect 16477 3163 16494 3180
rect 16517 3163 16534 3180
rect 16437 3163 16454 3180
rect 16557 3163 16574 3180
rect 16477 3163 16494 3180
rect 16437 3163 16454 3180
rect 16477 3163 16494 3180
rect 16597 3163 16614 3180
rect 16397 3163 16414 3180
rect 16477 3163 16494 3180
rect 16557 3163 16574 3180
rect 16517 3163 16534 3180
rect 16397 3163 16414 3180
rect 16317 3163 16334 3180
rect 16197 3163 16214 3180
rect 16357 3163 16374 3180
rect 16277 3163 16294 3180
rect 16277 3163 16294 3180
rect 16117 3163 16134 3180
rect 16157 3163 16174 3180
rect 16237 3163 16254 3180
rect 16157 3163 16174 3180
rect 16117 3163 16134 3180
rect 16197 3163 16214 3180
rect 16197 3163 16214 3180
rect 16317 3163 16334 3180
rect 16277 3163 16294 3180
rect 16237 3163 16254 3180
rect 16157 3163 16174 3180
rect 16157 3163 16174 3180
rect 16197 3163 16214 3180
rect 16157 3163 16174 3180
rect 16357 3163 16374 3180
rect 16237 3163 16254 3180
rect 16237 3163 16254 3180
rect 16317 3163 16334 3180
rect 16157 3163 16174 3180
rect 16357 3163 16374 3180
rect 16237 3163 16254 3180
rect 16357 3163 16374 3180
rect 16317 3163 16334 3180
rect 16277 3163 16294 3180
rect 16317 3163 16334 3180
rect 16117 3163 16134 3180
rect 16317 3163 16334 3180
rect 16357 3163 16374 3180
rect 16117 3163 16134 3180
rect 16117 3163 16134 3180
rect 16317 3163 16334 3180
rect 16117 3163 16134 3180
rect 16157 3163 16174 3180
rect 16237 3163 16254 3180
rect 16157 3163 16174 3180
rect 16197 3163 16214 3180
rect 16117 3163 16134 3180
rect 16277 3163 16294 3180
rect 16277 3163 16294 3180
rect 16357 3163 16374 3180
rect 16197 3163 16214 3180
rect 16357 3163 16374 3180
rect 16277 3163 16294 3180
rect 16197 3163 16214 3180
rect 16237 3163 16254 3180
rect 16237 3163 16254 3180
rect 16357 3163 16374 3180
rect 16117 3163 16134 3180
rect 16197 3163 16214 3180
rect 16317 3163 16334 3180
rect 16277 3163 16294 3180
rect 16037 3163 16054 3180
rect 15997 3163 16014 3180
rect 15957 3163 15974 3180
rect 15997 3163 16014 3180
rect 15877 3163 15894 3180
rect 15837 3163 15854 3180
rect 15877 3163 15894 3180
rect 15877 3163 15894 3180
rect 15837 3163 15854 3180
rect 15957 3163 15974 3180
rect 16077 3163 16094 3180
rect 15837 3163 15854 3180
rect 15917 3163 15934 3180
rect 15917 3163 15934 3180
rect 16037 3163 16054 3180
rect 15877 3163 15894 3180
rect 15957 3163 15974 3180
rect 15997 3163 16014 3180
rect 16037 3163 16054 3180
rect 16077 3163 16094 3180
rect 15957 3163 15974 3180
rect 16077 3163 16094 3180
rect 15837 3163 15854 3180
rect 15997 3163 16014 3180
rect 16077 3163 16094 3180
rect 15877 3163 15894 3180
rect 16037 3163 16054 3180
rect 15877 3163 15894 3180
rect 15917 3163 15934 3180
rect 15837 3163 15854 3180
rect 15917 3163 15934 3180
rect 15997 3163 16014 3180
rect 15837 3163 15854 3180
rect 15957 3163 15974 3180
rect 16077 3163 16094 3180
rect 15877 3163 15894 3180
rect 15837 3163 15854 3180
rect 15997 3163 16014 3180
rect 15957 3163 15974 3180
rect 15917 3163 15934 3180
rect 15877 3163 15894 3180
rect 16037 3163 16054 3180
rect 15917 3163 15934 3180
rect 16037 3163 16054 3180
rect 15997 3163 16014 3180
rect 15957 3163 15974 3180
rect 16077 3163 16094 3180
rect 16037 3163 16054 3180
rect 15917 3163 15934 3180
rect 15997 3163 16014 3180
rect 15837 3163 15854 3180
rect 16077 3163 16094 3180
rect 16077 3163 16094 3180
rect 15917 3163 15934 3180
rect 16037 3163 16054 3180
rect 15957 3163 15974 3180
rect 15757 3163 15774 3180
rect 15557 3163 15574 3180
rect 15637 3163 15654 3180
rect 15557 3163 15574 3180
rect 15717 3163 15734 3180
rect 15797 3163 15814 3180
rect 15677 3163 15694 3180
rect 15757 3163 15774 3180
rect 15717 3163 15734 3180
rect 15797 3163 15814 3180
rect 15557 3163 15574 3180
rect 15557 3163 15574 3180
rect 15637 3163 15654 3180
rect 15597 3163 15614 3180
rect 15757 3163 15774 3180
rect 15557 3163 15574 3180
rect 15797 3163 15814 3180
rect 15797 3163 15814 3180
rect 15677 3163 15694 3180
rect 15637 3163 15654 3180
rect 15597 3163 15614 3180
rect 15757 3163 15774 3180
rect 15797 3163 15814 3180
rect 15717 3163 15734 3180
rect 15677 3163 15694 3180
rect 15717 3163 15734 3180
rect 15677 3163 15694 3180
rect 15597 3163 15614 3180
rect 15597 3163 15614 3180
rect 15797 3163 15814 3180
rect 15717 3163 15734 3180
rect 15757 3163 15774 3180
rect 15757 3163 15774 3180
rect 15677 3163 15694 3180
rect 15717 3163 15734 3180
rect 15637 3163 15654 3180
rect 15757 3163 15774 3180
rect 15677 3163 15694 3180
rect 15717 3163 15734 3180
rect 15557 3163 15574 3180
rect 15797 3163 15814 3180
rect 15597 3163 15614 3180
rect 15637 3163 15654 3180
rect 15557 3163 15574 3180
rect 15597 3163 15614 3180
rect 15637 3163 15654 3180
rect 15797 3163 15814 3180
rect 15637 3163 15654 3180
rect 15677 3163 15694 3180
rect 15557 3163 15574 3180
rect 15637 3163 15654 3180
rect 15597 3163 15614 3180
rect 15597 3163 15614 3180
rect 15717 3163 15734 3180
rect 15757 3163 15774 3180
rect 15677 3163 15694 3180
rect 14562 2394 14579 2411
rect 14522 2394 14539 2411
rect 15082 2394 15099 2411
rect 14882 2394 14899 2411
rect 15402 2394 15419 2411
rect 15522 2394 15539 2411
rect 15042 2394 15059 2411
rect 14922 2394 14939 2411
rect 15562 2394 15579 2411
rect 15002 2394 15019 2411
rect 14882 2394 14899 2411
rect 15162 2394 15179 2411
rect 15362 2394 15379 2411
rect 14962 2394 14979 2411
rect 14962 2394 14979 2411
rect 15442 2394 15459 2411
rect 15122 2394 15139 2411
rect 14922 2394 14939 2411
rect 15322 2394 15339 2411
rect 15562 2394 15579 2411
rect 15522 2394 15539 2411
rect 15482 2394 15499 2411
rect 15442 2394 15459 2411
rect 15402 2394 15419 2411
rect 15362 2394 15379 2411
rect 15322 2394 15339 2411
rect 15242 2394 15259 2411
rect 15282 2394 15299 2411
rect 15282 2394 15299 2411
rect 15202 2394 15219 2411
rect 15162 2394 15179 2411
rect 15242 2394 15259 2411
rect 15122 2394 15139 2411
rect 15482 2394 15499 2411
rect 15082 2394 15099 2411
rect 15202 2394 15219 2411
rect 15042 2394 15059 2411
rect 15002 2394 15019 2411
rect 14482 2394 14499 2411
rect 14482 2394 14499 2411
rect 14442 2394 14459 2411
rect 14402 2394 14419 2411
rect 14682 2394 14699 2411
rect 14842 2394 14859 2411
rect 14802 2394 14819 2411
rect 14442 2394 14459 2411
rect 14762 2394 14779 2411
rect 14402 2394 14419 2411
rect 14642 2394 14659 2411
rect 14842 2394 14859 2411
rect 14602 2394 14619 2411
rect 14802 2394 14819 2411
rect 14762 2394 14779 2411
rect 14562 2394 14579 2411
rect 14722 2394 14739 2411
rect 14682 2394 14699 2411
rect 14642 2394 14659 2411
rect 14722 2394 14739 2411
rect 14602 2394 14619 2411
rect 14522 2394 14539 2411
rect 15842 2394 15859 2411
rect 16402 2394 16419 2411
rect 15882 2394 15899 2411
rect 15762 2394 15779 2411
rect 15922 2394 15939 2411
rect 15842 2394 15859 2411
rect 15882 2394 15899 2411
rect 15922 2394 15939 2411
rect 16682 2394 16699 2411
rect 15682 2394 15699 2411
rect 16242 2394 16259 2411
rect 16362 2394 16379 2411
rect 16202 2394 16219 2411
rect 16322 2394 16339 2411
rect 16642 2394 16659 2411
rect 16362 2394 16379 2411
rect 15722 2394 15739 2411
rect 16322 2394 16339 2411
rect 16602 2394 16619 2411
rect 16282 2394 16299 2411
rect 15682 2394 15699 2411
rect 16282 2394 16299 2411
rect 15642 2394 15659 2411
rect 16562 2394 16579 2411
rect 16522 2394 16539 2411
rect 15602 2394 15619 2411
rect 16242 2394 16259 2411
rect 16482 2394 16499 2411
rect 15642 2394 15659 2411
rect 16202 2394 16219 2411
rect 16162 2394 16179 2411
rect 15722 2394 15739 2411
rect 16402 2394 16419 2411
rect 16442 2394 16459 2411
rect 16162 2394 16179 2411
rect 16722 2394 16739 2411
rect 16682 2394 16699 2411
rect 16642 2394 16659 2411
rect 16602 2394 16619 2411
rect 16562 2394 16579 2411
rect 16522 2394 16539 2411
rect 15802 2394 15819 2411
rect 16482 2394 16499 2411
rect 16122 2394 16139 2411
rect 15602 2394 15619 2411
rect 16082 2394 16099 2411
rect 16042 2394 16059 2411
rect 16002 2394 16019 2411
rect 15802 2394 15819 2411
rect 15962 2394 15979 2411
rect 16082 2394 16099 2411
rect 15762 2394 15779 2411
rect 16042 2394 16059 2411
rect 16002 2394 16019 2411
rect 16442 2394 16459 2411
rect 16122 2394 16139 2411
rect 16722 2394 16739 2411
rect 15962 2394 15979 2411
rect 17402 2394 17419 2411
rect 17362 2394 17379 2411
rect 17322 2394 17339 2411
rect 17282 2394 17299 2411
rect 17242 2394 17259 2411
rect 16882 2394 16899 2411
rect 16842 2394 16859 2411
rect 18082 2394 18099 2411
rect 18042 2394 18059 2411
rect 17002 2394 17019 2411
rect 17002 2394 17019 2411
rect 16962 2394 16979 2411
rect 18002 2394 18019 2411
rect 17962 2394 17979 2411
rect 16802 2394 16819 2411
rect 17922 2394 17939 2411
rect 16962 2394 16979 2411
rect 17882 2394 17899 2411
rect 16842 2394 16859 2411
rect 16922 2394 16939 2411
rect 17842 2394 17859 2411
rect 17802 2394 17819 2411
rect 16922 2394 16939 2411
rect 17202 2394 17219 2411
rect 17762 2394 17779 2411
rect 17722 2394 17739 2411
rect 17682 2394 17699 2411
rect 17642 2394 17659 2411
rect 17602 2394 17619 2411
rect 16802 2394 16819 2411
rect 17562 2394 17579 2411
rect 17162 2394 17179 2411
rect 16882 2394 16899 2411
rect 18082 2394 18099 2411
rect 17122 2394 17139 2411
rect 17082 2394 17099 2411
rect 17042 2394 17059 2411
rect 18042 2394 18059 2411
rect 17122 2394 17139 2411
rect 18002 2394 18019 2411
rect 17082 2394 17099 2411
rect 17042 2394 17059 2411
rect 17482 2394 17499 2411
rect 17442 2394 17459 2411
rect 17522 2394 17539 2411
rect 17962 2394 17979 2411
rect 17522 2394 17539 2411
rect 17922 2394 17939 2411
rect 17882 2394 17899 2411
rect 17842 2394 17859 2411
rect 17802 2394 17819 2411
rect 17762 2394 17779 2411
rect 17722 2394 17739 2411
rect 17682 2394 17699 2411
rect 17642 2394 17659 2411
rect 17602 2394 17619 2411
rect 17562 2394 17579 2411
rect 17402 2394 17419 2411
rect 17362 2394 17379 2411
rect 17322 2394 17339 2411
rect 17282 2394 17299 2411
rect 17242 2394 17259 2411
rect 17202 2394 17219 2411
rect 17162 2394 17179 2411
rect 17482 2394 17499 2411
rect 17442 2394 17459 2411
rect -9412 2394 -9395 2411
rect -9412 2394 -9395 2411
rect -365 8582 -348 8599
rect -325 8582 -308 8599
rect -285 8582 -268 8599
rect -245 8582 -228 8599
rect -205 8582 -188 8599
rect -165 8582 -148 8599
rect -125 8582 -108 8599
rect -85 8582 -68 8599
rect -45 8582 -28 8599
rect -5 8582 13 8599
rect 36 8582 53 8599
rect 76 8582 93 8599
rect -1685 8582 -1668 8599
rect -1725 8582 -1708 8599
rect -1765 8582 -1748 8599
rect -1805 8582 -1788 8599
rect -1845 8582 -1828 8599
rect -1885 8582 -1868 8599
rect -1925 8582 -1908 8599
rect -1965 8582 -1948 8599
rect -2005 8582 -1988 8599
rect -2045 8582 -2028 8599
rect -2085 8582 -2068 8599
rect -2125 8582 -2108 8599
rect -2165 8582 -2148 8599
rect -2205 8582 -2188 8599
rect -965 8582 -948 8599
rect -1685 8582 -1668 8599
rect -1725 8582 -1708 8599
rect -1765 8582 -1748 8599
rect -1805 8582 -1788 8599
rect -1845 8582 -1828 8599
rect -1885 8582 -1868 8599
rect -1925 8582 -1908 8599
rect -1965 8582 -1948 8599
rect -2005 8582 -1988 8599
rect -2045 8582 -2028 8599
rect -2085 8582 -2068 8599
rect -2125 8582 -2108 8599
rect -2165 8582 -2148 8599
rect -2205 8582 -2188 8599
rect -925 8582 -908 8599
rect -2245 8582 -2228 8599
rect -2245 8582 -2228 8599
rect -885 8582 -868 8599
rect -845 8582 -828 8599
rect -805 8582 -788 8599
rect -765 8582 -748 8599
rect -725 8582 -708 8599
rect -685 8582 -668 8599
rect -645 8582 -628 8599
rect -605 8582 -588 8599
rect -565 8582 -548 8599
rect -525 8582 -508 8599
rect -485 8582 -468 8599
rect -445 8582 -428 8599
rect -405 8582 -388 8599
rect -3245 8582 -3228 8599
rect -2485 8582 -2468 8599
rect -2725 8582 -2708 8599
rect -2565 8582 -2548 8599
rect -2285 8582 -2268 8599
rect -3285 8582 -3268 8599
rect -2765 8582 -2748 8599
rect -2805 8582 -2788 8599
rect -2765 8582 -2748 8599
rect -3085 8582 -3068 8599
rect -2805 8582 -2788 8599
rect -2525 8582 -2508 8599
rect -3325 8582 -3308 8599
rect -3405 8582 -3388 8599
rect -3325 8582 -3308 8599
rect -2525 8582 -2508 8599
rect -2325 8582 -2308 8599
rect -2365 8582 -2348 8599
rect -2965 8582 -2948 8599
rect -3125 8582 -3108 8599
rect -2565 8582 -2548 8599
rect -2645 8582 -2628 8599
rect -3445 8582 -3428 8599
rect -2605 8582 -2588 8599
rect -3285 8582 -3268 8599
rect -2405 8582 -2388 8599
rect -2365 8582 -2348 8599
rect -2685 8582 -2668 8599
rect -2845 8582 -2828 8599
rect -3165 8582 -3148 8599
rect -2845 8582 -2828 8599
rect -2605 8582 -2588 8599
rect -3365 8582 -3348 8599
rect -2885 8582 -2868 8599
rect -2925 8582 -2908 8599
rect -3445 8582 -3428 8599
rect -2405 8582 -2388 8599
rect -2285 8582 -2268 8599
rect -3405 8582 -3388 8599
rect -3005 8582 -2988 8599
rect -2325 8582 -2308 8599
rect -2885 8582 -2868 8599
rect -2445 8582 -2428 8599
rect -2685 8582 -2668 8599
rect -2725 8582 -2708 8599
rect -2925 8582 -2908 8599
rect -3205 8582 -3188 8599
rect -3365 8582 -3348 8599
rect -2645 8582 -2628 8599
rect -2965 8582 -2948 8599
rect -3005 8582 -2988 8599
rect -3045 8582 -3028 8599
rect -3085 8582 -3068 8599
rect -2445 8582 -2428 8599
rect -3125 8582 -3108 8599
rect -3165 8582 -3148 8599
rect -3205 8582 -3188 8599
rect -3245 8582 -3228 8599
rect -3045 8582 -3028 8599
rect -2485 8582 -2468 8599
rect -3925 8582 -3908 8599
rect -4485 8582 -4468 8599
rect -4405 8582 -4388 8599
rect -3765 8582 -3748 8599
rect -4285 8582 -4268 8599
rect -4325 8582 -4308 8599
rect -3565 8582 -3548 8599
rect -4565 8582 -4548 8599
rect -3685 8582 -3668 8599
rect -3605 8582 -3588 8599
rect -3765 8582 -3748 8599
rect -3885 8582 -3868 8599
rect -4205 8582 -4188 8599
rect -3885 8582 -3868 8599
rect -4245 8582 -4228 8599
rect -3605 8582 -3588 8599
rect -3805 8582 -3788 8599
rect -3485 8582 -3468 8599
rect -4485 8582 -4468 8599
rect -3645 8582 -3628 8599
rect -4125 8582 -4108 8599
rect -3485 8582 -3468 8599
rect -3965 8582 -3948 8599
rect -3805 8582 -3788 8599
rect -3725 8582 -3708 8599
rect -4445 8582 -4428 8599
rect -4165 8582 -4148 8599
rect -3645 8582 -3628 8599
rect -4445 8582 -4428 8599
rect -4365 8582 -4348 8599
rect -4605 8582 -4588 8599
rect -4405 8582 -4388 8599
rect -3965 8582 -3948 8599
rect -4045 8582 -4028 8599
rect -4005 8582 -3988 8599
rect -3845 8582 -3828 8599
rect -4285 8582 -4268 8599
rect -4605 8582 -4588 8599
rect -4325 8582 -4308 8599
rect -3845 8582 -3828 8599
rect -4645 8582 -4628 8599
rect -3565 8582 -3548 8599
rect -4085 8582 -4068 8599
rect -4525 8582 -4508 8599
rect -4365 8582 -4348 8599
rect -4245 8582 -4228 8599
rect -3525 8582 -3508 8599
rect -4165 8582 -4148 8599
rect -4645 8582 -4628 8599
rect -3525 8582 -3508 8599
rect -4525 8582 -4508 8599
rect -3685 8582 -3668 8599
rect -4085 8582 -4068 8599
rect -4005 8582 -3988 8599
rect -4205 8582 -4188 8599
rect -3925 8582 -3908 8599
rect -3725 8582 -3708 8599
rect -4125 8582 -4108 8599
rect -4565 8582 -4548 8599
rect -4045 8582 -4028 8599
rect -5845 8582 -5828 8599
rect -5845 8582 -5828 8599
rect -5285 8582 -5268 8599
rect -4925 8582 -4908 8599
rect -5445 8582 -5428 8599
rect -5365 8582 -5348 8599
rect -5165 8582 -5148 8599
rect -5165 8582 -5148 8599
rect -4965 8582 -4948 8599
rect -5445 8582 -5428 8599
rect -5485 8582 -5468 8599
rect -5245 8582 -5228 8599
rect -5005 8582 -4988 8599
rect -5525 8582 -5508 8599
rect -4765 8582 -4748 8599
rect -4805 8582 -4788 8599
rect -5765 8582 -5748 8599
rect -5525 8582 -5508 8599
rect -5565 8582 -5548 8599
rect -5125 8582 -5108 8599
rect -5565 8582 -5548 8599
rect -5605 8582 -5588 8599
rect -4885 8582 -4868 8599
rect -5045 8582 -5028 8599
rect -5685 8582 -5668 8599
rect -5085 8582 -5068 8599
rect -5805 8582 -5788 8599
rect -5605 8582 -5588 8599
rect -5645 8582 -5628 8599
rect -5205 8582 -5188 8599
rect -5685 8582 -5668 8599
rect -4845 8582 -4828 8599
rect -4925 8582 -4908 8599
rect -5725 8582 -5708 8599
rect -4685 8582 -4668 8599
rect -5205 8582 -5188 8599
rect -5765 8582 -5748 8599
rect -4685 8582 -4668 8599
rect -5405 8582 -5388 8599
rect -4965 8582 -4948 8599
rect -4845 8582 -4828 8599
rect -5285 8582 -5268 8599
rect -5805 8582 -5788 8599
rect -5325 8582 -5308 8599
rect -4765 8582 -4748 8599
rect -4805 8582 -4788 8599
rect -5005 8582 -4988 8599
rect -4885 8582 -4868 8599
rect -5125 8582 -5108 8599
rect -5645 8582 -5628 8599
rect -5365 8582 -5348 8599
rect -5085 8582 -5068 8599
rect -5045 8582 -5028 8599
rect -4725 8582 -4708 8599
rect -5325 8582 -5308 8599
rect -5725 8582 -5708 8599
rect -4725 8582 -4708 8599
rect -5245 8582 -5228 8599
rect -5485 8582 -5468 8599
rect -5405 8582 -5388 8599
rect -6166 8582 -6149 8599
rect -6446 8582 -6429 8599
rect -6926 8582 -6909 8599
rect -6766 8582 -6749 8599
rect -6246 8582 -6229 8599
rect -5965 8582 -5948 8599
rect -6046 8582 -6029 8599
rect -6886 8582 -6869 8599
rect -6486 8582 -6469 8599
rect -6446 8582 -6429 8599
rect -6806 8582 -6789 8599
rect -6046 8582 -6029 8599
rect -5885 8582 -5868 8599
rect -6326 8582 -6309 8599
rect -6526 8582 -6509 8599
rect -6686 8582 -6669 8599
rect -6646 8582 -6629 8599
rect -6126 8582 -6109 8599
rect -6766 8582 -6749 8599
rect -6246 8582 -6229 8599
rect -6566 8582 -6549 8599
rect -6326 8582 -6309 8599
rect -5925 8582 -5908 8599
rect -6806 8582 -6789 8599
rect -6006 8582 -5989 8599
rect -6366 8582 -6349 8599
rect -7006 8582 -6989 8599
rect -6566 8582 -6549 8599
rect -6486 8582 -6469 8599
rect -6086 8582 -6069 8599
rect -6846 8582 -6829 8599
rect -6006 8582 -5989 8599
rect -5965 8582 -5948 8599
rect -6966 8582 -6949 8599
rect -6366 8582 -6349 8599
rect -6286 8582 -6269 8599
rect -6166 8582 -6149 8599
rect -6846 8582 -6829 8599
rect -6966 8582 -6949 8599
rect -6526 8582 -6509 8599
rect -6206 8582 -6189 8599
rect -6606 8582 -6589 8599
rect -6726 8582 -6709 8599
rect -7006 8582 -6989 8599
rect -6926 8582 -6909 8599
rect -6126 8582 -6109 8599
rect -6726 8582 -6709 8599
rect -5885 8582 -5868 8599
rect -5925 8582 -5908 8599
rect -6646 8582 -6629 8599
rect -6406 8582 -6389 8599
rect -6286 8582 -6269 8599
rect -6206 8582 -6189 8599
rect -6606 8582 -6589 8599
rect -6406 8582 -6389 8599
rect -6686 8582 -6669 8599
rect -6086 8582 -6069 8599
rect -6886 8582 -6869 8599
rect -7286 8582 -7269 8599
rect -7366 8582 -7349 8599
rect -7766 8582 -7749 8599
rect -7086 8582 -7069 8599
rect -8126 8582 -8109 8599
rect -7086 8582 -7069 8599
rect -7806 8582 -7789 8599
rect -7966 8582 -7949 8599
rect -7886 8582 -7869 8599
rect -7726 8582 -7709 8599
rect -7286 8582 -7269 8599
rect -7566 8582 -7549 8599
rect -7806 8582 -7789 8599
rect -7326 8582 -7309 8599
rect -7206 8582 -7189 8599
rect -8126 8582 -8109 8599
rect -8166 8582 -8149 8599
rect -7646 8582 -7629 8599
rect -7686 8582 -7669 8599
rect -7126 8582 -7109 8599
rect -7646 8582 -7629 8599
rect -8166 8582 -8149 8599
rect -7446 8582 -7429 8599
rect -8006 8582 -7989 8599
rect -7486 8582 -7469 8599
rect -7046 8582 -7029 8599
rect -7166 8582 -7149 8599
rect -7966 8582 -7949 8599
rect -7446 8582 -7429 8599
rect -8086 8582 -8069 8599
rect -8006 8582 -7989 8599
rect -7046 8582 -7029 8599
rect -7326 8582 -7309 8599
rect -7406 8582 -7389 8599
rect -8206 8582 -8189 8599
rect -7526 8582 -7509 8599
rect -7166 8582 -7149 8599
rect -7606 8582 -7589 8599
rect -7766 8582 -7749 8599
rect -7486 8582 -7469 8599
rect -8206 8582 -8189 8599
rect -7246 8582 -7229 8599
rect -8046 8582 -8029 8599
rect -7686 8582 -7669 8599
rect -7206 8582 -7189 8599
rect -7886 8582 -7869 8599
rect -7726 8582 -7709 8599
rect -7526 8582 -7509 8599
rect -7366 8582 -7349 8599
rect -7846 8582 -7829 8599
rect -7926 8582 -7909 8599
rect -7406 8582 -7389 8599
rect -7846 8582 -7829 8599
rect -7246 8582 -7229 8599
rect -7566 8582 -7549 8599
rect -7606 8582 -7589 8599
rect -8046 8582 -8029 8599
rect -7126 8582 -7109 8599
rect -8086 8582 -8069 8599
rect -7926 8582 -7909 8599
rect -8806 8582 -8789 8599
rect -8886 8582 -8869 8599
rect -8606 8582 -8589 8599
rect -8926 8582 -8909 8599
rect -9166 8582 -9149 8599
rect -8246 8582 -8229 8599
rect -8286 8582 -8269 8599
rect -8446 8582 -8429 8599
rect -8686 8582 -8669 8599
rect -8286 8582 -8269 8599
rect -8606 8582 -8589 8599
rect -8566 8582 -8549 8599
rect -8406 8582 -8389 8599
rect -9366 8582 -9349 8599
rect -8926 8582 -8909 8599
rect -8486 8582 -8469 8599
rect -8846 8582 -8829 8599
rect -9286 8582 -9269 8599
rect -8806 8582 -8789 8599
rect -8526 8582 -8509 8599
rect -8966 8582 -8949 8599
rect -8766 8582 -8749 8599
rect -9366 8582 -9349 8599
rect -9086 8582 -9069 8599
rect -8246 8582 -8229 8599
rect -8486 8582 -8469 8599
rect -9326 8582 -9309 8599
rect -8886 8582 -8869 8599
rect -8526 8582 -8509 8599
rect -9326 8582 -9309 8599
rect -9006 8582 -8989 8599
rect -9206 8582 -9189 8599
rect -9166 8582 -9149 8599
rect -8646 8582 -8629 8599
rect -8846 8582 -8829 8599
rect -9206 8582 -9189 8599
rect -8366 8582 -8349 8599
rect -9246 8582 -9229 8599
rect -8326 8582 -8309 8599
rect -9286 8582 -9269 8599
rect -8726 8582 -8709 8599
rect -9126 8582 -9109 8599
rect -9246 8582 -9229 8599
rect -8686 8582 -8669 8599
rect -9406 8582 -9389 8599
rect -8966 8582 -8949 8599
rect -9406 8582 -9389 8599
rect -9046 8582 -9029 8599
rect -8446 8582 -8429 8599
rect -8326 8582 -8309 8599
rect -8646 8582 -8629 8599
rect -9046 8582 -9029 8599
rect -8366 8582 -8349 8599
rect -8766 8582 -8749 8599
rect -9126 8582 -9109 8599
rect -8566 8582 -8549 8599
rect -8406 8582 -8389 8599
rect -9006 8582 -8989 8599
rect -9086 8582 -9069 8599
rect -8726 8582 -8709 8599
rect -10606 8582 -10589 8599
rect -10606 8582 -10589 8599
rect -10326 8582 -10309 8599
rect -10406 8582 -10389 8599
rect -10086 8582 -10069 8599
rect -10446 8582 -10429 8599
rect -10366 8582 -10349 8599
rect -10406 8582 -10389 8599
rect -10486 8582 -10469 8599
rect -9646 8582 -9629 8599
rect -10126 8582 -10109 8599
rect -9686 8582 -9669 8599
rect -10246 8582 -10229 8599
rect -9726 8582 -9709 8599
rect -10446 8582 -10429 8599
rect -10526 8582 -10509 8599
rect -9806 8582 -9789 8599
rect -9486 8582 -9469 8599
rect -9886 8582 -9869 8599
rect -10246 8582 -10229 8599
rect -10046 8582 -10029 8599
rect -9606 8582 -9589 8599
rect -10126 8582 -10109 8599
rect -10566 8582 -10549 8599
rect -10006 8582 -9989 8599
rect -9526 8582 -9509 8599
rect -9446 8582 -9429 8599
rect -9446 8582 -9429 8599
rect -10286 8582 -10269 8599
rect -10086 8582 -10069 8599
rect -9526 8582 -9509 8599
rect -10046 8582 -10029 8599
rect -9726 8582 -9709 8599
rect -10006 8582 -9989 8599
rect -9846 8582 -9829 8599
rect -10366 8582 -10349 8599
rect -10206 8582 -10189 8599
rect -10166 8582 -10149 8599
rect -9886 8582 -9869 8599
rect -9806 8582 -9789 8599
rect -9966 8582 -9949 8599
rect -9486 8582 -9469 8599
rect -9686 8582 -9669 8599
rect -10486 8582 -10469 8599
rect -9766 8582 -9749 8599
rect -9966 8582 -9949 8599
rect -10526 8582 -10509 8599
rect -9926 8582 -9909 8599
rect -9566 8582 -9549 8599
rect -10326 8582 -10309 8599
rect -9566 8582 -9549 8599
rect -9646 8582 -9629 8599
rect -10206 8582 -10189 8599
rect -10566 8582 -10549 8599
rect -9846 8582 -9829 8599
rect -9766 8582 -9749 8599
rect -10166 8582 -10149 8599
rect -10286 8582 -10269 8599
rect -9926 8582 -9909 8599
rect -9606 8582 -9589 8599
rect -10726 8582 -10709 8599
rect -11606 8582 -11589 8599
rect -11166 8582 -11149 8599
rect -10686 8582 -10669 8599
rect -10806 8582 -10789 8599
rect -11366 8582 -11349 8599
rect -11646 8582 -11629 8599
rect -10886 8582 -10869 8599
rect -11126 8582 -11109 8599
rect -11006 8582 -10989 8599
rect -10726 8582 -10709 8599
rect -11086 8582 -11069 8599
rect -11406 8582 -11389 8599
rect -11526 8582 -11509 8599
rect -11486 8582 -11469 8599
rect -11686 8582 -11669 8599
rect -11326 8582 -11309 8599
rect -11126 8582 -11109 8599
rect -11406 8582 -11389 8599
rect -11086 8582 -11069 8599
rect -10926 8582 -10909 8599
rect -11286 8582 -11269 8599
rect -11686 8582 -11669 8599
rect -11566 8582 -11549 8599
rect -11166 8582 -11149 8599
rect -10766 8582 -10749 8599
rect -11646 8582 -11629 8599
rect -10966 8582 -10949 8599
rect -11246 8582 -11229 8599
rect -11446 8582 -11429 8599
rect -11766 8582 -11749 8599
rect -10766 8582 -10749 8599
rect -11046 8582 -11029 8599
rect -11486 8582 -11469 8599
rect -11566 8582 -11549 8599
rect -11446 8582 -11429 8599
rect -11726 8582 -11709 8599
rect -11246 8582 -11229 8599
rect -11606 8582 -11589 8599
rect -11366 8582 -11349 8599
rect -11046 8582 -11029 8599
rect -10846 8582 -10829 8599
rect -10926 8582 -10909 8599
rect -11326 8582 -11309 8599
rect -10646 8582 -10629 8599
rect -10646 8582 -10629 8599
rect -10806 8582 -10789 8599
rect -11766 8582 -11749 8599
rect -11006 8582 -10989 8599
rect -11206 8582 -11189 8599
rect -11206 8582 -11189 8599
rect -10846 8582 -10829 8599
rect -11726 8582 -11709 8599
rect -10886 8582 -10869 8599
rect -11286 8582 -11269 8599
rect -10686 8582 -10669 8599
rect -11526 8582 -11509 8599
rect -10966 8582 -10949 8599
rect -12166 8582 -12149 8599
rect -12566 8582 -12549 8599
rect -12046 8582 -12029 8599
rect -12126 8582 -12109 8599
rect -12286 8582 -12269 8599
rect -12886 8582 -12869 8599
rect -12806 8582 -12789 8599
rect -12686 8582 -12669 8599
rect -11926 8582 -11909 8599
rect -12406 8582 -12389 8599
rect -12606 8582 -12589 8599
rect -12366 8582 -12349 8599
rect -12526 8582 -12509 8599
rect -12006 8582 -11989 8599
rect -12966 8582 -12949 8599
rect -12446 8582 -12429 8599
rect -11966 8582 -11949 8599
rect -12206 8582 -12189 8599
rect -12766 8582 -12749 8599
rect -12926 8582 -12909 8599
rect -12646 8582 -12629 8599
rect -12726 8582 -12709 8599
rect -11846 8582 -11829 8599
rect -11886 8582 -11869 8599
rect -12966 8582 -12949 8599
rect -11846 8582 -11829 8599
rect -11966 8582 -11949 8599
rect -12326 8582 -12309 8599
rect -12606 8582 -12589 8599
rect -12686 8582 -12669 8599
rect -12086 8582 -12069 8599
rect -12726 8582 -12709 8599
rect -12166 8582 -12149 8599
rect -12886 8582 -12869 8599
rect -12206 8582 -12189 8599
rect -11886 8582 -11869 8599
rect -12006 8582 -11989 8599
rect -12766 8582 -12749 8599
rect -12246 8582 -12229 8599
rect -12926 8582 -12909 8599
rect -12246 8582 -12229 8599
rect -12086 8582 -12069 8599
rect -12806 8582 -12789 8599
rect -12406 8582 -12389 8599
rect -12366 8582 -12349 8599
rect -12486 8582 -12469 8599
rect -12446 8582 -12429 8599
rect -12846 8582 -12829 8599
rect -12486 8582 -12469 8599
rect -11926 8582 -11909 8599
rect -12286 8582 -12269 8599
rect -12846 8582 -12829 8599
rect -12126 8582 -12109 8599
rect -11806 8582 -11789 8599
rect -12326 8582 -12309 8599
rect -12046 8582 -12029 8599
rect -11806 8582 -11789 8599
rect -12566 8582 -12549 8599
rect -12646 8582 -12629 8599
rect -12526 8582 -12509 8599
rect -13246 8582 -13229 8599
rect -13166 8582 -13149 8599
rect -13406 8582 -13389 8599
rect -13686 8582 -13669 8599
rect -13966 8582 -13949 8599
rect -13966 8582 -13949 8599
rect -13486 8582 -13469 8599
rect -14006 8582 -13989 8599
rect -14126 8582 -14109 8599
rect -14006 8582 -13989 8599
rect -13486 8582 -13469 8599
rect -13886 8582 -13869 8599
rect -13606 8582 -13589 8599
rect -13566 8582 -13549 8599
rect -14046 8582 -14029 8599
rect -13046 8582 -13029 8599
rect -13286 8582 -13269 8599
rect -13606 8582 -13589 8599
rect -13206 8582 -13189 8599
rect -13646 8582 -13629 8599
rect -13526 8582 -13509 8599
rect -13926 8582 -13909 8599
rect -13006 8582 -12989 8599
rect -13766 8582 -13749 8599
rect -13846 8582 -13829 8599
rect -13566 8582 -13549 8599
rect -13726 8582 -13709 8599
rect -13086 8582 -13069 8599
rect -14166 8582 -14149 8599
rect -13206 8582 -13189 8599
rect -13326 8582 -13309 8599
rect -13086 8582 -13069 8599
rect -13726 8582 -13709 8599
rect -13686 8582 -13669 8599
rect -13366 8582 -13349 8599
rect -13126 8582 -13109 8599
rect -13046 8582 -13029 8599
rect -13286 8582 -13269 8599
rect -13406 8582 -13389 8599
rect -13246 8582 -13229 8599
rect -14086 8582 -14069 8599
rect -13446 8582 -13429 8599
rect -13366 8582 -13349 8599
rect -14086 8582 -14069 8599
rect -14126 8582 -14109 8599
rect -14166 8582 -14149 8599
rect -13766 8582 -13749 8599
rect -13846 8582 -13829 8599
rect -13446 8582 -13429 8599
rect -13166 8582 -13149 8599
rect -13326 8582 -13309 8599
rect -13886 8582 -13869 8599
rect -13806 8582 -13789 8599
rect -13006 8582 -12989 8599
rect -13646 8582 -13629 8599
rect -13526 8582 -13509 8599
rect -13926 8582 -13909 8599
rect -14046 8582 -14029 8599
rect -13126 8582 -13109 8599
rect -13806 8582 -13789 8599
rect -15366 8582 -15349 8599
rect -15366 8582 -15349 8599
rect -15126 8582 -15109 8599
rect -14966 8582 -14949 8599
rect -14606 8582 -14589 8599
rect -15166 8582 -15149 8599
rect -15126 8582 -15109 8599
rect -15206 8582 -15189 8599
rect -14686 8582 -14669 8599
rect -15046 8582 -15029 8599
rect -14526 8582 -14509 8599
rect -15086 8582 -15069 8599
rect -14406 8582 -14389 8599
rect -14926 8582 -14909 8599
rect -14766 8582 -14749 8599
rect -14566 8582 -14549 8599
rect -14366 8582 -14349 8599
rect -15326 8582 -15309 8599
rect -14246 8582 -14229 8599
rect -15006 8582 -14989 8599
rect -15326 8582 -15309 8599
rect -14526 8582 -14509 8599
rect -14326 8582 -14309 8599
rect -14646 8582 -14629 8599
rect -15246 8582 -15229 8599
rect -14726 8582 -14709 8599
rect -14646 8582 -14629 8599
rect -14486 8582 -14469 8599
rect -15286 8582 -15269 8599
rect -14726 8582 -14709 8599
rect -14846 8582 -14829 8599
rect -14286 8582 -14269 8599
rect -15246 8582 -15229 8599
rect -14606 8582 -14589 8599
rect -14686 8582 -14669 8599
rect -15006 8582 -14989 8599
rect -14206 8582 -14189 8599
rect -14286 8582 -14269 8599
rect -15046 8582 -15029 8599
rect -14886 8582 -14869 8599
rect -14926 8582 -14909 8599
rect -15166 8582 -15149 8599
rect -15286 8582 -15269 8599
rect -14566 8582 -14549 8599
rect -14966 8582 -14949 8599
rect -14366 8582 -14349 8599
rect -15086 8582 -15069 8599
rect -14806 8582 -14789 8599
rect -14206 8582 -14189 8599
rect -14406 8582 -14389 8599
rect -14446 8582 -14429 8599
rect -14766 8582 -14749 8599
rect -14326 8582 -14309 8599
rect -14806 8582 -14789 8599
rect -14846 8582 -14829 8599
rect -14486 8582 -14469 8599
rect -14446 8582 -14429 8599
rect -14886 8582 -14869 8599
rect -14246 8582 -14229 8599
rect -15206 8582 -15189 8599
rect -15486 8582 -15469 8599
rect -15726 8582 -15709 8599
rect -15846 8582 -15829 8599
rect -16246 8582 -16229 8599
rect -16006 8582 -15989 8599
rect -15846 8582 -15829 8599
rect -15766 8582 -15749 8599
rect -15766 8582 -15749 8599
rect -16126 8582 -16109 8599
rect -16526 8582 -16509 8599
rect -16006 8582 -15989 8599
rect -16326 8582 -16309 8599
rect -15526 8582 -15509 8599
rect -16046 8582 -16029 8599
rect -16046 8582 -16029 8599
rect -15646 8582 -15629 8599
rect -15646 8582 -15629 8599
rect -15566 8582 -15549 8599
rect -15406 8582 -15389 8599
rect -15686 8582 -15669 8599
rect -16486 8582 -16469 8599
rect -16366 8582 -16349 8599
rect -15486 8582 -15469 8599
rect -15406 8582 -15389 8599
rect -15686 8582 -15669 8599
rect -15886 8582 -15869 8599
rect -15886 8582 -15869 8599
rect -15926 8582 -15909 8599
rect -16286 8582 -16269 8599
rect -16446 8582 -16429 8599
rect -15606 8582 -15589 8599
rect -15526 8582 -15509 8599
rect -16486 8582 -16469 8599
rect -15726 8582 -15709 8599
rect -16206 8582 -16189 8599
rect -16206 8582 -16189 8599
rect -15966 8582 -15949 8599
rect -15446 8582 -15429 8599
rect -15446 8582 -15429 8599
rect -16086 8582 -16069 8599
rect -16166 8582 -16149 8599
rect -16366 8582 -16349 8599
rect -16286 8582 -16269 8599
rect -16086 8582 -16069 8599
rect -16166 8582 -16149 8599
rect -15966 8582 -15949 8599
rect -16446 8582 -16429 8599
rect -16326 8582 -16309 8599
rect -16406 8582 -16389 8599
rect -16126 8582 -16109 8599
rect -15806 8582 -15789 8599
rect -15606 8582 -15589 8599
rect -16406 8582 -16389 8599
rect -16526 8582 -16509 8599
rect -15566 8582 -15549 8599
rect -16246 8582 -16229 8599
rect -15806 8582 -15789 8599
rect -15926 8582 -15909 8599
rect -17326 8582 -17309 8599
rect -17206 8582 -17189 8599
rect -17246 8582 -17229 8599
rect -16846 8582 -16829 8599
rect -17566 8582 -17549 8599
rect -16606 8582 -16589 8599
rect -16686 8582 -16669 8599
rect -17406 8582 -17389 8599
rect -16766 8582 -16749 8599
rect -17446 8582 -17429 8599
rect -17046 8582 -17029 8599
rect -16966 8582 -16949 8599
rect -16806 8582 -16789 8599
rect -17126 8582 -17109 8599
rect -16926 8582 -16909 8599
rect -17686 8582 -17669 8599
rect -17726 8582 -17709 8599
rect -17606 8582 -17589 8599
rect -16886 8582 -16869 8599
rect -17486 8582 -17469 8599
rect -16726 8582 -16709 8599
rect -17286 8582 -17269 8599
rect -16886 8582 -16869 8599
rect -17366 8582 -17349 8599
rect -17486 8582 -17469 8599
rect -17726 8582 -17709 8599
rect -16966 8582 -16949 8599
rect -16646 8582 -16629 8599
rect -17286 8582 -17269 8599
rect -17526 8582 -17509 8599
rect -17566 8582 -17549 8599
rect -17686 8582 -17669 8599
rect -17206 8582 -17189 8599
rect -16646 8582 -16629 8599
rect -17326 8582 -17309 8599
rect -17406 8582 -17389 8599
rect -17006 8582 -16989 8599
rect -17246 8582 -17229 8599
rect -16846 8582 -16829 8599
rect -16926 8582 -16909 8599
rect -17046 8582 -17029 8599
rect -17526 8582 -17509 8599
rect -17606 8582 -17589 8599
rect -16686 8582 -16669 8599
rect -17086 8582 -17069 8599
rect -17086 8582 -17069 8599
rect -17646 8582 -17629 8599
rect -16606 8582 -16589 8599
rect -17646 8582 -17629 8599
rect -16566 8582 -16549 8599
rect -16766 8582 -16749 8599
rect -17366 8582 -17349 8599
rect -17166 8582 -17149 8599
rect -16806 8582 -16789 8599
rect -17446 8582 -17429 8599
rect -17166 8582 -17149 8599
rect -17006 8582 -16989 8599
rect -16566 8582 -16549 8599
rect -17126 8582 -17109 8599
rect -16726 8582 -16709 8599
rect -17846 8582 -17829 8599
rect -18166 8582 -18149 8599
rect -18086 8582 -18069 8599
rect -18606 8582 -18589 8599
rect -18006 8582 -17989 8599
rect -18006 8582 -17989 8599
rect -18486 8582 -18469 8599
rect -18446 8582 -18429 8599
rect -17926 8582 -17909 8599
rect -18246 8582 -18229 8599
rect -18926 8582 -18909 8599
rect -18846 8582 -18829 8599
rect -18046 8582 -18029 8599
rect -18806 8582 -18789 8599
rect -18246 8582 -18229 8599
rect -17926 8582 -17909 8599
rect -18326 8582 -18309 8599
rect -18406 8582 -18389 8599
rect -18686 8582 -18669 8599
rect -18566 8582 -18549 8599
rect -18086 8582 -18069 8599
rect -17806 8582 -17789 8599
rect -18686 8582 -18669 8599
rect -18766 8582 -18749 8599
rect -18046 8582 -18029 8599
rect -17886 8582 -17869 8599
rect -18326 8582 -18309 8599
rect -18206 8582 -18189 8599
rect -18126 8582 -18109 8599
rect -18286 8582 -18269 8599
rect -18526 8582 -18509 8599
rect -18366 8582 -18349 8599
rect -18526 8582 -18509 8599
rect -18446 8582 -18429 8599
rect -18766 8582 -18749 8599
rect -17966 8582 -17949 8599
rect -18646 8582 -18629 8599
rect -17846 8582 -17829 8599
rect -18126 8582 -18109 8599
rect -18646 8582 -18629 8599
rect -18926 8582 -18909 8599
rect -18486 8582 -18469 8599
rect -18286 8582 -18269 8599
rect -18206 8582 -18189 8599
rect -18366 8582 -18349 8599
rect -17766 8582 -17749 8599
rect -18886 8582 -18869 8599
rect -18726 8582 -18709 8599
rect -17886 8582 -17869 8599
rect -18566 8582 -18549 8599
rect -18406 8582 -18389 8599
rect -18726 8582 -18709 8599
rect -18806 8582 -18789 8599
rect -17766 8582 -17749 8599
rect -17806 8582 -17789 8599
rect -18166 8582 -18149 8599
rect -18846 8582 -18829 8599
rect -18886 8582 -18869 8599
rect -17966 8582 -17949 8599
rect -18606 8582 -18589 8599
rect -14173 2394 -14156 2411
rect -14173 2394 -14156 2411
rect -11926 4652 -11909 4669
rect -11966 4652 -11949 4669
rect -11926 4652 -11909 4669
rect -12006 4652 -11989 4669
rect -12046 4652 -12029 4669
rect -11966 4652 -11949 4669
rect -12086 4652 -12069 4669
rect -12126 4652 -12109 4669
rect -12006 4652 -11989 4669
rect -12166 4652 -12149 4669
rect -12046 4652 -12029 4669
rect -12086 4652 -12069 4669
rect -11806 4652 -11789 4669
rect -12126 4652 -12109 4669
rect -12166 4652 -12149 4669
rect -12206 4652 -12189 4669
rect -11846 4652 -11829 4669
rect -12246 4652 -12229 4669
rect -12286 4652 -12269 4669
rect -12326 4652 -12309 4669
rect -11886 4652 -11869 4669
rect -12366 4652 -12349 4669
rect -12006 4652 -11989 4669
rect -12206 4652 -12189 4669
rect -12206 4652 -12189 4669
rect -12246 4652 -12229 4669
rect -12286 4652 -12269 4669
rect -12326 4652 -12309 4669
rect -11806 4652 -11789 4669
rect -12366 4652 -12349 4669
rect -11966 4652 -11949 4669
rect -11846 4652 -11829 4669
rect -11846 4652 -11829 4669
rect -11886 4652 -11869 4669
rect -11886 4652 -11869 4669
rect -12166 4652 -12149 4669
rect -12006 4652 -11989 4669
rect -11846 4652 -11829 4669
rect -12206 4652 -12189 4669
rect -11966 4652 -11949 4669
rect -12326 4652 -12309 4669
rect -12246 4652 -12229 4669
rect -12086 4652 -12069 4669
rect -12126 4652 -12109 4669
rect -12286 4652 -12269 4669
rect -11886 4652 -11869 4669
rect -12046 4652 -12029 4669
rect -12246 4652 -12229 4669
rect -12086 4652 -12069 4669
rect -11806 4652 -11789 4669
rect -12366 4652 -12349 4669
rect -12166 4652 -12149 4669
rect -12126 4652 -12109 4669
rect -11926 4652 -11909 4669
rect -12046 4652 -12029 4669
rect -12326 4652 -12309 4669
rect -11806 4652 -11789 4669
rect -12286 4652 -12269 4669
rect -11926 4652 -11909 4669
rect -12366 4652 -12349 4669
rect -12806 4652 -12789 4669
rect -12486 4652 -12469 4669
rect -12726 4652 -12709 4669
rect -12606 4652 -12589 4669
rect -12926 4652 -12909 4669
rect -12486 4652 -12469 4669
rect -12646 4652 -12629 4669
rect -12526 4652 -12509 4669
rect -12566 4652 -12549 4669
rect -12686 4652 -12669 4669
rect -12406 4652 -12389 4669
rect -12606 4652 -12589 4669
rect -12526 4652 -12509 4669
rect -12966 4652 -12949 4669
rect -12446 4652 -12429 4669
rect -12766 4652 -12749 4669
rect -12926 4652 -12909 4669
rect -12646 4652 -12629 4669
rect -12966 4652 -12949 4669
rect -12686 4652 -12669 4669
rect -12726 4652 -12709 4669
rect -12886 4652 -12869 4669
rect -12766 4652 -12749 4669
rect -12806 4652 -12789 4669
rect -12446 4652 -12429 4669
rect -12846 4652 -12829 4669
rect -12846 4652 -12829 4669
rect -12566 4652 -12549 4669
rect -12886 4652 -12869 4669
rect -12406 4652 -12389 4669
rect -12406 4652 -12389 4669
rect -12446 4652 -12429 4669
rect -12406 4652 -12389 4669
rect -12446 4652 -12429 4669
rect -12726 4652 -12709 4669
rect -12526 4652 -12509 4669
rect -12886 4652 -12869 4669
rect -12566 4652 -12549 4669
rect -12806 4652 -12789 4669
rect -12606 4652 -12589 4669
rect -12926 4652 -12909 4669
rect -12486 4652 -12469 4669
rect -12646 4652 -12629 4669
rect -12526 4652 -12509 4669
rect -12566 4652 -12549 4669
rect -12686 4652 -12669 4669
rect -12606 4652 -12589 4669
rect -12646 4652 -12629 4669
rect -12966 4652 -12949 4669
rect -12686 4652 -12669 4669
rect -12726 4652 -12709 4669
rect -12766 4652 -12749 4669
rect -12806 4652 -12789 4669
rect -12846 4652 -12829 4669
rect -12846 4652 -12829 4669
rect -12886 4652 -12869 4669
rect -12926 4652 -12909 4669
rect -12486 4652 -12469 4669
rect -12966 4652 -12949 4669
rect -12766 4652 -12749 4669
rect -13206 4652 -13189 4669
rect -13126 4652 -13109 4669
rect -13246 4652 -13229 4669
rect -13566 4652 -13549 4669
rect -13286 4652 -13269 4669
rect -13406 4652 -13389 4669
rect -13006 4652 -12989 4669
rect -13166 4652 -13149 4669
rect -13326 4652 -13309 4669
rect -13446 4652 -13429 4669
rect -13126 4652 -13109 4669
rect -13046 4652 -13029 4669
rect -13206 4652 -13189 4669
rect -13246 4652 -13229 4669
rect -13366 4652 -13349 4669
rect -13526 4652 -13509 4669
rect -13326 4652 -13309 4669
rect -13246 4652 -13229 4669
rect -13486 4652 -13469 4669
rect -13006 4652 -12989 4669
rect -13486 4652 -13469 4669
rect -13446 4652 -13429 4669
rect -13006 4652 -12989 4669
rect -13286 4652 -13269 4669
rect -13006 4652 -12989 4669
rect -13086 4652 -13069 4669
rect -13046 4652 -13029 4669
rect -13326 4652 -13309 4669
rect -13566 4652 -13549 4669
rect -13406 4652 -13389 4669
rect -13126 4652 -13109 4669
rect -13526 4652 -13509 4669
rect -13166 4652 -13149 4669
rect -13086 4652 -13069 4669
rect -13126 4652 -13109 4669
rect -13166 4652 -13149 4669
rect -13206 4652 -13189 4669
rect -13206 4652 -13189 4669
rect -13246 4652 -13229 4669
rect -13286 4652 -13269 4669
rect -13286 4652 -13269 4669
rect -13046 4652 -13029 4669
rect -13166 4652 -13149 4669
rect -13566 4652 -13549 4669
rect -13326 4652 -13309 4669
rect -13566 4652 -13549 4669
rect -13086 4652 -13069 4669
rect -13086 4652 -13069 4669
rect -13446 4652 -13429 4669
rect -13486 4652 -13469 4669
rect -13526 4652 -13509 4669
rect -13406 4652 -13389 4669
rect -13446 4652 -13429 4669
rect -13486 4652 -13469 4669
rect -13526 4652 -13509 4669
rect -13406 4652 -13389 4669
rect -13366 4652 -13349 4669
rect -13366 4652 -13349 4669
rect -13046 4652 -13029 4669
rect -13366 4652 -13349 4669
rect -13846 4652 -13829 4669
rect -14086 4652 -14069 4669
rect -13606 4652 -13589 4669
rect -14126 4652 -14109 4669
rect -13806 4652 -13789 4669
rect -14046 4652 -14029 4669
rect -13686 4652 -13669 4669
rect -13966 4652 -13949 4669
rect -14166 4652 -14149 4669
rect -14126 4652 -14109 4669
rect -13886 4652 -13869 4669
rect -13966 4652 -13949 4669
rect -13646 4652 -13629 4669
rect -14086 4652 -14069 4669
rect -13766 4652 -13749 4669
rect -13606 4652 -13589 4669
rect -13766 4652 -13749 4669
rect -13846 4652 -13829 4669
rect -13686 4652 -13669 4669
rect -13926 4652 -13909 4669
rect -13646 4652 -13629 4669
rect -14006 4652 -13989 4669
rect -13886 4652 -13869 4669
rect -13726 4652 -13709 4669
rect -14006 4652 -13989 4669
rect -13926 4652 -13909 4669
rect -14166 4652 -14149 4669
rect -13806 4652 -13789 4669
rect -13726 4652 -13709 4669
rect -14046 4652 -14029 4669
rect -13766 4652 -13749 4669
rect -13646 4652 -13629 4669
rect -14126 4652 -14109 4669
rect -14006 4652 -13989 4669
rect -13686 4652 -13669 4669
rect -13806 4652 -13789 4669
rect -13766 4652 -13749 4669
rect -14086 4652 -14069 4669
rect -14166 4652 -14149 4669
rect -14126 4652 -14109 4669
rect -13646 4652 -13629 4669
rect -13846 4652 -13829 4669
rect -14166 4652 -14149 4669
rect -13846 4652 -13829 4669
rect -13886 4652 -13869 4669
rect -13886 4652 -13869 4669
rect -13686 4652 -13669 4669
rect -13726 4652 -13709 4669
rect -13926 4652 -13909 4669
rect -13806 4652 -13789 4669
rect -13606 4652 -13589 4669
rect -13966 4652 -13949 4669
rect -13966 4652 -13949 4669
rect -13926 4652 -13909 4669
rect -14006 4652 -13989 4669
rect -13606 4652 -13589 4669
rect -13726 4652 -13709 4669
rect -14046 4652 -14029 4669
rect -14046 4652 -14029 4669
rect -14086 4652 -14069 4669
rect -10606 4652 -10589 4669
rect -10606 4652 -10589 4669
rect -10606 4652 -10589 4669
rect -10606 4652 -10589 4669
rect -10006 4652 -9989 4669
rect -10006 4652 -9989 4669
rect -10006 4652 -9989 4669
rect -10006 4652 -9989 4669
rect -9926 4652 -9909 4669
rect -9526 4652 -9509 4669
rect -9606 4652 -9589 4669
rect -9846 4652 -9829 4669
rect -9886 4652 -9869 4669
rect -9686 4652 -9669 4669
rect -9726 4652 -9709 4669
rect -9966 4652 -9949 4669
rect -9806 4652 -9789 4669
rect -9886 4652 -9869 4669
rect -9726 4652 -9709 4669
rect -9606 4652 -9589 4669
rect -9726 4652 -9709 4669
rect -9526 4652 -9509 4669
rect -9446 4652 -9429 4669
rect -9606 4652 -9589 4669
rect -9566 4652 -9549 4669
rect -9846 4652 -9829 4669
rect -9766 4652 -9749 4669
rect -9886 4652 -9869 4669
rect -9966 4652 -9949 4669
rect -9566 4652 -9549 4669
rect -9966 4652 -9949 4669
rect -9646 4652 -9629 4669
rect -9646 4652 -9629 4669
rect -9446 4652 -9429 4669
rect -9806 4652 -9789 4669
rect -9926 4652 -9909 4669
rect -9686 4652 -9669 4669
rect -9486 4652 -9469 4669
rect -9806 4652 -9789 4669
rect -9646 4652 -9629 4669
rect -9526 4652 -9509 4669
rect -9926 4652 -9909 4669
rect -9606 4652 -9589 4669
rect -9686 4652 -9669 4669
rect -9446 4652 -9429 4669
rect -9726 4652 -9709 4669
rect -9686 4652 -9669 4669
rect -9766 4652 -9749 4669
rect -9846 4652 -9829 4669
rect -9446 4652 -9429 4669
rect -9886 4652 -9869 4669
rect -9646 4652 -9629 4669
rect -9486 4652 -9469 4669
rect -9806 4652 -9789 4669
rect -9486 4652 -9469 4669
rect -9926 4652 -9909 4669
rect -9486 4652 -9469 4669
rect -9966 4652 -9949 4669
rect -9766 4652 -9749 4669
rect -9526 4652 -9509 4669
rect -9566 4652 -9549 4669
rect -9846 4652 -9829 4669
rect -9766 4652 -9749 4669
rect -9566 4652 -9549 4669
rect -10166 4652 -10149 4669
rect -10046 4652 -10029 4669
rect -10246 4652 -10229 4669
rect -10086 4652 -10069 4669
rect -10126 4652 -10109 4669
rect -10286 4652 -10269 4669
rect -10486 4652 -10469 4669
rect -10526 4652 -10509 4669
rect -10566 4652 -10549 4669
rect -10126 4652 -10109 4669
rect -10326 4652 -10309 4669
rect -10366 4652 -10349 4669
rect -10406 4652 -10389 4669
rect -10446 4652 -10429 4669
rect -10486 4652 -10469 4669
rect -10526 4652 -10509 4669
rect -10566 4652 -10549 4669
rect -10046 4652 -10029 4669
rect -10326 4652 -10309 4669
rect -10366 4652 -10349 4669
rect -10406 4652 -10389 4669
rect -10446 4652 -10429 4669
rect -10566 4652 -10549 4669
rect -10086 4652 -10069 4669
rect -10206 4652 -10189 4669
rect -10166 4652 -10149 4669
rect -10326 4652 -10309 4669
rect -10086 4652 -10069 4669
rect -10366 4652 -10349 4669
rect -10406 4652 -10389 4669
rect -10126 4652 -10109 4669
rect -10446 4652 -10429 4669
rect -10246 4652 -10229 4669
rect -10286 4652 -10269 4669
rect -10286 4652 -10269 4669
rect -10046 4652 -10029 4669
rect -10206 4652 -10189 4669
rect -10486 4652 -10469 4669
rect -10526 4652 -10509 4669
rect -10206 4652 -10189 4669
rect -10566 4652 -10549 4669
rect -10166 4652 -10149 4669
rect -10286 4652 -10269 4669
rect -10366 4652 -10349 4669
rect -10126 4652 -10109 4669
rect -10326 4652 -10309 4669
rect -10446 4652 -10429 4669
rect -10486 4652 -10469 4669
rect -10246 4652 -10229 4669
rect -10526 4652 -10509 4669
rect -10046 4652 -10029 4669
rect -10166 4652 -10149 4669
rect -10206 4652 -10189 4669
rect -10246 4652 -10229 4669
rect -10086 4652 -10069 4669
rect -10406 4652 -10389 4669
rect -11206 4652 -11189 4669
rect -11206 4652 -11189 4669
rect -11206 4652 -11189 4669
rect -11206 4652 -11189 4669
rect -11046 4652 -11029 4669
rect -10846 4652 -10829 4669
rect -11166 4652 -11149 4669
rect -11006 4652 -10989 4669
rect -10686 4652 -10669 4669
rect -10726 4652 -10709 4669
rect -10766 4652 -10749 4669
rect -10726 4652 -10709 4669
rect -10646 4652 -10629 4669
rect -11046 4652 -11029 4669
rect -10686 4652 -10669 4669
rect -10886 4652 -10869 4669
rect -10646 4652 -10629 4669
rect -10926 4652 -10909 4669
rect -10806 4652 -10789 4669
rect -11126 4652 -11109 4669
rect -11086 4652 -11069 4669
rect -10886 4652 -10869 4669
rect -11086 4652 -11069 4669
rect -10966 4652 -10949 4669
rect -11166 4652 -11149 4669
rect -11086 4652 -11069 4669
rect -10766 4652 -10749 4669
rect -10766 4652 -10749 4669
rect -11126 4652 -11109 4669
rect -10646 4652 -10629 4669
rect -10806 4652 -10789 4669
rect -11006 4652 -10989 4669
rect -11126 4652 -11109 4669
rect -10686 4652 -10669 4669
rect -10846 4652 -10829 4669
rect -10966 4652 -10949 4669
rect -10646 4652 -10629 4669
rect -10726 4652 -10709 4669
rect -10886 4652 -10869 4669
rect -10926 4652 -10909 4669
rect -11166 4652 -11149 4669
rect -10966 4652 -10949 4669
rect -10926 4652 -10909 4669
rect -10926 4652 -10909 4669
rect -11086 4652 -11069 4669
rect -10686 4652 -10669 4669
rect -10966 4652 -10949 4669
rect -10806 4652 -10789 4669
rect -11006 4652 -10989 4669
rect -10846 4652 -10829 4669
rect -10846 4652 -10829 4669
rect -11126 4652 -11109 4669
rect -10726 4652 -10709 4669
rect -11046 4652 -11029 4669
rect -11006 4652 -10989 4669
rect -10886 4652 -10869 4669
rect -10766 4652 -10749 4669
rect -11166 4652 -11149 4669
rect -11046 4652 -11029 4669
rect -10806 4652 -10789 4669
rect -11686 4652 -11669 4669
rect -11726 4652 -11709 4669
rect -11406 4652 -11389 4669
rect -11766 4652 -11749 4669
rect -11606 4652 -11589 4669
rect -11526 4652 -11509 4669
rect -11246 4652 -11229 4669
rect -11286 4652 -11269 4669
rect -11326 4652 -11309 4669
rect -11366 4652 -11349 4669
rect -11686 4652 -11669 4669
rect -11446 4652 -11429 4669
rect -11246 4652 -11229 4669
rect -11446 4652 -11429 4669
rect -11646 4652 -11629 4669
rect -11526 4652 -11509 4669
rect -11246 4652 -11229 4669
rect -11286 4652 -11269 4669
rect -11486 4652 -11469 4669
rect -11286 4652 -11269 4669
rect -11246 4652 -11229 4669
rect -11566 4652 -11549 4669
rect -11326 4652 -11309 4669
rect -11646 4652 -11629 4669
rect -11366 4652 -11349 4669
rect -11566 4652 -11549 4669
rect -11606 4652 -11589 4669
rect -11326 4652 -11309 4669
rect -11406 4652 -11389 4669
rect -11766 4652 -11749 4669
rect -11726 4652 -11709 4669
rect -11766 4652 -11749 4669
rect -11526 4652 -11509 4669
rect -11606 4652 -11589 4669
rect -11686 4652 -11669 4669
rect -11686 4652 -11669 4669
rect -11446 4652 -11429 4669
rect -11446 4652 -11429 4669
rect -11366 4652 -11349 4669
rect -11726 4652 -11709 4669
rect -11406 4652 -11389 4669
rect -11646 4652 -11629 4669
rect -11486 4652 -11469 4669
rect -11646 4652 -11629 4669
rect -11406 4652 -11389 4669
rect -11726 4652 -11709 4669
rect -11486 4652 -11469 4669
rect -11566 4652 -11549 4669
rect -11766 4652 -11749 4669
rect -11526 4652 -11509 4669
rect -11286 4652 -11269 4669
rect -11486 4652 -11469 4669
rect -11326 4652 -11309 4669
rect -11366 4652 -11349 4669
rect -11566 4652 -11549 4669
rect -11606 4652 -11589 4669
rect -16606 4652 -16589 4669
rect -16646 4652 -16629 4669
rect -16686 4652 -16669 4669
rect -16726 4652 -16709 4669
rect -16766 4652 -16749 4669
rect -16566 4652 -16549 4669
rect -16606 4652 -16589 4669
rect -16646 4652 -16629 4669
rect -16686 4652 -16669 4669
rect -16726 4652 -16709 4669
rect -16766 4652 -16749 4669
rect -16566 4652 -16549 4669
rect -17126 4652 -17109 4669
rect -16646 4652 -16629 4669
rect -16566 4652 -16549 4669
rect -16766 4652 -16749 4669
rect -16606 4652 -16589 4669
rect -16926 4652 -16909 4669
rect -17006 4652 -16989 4669
rect -16686 4652 -16669 4669
rect -16846 4652 -16829 4669
rect -17086 4652 -17069 4669
rect -16766 4652 -16749 4669
rect -16566 4652 -16549 4669
rect -16886 4652 -16869 4669
rect -16846 4652 -16829 4669
rect -16726 4652 -16709 4669
rect -16886 4652 -16869 4669
rect -16966 4652 -16949 4669
rect -17046 4652 -17029 4669
rect -16806 4652 -16789 4669
rect -16646 4652 -16629 4669
rect -17046 4652 -17029 4669
rect -17046 4652 -17029 4669
rect -17086 4652 -17069 4669
rect -17126 4652 -17109 4669
rect -16806 4652 -16789 4669
rect -17006 4652 -16989 4669
rect -16806 4652 -16789 4669
rect -16846 4652 -16829 4669
rect -16886 4652 -16869 4669
rect -16926 4652 -16909 4669
rect -16966 4652 -16949 4669
rect -17006 4652 -16989 4669
rect -17046 4652 -17029 4669
rect -17086 4652 -17069 4669
rect -17126 4652 -17109 4669
rect -16606 4652 -16589 4669
rect -16726 4652 -16709 4669
rect -16806 4652 -16789 4669
rect -16846 4652 -16829 4669
rect -16886 4652 -16869 4669
rect -16926 4652 -16909 4669
rect -16926 4652 -16909 4669
rect -17086 4652 -17069 4669
rect -16966 4652 -16949 4669
rect -16686 4652 -16669 4669
rect -17006 4652 -16989 4669
rect -17126 4652 -17109 4669
rect -16966 4652 -16949 4669
rect -17686 4652 -17669 4669
rect -17486 4652 -17469 4669
rect -17686 4652 -17669 4669
rect -17166 4652 -17149 4669
rect -17726 4652 -17709 4669
rect -17566 4652 -17549 4669
rect -17486 4652 -17469 4669
rect -17406 4652 -17389 4669
rect -17286 4652 -17269 4669
rect -17446 4652 -17429 4669
rect -17446 4652 -17429 4669
rect -17606 4652 -17589 4669
rect -17566 4652 -17549 4669
rect -17646 4652 -17629 4669
rect -17326 4652 -17309 4669
rect -17726 4652 -17709 4669
rect -17526 4652 -17509 4669
rect -17246 4652 -17229 4669
rect -17326 4652 -17309 4669
rect -17166 4652 -17149 4669
rect -17286 4652 -17269 4669
rect -17526 4652 -17509 4669
rect -17646 4652 -17629 4669
rect -17206 4652 -17189 4669
rect -17406 4652 -17389 4669
rect -17606 4652 -17589 4669
rect -17366 4652 -17349 4669
rect -17206 4652 -17189 4669
rect -17366 4652 -17349 4669
rect -17246 4652 -17229 4669
rect -17246 4652 -17229 4669
rect -17526 4652 -17509 4669
rect -17286 4652 -17269 4669
rect -17566 4652 -17549 4669
rect -17246 4652 -17229 4669
rect -17286 4652 -17269 4669
rect -17326 4652 -17309 4669
rect -17366 4652 -17349 4669
rect -17406 4652 -17389 4669
rect -17446 4652 -17429 4669
rect -17486 4652 -17469 4669
rect -17526 4652 -17509 4669
rect -17566 4652 -17549 4669
rect -17606 4652 -17589 4669
rect -17646 4652 -17629 4669
rect -17686 4652 -17669 4669
rect -17726 4652 -17709 4669
rect -17326 4652 -17309 4669
rect -17606 4652 -17589 4669
rect -17366 4652 -17349 4669
rect -17646 4652 -17629 4669
rect -17166 4652 -17149 4669
rect -17206 4652 -17189 4669
rect -17166 4652 -17149 4669
rect -17206 4652 -17189 4669
rect -17406 4652 -17389 4669
rect -17686 4652 -17669 4669
rect -17446 4652 -17429 4669
rect -17726 4652 -17709 4669
rect -17486 4652 -17469 4669
rect -17846 4652 -17829 4669
rect -17766 4652 -17749 4669
rect -17766 4652 -17749 4669
rect -17806 4652 -17789 4669
rect -17846 4652 -17829 4669
rect -18046 4652 -18029 4669
rect -17806 4652 -17789 4669
rect -17926 4652 -17909 4669
rect -17846 4652 -17829 4669
rect -17886 4652 -17869 4669
rect -18086 4652 -18069 4669
rect -18126 4652 -18109 4669
rect -18326 4652 -18309 4669
rect -18126 4652 -18109 4669
rect -17766 4652 -17749 4669
rect -18166 4652 -18149 4669
rect -18126 4652 -18109 4669
rect -18206 4652 -18189 4669
rect -18166 4652 -18149 4669
rect -17886 4652 -17869 4669
rect -18286 4652 -18269 4669
rect -18246 4652 -18229 4669
rect -17966 4652 -17949 4669
rect -18286 4652 -18269 4669
rect -17806 4652 -17789 4669
rect -18006 4652 -17989 4669
rect -18246 4652 -18229 4669
rect -18326 4652 -18309 4669
rect -17926 4652 -17909 4669
rect -18206 4652 -18189 4669
rect -18166 4652 -18149 4669
rect -17806 4652 -17789 4669
rect -17926 4652 -17909 4669
rect -18246 4652 -18229 4669
rect -17886 4652 -17869 4669
rect -18086 4652 -18069 4669
rect -18006 4652 -17989 4669
rect -18326 4652 -18309 4669
rect -18126 4652 -18109 4669
rect -17966 4652 -17949 4669
rect -18046 4652 -18029 4669
rect -17926 4652 -17909 4669
rect -17886 4652 -17869 4669
rect -18206 4652 -18189 4669
rect -17966 4652 -17949 4669
rect -18046 4652 -18029 4669
rect -18246 4652 -18229 4669
rect -18006 4652 -17989 4669
rect -18286 4652 -18269 4669
rect -17966 4652 -17949 4669
rect -17766 4652 -17749 4669
rect -18286 4652 -18269 4669
rect -18166 4652 -18149 4669
rect -18046 4652 -18029 4669
rect -18006 4652 -17989 4669
rect -18086 4652 -18069 4669
rect -17846 4652 -17829 4669
rect -18326 4652 -18309 4669
rect -18206 4652 -18189 4669
rect -18086 4652 -18069 4669
rect -18366 4652 -18349 4669
rect -18846 4652 -18829 4669
rect -18766 4652 -18749 4669
rect -18566 4652 -18549 4669
rect -18686 4652 -18669 4669
rect -18646 4652 -18629 4669
rect -18406 4652 -18389 4669
rect -18886 4652 -18869 4669
rect -18806 4652 -18789 4669
rect -18606 4652 -18589 4669
rect -18446 4652 -18429 4669
rect -18366 4652 -18349 4669
rect -18606 4652 -18589 4669
rect -18406 4652 -18389 4669
rect -18726 4652 -18709 4669
rect -18486 4652 -18469 4669
rect -18486 4652 -18469 4669
rect -18846 4652 -18829 4669
rect -18646 4652 -18629 4669
rect -18526 4652 -18509 4669
rect -18926 4652 -18909 4669
rect -18806 4652 -18789 4669
rect -18446 4652 -18429 4669
rect -18926 4652 -18909 4669
rect -18886 4652 -18869 4669
rect -18766 4652 -18749 4669
rect -18686 4652 -18669 4669
rect -18526 4652 -18509 4669
rect -18566 4652 -18549 4669
rect -18726 4652 -18709 4669
rect -18766 4652 -18749 4669
rect -18806 4652 -18789 4669
rect -18366 4652 -18349 4669
rect -18846 4652 -18829 4669
rect -18886 4652 -18869 4669
rect -18926 4652 -18909 4669
rect -18686 4652 -18669 4669
rect -18726 4652 -18709 4669
rect -18766 4652 -18749 4669
rect -18806 4652 -18789 4669
rect -18846 4652 -18829 4669
rect -18886 4652 -18869 4669
rect -18926 4652 -18909 4669
rect -18366 4652 -18349 4669
rect -18406 4652 -18389 4669
rect -18446 4652 -18429 4669
rect -18406 4652 -18389 4669
rect -18486 4652 -18469 4669
rect -18526 4652 -18509 4669
rect -18446 4652 -18429 4669
rect -18566 4652 -18549 4669
rect -18606 4652 -18589 4669
rect -18486 4652 -18469 4669
rect -18646 4652 -18629 4669
rect -18526 4652 -18509 4669
rect -18566 4652 -18549 4669
rect -18606 4652 -18589 4669
rect -18646 4652 -18629 4669
rect -18686 4652 -18669 4669
rect -18726 4652 -18709 4669
rect -15366 4652 -15349 4669
rect -15366 4652 -15349 4669
rect -15366 4652 -15349 4669
rect -15366 4652 -15349 4669
rect -14766 4652 -14749 4669
rect -14766 4652 -14749 4669
rect -14766 4652 -14749 4669
rect -14766 4652 -14749 4669
rect -14726 4652 -14709 4669
rect -14646 4652 -14629 4669
rect -14246 4652 -14229 4669
rect -14286 4652 -14269 4669
rect -14446 4652 -14429 4669
rect -14726 4652 -14709 4669
rect -14606 4652 -14589 4669
rect -14686 4652 -14669 4669
rect -14726 4652 -14709 4669
rect -14326 4652 -14309 4669
rect -14206 4652 -14189 4669
rect -14366 4652 -14349 4669
rect -14486 4652 -14469 4669
rect -14486 4652 -14469 4669
rect -14566 4652 -14549 4669
rect -14686 4652 -14669 4669
rect -14566 4652 -14549 4669
rect -14246 4652 -14229 4669
rect -14486 4652 -14469 4669
rect -14406 4652 -14389 4669
rect -14286 4652 -14269 4669
rect -14366 4652 -14349 4669
rect -14526 4652 -14509 4669
rect -14326 4652 -14309 4669
rect -14286 4652 -14269 4669
rect -14646 4652 -14629 4669
rect -14726 4652 -14709 4669
rect -14446 4652 -14429 4669
rect -14606 4652 -14589 4669
rect -14646 4652 -14629 4669
rect -14646 4652 -14629 4669
rect -14486 4652 -14469 4669
rect -14366 4652 -14349 4669
rect -14526 4652 -14509 4669
rect -14686 4652 -14669 4669
rect -14406 4652 -14389 4669
rect -14566 4652 -14549 4669
rect -14326 4652 -14309 4669
rect -14246 4652 -14229 4669
rect -14286 4652 -14269 4669
rect -14406 4652 -14389 4669
rect -14446 4652 -14429 4669
rect -14606 4652 -14589 4669
rect -14206 4652 -14189 4669
rect -14526 4652 -14509 4669
rect -14446 4652 -14429 4669
rect -14326 4652 -14309 4669
rect -14566 4652 -14549 4669
rect -14406 4652 -14389 4669
rect -14206 4652 -14189 4669
rect -14366 4652 -14349 4669
rect -14526 4652 -14509 4669
rect -14246 4652 -14229 4669
rect -14606 4652 -14589 4669
rect -14686 4652 -14669 4669
rect -14206 4652 -14189 4669
rect -15126 4652 -15109 4669
rect -15166 4652 -15149 4669
rect -15206 4652 -15189 4669
rect -15246 4652 -15229 4669
rect -15286 4652 -15269 4669
rect -15326 4652 -15309 4669
rect -14846 4652 -14829 4669
rect -15166 4652 -15149 4669
rect -15206 4652 -15189 4669
rect -14886 4652 -14869 4669
rect -14926 4652 -14909 4669
rect -14966 4652 -14949 4669
rect -15006 4652 -14989 4669
rect -15046 4652 -15029 4669
rect -15006 4652 -14989 4669
rect -14806 4652 -14789 4669
rect -14846 4652 -14829 4669
rect -14886 4652 -14869 4669
rect -14926 4652 -14909 4669
rect -14966 4652 -14949 4669
rect -15006 4652 -14989 4669
rect -15046 4652 -15029 4669
rect -15086 4652 -15069 4669
rect -15246 4652 -15229 4669
rect -14806 4652 -14789 4669
rect -15286 4652 -15269 4669
rect -14846 4652 -14829 4669
rect -15326 4652 -15309 4669
rect -15326 4652 -15309 4669
rect -15046 4652 -15029 4669
rect -15166 4652 -15149 4669
rect -15006 4652 -14989 4669
rect -15126 4652 -15109 4669
rect -15286 4652 -15269 4669
rect -15126 4652 -15109 4669
rect -14806 4652 -14789 4669
rect -15206 4652 -15189 4669
rect -15086 4652 -15069 4669
rect -15326 4652 -15309 4669
rect -14846 4652 -14829 4669
rect -15086 4652 -15069 4669
rect -15126 4652 -15109 4669
rect -15246 4652 -15229 4669
rect -14886 4652 -14869 4669
rect -14886 4652 -14869 4669
rect -15166 4652 -15149 4669
rect -14926 4652 -14909 4669
rect -14806 4652 -14789 4669
rect -15206 4652 -15189 4669
rect -14966 4652 -14949 4669
rect -15046 4652 -15029 4669
rect -14926 4652 -14909 4669
rect -15286 4652 -15269 4669
rect -15246 4652 -15229 4669
rect -15086 4652 -15069 4669
rect -14966 4652 -14949 4669
rect -15966 4652 -15949 4669
rect -15966 4652 -15949 4669
rect -15966 4652 -15949 4669
rect -15966 4652 -15949 4669
rect -15646 4652 -15629 4669
rect -15806 4652 -15789 4669
rect -15766 4652 -15749 4669
rect -15686 4652 -15669 4669
rect -15726 4652 -15709 4669
rect -15406 4652 -15389 4669
rect -15846 4652 -15829 4669
rect -15446 4652 -15429 4669
rect -15766 4652 -15749 4669
rect -15526 4652 -15509 4669
rect -15486 4652 -15469 4669
rect -15526 4652 -15509 4669
rect -15606 4652 -15589 4669
rect -15926 4652 -15909 4669
rect -15446 4652 -15429 4669
rect -15526 4652 -15509 4669
rect -15526 4652 -15509 4669
rect -15406 4652 -15389 4669
rect -15566 4652 -15549 4669
rect -15486 4652 -15469 4669
rect -15606 4652 -15589 4669
rect -15646 4652 -15629 4669
rect -15686 4652 -15669 4669
rect -15926 4652 -15909 4669
rect -15726 4652 -15709 4669
rect -15886 4652 -15869 4669
rect -15566 4652 -15549 4669
rect -15446 4652 -15429 4669
rect -15806 4652 -15789 4669
rect -15766 4652 -15749 4669
rect -15566 4652 -15549 4669
rect -15846 4652 -15829 4669
rect -15606 4652 -15589 4669
rect -15726 4652 -15709 4669
rect -15646 4652 -15629 4669
rect -15766 4652 -15749 4669
rect -15806 4652 -15789 4669
rect -15406 4652 -15389 4669
rect -15886 4652 -15869 4669
rect -15846 4652 -15829 4669
rect -15446 4652 -15429 4669
rect -15846 4652 -15829 4669
rect -15726 4652 -15709 4669
rect -15566 4652 -15549 4669
rect -15926 4652 -15909 4669
rect -15486 4652 -15469 4669
rect -15686 4652 -15669 4669
rect -15806 4652 -15789 4669
rect -15406 4652 -15389 4669
rect -15606 4652 -15589 4669
rect -15886 4652 -15869 4669
rect -15646 4652 -15629 4669
rect -15486 4652 -15469 4669
rect -15886 4652 -15869 4669
rect -15686 4652 -15669 4669
rect -15926 4652 -15909 4669
rect -16526 4652 -16509 4669
rect -16166 4652 -16149 4669
rect -16006 4652 -15989 4669
rect -16526 4652 -16509 4669
rect -16046 4652 -16029 4669
rect -16006 4652 -15989 4669
rect -16086 4652 -16069 4669
rect -16366 4652 -16349 4669
rect -16126 4652 -16109 4669
rect -16166 4652 -16149 4669
rect -16206 4652 -16189 4669
rect -16006 4652 -15989 4669
rect -16246 4652 -16229 4669
rect -16286 4652 -16269 4669
rect -16246 4652 -16229 4669
rect -16326 4652 -16309 4669
rect -16366 4652 -16349 4669
rect -16526 4652 -16509 4669
rect -16086 4652 -16069 4669
rect -16126 4652 -16109 4669
rect -16326 4652 -16309 4669
rect -16406 4652 -16389 4669
rect -16206 4652 -16189 4669
rect -16206 4652 -16189 4669
rect -16486 4652 -16469 4669
rect -16486 4652 -16469 4669
rect -16006 4652 -15989 4669
rect -16446 4652 -16429 4669
rect -16286 4652 -16269 4669
rect -16166 4652 -16149 4669
rect -16246 4652 -16229 4669
rect -16046 4652 -16029 4669
rect -16166 4652 -16149 4669
rect -16446 4652 -16429 4669
rect -16286 4652 -16269 4669
rect -16366 4652 -16349 4669
rect -16406 4652 -16389 4669
rect -16526 4652 -16509 4669
rect -16446 4652 -16429 4669
rect -16286 4652 -16269 4669
rect -16326 4652 -16309 4669
rect -16406 4652 -16389 4669
rect -16326 4652 -16309 4669
rect -16486 4652 -16469 4669
rect -16206 4652 -16189 4669
rect -16126 4652 -16109 4669
rect -16046 4652 -16029 4669
rect -16086 4652 -16069 4669
rect -16366 4652 -16349 4669
rect -16046 4652 -16029 4669
rect -16246 4652 -16229 4669
rect -16086 4652 -16069 4669
rect -16406 4652 -16389 4669
rect -16126 4652 -16109 4669
rect -16446 4652 -16429 4669
rect -16486 4652 -16469 4669
rect -18166 3163 -18149 3180
rect -18846 3163 -18829 3180
rect -18486 3163 -18469 3180
rect -18686 3163 -18669 3180
rect -18726 3163 -18709 3180
rect -18446 3163 -18429 3180
rect -18446 3163 -18429 3180
rect -18886 3163 -18869 3180
rect -18566 3163 -18549 3180
rect -18486 3163 -18469 3180
rect -18886 3163 -18869 3180
rect -18886 3163 -18869 3180
rect -18606 3163 -18589 3180
rect -18766 3163 -18749 3180
rect -18686 3163 -18669 3180
rect -18566 3163 -18549 3180
rect -18486 3163 -18469 3180
rect -18646 3163 -18629 3180
rect -18606 3163 -18589 3180
rect -18406 3163 -18389 3180
rect -18926 3163 -18909 3180
rect -18926 3163 -18909 3180
rect -18406 3163 -18389 3180
rect -18686 3163 -18669 3180
rect -18726 3163 -18709 3180
rect -18446 3163 -18429 3180
rect -18606 3163 -18589 3180
rect -18726 3163 -18709 3180
rect -18406 3163 -18389 3180
rect -18806 3163 -18789 3180
rect -18566 3163 -18549 3180
rect -18806 3163 -18789 3180
rect -18526 3163 -18509 3180
rect -18846 3163 -18829 3180
rect -18446 3163 -18429 3180
rect -18766 3163 -18749 3180
rect -18646 3163 -18629 3180
rect -18846 3163 -18829 3180
rect -18926 3163 -18909 3180
rect -18686 3163 -18669 3180
rect -18646 3163 -18629 3180
rect -18926 3163 -18909 3180
rect -18886 3163 -18869 3180
rect -18766 3163 -18749 3180
rect -18486 3163 -18469 3180
rect -18766 3163 -18749 3180
rect -18726 3163 -18709 3180
rect -18526 3163 -18509 3180
rect -18526 3163 -18509 3180
rect -18846 3163 -18829 3180
rect -18526 3163 -18509 3180
rect -18566 3163 -18549 3180
rect -18646 3163 -18629 3180
rect -18406 3163 -18389 3180
rect -18606 3163 -18589 3180
rect -18806 3163 -18789 3180
rect -18806 3163 -18789 3180
rect -14366 3163 -14349 3180
rect -14526 3163 -14509 3180
rect -14206 3163 -14189 3180
rect -14326 3163 -14309 3180
rect -14286 3163 -14269 3180
rect -14326 3163 -14309 3180
rect -14246 3163 -14229 3180
rect -14486 3163 -14469 3180
rect -14286 3163 -14269 3180
rect -14566 3163 -14549 3180
rect -14566 3163 -14549 3180
rect -14406 3163 -14389 3180
rect -14286 3163 -14269 3180
rect -14406 3163 -14389 3180
rect -14366 3163 -14349 3180
rect -14246 3163 -14229 3180
rect -14446 3163 -14429 3180
rect -14446 3163 -14429 3180
rect -14326 3163 -14309 3180
rect -14486 3163 -14469 3180
rect -14606 3163 -14589 3180
rect -14206 3163 -14189 3180
rect -14246 3163 -14229 3180
rect -14486 3163 -14469 3180
rect -14206 3163 -14189 3180
rect -14606 3163 -14589 3180
rect -14526 3163 -14509 3180
rect -14406 3163 -14389 3180
rect -14606 3163 -14589 3180
rect -14486 3163 -14469 3180
rect -14566 3163 -14549 3180
rect -14606 3163 -14589 3180
rect -14366 3163 -14349 3180
rect -14446 3163 -14429 3180
rect -14246 3163 -14229 3180
rect -14206 3163 -14189 3180
rect -14526 3163 -14509 3180
rect -14526 3163 -14509 3180
rect -14286 3163 -14269 3180
rect -14446 3163 -14429 3180
rect -14366 3163 -14349 3180
rect -14406 3163 -14389 3180
rect -14566 3163 -14549 3180
rect -14326 3163 -14309 3180
rect -15166 3163 -15149 3180
rect -15166 3163 -15149 3180
rect -15166 3163 -15149 3180
rect -15166 3163 -15149 3180
rect -15126 3163 -15109 3180
rect -14806 3163 -14789 3180
rect -15086 3163 -15069 3180
rect -14846 3163 -14829 3180
rect -15086 3163 -15069 3180
rect -14766 3163 -14749 3180
rect -15126 3163 -15109 3180
rect -14766 3163 -14749 3180
rect -14886 3163 -14869 3180
rect -14886 3163 -14869 3180
rect -14766 3163 -14749 3180
rect -15046 3163 -15029 3180
rect -14926 3163 -14909 3180
rect -14766 3163 -14749 3180
rect -14806 3163 -14789 3180
rect -15126 3163 -15109 3180
rect -14966 3163 -14949 3180
rect -15006 3163 -14989 3180
rect -15046 3163 -15029 3180
rect -14926 3163 -14909 3180
rect -15086 3163 -15069 3180
rect -14966 3163 -14949 3180
rect -14726 3163 -14709 3180
rect -14646 3163 -14629 3180
rect -14846 3163 -14829 3180
rect -15126 3163 -15109 3180
rect -14726 3163 -14709 3180
rect -14686 3163 -14669 3180
rect -14886 3163 -14869 3180
rect -14726 3163 -14709 3180
rect -14926 3163 -14909 3180
rect -14966 3163 -14949 3180
rect -15006 3163 -14989 3180
rect -15046 3163 -15029 3180
rect -15006 3163 -14989 3180
rect -14686 3163 -14669 3180
rect -14806 3163 -14789 3180
rect -14846 3163 -14829 3180
rect -14886 3163 -14869 3180
rect -14926 3163 -14909 3180
rect -14966 3163 -14949 3180
rect -15006 3163 -14989 3180
rect -15046 3163 -15029 3180
rect -14646 3163 -14629 3180
rect -14726 3163 -14709 3180
rect -15086 3163 -15069 3180
rect -14646 3163 -14629 3180
rect -14806 3163 -14789 3180
rect -14646 3163 -14629 3180
rect -14686 3163 -14669 3180
rect -14846 3163 -14829 3180
rect -14686 3163 -14669 3180
rect -15286 3163 -15269 3180
rect -15606 3163 -15589 3180
rect -15406 3163 -15389 3180
rect -15326 3163 -15309 3180
rect -15686 3163 -15669 3180
rect -15246 3163 -15229 3180
rect -15286 3163 -15269 3180
rect -15566 3163 -15549 3180
rect -15366 3163 -15349 3180
rect -15206 3163 -15189 3180
rect -15406 3163 -15389 3180
rect -15446 3163 -15429 3180
rect -15566 3163 -15549 3180
rect -15686 3163 -15669 3180
rect -15326 3163 -15309 3180
rect -15566 3163 -15549 3180
rect -15206 3163 -15189 3180
rect -15686 3163 -15669 3180
rect -15486 3163 -15469 3180
rect -15446 3163 -15429 3180
rect -15486 3163 -15469 3180
rect -15566 3163 -15549 3180
rect -15366 3163 -15349 3180
rect -15366 3163 -15349 3180
rect -15486 3163 -15469 3180
rect -15646 3163 -15629 3180
rect -15606 3163 -15589 3180
rect -15406 3163 -15389 3180
rect -15206 3163 -15189 3180
rect -15606 3163 -15589 3180
rect -15606 3163 -15589 3180
rect -15526 3163 -15509 3180
rect -15646 3163 -15629 3180
rect -15326 3163 -15309 3180
rect -15526 3163 -15509 3180
rect -15646 3163 -15629 3180
rect -15446 3163 -15429 3180
rect -15526 3163 -15509 3180
rect -15206 3163 -15189 3180
rect -15406 3163 -15389 3180
rect -15286 3163 -15269 3180
rect -15246 3163 -15229 3180
rect -15646 3163 -15629 3180
rect -15686 3163 -15669 3180
rect -15246 3163 -15229 3180
rect -15246 3163 -15229 3180
rect -15286 3163 -15269 3180
rect -15446 3163 -15429 3180
rect -15486 3163 -15469 3180
rect -15526 3163 -15509 3180
rect -15366 3163 -15349 3180
rect -15326 3163 -15309 3180
rect -16246 3163 -16229 3180
rect -16246 3163 -16229 3180
rect -16246 3163 -16229 3180
rect -16246 3163 -16229 3180
rect -15806 3163 -15789 3180
rect -16126 3163 -16109 3180
rect -15806 3163 -15789 3180
rect -15926 3163 -15909 3180
rect -16126 3163 -16109 3180
rect -16206 3163 -16189 3180
rect -16006 3163 -15989 3180
rect -15766 3163 -15749 3180
rect -15886 3163 -15869 3180
rect -16046 3163 -16029 3180
rect -15926 3163 -15909 3180
rect -15726 3163 -15709 3180
rect -15966 3163 -15949 3180
rect -15846 3163 -15829 3180
rect -16166 3163 -16149 3180
rect -15726 3163 -15709 3180
rect -15966 3163 -15949 3180
rect -16086 3163 -16069 3180
rect -16046 3163 -16029 3180
rect -16166 3163 -16149 3180
rect -16206 3163 -16189 3180
rect -15726 3163 -15709 3180
rect -16086 3163 -16069 3180
rect -15926 3163 -15909 3180
rect -16166 3163 -16149 3180
rect -15846 3163 -15829 3180
rect -15766 3163 -15749 3180
rect -16126 3163 -16109 3180
rect -16006 3163 -15989 3180
rect -16086 3163 -16069 3180
rect -15806 3163 -15789 3180
rect -15966 3163 -15949 3180
rect -16086 3163 -16069 3180
rect -15726 3163 -15709 3180
rect -16006 3163 -15989 3180
rect -16126 3163 -16109 3180
rect -16206 3163 -16189 3180
rect -15806 3163 -15789 3180
rect -15886 3163 -15869 3180
rect -15926 3163 -15909 3180
rect -15766 3163 -15749 3180
rect -15846 3163 -15829 3180
rect -15886 3163 -15869 3180
rect -16166 3163 -16149 3180
rect -16046 3163 -16029 3180
rect -16006 3163 -15989 3180
rect -16206 3163 -16189 3180
rect -15766 3163 -15749 3180
rect -15846 3163 -15829 3180
rect -15966 3163 -15949 3180
rect -16046 3163 -16029 3180
rect -15886 3163 -15869 3180
rect -16406 3163 -16389 3180
rect -16446 3163 -16429 3180
rect -16766 3163 -16749 3180
rect -16526 3163 -16509 3180
rect -16486 3163 -16469 3180
rect -16486 3163 -16469 3180
rect -16566 3163 -16549 3180
rect -16286 3163 -16269 3180
rect -16326 3163 -16309 3180
rect -16726 3163 -16709 3180
rect -16286 3163 -16269 3180
rect -16406 3163 -16389 3180
rect -16326 3163 -16309 3180
rect -16646 3163 -16629 3180
rect -16366 3163 -16349 3180
rect -16526 3163 -16509 3180
rect -16646 3163 -16629 3180
rect -16606 3163 -16589 3180
rect -16766 3163 -16749 3180
rect -16566 3163 -16549 3180
rect -16366 3163 -16349 3180
rect -16606 3163 -16589 3180
rect -16366 3163 -16349 3180
rect -16566 3163 -16549 3180
rect -16766 3163 -16749 3180
rect -16326 3163 -16309 3180
rect -16446 3163 -16429 3180
rect -16606 3163 -16589 3180
rect -16726 3163 -16709 3180
rect -16366 3163 -16349 3180
rect -16606 3163 -16589 3180
rect -16526 3163 -16509 3180
rect -16486 3163 -16469 3180
rect -16406 3163 -16389 3180
rect -16526 3163 -16509 3180
rect -16446 3163 -16429 3180
rect -16686 3163 -16669 3180
rect -16486 3163 -16469 3180
rect -16646 3163 -16629 3180
rect -16286 3163 -16269 3180
rect -16646 3163 -16629 3180
rect -16726 3163 -16709 3180
rect -16326 3163 -16309 3180
rect -16766 3163 -16749 3180
rect -16686 3163 -16669 3180
rect -16446 3163 -16429 3180
rect -16286 3163 -16269 3180
rect -16406 3163 -16389 3180
rect -16566 3163 -16549 3180
rect -16686 3163 -16669 3180
rect -16726 3163 -16709 3180
rect -16686 3163 -16669 3180
rect -16806 3163 -16789 3180
rect -17166 3163 -17149 3180
rect -17206 3163 -17189 3180
rect -17126 3163 -17109 3180
rect -17046 3163 -17029 3180
rect -16846 3163 -16829 3180
rect -17246 3163 -17229 3180
rect -16926 3163 -16909 3180
rect -17166 3163 -17149 3180
rect -17046 3163 -17029 3180
rect -16846 3163 -16829 3180
rect -17086 3163 -17069 3180
rect -17286 3163 -17269 3180
rect -17006 3163 -16989 3180
rect -17286 3163 -17269 3180
rect -16886 3163 -16869 3180
rect -17046 3163 -17029 3180
rect -17206 3163 -17189 3180
rect -17006 3163 -16989 3180
rect -16966 3163 -16949 3180
rect -17286 3163 -17269 3180
rect -16886 3163 -16869 3180
rect -17246 3163 -17229 3180
rect -16886 3163 -16869 3180
rect -17206 3163 -17189 3180
rect -16806 3163 -16789 3180
rect -17086 3163 -17069 3180
rect -17126 3163 -17109 3180
rect -16966 3163 -16949 3180
rect -17126 3163 -17109 3180
rect -16926 3163 -16909 3180
rect -16846 3163 -16829 3180
rect -17286 3163 -17269 3180
rect -17006 3163 -16989 3180
rect -16886 3163 -16869 3180
rect -16966 3163 -16949 3180
rect -17126 3163 -17109 3180
rect -16806 3163 -16789 3180
rect -16926 3163 -16909 3180
rect -17006 3163 -16989 3180
rect -16966 3163 -16949 3180
rect -17046 3163 -17029 3180
rect -17086 3163 -17069 3180
rect -17246 3163 -17229 3180
rect -17166 3163 -17149 3180
rect -16846 3163 -16829 3180
rect -17086 3163 -17069 3180
rect -16806 3163 -16789 3180
rect -16926 3163 -16909 3180
rect -17206 3163 -17189 3180
rect -17166 3163 -17149 3180
rect -17246 3163 -17229 3180
rect -17566 3163 -17549 3180
rect -17846 3163 -17829 3180
rect -17446 3163 -17429 3180
rect -17766 3163 -17749 3180
rect -17686 3163 -17669 3180
rect -17606 3163 -17589 3180
rect -17686 3163 -17669 3180
rect -17726 3163 -17709 3180
rect -17486 3163 -17469 3180
rect -17406 3163 -17389 3180
rect -17486 3163 -17469 3180
rect -17566 3163 -17549 3180
rect -17486 3163 -17469 3180
rect -17526 3163 -17509 3180
rect -17646 3163 -17629 3180
rect -17326 3163 -17309 3180
rect -17726 3163 -17709 3180
rect -17806 3163 -17789 3180
rect -17766 3163 -17749 3180
rect -17526 3163 -17509 3180
rect -17526 3163 -17509 3180
rect -17566 3163 -17549 3180
rect -17606 3163 -17589 3180
rect -17766 3163 -17749 3180
rect -17326 3163 -17309 3180
rect -17846 3163 -17829 3180
rect -17686 3163 -17669 3180
rect -17366 3163 -17349 3180
rect -17486 3163 -17469 3180
rect -17846 3163 -17829 3180
rect -17766 3163 -17749 3180
rect -17726 3163 -17709 3180
rect -17366 3163 -17349 3180
rect -17566 3163 -17549 3180
rect -17406 3163 -17389 3180
rect -17526 3163 -17509 3180
rect -17646 3163 -17629 3180
rect -17446 3163 -17429 3180
rect -17686 3163 -17669 3180
rect -17326 3163 -17309 3180
rect -17406 3163 -17389 3180
rect -17446 3163 -17429 3180
rect -17606 3163 -17589 3180
rect -17606 3163 -17589 3180
rect -17806 3163 -17789 3180
rect -17406 3163 -17389 3180
rect -17806 3163 -17789 3180
rect -17726 3163 -17709 3180
rect -17326 3163 -17309 3180
rect -17646 3163 -17629 3180
rect -17366 3163 -17349 3180
rect -17646 3163 -17629 3180
rect -17446 3163 -17429 3180
rect -17806 3163 -17789 3180
rect -17366 3163 -17349 3180
rect -17846 3163 -17829 3180
rect -18166 3163 -18149 3180
rect -17926 3163 -17909 3180
rect -17966 3163 -17949 3180
rect -18006 3163 -17989 3180
rect -17886 3163 -17869 3180
rect -18206 3163 -18189 3180
rect -17926 3163 -17909 3180
rect -18046 3163 -18029 3180
rect -18326 3163 -18309 3180
rect -18286 3163 -18269 3180
rect -18286 3163 -18269 3180
rect -18366 3163 -18349 3180
rect -18166 3163 -18149 3180
rect -18006 3163 -17989 3180
rect -18126 3163 -18109 3180
rect -18046 3163 -18029 3180
rect -18366 3163 -18349 3180
rect -17926 3163 -17909 3180
rect -18046 3163 -18029 3180
rect -18246 3163 -18229 3180
rect -18246 3163 -18229 3180
rect -17926 3163 -17909 3180
rect -18366 3163 -18349 3180
rect -18126 3163 -18109 3180
rect -18126 3163 -18109 3180
rect -17966 3163 -17949 3180
rect -18326 3163 -18309 3180
rect -18206 3163 -18189 3180
rect -18246 3163 -18229 3180
rect -18086 3163 -18069 3180
rect -17966 3163 -17949 3180
rect -18246 3163 -18229 3180
rect -17966 3163 -17949 3180
rect -18326 3163 -18309 3180
rect -18326 3163 -18309 3180
rect -17886 3163 -17869 3180
rect -18046 3163 -18029 3180
rect -18126 3163 -18109 3180
rect -18206 3163 -18189 3180
rect -18286 3163 -18269 3180
rect -17886 3163 -17869 3180
rect -18206 3163 -18189 3180
rect -18166 3163 -18149 3180
rect -18086 3163 -18069 3180
rect -18286 3163 -18269 3180
rect -17886 3163 -17869 3180
rect -18006 3163 -17989 3180
rect -18006 3163 -17989 3180
rect -18366 3163 -18349 3180
rect -18086 3163 -18069 3180
rect -18086 3163 -18069 3180
rect -16733 2394 -16716 2411
rect -17373 2394 -17356 2411
rect -16653 2394 -16636 2411
rect -16613 2394 -16596 2411
rect -17213 2394 -17196 2411
rect -17253 2394 -17236 2411
rect -16813 2394 -16796 2411
rect -17413 2394 -17396 2411
rect -16853 2394 -16836 2411
rect -17453 2394 -17436 2411
rect -16853 2394 -16836 2411
rect -17133 2394 -17116 2411
rect -17413 2394 -17396 2411
rect -17453 2394 -17436 2411
rect -17293 2394 -17276 2411
rect -16573 2394 -16556 2411
rect -16893 2394 -16876 2411
rect -17293 2394 -17276 2411
rect -16573 2394 -16556 2411
rect -16693 2394 -16676 2411
rect -17253 2394 -17236 2411
rect -16693 2394 -16676 2411
rect -16933 2394 -16916 2411
rect -17173 2394 -17156 2411
rect -16773 2394 -16756 2411
rect -17053 2394 -17036 2411
rect -16973 2394 -16956 2411
rect -17333 2394 -17316 2411
rect -17173 2394 -17156 2411
rect -16933 2394 -16916 2411
rect -17013 2394 -16996 2411
rect -17333 2394 -17316 2411
rect -17213 2394 -17196 2411
rect -17013 2394 -16996 2411
rect -16893 2394 -16876 2411
rect -17133 2394 -17116 2411
rect -17093 2394 -17076 2411
rect -17053 2394 -17036 2411
rect -16773 2394 -16756 2411
rect -16613 2394 -16596 2411
rect -16813 2394 -16796 2411
rect -16973 2394 -16956 2411
rect -16653 2394 -16636 2411
rect -17373 2394 -17356 2411
rect -16733 2394 -16716 2411
rect -17093 2394 -17076 2411
rect -15373 2394 -15356 2411
rect -15373 2394 -15356 2411
rect -16333 2394 -16316 2411
rect -16053 2394 -16036 2411
rect -15493 2394 -15476 2411
rect -15693 2394 -15676 2411
rect -16373 2394 -16356 2411
rect -15453 2394 -15436 2411
rect -15973 2394 -15956 2411
rect -15853 2394 -15836 2411
rect -16093 2394 -16076 2411
rect -15893 2394 -15876 2411
rect -15533 2394 -15516 2411
rect -16133 2394 -16116 2411
rect -15733 2394 -15716 2411
rect -16253 2394 -16236 2411
rect -15773 2394 -15756 2411
rect -15893 2394 -15876 2411
rect -16133 2394 -16116 2411
rect -15573 2394 -15556 2411
rect -16293 2394 -16276 2411
rect -15493 2394 -15476 2411
rect -16173 2394 -16156 2411
rect -16333 2394 -16316 2411
rect -15933 2394 -15916 2411
rect -16173 2394 -16156 2411
rect -15573 2394 -15556 2411
rect -15853 2394 -15836 2411
rect -16373 2394 -16356 2411
rect -16093 2394 -16076 2411
rect -15413 2394 -15396 2411
rect -15613 2394 -15596 2411
rect -15613 2394 -15596 2411
rect -16013 2394 -15996 2411
rect -16213 2394 -16196 2411
rect -15653 2394 -15636 2411
rect -15413 2394 -15396 2411
rect -15813 2394 -15796 2411
rect -15693 2394 -15676 2411
rect -15973 2394 -15956 2411
rect -15813 2394 -15796 2411
rect -15453 2394 -15436 2411
rect -15733 2394 -15716 2411
rect -16253 2394 -16236 2411
rect -15533 2394 -15516 2411
rect -15773 2394 -15756 2411
rect -16013 2394 -15996 2411
rect -15933 2394 -15916 2411
rect -16213 2394 -16196 2411
rect -16293 2394 -16276 2411
rect -15653 2394 -15636 2411
rect -16053 2394 -16036 2411
rect -16533 2394 -16516 2411
rect -16493 2394 -16476 2411
rect -16413 2394 -16396 2411
rect -16533 2394 -16516 2411
rect -16413 2394 -16396 2411
rect -16453 2394 -16436 2411
rect -16453 2394 -16436 2411
rect -16493 2394 -16476 2411
rect -15213 2394 -15196 2411
rect -14693 2394 -14676 2411
rect -15173 2394 -15156 2411
rect -14373 2394 -14356 2411
rect -14213 2394 -14196 2411
rect -14213 2394 -14196 2411
rect -14893 2394 -14876 2411
rect -15293 2394 -15276 2411
rect -14733 2394 -14716 2411
rect -14253 2394 -14236 2411
rect -14373 2394 -14356 2411
rect -14573 2394 -14556 2411
rect -15173 2394 -15156 2411
rect -14413 2394 -14396 2411
rect -15213 2394 -15196 2411
rect -14493 2394 -14476 2411
rect -14333 2394 -14316 2411
rect -14333 2394 -14316 2411
rect -14853 2394 -14836 2411
rect -15333 2394 -15316 2411
rect -15013 2394 -14996 2411
rect -15253 2394 -15236 2411
rect -14933 2394 -14916 2411
rect -14813 2394 -14796 2411
rect -14733 2394 -14716 2411
rect -14493 2394 -14476 2411
rect -14653 2394 -14636 2411
rect -15253 2394 -15236 2411
rect -14453 2394 -14436 2411
rect -14933 2394 -14916 2411
rect -15333 2394 -15316 2411
rect -15293 2394 -15276 2411
rect -14533 2394 -14516 2411
rect -14813 2394 -14796 2411
rect -14893 2394 -14876 2411
rect -15013 2394 -14996 2411
rect -15053 2394 -15036 2411
rect -15053 2394 -15036 2411
rect -14773 2394 -14756 2411
rect -14613 2394 -14596 2411
rect -14973 2394 -14956 2411
rect -14573 2394 -14556 2411
rect -14853 2394 -14836 2411
rect -14653 2394 -14636 2411
rect -14693 2394 -14676 2411
rect -14293 2394 -14276 2411
rect -15093 2394 -15076 2411
rect -15133 2394 -15116 2411
rect -15093 2394 -15076 2411
rect -14253 2394 -14236 2411
rect -14413 2394 -14396 2411
rect -14973 2394 -14956 2411
rect -14293 2394 -14276 2411
rect -15133 2394 -15116 2411
rect -14773 2394 -14756 2411
rect -14533 2394 -14516 2411
rect -14613 2394 -14596 2411
rect -14453 2394 -14436 2411
rect -10805 3163 -10788 3180
rect -10605 3163 -10588 3180
rect -10605 3163 -10588 3180
rect -10605 3163 -10588 3180
rect -10605 3163 -10588 3180
rect -10485 3163 -10468 3180
rect -10525 3163 -10508 3180
rect -10565 3163 -10548 3180
rect -10325 3163 -10308 3180
rect -10365 3163 -10348 3180
rect -10405 3163 -10388 3180
rect -10445 3163 -10428 3180
rect -10485 3163 -10468 3180
rect -10525 3163 -10508 3180
rect -10565 3163 -10548 3180
rect -10325 3163 -10308 3180
rect -10365 3163 -10348 3180
rect -10405 3163 -10388 3180
rect -10445 3163 -10428 3180
rect -10565 3163 -10548 3180
rect -10325 3163 -10308 3180
rect -10365 3163 -10348 3180
rect -10405 3163 -10388 3180
rect -10445 3163 -10428 3180
rect -10485 3163 -10468 3180
rect -10525 3163 -10508 3180
rect -10565 3163 -10548 3180
rect -10365 3163 -10348 3180
rect -10325 3163 -10308 3180
rect -10445 3163 -10428 3180
rect -10645 3163 -10628 3180
rect -10485 3163 -10468 3180
rect -10525 3163 -10508 3180
rect -10685 3163 -10668 3180
rect -10725 3163 -10708 3180
rect -10405 3163 -10388 3180
rect -10765 3163 -10748 3180
rect -11045 3163 -11028 3180
rect -11045 3163 -11028 3180
rect -11325 3163 -11308 3180
rect -11365 3163 -11348 3180
rect -11325 3163 -11308 3180
rect -11245 3163 -11228 3180
rect -11125 3163 -11108 3180
rect -10925 3163 -10908 3180
rect -10885 3163 -10868 3180
rect -11005 3163 -10988 3180
rect -11125 3163 -11108 3180
rect -11365 3163 -11348 3180
rect -11245 3163 -11228 3180
rect -11125 3163 -11108 3180
rect -11285 3163 -11268 3180
rect -10965 3163 -10948 3180
rect -11085 3163 -11068 3180
rect -10885 3163 -10868 3180
rect -10885 3163 -10868 3180
rect -10925 3163 -10908 3180
rect -11165 3163 -11148 3180
rect -10965 3163 -10948 3180
rect -10925 3163 -10908 3180
rect -10925 3163 -10908 3180
rect -11205 3163 -11188 3180
rect -11245 3163 -11228 3180
rect -11205 3163 -11188 3180
rect -11085 3163 -11068 3180
rect -11325 3163 -11308 3180
rect -11285 3163 -11268 3180
rect -10965 3163 -10948 3180
rect -11205 3163 -11188 3180
rect -11285 3163 -11268 3180
rect -11205 3163 -11188 3180
rect -11325 3163 -11308 3180
rect -11085 3163 -11068 3180
rect -11005 3163 -10988 3180
rect -11365 3163 -11348 3180
rect -10965 3163 -10948 3180
rect -11165 3163 -11148 3180
rect -11045 3163 -11028 3180
rect -11125 3163 -11108 3180
rect -11285 3163 -11268 3180
rect -11365 3163 -11348 3180
rect -11045 3163 -11028 3180
rect -11165 3163 -11148 3180
rect -11245 3163 -11228 3180
rect -11005 3163 -10988 3180
rect -11005 3163 -10988 3180
rect -10885 3163 -10868 3180
rect -11085 3163 -11068 3180
rect -11165 3163 -11148 3180
rect -11925 3163 -11908 3180
rect -11925 3163 -11908 3180
rect -11925 3163 -11908 3180
rect -11925 3163 -11908 3180
rect -11765 3163 -11748 3180
rect -11525 3163 -11508 3180
rect -11605 3163 -11588 3180
rect -11685 3163 -11668 3180
rect -11685 3163 -11668 3180
rect -11445 3163 -11428 3180
rect -11445 3163 -11428 3180
rect -11805 3163 -11788 3180
rect -11725 3163 -11708 3180
rect -11445 3163 -11428 3180
rect -11805 3163 -11788 3180
rect -11405 3163 -11388 3180
rect -11845 3163 -11828 3180
rect -11765 3163 -11748 3180
rect -11645 3163 -11628 3180
rect -11845 3163 -11828 3180
rect -11485 3163 -11468 3180
rect -11485 3163 -11468 3180
rect -11525 3163 -11508 3180
rect -11645 3163 -11628 3180
rect -11405 3163 -11388 3180
rect -11805 3163 -11788 3180
rect -11845 3163 -11828 3180
rect -11725 3163 -11708 3180
rect -11885 3163 -11868 3180
rect -11485 3163 -11468 3180
rect -11885 3163 -11868 3180
rect -11605 3163 -11588 3180
rect -11565 3163 -11548 3180
rect -11445 3163 -11428 3180
rect -11765 3163 -11748 3180
rect -11525 3163 -11508 3180
rect -11885 3163 -11868 3180
rect -11485 3163 -11468 3180
rect -11565 3163 -11548 3180
rect -11645 3163 -11628 3180
rect -11685 3163 -11668 3180
rect -11565 3163 -11548 3180
rect -11605 3163 -11588 3180
rect -11805 3163 -11788 3180
rect -11885 3163 -11868 3180
rect -11725 3163 -11708 3180
rect -11645 3163 -11628 3180
rect -11725 3163 -11708 3180
rect -11565 3163 -11548 3180
rect -11605 3163 -11588 3180
rect -11405 3163 -11388 3180
rect -11525 3163 -11508 3180
rect -11765 3163 -11748 3180
rect -11685 3163 -11668 3180
rect -11845 3163 -11828 3180
rect -11405 3163 -11388 3180
rect -12125 3163 -12108 3180
rect -12125 3163 -12108 3180
rect -12125 3163 -12108 3180
rect -12325 3163 -12308 3180
rect -12285 3163 -12268 3180
rect -12285 3163 -12268 3180
rect -12045 3163 -12028 3180
rect -12245 3163 -12228 3180
rect -12245 3163 -12228 3180
rect -12045 3163 -12028 3180
rect -12445 3163 -12428 3180
rect -12365 3163 -12348 3180
rect -12365 3163 -12348 3180
rect -12125 3163 -12108 3180
rect -12245 3163 -12228 3180
rect -12245 3163 -12228 3180
rect -12325 3163 -12308 3180
rect -12405 3163 -12388 3180
rect -12325 3163 -12308 3180
rect -12405 3163 -12388 3180
rect -12085 3163 -12068 3180
rect -12205 3163 -12188 3180
rect -12445 3163 -12428 3180
rect -12085 3163 -12068 3180
rect -12405 3163 -12388 3180
rect -12405 3163 -12388 3180
rect -12165 3163 -12148 3180
rect -12045 3163 -12028 3180
rect -12445 3163 -12428 3180
rect -12085 3163 -12068 3180
rect -12365 3163 -12348 3180
rect -11965 3163 -11948 3180
rect -12005 3163 -11988 3180
rect -12005 3163 -11988 3180
rect -12285 3163 -12268 3180
rect -11965 3163 -11948 3180
rect -12005 3163 -11988 3180
rect -12285 3163 -12268 3180
rect -12165 3163 -12148 3180
rect -12165 3163 -12148 3180
rect -12205 3163 -12188 3180
rect -12445 3163 -12428 3180
rect -12365 3163 -12348 3180
rect -11965 3163 -11948 3180
rect -12005 3163 -11988 3180
rect -12045 3163 -12028 3180
rect -12165 3163 -12148 3180
rect -12085 3163 -12068 3180
rect -11965 3163 -11948 3180
rect -12205 3163 -12188 3180
rect -12205 3163 -12188 3180
rect -12325 3163 -12308 3180
rect -13006 3163 -12989 3180
rect -13006 3163 -12989 3180
rect -13006 3163 -12989 3180
rect -13006 3163 -12989 3180
rect -12766 3163 -12749 3180
rect -12806 3163 -12789 3180
rect -12486 3163 -12469 3180
rect -12726 3163 -12709 3180
rect -12966 3163 -12949 3180
rect -12686 3163 -12669 3180
rect -12606 3163 -12589 3180
rect -12926 3163 -12909 3180
rect -12486 3163 -12469 3180
rect -12646 3163 -12629 3180
rect -12526 3163 -12509 3180
rect -12566 3163 -12549 3180
rect -12686 3163 -12669 3180
rect -12606 3163 -12589 3180
rect -12526 3163 -12509 3180
rect -12966 3163 -12949 3180
rect -12766 3163 -12749 3180
rect -12926 3163 -12909 3180
rect -12726 3163 -12709 3180
rect -12646 3163 -12629 3180
rect -12766 3163 -12749 3180
rect -12966 3163 -12949 3180
rect -12966 3163 -12949 3180
rect -12686 3163 -12669 3180
rect -12726 3163 -12709 3180
rect -12886 3163 -12869 3180
rect -12766 3163 -12749 3180
rect -12806 3163 -12789 3180
rect -12846 3163 -12829 3180
rect -12846 3163 -12829 3180
rect -12846 3163 -12829 3180
rect -12566 3163 -12549 3180
rect -12886 3163 -12869 3180
rect -12886 3163 -12869 3180
rect -12846 3163 -12829 3180
rect -12486 3163 -12469 3180
rect -12806 3163 -12789 3180
rect -12726 3163 -12709 3180
rect -12526 3163 -12509 3180
rect -12886 3163 -12869 3180
rect -12566 3163 -12549 3180
rect -12806 3163 -12789 3180
rect -12606 3163 -12589 3180
rect -12926 3163 -12909 3180
rect -12486 3163 -12469 3180
rect -12646 3163 -12629 3180
rect -12926 3163 -12909 3180
rect -12526 3163 -12509 3180
rect -12566 3163 -12549 3180
rect -12686 3163 -12669 3180
rect -12606 3163 -12589 3180
rect -12646 3163 -12629 3180
rect -13286 3163 -13269 3180
rect -13086 3163 -13069 3180
rect -13486 3163 -13469 3180
rect -13046 3163 -13029 3180
rect -13206 3163 -13189 3180
rect -13046 3163 -13029 3180
rect -13166 3163 -13149 3180
rect -13046 3163 -13029 3180
rect -13166 3163 -13149 3180
rect -13526 3163 -13509 3180
rect -13126 3163 -13109 3180
rect -13126 3163 -13109 3180
rect -13246 3163 -13229 3180
rect -13326 3163 -13309 3180
rect -13166 3163 -13149 3180
rect -13406 3163 -13389 3180
rect -13086 3163 -13069 3180
rect -13326 3163 -13309 3180
rect -13086 3163 -13069 3180
rect -13446 3163 -13429 3180
rect -13486 3163 -13469 3180
rect -13326 3163 -13309 3180
rect -13486 3163 -13469 3180
rect -13206 3163 -13189 3180
rect -13126 3163 -13109 3180
rect -13206 3163 -13189 3180
rect -13526 3163 -13509 3180
rect -13406 3163 -13389 3180
rect -13286 3163 -13269 3180
rect -13446 3163 -13429 3180
rect -13246 3163 -13229 3180
rect -13326 3163 -13309 3180
rect -13526 3163 -13509 3180
rect -13486 3163 -13469 3180
rect -13446 3163 -13429 3180
rect -13086 3163 -13069 3180
rect -13526 3163 -13509 3180
rect -13246 3163 -13229 3180
rect -13246 3163 -13229 3180
rect -13406 3163 -13389 3180
rect -13206 3163 -13189 3180
rect -13286 3163 -13269 3180
rect -13166 3163 -13149 3180
rect -13286 3163 -13269 3180
rect -13366 3163 -13349 3180
rect -13126 3163 -13109 3180
rect -13366 3163 -13349 3180
rect -13366 3163 -13349 3180
rect -13406 3163 -13389 3180
rect -13446 3163 -13429 3180
rect -13046 3163 -13029 3180
rect -13366 3163 -13349 3180
rect -14086 3163 -14069 3180
rect -14086 3163 -14069 3180
rect -14086 3163 -14069 3180
rect -14086 3163 -14069 3180
rect -13726 3163 -13709 3180
rect -13566 3163 -13549 3180
rect -13766 3163 -13749 3180
rect -13966 3163 -13949 3180
rect -13926 3163 -13909 3180
rect -13646 3163 -13629 3180
rect -13566 3163 -13549 3180
rect -13686 3163 -13669 3180
rect -13966 3163 -13949 3180
rect -13646 3163 -13629 3180
rect -13646 3163 -13629 3180
rect -13646 3163 -13629 3180
rect -13566 3163 -13549 3180
rect -13846 3163 -13829 3180
rect -13966 3163 -13949 3180
rect -13686 3163 -13669 3180
rect -14046 3163 -14029 3180
rect -14006 3163 -13989 3180
rect -13806 3163 -13789 3180
rect -13766 3163 -13749 3180
rect -13846 3163 -13829 3180
rect -13846 3163 -13829 3180
rect -13926 3163 -13909 3180
rect -13926 3163 -13909 3180
rect -13886 3163 -13869 3180
rect -14006 3163 -13989 3180
rect -13606 3163 -13589 3180
rect -13886 3163 -13869 3180
rect -13806 3163 -13789 3180
rect -13886 3163 -13869 3180
rect -13566 3163 -13549 3180
rect -13966 3163 -13949 3180
rect -13686 3163 -13669 3180
rect -13686 3163 -13669 3180
rect -13726 3163 -13709 3180
rect -14046 3163 -14029 3180
rect -13766 3163 -13749 3180
rect -13726 3163 -13709 3180
rect -13606 3163 -13589 3180
rect -13726 3163 -13709 3180
rect -14006 3163 -13989 3180
rect -13926 3163 -13909 3180
rect -13886 3163 -13869 3180
rect -13806 3163 -13789 3180
rect -13806 3163 -13789 3180
rect -13846 3163 -13829 3180
rect -14046 3163 -14029 3180
rect -14046 3163 -14029 3180
rect -14006 3163 -13989 3180
rect -13766 3163 -13749 3180
rect -13606 3163 -13589 3180
rect -13606 3163 -13589 3180
rect -9765 3163 -9748 3180
rect -9765 3163 -9748 3180
rect -9765 3163 -9748 3180
rect -14126 3163 -14109 3180
rect -9765 3163 -9748 3180
rect -14126 3163 -14109 3180
rect -9685 3163 -9668 3180
rect -9605 3163 -9588 3180
rect -9725 3163 -9708 3180
rect -9565 3163 -9548 3180
rect -9485 3163 -9468 3180
rect -9605 3163 -9588 3180
rect -14166 3163 -14149 3180
rect -9645 3163 -9628 3180
rect -9485 3163 -9468 3180
rect -9525 3163 -9508 3180
rect -9565 3163 -9548 3180
rect -9445 3163 -9428 3180
rect -9565 3163 -9548 3180
rect -9525 3163 -9508 3180
rect -9485 3163 -9468 3180
rect -9565 3163 -9548 3180
rect -9445 3163 -9428 3180
rect -9485 3163 -9468 3180
rect -9645 3163 -9628 3180
rect -9605 3163 -9588 3180
rect -9445 3163 -9428 3180
rect -9725 3163 -9708 3180
rect -9725 3163 -9708 3180
rect -9445 3163 -9428 3180
rect -9685 3163 -9668 3180
rect -14166 3163 -14149 3180
rect -9725 3163 -9708 3180
rect -9645 3163 -9628 3180
rect -9645 3163 -9628 3180
rect -14166 3163 -14149 3180
rect -9525 3163 -9508 3180
rect -9525 3163 -9508 3180
rect -9605 3163 -9588 3180
rect -9685 3163 -9668 3180
rect -9685 3163 -9668 3180
rect -10285 3163 -10268 3180
rect -9845 3163 -9828 3180
rect -14126 3163 -14109 3180
rect -10285 3163 -10268 3180
rect -14166 3163 -14149 3180
rect -10005 3163 -9988 3180
rect -10005 3163 -9988 3180
rect -10005 3163 -9988 3180
rect -14126 3163 -14109 3180
rect -10005 3163 -9988 3180
rect -10045 3163 -10028 3180
rect -9965 3163 -9948 3180
rect -10125 3163 -10108 3180
rect -9965 3163 -9948 3180
rect -9805 3163 -9788 3180
rect -10285 3163 -10268 3180
rect -10125 3163 -10108 3180
rect -9885 3163 -9868 3180
rect -10045 3163 -10028 3180
rect -10205 3163 -10188 3180
rect -9925 3163 -9908 3180
rect -9925 3163 -9908 3180
rect -10245 3163 -10228 3180
rect -10085 3163 -10068 3180
rect -9925 3163 -9908 3180
rect -10245 3163 -10228 3180
rect -10165 3163 -10148 3180
rect -9965 3163 -9948 3180
rect -9885 3163 -9868 3180
rect -9805 3163 -9788 3180
rect -10125 3163 -10108 3180
rect -10085 3163 -10068 3180
rect -10045 3163 -10028 3180
rect -10085 3163 -10068 3180
rect -10245 3163 -10228 3180
rect -10285 3163 -10268 3180
rect -10165 3163 -10148 3180
rect -10205 3163 -10188 3180
rect -9805 3163 -9788 3180
rect -9925 3163 -9908 3180
rect -10205 3163 -10188 3180
rect -10205 3163 -10188 3180
rect -9885 3163 -9868 3180
rect -9845 3163 -9828 3180
rect -10245 3163 -10228 3180
rect -10125 3163 -10108 3180
rect -10045 3163 -10028 3180
rect -9885 3163 -9868 3180
rect -10085 3163 -10068 3180
rect -9805 3163 -9788 3180
rect -9845 3163 -9828 3180
rect -10165 3163 -10148 3180
rect -9965 3163 -9948 3180
rect -10165 3163 -10148 3180
rect -9845 3163 -9828 3180
rect -10845 3163 -10828 3180
rect -10845 3163 -10828 3180
rect -10845 3163 -10828 3180
rect -10845 3163 -10828 3180
rect -10805 3163 -10788 3180
rect -10765 3163 -10748 3180
rect -10765 3163 -10748 3180
rect -10645 3163 -10628 3180
rect -10805 3163 -10788 3180
rect -10685 3163 -10668 3180
rect -10725 3163 -10708 3180
rect -10645 3163 -10628 3180
rect -10725 3163 -10708 3180
rect -10685 3163 -10668 3180
rect -10805 3163 -10788 3180
rect -10645 3163 -10628 3180
rect -10685 3163 -10668 3180
rect -10725 3163 -10708 3180
rect -10765 3163 -10748 3180
rect -13133 2394 -13116 2411
rect -13053 2394 -13036 2411
rect -13013 2394 -12996 2411
rect -13733 2394 -13716 2411
rect -13573 2394 -13556 2411
rect -14093 2394 -14076 2411
rect -13173 2394 -13156 2411
rect -13973 2394 -13956 2411
rect -13213 2394 -13196 2411
rect -14013 2394 -13996 2411
rect -13253 2394 -13236 2411
rect -13293 2394 -13276 2411
rect -13413 2394 -13396 2411
rect -13773 2394 -13756 2411
rect -14133 2394 -14116 2411
rect -14053 2394 -14036 2411
rect -13613 2394 -13596 2411
rect -13333 2394 -13316 2411
rect -13453 2394 -13436 2411
rect -13813 2394 -13796 2411
rect -13373 2394 -13356 2411
rect -13893 2394 -13876 2411
rect -14093 2394 -14076 2411
rect -13493 2394 -13476 2411
rect -14133 2394 -14116 2411
rect -13533 2394 -13516 2411
rect -13653 2394 -13636 2411
rect -14013 2394 -13996 2411
rect -13853 2394 -13836 2411
rect -13573 2394 -13556 2411
rect -13933 2394 -13916 2411
rect -13173 2394 -13156 2411
rect -13933 2394 -13916 2411
rect -13213 2394 -13196 2411
rect -13613 2394 -13596 2411
rect -13253 2394 -13236 2411
rect -13653 2394 -13636 2411
rect -13293 2394 -13276 2411
rect -13693 2394 -13676 2411
rect -13333 2394 -13316 2411
rect -13693 2394 -13676 2411
rect -14053 2394 -14036 2411
rect -13893 2394 -13876 2411
rect -13373 2394 -13356 2411
rect -13733 2394 -13716 2411
rect -13853 2394 -13836 2411
rect -13413 2394 -13396 2411
rect -13773 2394 -13756 2411
rect -13973 2394 -13956 2411
rect -13453 2394 -13436 2411
rect -13813 2394 -13796 2411
rect -13493 2394 -13476 2411
rect -13533 2394 -13516 2411
rect -13053 2394 -13036 2411
rect -13093 2394 -13076 2411
rect -13013 2394 -12996 2411
rect -13133 2394 -13116 2411
rect -13093 2394 -13076 2411
rect -12733 2394 -12716 2411
rect -12453 2394 -12436 2411
rect -12493 2394 -12476 2411
rect -12253 2394 -12236 2411
rect -12893 2394 -12876 2411
rect -12213 2394 -12196 2411
rect -12253 2394 -12236 2411
rect -12773 2394 -12756 2411
rect -12293 2394 -12276 2411
rect -12613 2394 -12596 2411
rect -12933 2394 -12916 2411
rect -12373 2394 -12356 2411
rect -11813 2394 -11796 2411
rect -11813 2394 -11796 2411
rect -11853 2394 -11836 2411
rect -11973 2394 -11956 2411
rect -12013 2394 -11996 2411
rect -12053 2394 -12036 2411
rect -11853 2394 -11836 2411
rect -11933 2394 -11916 2411
rect -11973 2394 -11956 2411
rect -12013 2394 -11996 2411
rect -12053 2394 -12036 2411
rect -11933 2394 -11916 2411
rect -11893 2394 -11876 2411
rect -11893 2394 -11876 2411
rect -12693 2394 -12676 2411
rect -12333 2394 -12316 2411
rect -12613 2394 -12596 2411
rect -12693 2394 -12676 2411
rect -12653 2394 -12636 2411
rect -12573 2394 -12556 2411
rect -12093 2394 -12076 2411
rect -12653 2394 -12636 2411
rect -12493 2394 -12476 2411
rect -12773 2394 -12756 2411
rect -12413 2394 -12396 2411
rect -12533 2394 -12516 2411
rect -12813 2394 -12796 2411
rect -12933 2394 -12916 2411
rect -12533 2394 -12516 2411
rect -12333 2394 -12316 2411
rect -12973 2394 -12956 2411
rect -12853 2394 -12836 2411
rect -12813 2394 -12796 2411
rect -12853 2394 -12836 2411
rect -12973 2394 -12956 2411
rect -12133 2394 -12116 2411
rect -12173 2394 -12156 2411
rect -12573 2394 -12556 2411
rect -12413 2394 -12396 2411
rect -12093 2394 -12076 2411
rect -12453 2394 -12436 2411
rect -12893 2394 -12876 2411
rect -12293 2394 -12276 2411
rect -12173 2394 -12156 2411
rect -12373 2394 -12356 2411
rect -12133 2394 -12116 2411
rect -12213 2394 -12196 2411
rect -12733 2394 -12716 2411
rect -10612 2394 -10595 2411
rect -10612 2394 -10595 2411
rect -10692 2394 -10675 2411
rect -10652 2394 -10635 2411
rect -10652 2394 -10635 2411
rect -10692 2394 -10675 2411
rect -10732 2394 -10715 2411
rect -10772 2394 -10755 2411
rect -10812 2394 -10795 2411
rect -10852 2394 -10835 2411
rect -11613 2394 -11596 2411
rect -11653 2394 -11636 2411
rect -11693 2394 -11676 2411
rect -11253 2394 -11236 2411
rect -11733 2394 -11716 2411
rect -11773 2394 -11756 2411
rect -11053 2394 -11036 2411
rect -11573 2394 -11556 2411
rect -11413 2394 -11396 2411
rect -11093 2394 -11076 2411
rect -11613 2394 -11596 2411
rect -11533 2394 -11516 2411
rect -11333 2394 -11316 2411
rect -11013 2394 -10996 2411
rect -11293 2394 -11276 2411
rect -11133 2394 -11116 2411
rect -11453 2394 -11436 2411
rect -11013 2394 -10996 2411
rect -11573 2394 -11556 2411
rect -11653 2394 -11636 2411
rect -11173 2394 -11156 2411
rect -11053 2394 -11036 2411
rect -11093 2394 -11076 2411
rect -11213 2394 -11196 2411
rect -11133 2394 -11116 2411
rect -11693 2394 -11676 2411
rect -11173 2394 -11156 2411
rect -11493 2394 -11476 2411
rect -11213 2394 -11196 2411
rect -11253 2394 -11236 2411
rect -11493 2394 -11476 2411
rect -11733 2394 -11716 2411
rect -11453 2394 -11436 2411
rect -11293 2394 -11276 2411
rect -11333 2394 -11316 2411
rect -11373 2394 -11356 2411
rect -11373 2394 -11356 2411
rect -11773 2394 -11756 2411
rect -11413 2394 -11396 2411
rect -11533 2394 -11516 2411
rect -10892 2394 -10875 2411
rect -10932 2394 -10915 2411
rect -10972 2394 -10955 2411
rect -10732 2394 -10715 2411
rect -10772 2394 -10755 2411
rect -10812 2394 -10795 2411
rect -10852 2394 -10835 2411
rect -10892 2394 -10875 2411
rect -10932 2394 -10915 2411
rect -10972 2394 -10955 2411
rect -9932 2394 -9915 2411
rect -9972 2394 -9955 2411
rect -10252 2394 -10235 2411
rect -10412 2394 -10395 2411
rect -9532 2394 -9515 2411
rect -10012 2394 -9995 2411
rect -10092 2394 -10075 2411
rect -10292 2394 -10275 2411
rect -10052 2394 -10035 2411
rect -10572 2394 -10555 2411
rect -10012 2394 -9995 2411
rect -10532 2394 -10515 2411
rect -9492 2394 -9475 2411
rect -10332 2394 -10315 2411
rect -10572 2394 -10555 2411
rect -9572 2394 -9555 2411
rect -10092 2394 -10075 2411
rect -10532 2394 -10515 2411
rect -10132 2394 -10115 2411
rect -10492 2394 -10475 2411
rect -9612 2394 -9595 2411
rect -9652 2394 -9635 2411
rect -9692 2394 -9675 2411
rect -9732 2394 -9715 2411
rect -9452 2394 -9435 2411
rect -9732 2394 -9715 2411
rect -9492 2394 -9475 2411
rect -9772 2394 -9755 2411
rect -9812 2394 -9795 2411
rect -9852 2394 -9835 2411
rect -9892 2394 -9875 2411
rect -9532 2394 -9515 2411
rect -9572 2394 -9555 2411
rect -9612 2394 -9595 2411
rect -9772 2394 -9755 2411
rect -10172 2394 -10155 2411
rect -9812 2394 -9795 2411
rect -10172 2394 -10155 2411
rect -9852 2394 -9835 2411
rect -10212 2394 -10195 2411
rect -10372 2394 -10355 2411
rect -10252 2394 -10235 2411
rect -9892 2394 -9875 2411
rect -9932 2394 -9915 2411
rect -9652 2394 -9635 2411
rect -10292 2394 -10275 2411
rect -9452 2394 -9435 2411
rect -10332 2394 -10315 2411
rect -10212 2394 -10195 2411
rect -9692 2394 -9675 2411
rect -10452 2394 -10435 2411
rect -10052 2394 -10035 2411
rect -9972 2394 -9955 2411
rect -10492 2394 -10475 2411
rect -10372 2394 -10355 2411
rect -10452 2394 -10435 2411
rect -10132 2394 -10115 2411
rect -10412 2394 -10395 2411
rect -4652 2394 -4635 2411
rect -4652 2394 -4635 2411
rect -2805 4652 -2788 4669
rect -2365 4652 -2348 4669
rect -2405 4652 -2388 4669
rect -2445 4652 -2428 4669
rect -2485 4652 -2468 4669
rect -2725 4652 -2708 4669
rect -2805 4652 -2788 4669
rect -2525 4652 -2508 4669
rect -2565 4652 -2548 4669
rect -2605 4652 -2588 4669
rect -2845 4652 -2828 4669
rect -2365 4652 -2348 4669
rect -2405 4652 -2388 4669
rect -2445 4652 -2428 4669
rect -2485 4652 -2468 4669
rect -2525 4652 -2508 4669
rect -2565 4652 -2548 4669
rect -2605 4652 -2588 4669
rect -2325 4652 -2308 4669
rect -2285 4652 -2268 4669
rect -2285 4652 -2268 4669
rect -2325 4652 -2308 4669
rect -2285 4652 -2268 4669
rect -2365 4652 -2348 4669
rect -2325 4652 -2308 4669
rect -2405 4652 -2388 4669
rect -2685 4652 -2668 4669
rect -2445 4652 -2428 4669
rect -2725 4652 -2708 4669
rect -2485 4652 -2468 4669
rect -2365 4652 -2348 4669
rect -2525 4652 -2508 4669
rect -2645 4652 -2628 4669
rect -2565 4652 -2548 4669
rect -2405 4652 -2388 4669
rect -2605 4652 -2588 4669
rect -2845 4652 -2828 4669
rect -2645 4652 -2628 4669
rect -2445 4652 -2428 4669
rect -2685 4652 -2668 4669
rect -2725 4652 -2708 4669
rect -2765 4652 -2748 4669
rect -2805 4652 -2788 4669
rect -2845 4652 -2828 4669
rect -2605 4652 -2588 4669
rect -2485 4652 -2468 4669
rect -2565 4652 -2548 4669
rect -2765 4652 -2748 4669
rect -2645 4652 -2628 4669
rect -2685 4652 -2668 4669
rect -2725 4652 -2708 4669
rect -2765 4652 -2748 4669
rect -2805 4652 -2788 4669
rect -2845 4652 -2828 4669
rect -2765 4652 -2748 4669
rect -2645 4652 -2628 4669
rect -2285 4652 -2268 4669
rect -2325 4652 -2308 4669
rect -2525 4652 -2508 4669
rect -2685 4652 -2668 4669
rect -2885 4652 -2868 4669
rect -2925 4652 -2908 4669
rect -3405 4652 -3388 4669
rect -3005 4652 -2988 4669
rect -2885 4652 -2868 4669
rect -2925 4652 -2908 4669
rect -3365 4652 -3348 4669
rect -2965 4652 -2948 4669
rect -3005 4652 -2988 4669
rect -3045 4652 -3028 4669
rect -3085 4652 -3068 4669
rect -3125 4652 -3108 4669
rect -3165 4652 -3148 4669
rect -3205 4652 -3188 4669
rect -3245 4652 -3228 4669
rect -3285 4652 -3268 4669
rect -3325 4652 -3308 4669
rect -3365 4652 -3348 4669
rect -3405 4652 -3388 4669
rect -3445 4652 -3428 4669
rect -2965 4652 -2948 4669
rect -3045 4652 -3028 4669
rect -3085 4652 -3068 4669
rect -3125 4652 -3108 4669
rect -3445 4652 -3428 4669
rect -3165 4652 -3148 4669
rect -3205 4652 -3188 4669
rect -3245 4652 -3228 4669
rect -3285 4652 -3268 4669
rect -2965 4652 -2948 4669
rect -3005 4652 -2988 4669
rect -3045 4652 -3028 4669
rect -3085 4652 -3068 4669
rect -3125 4652 -3108 4669
rect -3165 4652 -3148 4669
rect -3205 4652 -3188 4669
rect -3245 4652 -3228 4669
rect -3285 4652 -3268 4669
rect -3325 4652 -3308 4669
rect -3365 4652 -3348 4669
rect -3405 4652 -3388 4669
rect -3445 4652 -3428 4669
rect -3045 4652 -3028 4669
rect -3085 4652 -3068 4669
rect -3125 4652 -3108 4669
rect -3165 4652 -3148 4669
rect -3205 4652 -3188 4669
rect -3245 4652 -3228 4669
rect -3285 4652 -3268 4669
rect -3325 4652 -3308 4669
rect -3365 4652 -3348 4669
rect -3405 4652 -3388 4669
rect -3445 4652 -3428 4669
rect -2885 4652 -2868 4669
rect -2925 4652 -2908 4669
rect -2965 4652 -2948 4669
rect -3005 4652 -2988 4669
rect -2885 4652 -2868 4669
rect -2925 4652 -2908 4669
rect -3325 4652 -3308 4669
rect -3885 4652 -3868 4669
rect -3925 4652 -3908 4669
rect -3485 4652 -3468 4669
rect -3925 4652 -3908 4669
rect -3925 4652 -3908 4669
rect -4045 4652 -4028 4669
rect -3565 4652 -3548 4669
rect -3485 4652 -3468 4669
rect -3485 4652 -3468 4669
rect -3525 4652 -3508 4669
rect -3845 4652 -3828 4669
rect -3525 4652 -3508 4669
rect -3565 4652 -3548 4669
rect -4045 4652 -4028 4669
rect -3605 4652 -3588 4669
rect -3645 4652 -3628 4669
rect -3885 4652 -3868 4669
rect -3605 4652 -3588 4669
rect -3685 4652 -3668 4669
rect -3725 4652 -3708 4669
rect -3765 4652 -3748 4669
rect -3885 4652 -3868 4669
rect -3805 4652 -3788 4669
rect -3965 4652 -3948 4669
rect -3925 4652 -3908 4669
rect -3845 4652 -3828 4669
rect -3965 4652 -3948 4669
rect -4005 4652 -3988 4669
rect -4005 4652 -3988 4669
rect -3725 4652 -3708 4669
rect -4045 4652 -4028 4669
rect -4005 4652 -3988 4669
rect -3565 4652 -3548 4669
rect -3645 4652 -3628 4669
rect -4045 4652 -4028 4669
rect -3605 4652 -3588 4669
rect -3685 4652 -3668 4669
rect -3565 4652 -3548 4669
rect -3645 4652 -3628 4669
rect -3765 4652 -3748 4669
rect -3965 4652 -3948 4669
rect -3725 4652 -3708 4669
rect -3805 4652 -3788 4669
rect -3845 4652 -3828 4669
rect -4005 4652 -3988 4669
rect -3525 4652 -3508 4669
rect -3765 4652 -3748 4669
rect -3485 4652 -3468 4669
rect -3805 4652 -3788 4669
rect -3845 4652 -3828 4669
rect -3525 4652 -3508 4669
rect -3685 4652 -3668 4669
rect -3605 4652 -3588 4669
rect -3885 4652 -3868 4669
rect -3725 4652 -3708 4669
rect -3645 4652 -3628 4669
rect -3805 4652 -3788 4669
rect -3765 4652 -3748 4669
rect -3965 4652 -3948 4669
rect -3685 4652 -3668 4669
rect -4565 4652 -4548 4669
rect -4085 4652 -4068 4669
rect -4605 4652 -4588 4669
rect -4525 4652 -4508 4669
rect -4645 4652 -4628 4669
rect -4285 4652 -4268 4669
rect -4565 4652 -4548 4669
rect -4165 4652 -4148 4669
rect -4605 4652 -4588 4669
rect -4325 4652 -4308 4669
rect -4645 4652 -4628 4669
rect -4365 4652 -4348 4669
rect -4205 4652 -4188 4669
rect -4405 4652 -4388 4669
rect -4125 4652 -4108 4669
rect -4445 4652 -4428 4669
rect -4245 4652 -4228 4669
rect -4085 4652 -4068 4669
rect -4125 4652 -4108 4669
rect -4165 4652 -4148 4669
rect -4205 4652 -4188 4669
rect -4245 4652 -4228 4669
rect -4285 4652 -4268 4669
rect -4325 4652 -4308 4669
rect -4365 4652 -4348 4669
rect -4405 4652 -4388 4669
rect -4445 4652 -4428 4669
rect -4525 4652 -4508 4669
rect -4485 4652 -4468 4669
rect -4485 4652 -4468 4669
rect -4605 4652 -4588 4669
rect -4645 4652 -4628 4669
rect -4525 4652 -4508 4669
rect -4325 4652 -4308 4669
rect -4205 4652 -4188 4669
rect -4645 4652 -4628 4669
rect -4125 4652 -4108 4669
rect -4285 4652 -4268 4669
rect -4365 4652 -4348 4669
rect -4445 4652 -4428 4669
rect -4085 4652 -4068 4669
rect -4165 4652 -4148 4669
rect -4405 4652 -4388 4669
rect -4565 4652 -4548 4669
rect -4365 4652 -4348 4669
rect -4245 4652 -4228 4669
rect -4565 4652 -4548 4669
rect -4245 4652 -4228 4669
rect -4445 4652 -4428 4669
rect -4165 4652 -4148 4669
rect -4605 4652 -4588 4669
rect -4325 4652 -4308 4669
rect -4525 4652 -4508 4669
rect -4085 4652 -4068 4669
rect -4205 4652 -4188 4669
rect -4125 4652 -4108 4669
rect -4485 4652 -4468 4669
rect -4285 4652 -4268 4669
rect -4485 4652 -4468 4669
rect -4405 4652 -4388 4669
rect -925 4652 -908 4669
rect -885 4652 -868 4669
rect -845 4652 -828 4669
rect -805 4652 -788 4669
rect -765 4652 -748 4669
rect -725 4652 -708 4669
rect -685 4652 -668 4669
rect -645 4652 -628 4669
rect -605 4652 -588 4669
rect -565 4652 -548 4669
rect -525 4652 -508 4669
rect -485 4652 -468 4669
rect -885 4652 -868 4669
rect -965 4652 -948 4669
rect -845 4652 -828 4669
rect -805 4652 -788 4669
rect -765 4652 -748 4669
rect -725 4652 -708 4669
rect -685 4652 -668 4669
rect -645 4652 -628 4669
rect -605 4652 -588 4669
rect -565 4652 -548 4669
rect -525 4652 -508 4669
rect -485 4652 -468 4669
rect -445 4652 -428 4669
rect -405 4652 -388 4669
rect -365 4652 -348 4669
rect -325 4652 -308 4669
rect -285 4652 -268 4669
rect -245 4652 -228 4669
rect -205 4652 -188 4669
rect -165 4652 -148 4669
rect -125 4652 -108 4669
rect -85 4652 -68 4669
rect -45 4652 -28 4669
rect -5 4652 13 4669
rect 36 4652 53 4669
rect 76 4652 93 4669
rect -965 4652 -948 4669
rect -925 4652 -908 4669
rect -445 4652 -428 4669
rect -405 4652 -388 4669
rect -365 4652 -348 4669
rect -325 4652 -308 4669
rect -285 4652 -268 4669
rect -245 4652 -228 4669
rect -205 4652 -188 4669
rect -165 4652 -148 4669
rect -125 4652 -108 4669
rect -85 4652 -68 4669
rect -45 4652 -28 4669
rect -5 4652 13 4669
rect 36 4652 53 4669
rect 76 4652 93 4669
rect -1965 4652 -1948 4669
rect -2005 4652 -1988 4669
rect -2045 4652 -2028 4669
rect -2085 4652 -2068 4669
rect -2125 4652 -2108 4669
rect -2165 4652 -2148 4669
rect -2205 4652 -2188 4669
rect -2245 4652 -2228 4669
rect -1685 4652 -1668 4669
rect -1725 4652 -1708 4669
rect -1765 4652 -1748 4669
rect -1805 4652 -1788 4669
rect -1845 4652 -1828 4669
rect -1885 4652 -1868 4669
rect -1925 4652 -1908 4669
rect -1965 4652 -1948 4669
rect -2005 4652 -1988 4669
rect -2045 4652 -2028 4669
rect -2085 4652 -2068 4669
rect -2125 4652 -2108 4669
rect -2165 4652 -2148 4669
rect -2205 4652 -2188 4669
rect -2205 4652 -2188 4669
rect -1765 4652 -1748 4669
rect -1805 4652 -1788 4669
rect -1845 4652 -1828 4669
rect -1885 4652 -1868 4669
rect -1925 4652 -1908 4669
rect -1965 4652 -1948 4669
rect -2005 4652 -1988 4669
rect -2045 4652 -2028 4669
rect -2085 4652 -2068 4669
rect -2125 4652 -2108 4669
rect -2205 4652 -2188 4669
rect -2165 4652 -2148 4669
rect -2245 4652 -2228 4669
rect -1685 4652 -1668 4669
rect -1725 4652 -1708 4669
rect -2245 4652 -2228 4669
rect -2245 4652 -2228 4669
rect -1685 4652 -1668 4669
rect -1725 4652 -1708 4669
rect -1765 4652 -1748 4669
rect -1805 4652 -1788 4669
rect -1845 4652 -1828 4669
rect -1885 4652 -1868 4669
rect -1925 4652 -1908 4669
rect -1685 4652 -1668 4669
rect -1725 4652 -1708 4669
rect -1765 4652 -1748 4669
rect -1805 4652 -1788 4669
rect -1845 4652 -1828 4669
rect -1885 4652 -1868 4669
rect -1925 4652 -1908 4669
rect -1965 4652 -1948 4669
rect -2005 4652 -1988 4669
rect -2045 4652 -2028 4669
rect -2085 4652 -2068 4669
rect -2125 4652 -2108 4669
rect -2165 4652 -2148 4669
rect -7326 4652 -7309 4669
rect -7206 4652 -7189 4669
rect -7606 4652 -7589 4669
rect -7406 4652 -7389 4669
rect -7126 4652 -7109 4669
rect -7446 4652 -7429 4669
rect -7446 4652 -7429 4669
rect -7486 4652 -7469 4669
rect -7166 4652 -7149 4669
rect -7446 4652 -7429 4669
rect -7486 4652 -7469 4669
rect -7046 4652 -7029 4669
rect -7326 4652 -7309 4669
rect -7406 4652 -7389 4669
rect -7526 4652 -7509 4669
rect -7526 4652 -7509 4669
rect -7486 4652 -7469 4669
rect -7246 4652 -7229 4669
rect -7566 4652 -7549 4669
rect -7406 4652 -7389 4669
rect -7526 4652 -7509 4669
rect -7526 4652 -7509 4669
rect -7606 4652 -7589 4669
rect -7246 4652 -7229 4669
rect -7566 4652 -7549 4669
rect -7606 4652 -7589 4669
rect -7126 4652 -7109 4669
rect -7286 4652 -7269 4669
rect -7606 4652 -7589 4669
rect -7566 4652 -7549 4669
rect -7246 4652 -7229 4669
rect -7166 4652 -7149 4669
rect -7366 4652 -7349 4669
rect -7446 4652 -7429 4669
rect -7046 4652 -7029 4669
rect -7406 4652 -7389 4669
rect -7566 4652 -7549 4669
rect -7326 4652 -7309 4669
rect -7286 4652 -7269 4669
rect -7366 4652 -7349 4669
rect -7206 4652 -7189 4669
rect -7086 4652 -7069 4669
rect -7326 4652 -7309 4669
rect -7086 4652 -7069 4669
rect -7126 4652 -7109 4669
rect -7286 4652 -7269 4669
rect -7486 4652 -7469 4669
rect -7366 4652 -7349 4669
rect -7366 4652 -7349 4669
rect -7046 4652 -7029 4669
rect -7206 4652 -7189 4669
rect -7166 4652 -7149 4669
rect -7246 4652 -7229 4669
rect -7086 4652 -7069 4669
rect -7046 4652 -7029 4669
rect -7286 4652 -7269 4669
rect -7086 4652 -7069 4669
rect -7126 4652 -7109 4669
rect -7166 4652 -7149 4669
rect -7206 4652 -7189 4669
rect -8166 4652 -8149 4669
rect -8206 4652 -8189 4669
rect -8126 4652 -8109 4669
rect -8126 4652 -8109 4669
rect -8046 4652 -8029 4669
rect -7646 4652 -7629 4669
rect -8086 4652 -8069 4669
rect -7686 4652 -7669 4669
rect -8086 4652 -8069 4669
rect -8166 4652 -8149 4669
rect -7726 4652 -7709 4669
rect -8006 4652 -7989 4669
rect -7766 4652 -7749 4669
rect -7806 4652 -7789 4669
rect -8206 4652 -8189 4669
rect -7646 4652 -7629 4669
rect -8006 4652 -7989 4669
rect -7966 4652 -7949 4669
rect -7686 4652 -7669 4669
rect -7726 4652 -7709 4669
rect -7766 4652 -7749 4669
rect -7846 4652 -7829 4669
rect -7806 4652 -7789 4669
rect -8046 4652 -8029 4669
rect -7846 4652 -7829 4669
rect -7886 4652 -7869 4669
rect -7886 4652 -7869 4669
rect -7926 4652 -7909 4669
rect -7926 4652 -7909 4669
rect -7966 4652 -7949 4669
rect -8046 4652 -8029 4669
rect -7926 4652 -7909 4669
rect -7766 4652 -7749 4669
rect -7966 4652 -7949 4669
rect -7806 4652 -7789 4669
rect -7646 4652 -7629 4669
rect -7686 4652 -7669 4669
rect -7646 4652 -7629 4669
rect -7966 4652 -7949 4669
rect -8086 4652 -8069 4669
rect -7766 4652 -7749 4669
rect -8206 4652 -8189 4669
rect -8046 4652 -8029 4669
rect -7686 4652 -7669 4669
rect -7886 4652 -7869 4669
rect -7926 4652 -7909 4669
rect -8166 4652 -8149 4669
rect -8086 4652 -8069 4669
rect -7846 4652 -7829 4669
rect -7726 4652 -7709 4669
rect -8166 4652 -8149 4669
rect -7846 4652 -7829 4669
rect -7726 4652 -7709 4669
rect -7886 4652 -7869 4669
rect -8206 4652 -8189 4669
rect -7806 4652 -7789 4669
rect -8126 4652 -8109 4669
rect -8006 4652 -7989 4669
rect -8006 4652 -7989 4669
rect -8126 4652 -8109 4669
rect -8646 4652 -8629 4669
rect -8406 4652 -8389 4669
rect -8366 4652 -8349 4669
rect -8286 4652 -8269 4669
rect -8406 4652 -8389 4669
rect -8486 4652 -8469 4669
rect -8526 4652 -8509 4669
rect -8446 4652 -8429 4669
rect -8606 4652 -8589 4669
rect -8486 4652 -8469 4669
rect -8526 4652 -8509 4669
rect -8246 4652 -8229 4669
rect -8526 4652 -8509 4669
rect -8446 4652 -8429 4669
rect -8566 4652 -8549 4669
rect -8686 4652 -8669 4669
rect -8766 4652 -8749 4669
rect -8606 4652 -8589 4669
rect -8766 4652 -8749 4669
rect -8646 4652 -8629 4669
rect -8726 4652 -8709 4669
rect -8806 4652 -8789 4669
rect -8686 4652 -8669 4669
rect -8446 4652 -8429 4669
rect -8726 4652 -8709 4669
rect -8286 4652 -8269 4669
rect -8606 4652 -8589 4669
rect -8766 4652 -8749 4669
rect -8646 4652 -8629 4669
rect -8806 4652 -8789 4669
rect -8406 4652 -8389 4669
rect -8726 4652 -8709 4669
rect -8806 4652 -8789 4669
rect -8326 4652 -8309 4669
rect -8406 4652 -8389 4669
rect -8526 4652 -8509 4669
rect -8366 4652 -8349 4669
rect -8326 4652 -8309 4669
rect -8246 4652 -8229 4669
rect -8446 4652 -8429 4669
rect -8246 4652 -8229 4669
rect -8566 4652 -8549 4669
rect -8566 4652 -8549 4669
rect -8486 4652 -8469 4669
rect -8646 4652 -8629 4669
rect -8286 4652 -8269 4669
rect -8606 4652 -8589 4669
rect -8566 4652 -8549 4669
rect -8686 4652 -8669 4669
rect -8806 4652 -8789 4669
rect -8326 4652 -8309 4669
rect -8766 4652 -8749 4669
rect -8486 4652 -8469 4669
rect -8726 4652 -8709 4669
rect -8246 4652 -8229 4669
rect -8366 4652 -8349 4669
rect -8366 4652 -8349 4669
rect -8286 4652 -8269 4669
rect -8686 4652 -8669 4669
rect -8326 4652 -8309 4669
rect -8926 4652 -8909 4669
rect -9166 4652 -9149 4669
rect -8846 4652 -8829 4669
rect -9366 4652 -9349 4669
rect -8846 4652 -8829 4669
rect -9246 4652 -9229 4669
rect -8886 4652 -8869 4669
rect -8886 4652 -8869 4669
rect -8926 4652 -8909 4669
rect -9086 4652 -9069 4669
rect -8966 4652 -8949 4669
rect -9326 4652 -9309 4669
rect -9006 4652 -8989 4669
rect -8846 4652 -8829 4669
rect -8886 4652 -8869 4669
rect -8966 4652 -8949 4669
rect -9406 4652 -9389 4669
rect -9326 4652 -9309 4669
rect -9166 4652 -9149 4669
rect -8926 4652 -8909 4669
rect -9046 4652 -9029 4669
rect -8966 4652 -8949 4669
rect -9086 4652 -9069 4669
rect -9006 4652 -8989 4669
rect -9206 4652 -9189 4669
rect -8966 4652 -8949 4669
rect -9126 4652 -9109 4669
rect -9406 4652 -9389 4669
rect -9366 4652 -9349 4669
rect -9046 4652 -9029 4669
rect -8886 4652 -8869 4669
rect -8846 4652 -8829 4669
rect -9006 4652 -8989 4669
rect -9286 4652 -9269 4669
rect -9246 4652 -9229 4669
rect -9246 4652 -9229 4669
rect -9126 4652 -9109 4669
rect -9366 4652 -9349 4669
rect -9166 4652 -9149 4669
rect -9366 4652 -9349 4669
rect -9406 4652 -9389 4669
rect -9206 4652 -9189 4669
rect -9286 4652 -9269 4669
rect -9286 4652 -9269 4669
rect -9406 4652 -9389 4669
rect -9086 4652 -9069 4669
rect -9126 4652 -9109 4669
rect -9326 4652 -9309 4669
rect -9166 4652 -9149 4669
rect -9206 4652 -9189 4669
rect -9086 4652 -9069 4669
rect -9326 4652 -9309 4669
rect -9046 4652 -9029 4669
rect -9046 4652 -9029 4669
rect -9006 4652 -8989 4669
rect -9126 4652 -9109 4669
rect -9206 4652 -9189 4669
rect -8926 4652 -8909 4669
rect -9246 4652 -9229 4669
rect -9286 4652 -9269 4669
rect -5845 4652 -5828 4669
rect -5845 4652 -5828 4669
rect -5845 4652 -5828 4669
rect -5845 4652 -5828 4669
rect -5245 4652 -5228 4669
rect -5245 4652 -5228 4669
rect -5245 4652 -5228 4669
rect -5245 4652 -5228 4669
rect -4725 4652 -4708 4669
rect -4845 4652 -4828 4669
rect -4765 4652 -4748 4669
rect -4885 4652 -4868 4669
rect -5125 4652 -5108 4669
rect -4805 4652 -4788 4669
rect -4885 4652 -4868 4669
rect -4805 4652 -4788 4669
rect -4765 4652 -4748 4669
rect -4845 4652 -4828 4669
rect -4845 4652 -4828 4669
rect -5085 4652 -5068 4669
rect -4685 4652 -4668 4669
rect -4885 4652 -4868 4669
rect -4685 4652 -4668 4669
rect -4925 4652 -4908 4669
rect -4965 4652 -4948 4669
rect -5005 4652 -4988 4669
rect -5045 4652 -5028 4669
rect -4885 4652 -4868 4669
rect -5085 4652 -5068 4669
rect -5125 4652 -5108 4669
rect -4725 4652 -4708 4669
rect -5165 4652 -5148 4669
rect -5205 4652 -5188 4669
rect -5085 4652 -5068 4669
rect -4925 4652 -4908 4669
rect -4725 4652 -4708 4669
rect -4965 4652 -4948 4669
rect -4725 4652 -4708 4669
rect -4965 4652 -4948 4669
rect -5045 4652 -5028 4669
rect -4925 4652 -4908 4669
rect -4805 4652 -4788 4669
rect -5125 4652 -5108 4669
rect -5165 4652 -5148 4669
rect -4765 4652 -4748 4669
rect -5005 4652 -4988 4669
rect -4765 4652 -4748 4669
rect -5005 4652 -4988 4669
rect -4685 4652 -4668 4669
rect -5205 4652 -5188 4669
rect -5165 4652 -5148 4669
rect -4925 4652 -4908 4669
rect -4965 4652 -4948 4669
rect -4805 4652 -4788 4669
rect -5005 4652 -4988 4669
rect -5045 4652 -5028 4669
rect -5085 4652 -5068 4669
rect -5125 4652 -5108 4669
rect -5045 4652 -5028 4669
rect -5165 4652 -5148 4669
rect -5205 4652 -5188 4669
rect -5205 4652 -5188 4669
rect -4845 4652 -4828 4669
rect -4685 4652 -4668 4669
rect -5725 4652 -5708 4669
rect -5765 4652 -5748 4669
rect -5805 4652 -5788 4669
rect -5725 4652 -5708 4669
rect -5645 4652 -5628 4669
rect -5285 4652 -5268 4669
rect -5725 4652 -5708 4669
rect -5685 4652 -5668 4669
rect -5285 4652 -5268 4669
rect -5325 4652 -5308 4669
rect -5365 4652 -5348 4669
rect -5405 4652 -5388 4669
rect -5445 4652 -5428 4669
rect -5485 4652 -5468 4669
rect -5525 4652 -5508 4669
rect -5565 4652 -5548 4669
rect -5605 4652 -5588 4669
rect -5645 4652 -5628 4669
rect -5685 4652 -5668 4669
rect -5285 4652 -5268 4669
rect -5765 4652 -5748 4669
rect -5325 4652 -5308 4669
rect -5365 4652 -5348 4669
rect -5805 4652 -5788 4669
rect -5405 4652 -5388 4669
rect -5445 4652 -5428 4669
rect -5485 4652 -5468 4669
rect -5405 4652 -5388 4669
rect -5525 4652 -5508 4669
rect -5285 4652 -5268 4669
rect -5565 4652 -5548 4669
rect -5325 4652 -5308 4669
rect -5365 4652 -5348 4669
rect -5605 4652 -5588 4669
rect -5325 4652 -5308 4669
rect -5405 4652 -5388 4669
rect -5645 4652 -5628 4669
rect -5365 4652 -5348 4669
rect -5445 4652 -5428 4669
rect -5645 4652 -5628 4669
rect -5685 4652 -5668 4669
rect -5725 4652 -5708 4669
rect -5765 4652 -5748 4669
rect -5805 4652 -5788 4669
rect -5805 4652 -5788 4669
rect -5485 4652 -5468 4669
rect -5445 4652 -5428 4669
rect -5485 4652 -5468 4669
rect -5525 4652 -5508 4669
rect -5525 4652 -5508 4669
rect -5565 4652 -5548 4669
rect -5565 4652 -5548 4669
rect -5605 4652 -5588 4669
rect -5685 4652 -5668 4669
rect -5605 4652 -5588 4669
rect -5765 4652 -5748 4669
rect -6446 4652 -6429 4669
rect -6446 4652 -6429 4669
rect -6446 4652 -6429 4669
rect -6446 4652 -6429 4669
rect -6406 4652 -6389 4669
rect -6086 4652 -6069 4669
rect -6086 4652 -6069 4669
rect -6246 4652 -6229 4669
rect -5885 4652 -5868 4669
rect -5885 4652 -5868 4669
rect -5925 4652 -5908 4669
rect -5965 4652 -5948 4669
rect -5925 4652 -5908 4669
rect -6006 4652 -5989 4669
rect -6086 4652 -6069 4669
rect -6126 4652 -6109 4669
rect -6166 4652 -6149 4669
rect -6286 4652 -6269 4669
rect -5885 4652 -5868 4669
rect -6206 4652 -6189 4669
rect -6326 4652 -6309 4669
rect -6006 4652 -5989 4669
rect -6046 4652 -6029 4669
rect -6086 4652 -6069 4669
rect -6006 4652 -5989 4669
rect -6126 4652 -6109 4669
rect -6166 4652 -6149 4669
rect -6206 4652 -6189 4669
rect -6246 4652 -6229 4669
rect -6286 4652 -6269 4669
rect -6326 4652 -6309 4669
rect -6366 4652 -6349 4669
rect -6406 4652 -6389 4669
rect -6166 4652 -6149 4669
rect -6206 4652 -6189 4669
rect -6246 4652 -6229 4669
rect -6206 4652 -6189 4669
rect -6326 4652 -6309 4669
rect -5925 4652 -5908 4669
rect -6006 4652 -5989 4669
rect -6126 4652 -6109 4669
rect -6126 4652 -6109 4669
rect -6366 4652 -6349 4669
rect -6406 4652 -6389 4669
rect -6286 4652 -6269 4669
rect -5965 4652 -5948 4669
rect -6166 4652 -6149 4669
rect -6246 4652 -6229 4669
rect -6326 4652 -6309 4669
rect -5965 4652 -5948 4669
rect -6286 4652 -6269 4669
rect -6046 4652 -6029 4669
rect -6046 4652 -6029 4669
rect -6366 4652 -6349 4669
rect -6366 4652 -6349 4669
rect -5885 4652 -5868 4669
rect -6046 4652 -6029 4669
rect -6406 4652 -6389 4669
rect -5965 4652 -5948 4669
rect -5925 4652 -5908 4669
rect -6646 4652 -6629 4669
rect -7006 4652 -6989 4669
rect -6526 4652 -6509 4669
rect -7006 4652 -6989 4669
rect -6886 4652 -6869 4669
rect -6886 4652 -6869 4669
rect -6486 4652 -6469 4669
rect -6806 4652 -6789 4669
rect -6526 4652 -6509 4669
rect -6766 4652 -6749 4669
rect -6566 4652 -6549 4669
rect -6566 4652 -6549 4669
rect -6486 4652 -6469 4669
rect -6966 4652 -6949 4669
rect -6606 4652 -6589 4669
rect -6926 4652 -6909 4669
rect -6646 4652 -6629 4669
rect -6606 4652 -6589 4669
rect -6926 4652 -6909 4669
rect -6486 4652 -6469 4669
rect -6926 4652 -6909 4669
rect -6966 4652 -6949 4669
rect -6766 4652 -6749 4669
rect -6806 4652 -6789 4669
rect -6846 4652 -6829 4669
rect -6886 4652 -6869 4669
rect -6926 4652 -6909 4669
rect -6966 4652 -6949 4669
rect -7006 4652 -6989 4669
rect -6646 4652 -6629 4669
rect -6486 4652 -6469 4669
rect -6526 4652 -6509 4669
rect -6566 4652 -6549 4669
rect -6606 4652 -6589 4669
rect -6646 4652 -6629 4669
rect -6686 4652 -6669 4669
rect -6526 4652 -6509 4669
rect -6566 4652 -6549 4669
rect -6686 4652 -6669 4669
rect -6726 4652 -6709 4669
rect -6606 4652 -6589 4669
rect -6766 4652 -6749 4669
rect -6686 4652 -6669 4669
rect -6806 4652 -6789 4669
rect -6846 4652 -6829 4669
rect -6966 4652 -6949 4669
rect -6846 4652 -6829 4669
rect -6726 4652 -6709 4669
rect -6686 4652 -6669 4669
rect -6886 4652 -6869 4669
rect -6726 4652 -6709 4669
rect -7006 4652 -6989 4669
rect -6726 4652 -6709 4669
rect -6766 4652 -6749 4669
rect -6806 4652 -6789 4669
rect -6846 4652 -6829 4669
rect -8525 3163 -8508 3180
rect -8485 3163 -8468 3180
rect -8445 3163 -8428 3180
rect -8645 3163 -8628 3180
rect -8565 3163 -8548 3180
rect -8565 3163 -8548 3180
rect -8405 3163 -8388 3180
rect -8445 3163 -8428 3180
rect -8645 3163 -8628 3180
rect -8365 3163 -8348 3180
rect -8245 3163 -8228 3180
rect -8245 3163 -8228 3180
rect -8605 3163 -8588 3180
rect -8165 3163 -8148 3180
rect -8445 3163 -8428 3180
rect -8285 3163 -8268 3180
rect -8485 3163 -8468 3180
rect -8245 3163 -8228 3180
rect -8165 3163 -8148 3180
rect -8645 3163 -8628 3180
rect -8565 3163 -8548 3180
rect -8365 3163 -8348 3180
rect -9165 3163 -9148 3180
rect -9085 3163 -9068 3180
rect -9205 3163 -9188 3180
rect -9125 3163 -9108 3180
rect -9005 3163 -8988 3180
rect -8725 3163 -8708 3180
rect -9005 3163 -8988 3180
rect -8925 3163 -8908 3180
rect -8805 3163 -8788 3180
rect -8885 3163 -8868 3180
rect -8845 3163 -8828 3180
rect -9125 3163 -9108 3180
rect -9165 3163 -9148 3180
rect -8885 3163 -8868 3180
rect -8765 3163 -8748 3180
rect -8725 3163 -8708 3180
rect -9005 3163 -8988 3180
rect -8805 3163 -8788 3180
rect -8725 3163 -8708 3180
rect -8885 3163 -8868 3180
rect -8965 3163 -8948 3180
rect -9045 3163 -9028 3180
rect -8765 3163 -8748 3180
rect -8845 3163 -8828 3180
rect -8805 3163 -8788 3180
rect -8925 3163 -8908 3180
rect -8845 3163 -8828 3180
rect -8845 3163 -8828 3180
rect -8925 3163 -8908 3180
rect -8925 3163 -8908 3180
rect -9045 3163 -9028 3180
rect -9045 3163 -9028 3180
rect -8805 3163 -8788 3180
rect -8965 3163 -8948 3180
rect -8765 3163 -8748 3180
rect -9085 3163 -9068 3180
rect -9125 3163 -9108 3180
rect -9005 3163 -8988 3180
rect -9165 3163 -9148 3180
rect -9205 3163 -9188 3180
rect -9205 3163 -9188 3180
rect -9165 3163 -9148 3180
rect -9085 3163 -9068 3180
rect -8965 3163 -8948 3180
rect -9085 3163 -9068 3180
rect -8765 3163 -8748 3180
rect -9125 3163 -9108 3180
rect -8965 3163 -8948 3180
rect -9045 3163 -9028 3180
rect -8725 3163 -8708 3180
rect -8885 3163 -8868 3180
rect -9205 3163 -9188 3180
rect -9245 3163 -9228 3180
rect -9365 3163 -9348 3180
rect -9285 3163 -9268 3180
rect -9325 3163 -9308 3180
rect -9365 3163 -9348 3180
rect -9285 3163 -9268 3180
rect -9405 3163 -9388 3180
rect -9405 3163 -9388 3180
rect -9285 3163 -9268 3180
rect -9245 3163 -9228 3180
rect -9325 3163 -9308 3180
rect -9325 3163 -9308 3180
rect -9365 3163 -9348 3180
rect -9405 3163 -9388 3180
rect -9245 3163 -9228 3180
rect -9405 3163 -9388 3180
rect -9365 3163 -9348 3180
rect -9285 3163 -9268 3180
rect -9325 3163 -9308 3180
rect -9245 3163 -9228 3180
rect -4885 3163 -4868 3180
rect -4725 3163 -4708 3180
rect -4725 3163 -4708 3180
rect -4725 3163 -4708 3180
rect -4845 3163 -4828 3180
rect -4725 3163 -4708 3180
rect -4765 3163 -4748 3180
rect -4805 3163 -4788 3180
rect -4885 3163 -4868 3180
rect -4765 3163 -4748 3180
rect -4765 3163 -4748 3180
rect -4805 3163 -4788 3180
rect -4685 3163 -4668 3180
rect -4805 3163 -4788 3180
rect -4885 3163 -4868 3180
rect -4805 3163 -4788 3180
rect -4845 3163 -4828 3180
rect -4685 3163 -4668 3180
rect -4765 3163 -4748 3180
rect -4845 3163 -4828 3180
rect -4845 3163 -4828 3180
rect -4685 3163 -4668 3180
rect -4885 3163 -4868 3180
rect -4685 3163 -4668 3180
rect -5445 3163 -5428 3180
rect -5445 3163 -5428 3180
rect -5445 3163 -5428 3180
rect -5445 3163 -5428 3180
rect -5405 3163 -5388 3180
rect -5085 3163 -5068 3180
rect -5125 3163 -5108 3180
rect -5165 3163 -5148 3180
rect -5205 3163 -5188 3180
rect -5085 3163 -5068 3180
rect -5285 3163 -5268 3180
rect -4925 3163 -4908 3180
rect -4965 3163 -4948 3180
rect -4965 3163 -4948 3180
rect -5045 3163 -5028 3180
rect -5325 3163 -5308 3180
rect -4925 3163 -4908 3180
rect -5285 3163 -5268 3180
rect -5365 3163 -5348 3180
rect -5125 3163 -5108 3180
rect -5165 3163 -5148 3180
rect -5325 3163 -5308 3180
rect -5005 3163 -4988 3180
rect -5405 3163 -5388 3180
rect -5125 3163 -5108 3180
rect -5005 3163 -4988 3180
rect -5285 3163 -5268 3180
rect -5325 3163 -5308 3180
rect -5245 3163 -5228 3180
rect -5205 3163 -5188 3180
rect -5165 3163 -5148 3180
rect -4925 3163 -4908 3180
rect -4965 3163 -4948 3180
rect -5245 3163 -5228 3180
rect -5005 3163 -4988 3180
rect -5365 3163 -5348 3180
rect -5045 3163 -5028 3180
rect -5085 3163 -5068 3180
rect -5365 3163 -5348 3180
rect -5125 3163 -5108 3180
rect -4965 3163 -4948 3180
rect -5045 3163 -5028 3180
rect -5285 3163 -5268 3180
rect -5165 3163 -5148 3180
rect -5205 3163 -5188 3180
rect -5325 3163 -5308 3180
rect -5205 3163 -5188 3180
rect -5245 3163 -5228 3180
rect -5365 3163 -5348 3180
rect -5405 3163 -5388 3180
rect -5085 3163 -5068 3180
rect -5405 3163 -5388 3180
rect -5005 3163 -4988 3180
rect -5045 3163 -5028 3180
rect -5245 3163 -5228 3180
rect -4925 3163 -4908 3180
rect -5645 3163 -5628 3180
rect -5845 3163 -5828 3180
rect -5925 3163 -5908 3180
rect -5805 3163 -5788 3180
rect -5845 3163 -5828 3180
rect -5525 3163 -5508 3180
rect -5565 3163 -5548 3180
rect -5885 3163 -5868 3180
rect -5685 3163 -5668 3180
rect -5485 3163 -5468 3180
rect -5605 3163 -5588 3180
rect -5645 3163 -5628 3180
rect -5965 3163 -5948 3180
rect -5765 3163 -5748 3180
rect -5485 3163 -5468 3180
rect -5605 3163 -5588 3180
rect -5965 3163 -5948 3180
rect -5925 3163 -5908 3180
rect -5685 3163 -5668 3180
rect -5685 3163 -5668 3180
rect -5525 3163 -5508 3180
rect -5845 3163 -5828 3180
rect -5645 3163 -5628 3180
rect -5805 3163 -5788 3180
rect -5565 3163 -5548 3180
rect -5685 3163 -5668 3180
rect -5885 3163 -5868 3180
rect -5725 3163 -5708 3180
rect -5605 3163 -5588 3180
rect -5765 3163 -5748 3180
rect -5765 3163 -5748 3180
rect -5965 3163 -5948 3180
rect -5725 3163 -5708 3180
rect -5805 3163 -5788 3180
rect -5525 3163 -5508 3180
rect -5925 3163 -5908 3180
rect -5885 3163 -5868 3180
rect -5765 3163 -5748 3180
rect -5725 3163 -5708 3180
rect -5485 3163 -5468 3180
rect -5845 3163 -5828 3180
rect -5525 3163 -5508 3180
rect -5805 3163 -5788 3180
rect -5965 3163 -5948 3180
rect -5565 3163 -5548 3180
rect -5925 3163 -5908 3180
rect -5485 3163 -5468 3180
rect -5725 3163 -5708 3180
rect -5605 3163 -5588 3180
rect -5885 3163 -5868 3180
rect -5645 3163 -5628 3180
rect -5565 3163 -5548 3180
rect -6525 3163 -6508 3180
rect -6525 3163 -6508 3180
rect -6525 3163 -6508 3180
rect -6525 3163 -6508 3180
rect -6165 3163 -6148 3180
rect -6285 3163 -6268 3180
rect -6205 3163 -6188 3180
rect -6325 3163 -6308 3180
rect -6005 3163 -5988 3180
rect -6045 3163 -6028 3180
rect -6085 3163 -6068 3180
rect -6005 3163 -5988 3180
rect -6125 3163 -6108 3180
rect -6165 3163 -6148 3180
rect -6205 3163 -6188 3180
rect -6245 3163 -6228 3180
rect -6285 3163 -6268 3180
rect -6325 3163 -6308 3180
rect -6365 3163 -6348 3180
rect -6405 3163 -6388 3180
rect -6165 3163 -6148 3180
rect -6205 3163 -6188 3180
rect -6245 3163 -6228 3180
rect -6485 3163 -6468 3180
rect -6205 3163 -6188 3180
rect -6325 3163 -6308 3180
rect -6005 3163 -5988 3180
rect -6005 3163 -5988 3180
rect -6125 3163 -6108 3180
rect -6125 3163 -6108 3180
rect -6365 3163 -6348 3180
rect -6405 3163 -6388 3180
rect -6285 3163 -6268 3180
rect -6085 3163 -6068 3180
rect -6165 3163 -6148 3180
rect -6245 3163 -6228 3180
rect -6325 3163 -6308 3180
rect -6285 3163 -6268 3180
rect -6045 3163 -6028 3180
rect -6045 3163 -6028 3180
rect -6365 3163 -6348 3180
rect -6365 3163 -6348 3180
rect -6485 3163 -6468 3180
rect -6045 3163 -6028 3180
rect -6405 3163 -6388 3180
rect -6125 3163 -6108 3180
rect -6405 3163 -6388 3180
rect -6085 3163 -6068 3180
rect -6445 3163 -6428 3180
rect -6445 3163 -6428 3180
rect -6445 3163 -6428 3180
rect -6085 3163 -6068 3180
rect -6445 3163 -6428 3180
rect -6245 3163 -6228 3180
rect -6485 3163 -6468 3180
rect -6485 3163 -6468 3180
rect -6685 3163 -6668 3180
rect -7045 3163 -7028 3180
rect -6965 3163 -6948 3180
rect -6565 3163 -6548 3180
rect -6565 3163 -6548 3180
rect -6965 3163 -6948 3180
rect -6845 3163 -6828 3180
rect -6605 3163 -6588 3180
rect -7005 3163 -6988 3180
rect -6765 3163 -6748 3180
rect -7045 3163 -7028 3180
rect -6765 3163 -6748 3180
rect -6965 3163 -6948 3180
rect -6645 3163 -6628 3180
rect -6605 3163 -6588 3180
rect -6925 3163 -6908 3180
rect -6645 3163 -6628 3180
rect -6685 3163 -6668 3180
rect -6805 3163 -6788 3180
rect -6885 3163 -6868 3180
rect -6925 3163 -6908 3180
rect -6925 3163 -6908 3180
rect -6725 3163 -6708 3180
rect -7045 3163 -7028 3180
rect -7005 3163 -6988 3180
rect -6725 3163 -6708 3180
rect -6565 3163 -6548 3180
rect -6765 3163 -6748 3180
rect -6805 3163 -6788 3180
rect -6925 3163 -6908 3180
rect -6845 3163 -6828 3180
rect -7045 3163 -7028 3180
rect -6685 3163 -6668 3180
rect -6885 3163 -6868 3180
rect -6645 3163 -6628 3180
rect -6725 3163 -6708 3180
rect -6605 3163 -6588 3180
rect -6765 3163 -6748 3180
rect -6685 3163 -6668 3180
rect -6645 3163 -6628 3180
rect -6805 3163 -6788 3180
rect -6845 3163 -6828 3180
rect -6965 3163 -6948 3180
rect -6845 3163 -6828 3180
rect -6725 3163 -6708 3180
rect -7005 3163 -6988 3180
rect -6605 3163 -6588 3180
rect -6805 3163 -6788 3180
rect -7005 3163 -6988 3180
rect -6885 3163 -6868 3180
rect -6885 3163 -6868 3180
rect -6565 3163 -6548 3180
rect -7605 3163 -7588 3180
rect -7605 3163 -7588 3180
rect -7605 3163 -7588 3180
rect -7605 3163 -7588 3180
rect -7165 3163 -7148 3180
rect -7445 3163 -7428 3180
rect -7485 3163 -7468 3180
rect -7325 3163 -7308 3180
rect -7405 3163 -7388 3180
rect -7525 3163 -7508 3180
rect -7525 3163 -7508 3180
rect -7485 3163 -7468 3180
rect -7245 3163 -7228 3180
rect -7565 3163 -7548 3180
rect -7405 3163 -7388 3180
rect -7525 3163 -7508 3180
rect -7525 3163 -7508 3180
rect -7125 3163 -7108 3180
rect -7245 3163 -7228 3180
rect -7565 3163 -7548 3180
rect -7445 3163 -7428 3180
rect -7125 3163 -7108 3180
rect -7285 3163 -7268 3180
rect -7445 3163 -7428 3180
rect -7565 3163 -7548 3180
rect -7245 3163 -7228 3180
rect -7165 3163 -7148 3180
rect -7365 3163 -7348 3180
rect -7445 3163 -7428 3180
rect -7405 3163 -7388 3180
rect -7565 3163 -7548 3180
rect -7325 3163 -7308 3180
rect -7285 3163 -7268 3180
rect -7365 3163 -7348 3180
rect -7205 3163 -7188 3180
rect -7085 3163 -7068 3180
rect -7325 3163 -7308 3180
rect -7085 3163 -7068 3180
rect -7125 3163 -7108 3180
rect -7285 3163 -7268 3180
rect -7485 3163 -7468 3180
rect -7365 3163 -7348 3180
rect -7365 3163 -7348 3180
rect -7205 3163 -7188 3180
rect -7165 3163 -7148 3180
rect -7245 3163 -7228 3180
rect -7085 3163 -7068 3180
rect -7285 3163 -7268 3180
rect -7085 3163 -7068 3180
rect -7125 3163 -7108 3180
rect -7165 3163 -7148 3180
rect -7205 3163 -7188 3180
rect -7325 3163 -7308 3180
rect -7205 3163 -7188 3180
rect -7485 3163 -7468 3180
rect -7405 3163 -7388 3180
rect -7765 3163 -7748 3180
rect -7645 3163 -7628 3180
rect -7845 3163 -7828 3180
rect -7965 3163 -7948 3180
rect -8045 3163 -8028 3180
rect -8005 3163 -7988 3180
rect -7685 3163 -7668 3180
rect -7725 3163 -7708 3180
rect -8125 3163 -8108 3180
rect -7805 3163 -7788 3180
rect -7925 3163 -7908 3180
rect -7885 3163 -7868 3180
rect -7685 3163 -7668 3180
rect -7925 3163 -7908 3180
rect -8085 3163 -8068 3180
rect -8085 3163 -8068 3180
rect -7725 3163 -7708 3180
rect -8045 3163 -8028 3180
rect -7845 3163 -7828 3180
rect -7965 3163 -7948 3180
rect -7725 3163 -7708 3180
rect -7805 3163 -7788 3180
rect -7765 3163 -7748 3180
rect -7845 3163 -7828 3180
rect -8125 3163 -8108 3180
rect -7845 3163 -7828 3180
rect -7885 3163 -7868 3180
rect -8045 3163 -8028 3180
rect -8085 3163 -8068 3180
rect -7725 3163 -7708 3180
rect -7645 3163 -7628 3180
rect -7885 3163 -7868 3180
rect -7685 3163 -7668 3180
rect -7805 3163 -7788 3180
rect -8005 3163 -7988 3180
rect -7885 3163 -7868 3180
rect -7965 3163 -7948 3180
rect -7805 3163 -7788 3180
rect -7925 3163 -7908 3180
rect -8125 3163 -8108 3180
rect -8005 3163 -7988 3180
rect -7685 3163 -7668 3180
rect -7925 3163 -7908 3180
rect -8005 3163 -7988 3180
rect -8125 3163 -8108 3180
rect -7645 3163 -7628 3180
rect -8045 3163 -8028 3180
rect -7965 3163 -7948 3180
rect -7765 3163 -7748 3180
rect -8085 3163 -8068 3180
rect -7645 3163 -7628 3180
rect -7765 3163 -7748 3180
rect -8685 3163 -8668 3180
rect -8685 3163 -8668 3180
rect -8685 3163 -8668 3180
rect -8685 3163 -8668 3180
rect -8205 3163 -8188 3180
rect -8285 3163 -8268 3180
rect -8605 3163 -8588 3180
rect -8365 3163 -8348 3180
rect -8525 3163 -8508 3180
rect -8485 3163 -8468 3180
rect -8645 3163 -8628 3180
rect -8285 3163 -8268 3180
rect -8205 3163 -8188 3180
rect -8405 3163 -8388 3180
rect -8445 3163 -8428 3180
rect -8285 3163 -8268 3180
rect -8165 3163 -8148 3180
rect -8605 3163 -8588 3180
rect -8325 3163 -8308 3180
rect -8325 3163 -8308 3180
rect -8405 3163 -8388 3180
rect -8565 3163 -8548 3180
rect -8525 3163 -8508 3180
rect -8365 3163 -8348 3180
rect -8485 3163 -8468 3180
rect -8325 3163 -8308 3180
rect -8405 3163 -8388 3180
rect -8165 3163 -8148 3180
rect -8525 3163 -8508 3180
rect -8205 3163 -8188 3180
rect -8245 3163 -8228 3180
rect -8325 3163 -8308 3180
rect -8605 3163 -8588 3180
rect -8205 3163 -8188 3180
rect -8612 2394 -8595 2411
rect -9292 2394 -9275 2411
rect -8492 2394 -8475 2411
rect -9332 2394 -9315 2411
rect -9372 2394 -9355 2411
rect -8772 2394 -8755 2411
rect -8572 2394 -8555 2411
rect -8812 2394 -8795 2411
rect -9372 2394 -9355 2411
rect -9012 2394 -8995 2411
rect -9052 2394 -9035 2411
rect -9092 2394 -9075 2411
rect -9132 2394 -9115 2411
rect -9172 2394 -9155 2411
rect -9212 2394 -9195 2411
rect -9252 2394 -9235 2411
rect -8852 2394 -8835 2411
rect -8892 2394 -8875 2411
rect -8932 2394 -8915 2411
rect -8972 2394 -8955 2411
rect -9012 2394 -8995 2411
rect -9052 2394 -9035 2411
rect -9092 2394 -9075 2411
rect -9132 2394 -9115 2411
rect -9172 2394 -9155 2411
rect -9212 2394 -9195 2411
rect -9252 2394 -9235 2411
rect -8852 2394 -8835 2411
rect -8892 2394 -8875 2411
rect -8772 2394 -8755 2411
rect -8972 2394 -8955 2411
rect -8372 2394 -8355 2411
rect -8692 2394 -8675 2411
rect -8652 2394 -8635 2411
rect -8652 2394 -8635 2411
rect -8412 2394 -8395 2411
rect -8252 2394 -8235 2411
rect -8292 2394 -8275 2411
rect -9292 2394 -9275 2411
rect -8332 2394 -8315 2411
rect -8252 2394 -8235 2411
rect -9332 2394 -9315 2411
rect -8732 2394 -8715 2411
rect -8532 2394 -8515 2411
rect -8532 2394 -8515 2411
rect -8732 2394 -8715 2411
rect -8332 2394 -8315 2411
rect -8492 2394 -8475 2411
rect -8292 2394 -8275 2411
rect -8692 2394 -8675 2411
rect -8612 2394 -8595 2411
rect -8452 2394 -8435 2411
rect -8372 2394 -8355 2411
rect -8452 2394 -8435 2411
rect -8932 2394 -8915 2411
rect -8412 2394 -8395 2411
rect -8812 2394 -8795 2411
rect -8572 2394 -8555 2411
rect -7932 2394 -7915 2411
rect -7612 2394 -7595 2411
rect -7772 2394 -7755 2411
rect -7852 2394 -7835 2411
rect -7732 2394 -7715 2411
rect -7092 2394 -7075 2411
rect -7972 2394 -7955 2411
rect -8052 2394 -8035 2411
rect -8172 2394 -8155 2411
rect -8052 2394 -8035 2411
rect -7772 2394 -7755 2411
rect -7492 2394 -7475 2411
rect -7852 2394 -7835 2411
rect -7932 2394 -7915 2411
rect -8172 2394 -8155 2411
rect -7332 2394 -7315 2411
rect -7652 2394 -7635 2411
rect -7572 2394 -7555 2411
rect -8012 2394 -7995 2411
rect -7692 2394 -7675 2411
rect -7572 2394 -7555 2411
rect -7132 2394 -7115 2411
rect -7372 2394 -7355 2411
rect -7732 2394 -7715 2411
rect -7652 2394 -7635 2411
rect -7972 2394 -7955 2411
rect -8012 2394 -7995 2411
rect -7332 2394 -7315 2411
rect -7612 2394 -7595 2411
rect -8132 2394 -8115 2411
rect -7452 2394 -7435 2411
rect -7372 2394 -7355 2411
rect -7172 2394 -7155 2411
rect -7292 2394 -7275 2411
rect -7412 2394 -7395 2411
rect -7052 2394 -7035 2411
rect -7532 2394 -7515 2411
rect -7052 2394 -7035 2411
rect -7452 2394 -7435 2411
rect -7092 2394 -7075 2411
rect -7212 2394 -7195 2411
rect -7412 2394 -7395 2411
rect -7252 2394 -7235 2411
rect -7132 2394 -7115 2411
rect -7692 2394 -7675 2411
rect -7172 2394 -7155 2411
rect -7492 2394 -7475 2411
rect -7212 2394 -7195 2411
rect -7292 2394 -7275 2411
rect -7252 2394 -7235 2411
rect -7532 2394 -7515 2411
rect -8092 2394 -8075 2411
rect -8212 2394 -8195 2411
rect -8092 2394 -8075 2411
rect -7892 2394 -7875 2411
rect -7892 2394 -7875 2411
rect -8212 2394 -8195 2411
rect -7812 2394 -7795 2411
rect -7812 2394 -7795 2411
rect -8132 2394 -8115 2411
rect -5852 2394 -5835 2411
rect -5852 2394 -5835 2411
rect -6812 2394 -6795 2411
rect -6852 2394 -6835 2411
rect -6892 2394 -6875 2411
rect -6932 2394 -6915 2411
rect -6932 2394 -6915 2411
rect -6772 2394 -6755 2411
rect -6972 2394 -6955 2411
rect -7012 2394 -6995 2411
rect -6692 2394 -6675 2411
rect -6732 2394 -6715 2411
rect -6972 2394 -6955 2411
rect -6372 2394 -6355 2411
rect -6132 2394 -6115 2411
rect -6412 2394 -6395 2411
rect -6332 2394 -6315 2411
rect -5892 2394 -5875 2411
rect -5892 2394 -5875 2411
rect -6412 2394 -6395 2411
rect -6572 2394 -6555 2411
rect -6292 2394 -6275 2411
rect -6292 2394 -6275 2411
rect -6372 2394 -6355 2411
rect -5932 2394 -5915 2411
rect -6452 2394 -6435 2411
rect -6052 2394 -6035 2411
rect -6092 2394 -6075 2411
rect -6452 2394 -6435 2411
rect -6332 2394 -6315 2411
rect -6172 2394 -6155 2411
rect -6492 2394 -6475 2411
rect -6772 2394 -6755 2411
rect -6892 2394 -6875 2411
rect -6532 2394 -6515 2411
rect -6132 2394 -6115 2411
rect -6492 2394 -6475 2411
rect -6652 2394 -6635 2411
rect -6652 2394 -6635 2411
rect -6572 2394 -6555 2411
rect -6212 2394 -6195 2411
rect -6172 2394 -6155 2411
rect -5932 2394 -5915 2411
rect -5972 2394 -5955 2411
rect -6612 2394 -6595 2411
rect -6052 2394 -6035 2411
rect -6092 2394 -6075 2411
rect -6212 2394 -6195 2411
rect -6012 2394 -5995 2411
rect -6612 2394 -6595 2411
rect -6012 2394 -5995 2411
rect -6252 2394 -6235 2411
rect -6252 2394 -6235 2411
rect -5972 2394 -5955 2411
rect -6532 2394 -6515 2411
rect -6812 2394 -6795 2411
rect -6692 2394 -6675 2411
rect -6852 2394 -6835 2411
rect -6732 2394 -6715 2411
rect -7012 2394 -6995 2411
rect -5052 2394 -5035 2411
rect -5092 2394 -5075 2411
rect -5172 2394 -5155 2411
rect -5132 2394 -5115 2411
rect -5172 2394 -5155 2411
rect -5212 2394 -5195 2411
rect -5252 2394 -5235 2411
rect -5292 2394 -5275 2411
rect -5332 2394 -5315 2411
rect -5372 2394 -5355 2411
rect -5412 2394 -5395 2411
rect -5452 2394 -5435 2411
rect -5492 2394 -5475 2411
rect -5532 2394 -5515 2411
rect -5572 2394 -5555 2411
rect -5212 2394 -5195 2411
rect -5772 2394 -5755 2411
rect -5732 2394 -5715 2411
rect -4732 2394 -4715 2411
rect -5252 2394 -5235 2411
rect -5412 2394 -5395 2411
rect -5292 2394 -5275 2411
rect -5612 2394 -5595 2411
rect -5332 2394 -5315 2411
rect -5452 2394 -5435 2411
rect -5692 2394 -5675 2411
rect -4772 2394 -4755 2411
rect -5492 2394 -5475 2411
rect -5532 2394 -5515 2411
rect -5092 2394 -5075 2411
rect -5612 2394 -5595 2411
rect -5652 2394 -5635 2411
rect -5692 2394 -5675 2411
rect -5732 2394 -5715 2411
rect -5572 2394 -5555 2411
rect -5772 2394 -5755 2411
rect -5812 2394 -5795 2411
rect -4852 2394 -4835 2411
rect -4892 2394 -4875 2411
rect -5132 2394 -5115 2411
rect -4932 2394 -4915 2411
rect -4692 2394 -4675 2411
rect -5652 2394 -5635 2411
rect -4692 2394 -4675 2411
rect -4812 2394 -4795 2411
rect -5812 2394 -5795 2411
rect -5012 2394 -4995 2411
rect -4732 2394 -4715 2411
rect -5052 2394 -5035 2411
rect -4772 2394 -4755 2411
rect -4812 2394 -4795 2411
rect -4852 2394 -4835 2411
rect -4892 2394 -4875 2411
rect -4932 2394 -4915 2411
rect -4972 2394 -4955 2411
rect -4972 2394 -4955 2411
rect -5012 2394 -4995 2411
rect -5372 2394 -5355 2411
rect -2965 3163 -2948 3180
rect -3445 3163 -3428 3180
rect -3325 3163 -3308 3180
rect -3365 3163 -3348 3180
rect -3405 3163 -3388 3180
rect -3445 3163 -3428 3180
rect -3365 3163 -3348 3180
rect 36 3163 53 3180
rect -3365 3163 -3348 3180
rect -3765 3163 -3748 3180
rect -3685 3163 -3668 3180
rect -3685 3163 -3668 3180
rect -3405 3163 -3388 3180
rect -3605 3163 -3588 3180
rect -3445 3163 -3428 3180
rect -3445 3163 -3428 3180
rect -3725 3163 -3708 3180
rect -3325 3163 -3308 3180
rect -3405 3163 -3388 3180
rect -3325 3163 -3308 3180
rect -165 3163 -148 3180
rect -325 3163 -308 3180
rect -405 3163 -388 3180
rect -525 3163 -508 3180
rect -445 3163 -428 3180
rect -125 3163 -108 3180
rect -205 3163 -188 3180
rect -85 3163 -68 3180
rect -405 3163 -388 3180
rect -125 3163 -108 3180
rect -445 3163 -428 3180
rect -285 3163 -268 3180
rect -405 3163 -388 3180
rect -445 3163 -428 3180
rect -365 3163 -348 3180
rect -325 3163 -308 3180
rect -85 3163 -68 3180
rect -405 3163 -388 3180
rect -485 3163 -468 3180
rect -45 3163 -28 3180
rect -445 3163 -428 3180
rect -45 3163 -28 3180
rect -565 3163 -548 3180
rect -245 3163 -228 3180
rect -245 3163 -228 3180
rect -565 3163 -548 3180
rect -245 3163 -228 3180
rect -205 3163 -188 3180
rect -165 3163 -148 3180
rect -565 3163 -548 3180
rect -565 3163 -548 3180
rect -205 3163 -188 3180
rect -485 3163 -468 3180
rect -325 3163 -308 3180
rect -365 3163 -348 3180
rect -245 3163 -228 3180
rect -125 3163 -108 3180
rect -365 3163 -348 3180
rect -525 3163 -508 3180
rect -525 3163 -508 3180
rect -285 3163 -268 3180
rect -85 3163 -68 3180
rect -485 3163 -468 3180
rect -45 3163 -28 3180
rect -45 3163 -28 3180
rect -325 3163 -308 3180
rect -525 3163 -508 3180
rect -125 3163 -108 3180
rect -205 3163 -188 3180
rect -165 3163 -148 3180
rect -85 3163 -68 3180
rect -365 3163 -348 3180
rect -285 3163 -268 3180
rect -485 3163 -468 3180
rect -165 3163 -148 3180
rect -285 3163 -268 3180
rect -685 3163 -668 3180
rect -1005 3163 -988 3180
rect -685 3163 -668 3180
rect -685 3163 -668 3180
rect -1005 3163 -988 3180
rect -885 3163 -868 3180
rect -765 3163 -748 3180
rect -1045 3163 -1028 3180
rect -845 3163 -828 3180
rect -605 3163 -588 3180
rect -885 3163 -868 3180
rect -725 3163 -708 3180
rect -965 3163 -948 3180
rect -805 3163 -788 3180
rect -1045 3163 -1028 3180
rect -1085 3163 -1068 3180
rect -605 3163 -588 3180
rect -645 3163 -628 3180
rect -845 3163 -828 3180
rect -1085 3163 -1068 3180
rect -1085 3163 -1068 3180
rect -725 3163 -708 3180
rect -925 3163 -908 3180
rect -725 3163 -708 3180
rect -605 3163 -588 3180
rect -925 3163 -908 3180
rect -685 3163 -668 3180
rect -965 3163 -948 3180
rect -925 3163 -908 3180
rect -725 3163 -708 3180
rect -645 3163 -628 3180
rect -885 3163 -868 3180
rect -845 3163 -828 3180
rect -845 3163 -828 3180
rect -765 3163 -748 3180
rect -925 3163 -908 3180
rect -805 3163 -788 3180
rect -765 3163 -748 3180
rect -885 3163 -868 3180
rect -605 3163 -588 3180
rect -645 3163 -628 3180
rect -965 3163 -948 3180
rect -1045 3163 -1028 3180
rect -1005 3163 -988 3180
rect -965 3163 -948 3180
rect -645 3163 -628 3180
rect -805 3163 -788 3180
rect -1005 3163 -988 3180
rect -1045 3163 -1028 3180
rect -1085 3163 -1068 3180
rect -765 3163 -748 3180
rect -805 3163 -788 3180
rect -1645 3163 -1628 3180
rect -1325 3163 -1308 3180
rect -1485 3163 -1468 3180
rect -1205 3163 -1188 3180
rect -1245 3163 -1228 3180
rect -1565 3163 -1548 3180
rect -1405 3163 -1388 3180
rect -1525 3163 -1508 3180
rect -1485 3163 -1468 3180
rect -1485 3163 -1468 3180
rect -1325 3163 -1308 3180
rect -1125 3163 -1108 3180
rect -1445 3163 -1428 3180
rect -1645 3163 -1628 3180
rect -1325 3163 -1308 3180
rect -1605 3163 -1588 3180
rect -1365 3163 -1348 3180
rect -1565 3163 -1548 3180
rect -1405 3163 -1388 3180
rect -1245 3163 -1228 3180
rect -1205 3163 -1188 3180
rect -1285 3163 -1268 3180
rect -1525 3163 -1508 3180
rect -1645 3163 -1628 3180
rect -1605 3163 -1588 3180
rect -1525 3163 -1508 3180
rect -1205 3163 -1188 3180
rect -1525 3163 -1508 3180
rect -1325 3163 -1308 3180
rect -1285 3163 -1268 3180
rect -1165 3163 -1148 3180
rect -1565 3163 -1548 3180
rect -1565 3163 -1548 3180
rect -1245 3163 -1228 3180
rect -1285 3163 -1268 3180
rect -1445 3163 -1428 3180
rect -1285 3163 -1268 3180
rect -1205 3163 -1188 3180
rect -1605 3163 -1588 3180
rect -1405 3163 -1388 3180
rect -1365 3163 -1348 3180
rect -1125 3163 -1108 3180
rect -1365 3163 -1348 3180
rect -1165 3163 -1148 3180
rect -1245 3163 -1228 3180
rect -1605 3163 -1588 3180
rect -1125 3163 -1108 3180
rect -1485 3163 -1468 3180
rect -1405 3163 -1388 3180
rect -1365 3163 -1348 3180
rect -1125 3163 -1108 3180
rect -1445 3163 -1428 3180
rect -1445 3163 -1428 3180
rect -1165 3163 -1148 3180
rect -1645 3163 -1628 3180
rect -1165 3163 -1148 3180
rect -3645 3163 -3628 3180
rect -3325 3163 -3308 3180
rect -3365 3163 -3348 3180
rect -3525 3163 -3508 3180
rect -3405 3163 -3388 3180
rect -3805 3163 -3788 3180
rect -3485 3163 -3468 3180
rect -3565 3163 -3548 3180
rect -3485 3163 -3468 3180
rect -3485 3163 -3468 3180
rect -3525 3163 -3508 3180
rect -3525 3163 -3508 3180
rect -3565 3163 -3548 3180
rect -3605 3163 -3588 3180
rect -3645 3163 -3628 3180
rect -3605 3163 -3588 3180
rect -3685 3163 -3668 3180
rect -3725 3163 -3708 3180
rect -3765 3163 -3748 3180
rect -3805 3163 -3788 3180
rect -3725 3163 -3708 3180
rect -3565 3163 -3548 3180
rect -3645 3163 -3628 3180
rect -3605 3163 -3588 3180
rect -3685 3163 -3668 3180
rect -3565 3163 -3548 3180
rect -3645 3163 -3628 3180
rect -3765 3163 -3748 3180
rect -3725 3163 -3708 3180
rect -3805 3163 -3788 3180
rect -3525 3163 -3508 3180
rect -3765 3163 -3748 3180
rect -3485 3163 -3468 3180
rect -3805 3163 -3788 3180
rect -4365 3163 -4348 3180
rect -4365 3163 -4348 3180
rect -4365 3163 -4348 3180
rect -4365 3163 -4348 3180
rect -4325 3163 -4308 3180
rect -3885 3163 -3868 3180
rect -4205 3163 -4188 3180
rect -4125 3163 -4108 3180
rect -4245 3163 -4228 3180
rect -4085 3163 -4068 3180
rect -4125 3163 -4108 3180
rect -4165 3163 -4148 3180
rect -4205 3163 -4188 3180
rect -4245 3163 -4228 3180
rect -4285 3163 -4268 3180
rect -4325 3163 -4308 3180
rect -4085 3163 -4068 3180
rect -4325 3163 -4308 3180
rect -4205 3163 -4188 3180
rect -4125 3163 -4108 3180
rect -4285 3163 -4268 3180
rect -4285 3163 -4268 3180
rect -4085 3163 -4068 3180
rect -4165 3163 -4148 3180
rect -4165 3163 -4148 3180
rect -4245 3163 -4228 3180
rect -4245 3163 -4228 3180
rect -4165 3163 -4148 3180
rect -4325 3163 -4308 3180
rect -4085 3163 -4068 3180
rect -4205 3163 -4188 3180
rect -4125 3163 -4108 3180
rect -4285 3163 -4268 3180
rect -3885 3163 -3868 3180
rect -3925 3163 -3908 3180
rect -3925 3163 -3908 3180
rect -3925 3163 -3908 3180
rect -4045 3163 -4028 3180
rect -3845 3163 -3828 3180
rect -4045 3163 -4028 3180
rect -3965 3163 -3948 3180
rect -3885 3163 -3868 3180
rect -3885 3163 -3868 3180
rect -3965 3163 -3948 3180
rect -3925 3163 -3908 3180
rect -3845 3163 -3828 3180
rect -3965 3163 -3948 3180
rect -4005 3163 -3988 3180
rect -4005 3163 -3988 3180
rect -4045 3163 -4028 3180
rect -4005 3163 -3988 3180
rect -4045 3163 -4028 3180
rect -3965 3163 -3948 3180
rect -3845 3163 -3828 3180
rect -4005 3163 -3988 3180
rect -3845 3163 -3828 3180
rect -4405 3163 -4388 3180
rect -4565 3163 -4548 3180
rect -4565 3163 -4548 3180
rect -4445 3163 -4428 3180
rect -4565 3163 -4548 3180
rect -4405 3163 -4388 3180
rect -4445 3163 -4428 3180
rect -4445 3163 -4428 3180
rect -4605 3163 -4588 3180
rect -4525 3163 -4508 3180
rect -4525 3163 -4508 3180
rect -4485 3163 -4468 3180
rect -4485 3163 -4468 3180
rect -4485 3163 -4468 3180
rect -4405 3163 -4388 3180
rect -4485 3163 -4468 3180
rect -4605 3163 -4588 3180
rect -4645 3163 -4628 3180
rect -4525 3163 -4508 3180
rect -4605 3163 -4588 3180
rect -4605 3163 -4588 3180
rect -4645 3163 -4628 3180
rect -4525 3163 -4508 3180
rect -4645 3163 -4628 3180
rect -4645 3163 -4628 3180
rect -4445 3163 -4428 3180
rect -4565 3163 -4548 3180
rect -4405 3163 -4388 3180
rect -1965 3163 -1948 3180
rect -2005 3163 -1988 3180
rect -2045 3163 -2028 3180
rect -2085 3163 -2068 3180
rect -2125 3163 -2108 3180
rect -2165 3163 -2148 3180
rect -2205 3163 -2188 3180
rect -1685 3163 -1668 3180
rect -1725 3163 -1708 3180
rect -1765 3163 -1748 3180
rect -1805 3163 -1788 3180
rect -1845 3163 -1828 3180
rect -1885 3163 -1868 3180
rect -1925 3163 -1908 3180
rect -1965 3163 -1948 3180
rect -2005 3163 -1988 3180
rect -2045 3163 -2028 3180
rect -2085 3163 -2068 3180
rect -2125 3163 -2108 3180
rect -2165 3163 -2148 3180
rect -2205 3163 -2188 3180
rect -2205 3163 -2188 3180
rect -1765 3163 -1748 3180
rect -1805 3163 -1788 3180
rect -1845 3163 -1828 3180
rect -1885 3163 -1868 3180
rect -1925 3163 -1908 3180
rect -1965 3163 -1948 3180
rect -2005 3163 -1988 3180
rect -2045 3163 -2028 3180
rect -2085 3163 -2068 3180
rect -2125 3163 -2108 3180
rect -2205 3163 -2188 3180
rect -2165 3163 -2148 3180
rect -1685 3163 -1668 3180
rect -1725 3163 -1708 3180
rect -1685 3163 -1668 3180
rect -1725 3163 -1708 3180
rect -1765 3163 -1748 3180
rect -1805 3163 -1788 3180
rect -1845 3163 -1828 3180
rect -1885 3163 -1868 3180
rect -1925 3163 -1908 3180
rect -1685 3163 -1668 3180
rect -1725 3163 -1708 3180
rect -1765 3163 -1748 3180
rect -1805 3163 -1788 3180
rect -1845 3163 -1828 3180
rect -1885 3163 -1868 3180
rect -1925 3163 -1908 3180
rect -1965 3163 -1948 3180
rect -2005 3163 -1988 3180
rect -2045 3163 -2028 3180
rect -2085 3163 -2068 3180
rect -2125 3163 -2108 3180
rect -2165 3163 -2148 3180
rect -2565 3163 -2548 3180
rect -2285 3163 -2268 3180
rect -2485 3163 -2468 3180
rect -2285 3163 -2268 3180
rect -2605 3163 -2588 3180
rect -2325 3163 -2308 3180
rect -2405 3163 -2388 3180
rect -2285 3163 -2268 3180
rect -2725 3163 -2708 3180
rect -2365 3163 -2348 3180
rect -2365 3163 -2348 3180
rect -2325 3163 -2308 3180
rect -2365 3163 -2348 3180
rect -2405 3163 -2388 3180
rect -2405 3163 -2388 3180
rect -2685 3163 -2668 3180
rect -2445 3163 -2428 3180
rect -2445 3163 -2428 3180
rect -2445 3163 -2428 3180
rect -2725 3163 -2708 3180
rect -2245 3163 -2228 3180
rect -2485 3163 -2468 3180
rect -2485 3163 -2468 3180
rect -2365 3163 -2348 3180
rect -2525 3163 -2508 3180
rect -2525 3163 -2508 3180
rect -2525 3163 -2508 3180
rect -2645 3163 -2628 3180
rect -2245 3163 -2228 3180
rect -2565 3163 -2548 3180
rect -2565 3163 -2548 3180
rect -2405 3163 -2388 3180
rect -2245 3163 -2228 3180
rect -2605 3163 -2588 3180
rect -2605 3163 -2588 3180
rect -2245 3163 -2228 3180
rect -2645 3163 -2628 3180
rect -2325 3163 -2308 3180
rect -2445 3163 -2428 3180
rect -2685 3163 -2668 3180
rect -2725 3163 -2708 3180
rect -2605 3163 -2588 3180
rect -2485 3163 -2468 3180
rect -2565 3163 -2548 3180
rect -2645 3163 -2628 3180
rect -2685 3163 -2668 3180
rect -2725 3163 -2708 3180
rect -2645 3163 -2628 3180
rect -2285 3163 -2268 3180
rect -2325 3163 -2308 3180
rect -2525 3163 -2508 3180
rect -2685 3163 -2668 3180
rect -3005 3163 -2988 3180
rect -3045 3163 -3028 3180
rect -2845 3163 -2828 3180
rect -3085 3163 -3068 3180
rect -3125 3163 -3108 3180
rect -3165 3163 -3148 3180
rect -3205 3163 -3188 3180
rect -3245 3163 -3228 3180
rect -3285 3163 -3268 3180
rect -3045 3163 -3028 3180
rect -3085 3163 -3068 3180
rect -3125 3163 -3108 3180
rect -3165 3163 -3148 3180
rect -3205 3163 -3188 3180
rect -2885 3163 -2868 3180
rect -3245 3163 -3228 3180
rect -2925 3163 -2908 3180
rect -3285 3163 -3268 3180
rect -3005 3163 -2988 3180
rect -2885 3163 -2868 3180
rect -2925 3163 -2908 3180
rect -2885 3163 -2868 3180
rect -2965 3163 -2948 3180
rect -2925 3163 -2908 3180
rect -3005 3163 -2988 3180
rect -2965 3163 -2948 3180
rect -3045 3163 -3028 3180
rect -3005 3163 -2988 3180
rect -3085 3163 -3068 3180
rect -2885 3163 -2868 3180
rect -3125 3163 -3108 3180
rect -2925 3163 -2908 3180
rect -3165 3163 -3148 3180
rect -3205 3163 -3188 3180
rect -2805 3163 -2788 3180
rect 76 3163 93 3180
rect -2845 3163 -2828 3180
rect -3245 3163 -3228 3180
rect 76 3163 93 3180
rect -3285 3163 -3268 3180
rect -2765 3163 -2748 3180
rect -2805 3163 -2788 3180
rect -5 3163 13 3180
rect -2845 3163 -2828 3180
rect 36 3163 53 3180
rect -2965 3163 -2948 3180
rect 76 3163 93 3180
rect -3045 3163 -3028 3180
rect -5 3163 13 3180
rect -3085 3163 -3068 3180
rect -2765 3163 -2748 3180
rect 36 3163 53 3180
rect -3125 3163 -3108 3180
rect -5 3163 13 3180
rect -2805 3163 -2788 3180
rect -2765 3163 -2748 3180
rect -2805 3163 -2788 3180
rect -2845 3163 -2828 3180
rect -2765 3163 -2748 3180
rect -5 3163 13 3180
rect 36 3163 53 3180
rect -3165 3163 -3148 3180
rect -3205 3163 -3188 3180
rect -3245 3163 -3228 3180
rect -3285 3163 -3268 3180
rect 76 3163 93 3180
rect -4572 2394 -4555 2411
rect -4612 2394 -4595 2411
rect -4452 2394 -4435 2411
rect -4332 2394 -4315 2411
rect -4492 2394 -4475 2411
rect -4532 2394 -4515 2411
rect -4372 2394 -4355 2411
rect -4252 2394 -4235 2411
rect -4132 2394 -4115 2411
rect -4412 2394 -4395 2411
rect -4212 2394 -4195 2411
rect -4572 2394 -4555 2411
rect -3492 2394 -3475 2411
rect -3532 2394 -3515 2411
rect -4292 2394 -4275 2411
rect -3572 2394 -3555 2411
rect -4372 2394 -4355 2411
rect -3612 2394 -3595 2411
rect -4172 2394 -4155 2411
rect -4292 2394 -4275 2411
rect -3652 2394 -3635 2411
rect -4412 2394 -4395 2411
rect -3692 2394 -3675 2411
rect -4612 2394 -4595 2411
rect -3732 2394 -3715 2411
rect -4332 2394 -4315 2411
rect -3772 2394 -3755 2411
rect -3812 2394 -3795 2411
rect -3852 2394 -3835 2411
rect -3892 2394 -3875 2411
rect -3932 2394 -3915 2411
rect -3972 2394 -3955 2411
rect -4012 2394 -3995 2411
rect -4052 2394 -4035 2411
rect -4092 2394 -4075 2411
rect -4132 2394 -4115 2411
rect -4172 2394 -4155 2411
rect -3492 2394 -3475 2411
rect -3532 2394 -3515 2411
rect -3572 2394 -3555 2411
rect -3612 2394 -3595 2411
rect -3652 2394 -3635 2411
rect -3692 2394 -3675 2411
rect -3732 2394 -3715 2411
rect -4452 2394 -4435 2411
rect -3772 2394 -3755 2411
rect -3812 2394 -3795 2411
rect -4492 2394 -4475 2411
rect -4052 2394 -4035 2411
rect -4212 2394 -4195 2411
rect -3852 2394 -3835 2411
rect -4012 2394 -3995 2411
rect -3892 2394 -3875 2411
rect -4252 2394 -4235 2411
rect -3932 2394 -3915 2411
rect -4092 2394 -4075 2411
rect -3972 2394 -3955 2411
rect -4532 2394 -4515 2411
rect -3372 2394 -3355 2411
rect -2492 2394 -2475 2411
rect -3412 2394 -3395 2411
rect -2532 2394 -2515 2411
rect -2572 2394 -2555 2411
rect -2612 2394 -2595 2411
rect -2652 2394 -2635 2411
rect -2292 2394 -2275 2411
rect -2332 2394 -2315 2411
rect -2292 2394 -2275 2411
rect -2332 2394 -2315 2411
rect -2692 2394 -2675 2411
rect -2732 2394 -2715 2411
rect -2772 2394 -2755 2411
rect -2812 2394 -2795 2411
rect -2492 2394 -2475 2411
rect -2852 2394 -2835 2411
rect -2892 2394 -2875 2411
rect -2532 2394 -2515 2411
rect -2932 2394 -2915 2411
rect -2972 2394 -2955 2411
rect -3452 2394 -3435 2411
rect -3052 2394 -3035 2411
rect -3012 2394 -2995 2411
rect -3012 2394 -2995 2411
rect -2452 2394 -2435 2411
rect -2412 2394 -2395 2411
rect -2372 2394 -2355 2411
rect -2452 2394 -2435 2411
rect -2412 2394 -2395 2411
rect -2372 2394 -2355 2411
rect -3092 2394 -3075 2411
rect -2612 2394 -2595 2411
rect -3132 2394 -3115 2411
rect -3052 2394 -3035 2411
rect -3172 2394 -3155 2411
rect -2812 2394 -2795 2411
rect -3212 2394 -3195 2411
rect -3092 2394 -3075 2411
rect -3252 2394 -3235 2411
rect -3452 2394 -3435 2411
rect -2692 2394 -2675 2411
rect -3292 2394 -3275 2411
rect -3132 2394 -3115 2411
rect -3332 2394 -3315 2411
rect -2852 2394 -2835 2411
rect -3172 2394 -3155 2411
rect -2572 2394 -2555 2411
rect -3212 2394 -3195 2411
rect -2892 2394 -2875 2411
rect -3252 2394 -3235 2411
rect -2732 2394 -2715 2411
rect -3292 2394 -3275 2411
rect -2932 2394 -2915 2411
rect -3332 2394 -3315 2411
rect -2652 2394 -2635 2411
rect -3372 2394 -3355 2411
rect -2972 2394 -2955 2411
rect -3412 2394 -3395 2411
rect -2772 2394 -2755 2411
rect -1092 2394 -1075 2411
rect -1092 2394 -1075 2411
rect -1412 2394 -1395 2411
rect -1452 2394 -1435 2411
rect -1892 2394 -1875 2411
rect -2052 2394 -2035 2411
rect -1292 2394 -1275 2411
rect -2092 2394 -2075 2411
rect -1332 2394 -1315 2411
rect -2132 2394 -2115 2411
rect -1372 2394 -1355 2411
rect -2172 2394 -2155 2411
rect -1492 2394 -1475 2411
rect -1532 2394 -1515 2411
rect -1572 2394 -1555 2411
rect -1612 2394 -1595 2411
rect -1652 2394 -1635 2411
rect -1692 2394 -1675 2411
rect -1732 2394 -1715 2411
rect -1772 2394 -1755 2411
rect -1812 2394 -1795 2411
rect -1852 2394 -1835 2411
rect -1892 2394 -1875 2411
rect -1932 2394 -1915 2411
rect -1972 2394 -1955 2411
rect -2012 2394 -1995 2411
rect -2052 2394 -2035 2411
rect -2092 2394 -2075 2411
rect -2132 2394 -2115 2411
rect -2172 2394 -2155 2411
rect -2212 2394 -2195 2411
rect -2252 2394 -2235 2411
rect -1412 2394 -1395 2411
rect -2212 2394 -2195 2411
rect -1452 2394 -1435 2411
rect -2252 2394 -2235 2411
rect -1492 2394 -1475 2411
rect -1532 2394 -1515 2411
rect -1572 2394 -1555 2411
rect -1612 2394 -1595 2411
rect -1972 2394 -1955 2411
rect -1652 2394 -1635 2411
rect -1932 2394 -1915 2411
rect -1692 2394 -1675 2411
rect -2012 2394 -1995 2411
rect -1732 2394 -1715 2411
rect -1292 2394 -1275 2411
rect -1772 2394 -1755 2411
rect -1332 2394 -1315 2411
rect -1812 2394 -1795 2411
rect -1372 2394 -1355 2411
rect -1852 2394 -1835 2411
rect -1212 2394 -1195 2411
rect -1252 2394 -1235 2411
rect -1132 2394 -1115 2411
rect -1132 2394 -1115 2411
rect -1172 2394 -1155 2411
rect -1212 2394 -1195 2411
rect -1252 2394 -1235 2411
rect -1172 2394 -1155 2411
rect -492 2394 -475 2411
rect -532 2394 -515 2411
rect -572 2394 -555 2411
rect -612 2394 -595 2411
rect -652 2394 -635 2411
rect -692 2394 -675 2411
rect -732 2394 -715 2411
rect -892 2394 -875 2411
rect -932 2394 -915 2411
rect -972 2394 -955 2411
rect -1012 2394 -995 2411
rect -1052 2394 -1035 2411
rect -932 2394 -915 2411
rect -972 2394 -955 2411
rect -1012 2394 -995 2411
rect -1052 2394 -1035 2411
rect -812 2394 -795 2411
rect -252 2394 -235 2411
rect -292 2394 -275 2411
rect -332 2394 -315 2411
rect -372 2394 -355 2411
rect -412 2394 -395 2411
rect -732 2394 -715 2411
rect -852 2394 -835 2411
rect -772 2394 -755 2411
rect -212 2394 -195 2411
rect -252 2394 -235 2411
rect -292 2394 -275 2411
rect -332 2394 -315 2411
rect -372 2394 -355 2411
rect -772 2394 -755 2411
rect -412 2394 -395 2411
rect -452 2394 -435 2411
rect -212 2394 -195 2411
rect -452 2394 -435 2411
rect -492 2394 -475 2411
rect -532 2394 -515 2411
rect -572 2394 -555 2411
rect -612 2394 -595 2411
rect -652 2394 -635 2411
rect -692 2394 -675 2411
rect -812 2394 -795 2411
rect -852 2394 -835 2411
rect -892 2394 -875 2411
<< l125d44 >>
rect -711 3435 -687 3921
rect 1342 3435 1366 3921
<< l67d44 >>
rect 18616 8582 18633 8599
rect 18616 8582 18633 8599
rect 18976 8582 18993 8599
rect 18936 8582 18953 8599
rect 18896 8582 18913 8599
rect 18856 8582 18873 8599
rect 18816 8582 18833 8599
rect 18776 8582 18793 8599
rect 18736 8582 18753 8599
rect 19136 8582 19153 8599
rect 19096 8582 19113 8599
rect 19056 8582 19073 8599
rect 19016 8582 19033 8599
rect 18976 8582 18993 8599
rect 18936 8582 18953 8599
rect 18896 8582 18913 8599
rect 18856 8582 18873 8599
rect 18816 8582 18833 8599
rect 18776 8582 18793 8599
rect 18736 8582 18753 8599
rect 19136 8582 19153 8599
rect 19096 8582 19113 8599
rect 19056 8582 19073 8599
rect 19016 8582 19033 8599
rect 18696 8582 18713 8599
rect 18656 8582 18673 8599
rect 18696 8582 18713 8599
rect 18656 8582 18673 8599
rect 18296 8582 18313 8599
rect 18336 8582 18353 8599
rect 18576 8582 18593 8599
rect 18536 8582 18553 8599
rect 18256 8582 18273 8599
rect 18496 8582 18513 8599
rect 18216 8582 18233 8599
rect 18176 8582 18193 8599
rect 18136 8582 18153 8599
rect 18096 8582 18113 8599
rect 18456 8582 18473 8599
rect 18416 8582 18433 8599
rect 18376 8582 18393 8599
rect 18576 8582 18593 8599
rect 18536 8582 18553 8599
rect 18496 8582 18513 8599
rect 18456 8582 18473 8599
rect 18416 8582 18433 8599
rect 18376 8582 18393 8599
rect 18336 8582 18353 8599
rect 18296 8582 18313 8599
rect 18256 8582 18273 8599
rect 18216 8582 18233 8599
rect 18176 8582 18193 8599
rect 18136 8582 18153 8599
rect 18096 8582 18113 8599
rect 17976 8582 17993 8599
rect 18016 8582 18033 8599
rect 18056 8582 18073 8599
rect 18016 8582 18033 8599
rect 18056 8582 18073 8599
rect 17976 8582 17993 8599
rect 16936 8582 16953 8599
rect 16896 8582 16913 8599
rect 16856 8582 16873 8599
rect 16976 8582 16993 8599
rect 16816 8582 16833 8599
rect 16936 8582 16953 8599
rect 17176 8582 17193 8599
rect 17176 8582 17193 8599
rect 17056 8582 17073 8599
rect 17136 8582 17153 8599
rect 17216 8582 17233 8599
rect 17096 8582 17113 8599
rect 17016 8582 17033 8599
rect 17056 8582 17073 8599
rect 17936 8582 17953 8599
rect 17416 8582 17433 8599
rect 16896 8582 16913 8599
rect 17376 8582 17393 8599
rect 17656 8582 17673 8599
rect 17336 8582 17353 8599
rect 17896 8582 17913 8599
rect 17296 8582 17313 8599
rect 17856 8582 17873 8599
rect 17136 8582 17153 8599
rect 17616 8582 17633 8599
rect 17856 8582 17873 8599
rect 16776 8582 16793 8599
rect 17576 8582 17593 8599
rect 17816 8582 17833 8599
rect 17816 8582 17833 8599
rect 17776 8582 17793 8599
rect 17096 8582 17113 8599
rect 17736 8582 17753 8599
rect 16856 8582 16873 8599
rect 17696 8582 17713 8599
rect 17656 8582 17673 8599
rect 17936 8582 17953 8599
rect 17616 8582 17633 8599
rect 17576 8582 17593 8599
rect 17216 8582 17233 8599
rect 17256 8582 17273 8599
rect 17256 8582 17273 8599
rect 17016 8582 17033 8599
rect 17776 8582 17793 8599
rect 17536 8582 17553 8599
rect 17496 8582 17513 8599
rect 17536 8582 17553 8599
rect 17456 8582 17473 8599
rect 17416 8582 17433 8599
rect 17496 8582 17513 8599
rect 17376 8582 17393 8599
rect 17336 8582 17353 8599
rect 17456 8582 17473 8599
rect 17296 8582 17313 8599
rect 16816 8582 16833 8599
rect 16776 8582 16793 8599
rect 17736 8582 17753 8599
rect 16976 8582 16993 8599
rect 17896 8582 17913 8599
rect 17696 8582 17713 8599
rect 15576 8582 15593 8599
rect 15576 8582 15593 8599
rect 16696 8582 16713 8599
rect 16256 8582 16273 8599
rect 16656 8582 16673 8599
rect 16616 8582 16633 8599
rect 16616 8582 16633 8599
rect 16216 8582 16233 8599
rect 16576 8582 16593 8599
rect 16456 8582 16473 8599
rect 16536 8582 16553 8599
rect 16656 8582 16673 8599
rect 16496 8582 16513 8599
rect 16176 8582 16193 8599
rect 16456 8582 16473 8599
rect 16696 8582 16713 8599
rect 16416 8582 16433 8599
rect 16136 8582 16153 8599
rect 15696 8582 15713 8599
rect 15816 8582 15833 8599
rect 15896 8582 15913 8599
rect 15776 8582 15793 8599
rect 15736 8582 15753 8599
rect 15656 8582 15673 8599
rect 15696 8582 15713 8599
rect 15816 8582 15833 8599
rect 15656 8582 15673 8599
rect 15856 8582 15873 8599
rect 15856 8582 15873 8599
rect 15736 8582 15753 8599
rect 15896 8582 15913 8599
rect 15776 8582 15793 8599
rect 16016 8582 16033 8599
rect 15976 8582 15993 8599
rect 15616 8582 15633 8599
rect 15936 8582 15953 8599
rect 16056 8582 16073 8599
rect 16016 8582 16033 8599
rect 15976 8582 15993 8599
rect 15936 8582 15953 8599
rect 16056 8582 16073 8599
rect 15616 8582 15633 8599
rect 16096 8582 16113 8599
rect 16096 8582 16113 8599
rect 16376 8582 16393 8599
rect 16336 8582 16353 8599
rect 16256 8582 16273 8599
rect 16536 8582 16553 8599
rect 16216 8582 16233 8599
rect 16336 8582 16353 8599
rect 16296 8582 16313 8599
rect 16176 8582 16193 8599
rect 16416 8582 16433 8599
rect 16576 8582 16593 8599
rect 16136 8582 16153 8599
rect 16296 8582 16313 8599
rect 16736 8582 16753 8599
rect 16496 8582 16513 8599
rect 16376 8582 16393 8599
rect 16736 8582 16753 8599
rect 15216 8582 15233 8599
rect 14416 8582 14433 8599
rect 15496 8582 15513 8599
rect 15056 8582 15073 8599
rect 14856 8582 14873 8599
rect 14816 8582 14833 8599
rect 15496 8582 15513 8599
rect 15176 8582 15193 8599
rect 15536 8582 15553 8599
rect 14776 8582 14793 8599
rect 15456 8582 15473 8599
rect 15016 8582 15033 8599
rect 15016 8582 15033 8599
rect 14736 8582 14753 8599
rect 15136 8582 15153 8599
rect 15336 8582 15353 8599
rect 15176 8582 15193 8599
rect 14696 8582 14713 8599
rect 15416 8582 15433 8599
rect 15256 8582 15273 8599
rect 15416 8582 15433 8599
rect 14656 8582 14673 8599
rect 14976 8582 14993 8599
rect 15456 8582 15473 8599
rect 15136 8582 15153 8599
rect 14616 8582 14633 8599
rect 14976 8582 14993 8599
rect 14656 8582 14673 8599
rect 15376 8582 15393 8599
rect 14576 8582 14593 8599
rect 15096 8582 15113 8599
rect 15536 8582 15553 8599
rect 14896 8582 14913 8599
rect 14536 8582 14553 8599
rect 14896 8582 14913 8599
rect 15336 8582 15353 8599
rect 14496 8582 14513 8599
rect 14616 8582 14633 8599
rect 14456 8582 14473 8599
rect 14936 8582 14953 8599
rect 14416 8582 14433 8599
rect 15056 8582 15073 8599
rect 14816 8582 14833 8599
rect 14576 8582 14593 8599
rect 14776 8582 14793 8599
rect 15376 8582 15393 8599
rect 14736 8582 14753 8599
rect 14856 8582 14873 8599
rect 14696 8582 14713 8599
rect 14536 8582 14553 8599
rect 15296 8582 15313 8599
rect 15216 8582 15233 8599
rect 15256 8582 15273 8599
rect 14496 8582 14513 8599
rect 15096 8582 15113 8599
rect 15296 8582 15313 8599
rect 14936 8582 14953 8599
rect 14456 8582 14473 8599
rect 13496 8582 13513 8599
rect 14336 8582 14353 8599
rect 13496 8582 13513 8599
rect 13976 8582 13993 8599
rect 13456 8582 13473 8599
rect 14016 8582 14033 8599
rect 13416 8582 13433 8599
rect 14256 8582 14273 8599
rect 13736 8582 13753 8599
rect 14216 8582 14233 8599
rect 13376 8582 13393 8599
rect 13936 8582 13953 8599
rect 13336 8582 13353 8599
rect 14176 8582 14193 8599
rect 13616 8582 13633 8599
rect 13896 8582 13913 8599
rect 13296 8582 13313 8599
rect 13856 8582 13873 8599
rect 13256 8582 13273 8599
rect 13816 8582 13833 8599
rect 13456 8582 13473 8599
rect 13776 8582 13793 8599
rect 13216 8582 13233 8599
rect 14136 8582 14153 8599
rect 13216 8582 13233 8599
rect 13696 8582 13713 8599
rect 14096 8582 14113 8599
rect 13736 8582 13753 8599
rect 13416 8582 13433 8599
rect 14056 8582 14073 8599
rect 13656 8582 13673 8599
rect 13576 8582 13593 8599
rect 14256 8582 14273 8599
rect 13376 8582 13393 8599
rect 14216 8582 14233 8599
rect 14176 8582 14193 8599
rect 14136 8582 14153 8599
rect 14096 8582 14113 8599
rect 14056 8582 14073 8599
rect 14016 8582 14033 8599
rect 13976 8582 13993 8599
rect 13936 8582 13953 8599
rect 13896 8582 13913 8599
rect 13856 8582 13873 8599
rect 13816 8582 13833 8599
rect 13776 8582 13793 8599
rect 13656 8582 13673 8599
rect 13336 8582 13353 8599
rect 13576 8582 13593 8599
rect 13616 8582 13633 8599
rect 13536 8582 13553 8599
rect 14296 8582 14313 8599
rect 13296 8582 13313 8599
rect 14296 8582 14313 8599
rect 13536 8582 13553 8599
rect 14376 8582 14393 8599
rect 13696 8582 13713 8599
rect 14336 8582 14353 8599
rect 13256 8582 13273 8599
rect 14376 8582 14393 8599
rect 13176 8582 13193 8599
rect 12096 8582 12113 8599
rect 12456 8582 12473 8599
rect 12496 8582 12513 8599
rect 12256 8582 12273 8599
rect 12296 8582 12313 8599
rect 13056 8582 13073 8599
rect 12536 8582 12553 8599
rect 12176 8582 12193 8599
rect 12056 8582 12073 8599
rect 12576 8582 12593 8599
rect 12096 8582 12113 8599
rect 13016 8582 13033 8599
rect 13056 8582 13073 8599
rect 13096 8582 13113 8599
rect 12536 8582 12553 8599
rect 12256 8582 12273 8599
rect 13016 8582 13033 8599
rect 13136 8582 13153 8599
rect 12496 8582 12513 8599
rect 12976 8582 12993 8599
rect 12696 8582 12713 8599
rect 12136 8582 12153 8599
rect 12856 8582 12873 8599
rect 12976 8582 12993 8599
rect 12816 8582 12833 8599
rect 12056 8582 12073 8599
rect 13136 8582 13153 8599
rect 12216 8582 12233 8599
rect 12856 8582 12873 8599
rect 12216 8582 12233 8599
rect 12736 8582 12753 8599
rect 12176 8582 12193 8599
rect 12016 8582 12033 8599
rect 12656 8582 12673 8599
rect 12816 8582 12833 8599
rect 12416 8582 12433 8599
rect 12336 8582 12353 8599
rect 13096 8582 13113 8599
rect 12896 8582 12913 8599
rect 12376 8582 12393 8599
rect 12776 8582 12793 8599
rect 12936 8582 12953 8599
rect 12776 8582 12793 8599
rect 12656 8582 12673 8599
rect 12456 8582 12473 8599
rect 12336 8582 12353 8599
rect 12136 8582 12153 8599
rect 13176 8582 13193 8599
rect 12376 8582 12393 8599
rect 12616 8582 12633 8599
rect 12696 8582 12713 8599
rect 12616 8582 12633 8599
rect 12416 8582 12433 8599
rect 12016 8582 12033 8599
rect 12736 8582 12753 8599
rect 12576 8582 12593 8599
rect 12896 8582 12913 8599
rect 12296 8582 12313 8599
rect 12936 8582 12953 8599
rect 10816 8582 10833 8599
rect 10816 8582 10833 8599
rect 11296 8582 11313 8599
rect 11136 8582 11153 8599
rect 11616 8582 11633 8599
rect 11496 8582 11513 8599
rect 11856 8582 11873 8599
rect 11456 8582 11473 8599
rect 10896 8582 10913 8599
rect 11376 8582 11393 8599
rect 11136 8582 11153 8599
rect 11776 8582 11793 8599
rect 10976 8582 10993 8599
rect 11576 8582 11593 8599
rect 11816 8582 11833 8599
rect 11976 8582 11993 8599
rect 11816 8582 11833 8599
rect 11736 8582 11753 8599
rect 11856 8582 11873 8599
rect 10896 8582 10913 8599
rect 11656 8582 11673 8599
rect 10936 8582 10953 8599
rect 10856 8582 10873 8599
rect 11176 8582 11193 8599
rect 11336 8582 11353 8599
rect 11376 8582 11393 8599
rect 10936 8582 10953 8599
rect 11296 8582 11313 8599
rect 11056 8582 11073 8599
rect 11456 8582 11473 8599
rect 11216 8582 11233 8599
rect 11016 8582 11033 8599
rect 11256 8582 11273 8599
rect 11936 8582 11953 8599
rect 10856 8582 10873 8599
rect 11896 8582 11913 8599
rect 11416 8582 11433 8599
rect 11336 8582 11353 8599
rect 11096 8582 11113 8599
rect 11576 8582 11593 8599
rect 11016 8582 11033 8599
rect 11216 8582 11233 8599
rect 11976 8582 11993 8599
rect 11616 8582 11633 8599
rect 11056 8582 11073 8599
rect 11096 8582 11113 8599
rect 11776 8582 11793 8599
rect 11656 8582 11673 8599
rect 10976 8582 10993 8599
rect 11256 8582 11273 8599
rect 11536 8582 11553 8599
rect 11696 8582 11713 8599
rect 11936 8582 11953 8599
rect 11536 8582 11553 8599
rect 11696 8582 11713 8599
rect 11176 8582 11193 8599
rect 11736 8582 11753 8599
rect 11896 8582 11913 8599
rect 11496 8582 11513 8599
rect 11416 8582 11433 8599
rect 9696 8582 9713 8599
rect 9856 8582 9873 8599
rect 10576 8582 10593 8599
rect 9696 8582 9713 8599
rect 9856 8582 9873 8599
rect 10496 8582 10513 8599
rect 10256 8582 10273 8599
rect 10656 8582 10673 8599
rect 10216 8582 10233 8599
rect 9656 8582 9673 8599
rect 9896 8582 9913 8599
rect 10616 8582 10633 8599
rect 10256 8582 10273 8599
rect 10456 8582 10473 8599
rect 10056 8582 10073 8599
rect 10416 8582 10433 8599
rect 10456 8582 10473 8599
rect 10096 8582 10113 8599
rect 10296 8582 10313 8599
rect 10416 8582 10433 8599
rect 9816 8582 9833 8599
rect 10376 8582 10393 8599
rect 9656 8582 9673 8599
rect 10536 8582 10553 8599
rect 10136 8582 10153 8599
rect 10776 8582 10793 8599
rect 10336 8582 10353 8599
rect 10376 8582 10393 8599
rect 10696 8582 10713 8599
rect 9936 8582 9953 8599
rect 9896 8582 9913 8599
rect 10336 8582 10353 8599
rect 10176 8582 10193 8599
rect 10656 8582 10673 8599
rect 9776 8582 9793 8599
rect 9976 8582 9993 8599
rect 10216 8582 10233 8599
rect 10776 8582 10793 8599
rect 10576 8582 10593 8599
rect 10296 8582 10313 8599
rect 10736 8582 10753 8599
rect 10136 8582 10153 8599
rect 10736 8582 10753 8599
rect 10616 8582 10633 8599
rect 10096 8582 10113 8599
rect 9816 8582 9833 8599
rect 10016 8582 10033 8599
rect 10536 8582 10553 8599
rect 9736 8582 9753 8599
rect 10056 8582 10073 8599
rect 9976 8582 9993 8599
rect 10496 8582 10513 8599
rect 9736 8582 9753 8599
rect 10176 8582 10193 8599
rect 9936 8582 9953 8599
rect 10016 8582 10033 8599
rect 10696 8582 10713 8599
rect 9776 8582 9793 8599
rect 9336 8582 9353 8599
rect 9496 8582 9513 8599
rect 9256 8582 9273 8599
rect 9456 8582 9473 8599
rect 8616 8582 8633 8599
rect 8536 8582 8553 8599
rect 9056 8582 9073 8599
rect 8536 8582 8553 8599
rect 9296 8582 9313 8599
rect 8496 8582 8513 8599
rect 8576 8582 8593 8599
rect 8776 8582 8793 8599
rect 8456 8582 8473 8599
rect 8616 8582 8633 8599
rect 9336 8582 9353 8599
rect 8736 8582 8753 8599
rect 9016 8582 9033 8599
rect 9136 8582 9153 8599
rect 8696 8582 8713 8599
rect 9256 8582 9273 8599
rect 8656 8582 8673 8599
rect 8896 8582 8913 8599
rect 9216 8582 9233 8599
rect 8976 8582 8993 8599
rect 9216 8582 9233 8599
rect 8856 8582 8873 8599
rect 8576 8582 8593 8599
rect 9376 8582 9393 8599
rect 8936 8582 8953 8599
rect 8896 8582 8913 8599
rect 9176 8582 9193 8599
rect 9176 8582 9193 8599
rect 8816 8582 8833 8599
rect 9136 8582 9153 8599
rect 9096 8582 9113 8599
rect 8776 8582 8793 8599
rect 8496 8582 8513 8599
rect 8856 8582 8873 8599
rect 9416 8582 9433 8599
rect 9056 8582 9073 8599
rect 8736 8582 8753 8599
rect 9016 8582 9033 8599
rect 8696 8582 8713 8599
rect 9296 8582 9313 8599
rect 8976 8582 8993 8599
rect 8816 8582 8833 8599
rect 8936 8582 8953 8599
rect 8656 8582 8673 8599
rect 9616 8582 9633 8599
rect 9576 8582 9593 8599
rect 9376 8582 9393 8599
rect 9536 8582 9553 8599
rect 9416 8582 9433 8599
rect 9496 8582 9513 8599
rect 9456 8582 9473 8599
rect 9096 8582 9113 8599
rect 9616 8582 9633 8599
rect 8456 8582 8473 8599
rect 9576 8582 9593 8599
rect 9536 8582 9553 8599
rect 7615 8582 7632 8599
rect 8335 8582 8352 8599
rect 7655 8582 7672 8599
rect 8095 8582 8112 8599
rect 7815 8582 7832 8599
rect 7695 8582 7712 8599
rect 7575 8582 7592 8599
rect 7975 8582 7992 8599
rect 7655 8582 7672 8599
rect 8055 8582 8072 8599
rect 7975 8582 7992 8599
rect 7535 8582 7552 8599
rect 8015 8582 8032 8599
rect 8135 8582 8152 8599
rect 7255 8582 7272 8599
rect 8295 8582 8312 8599
rect 7775 8582 7792 8599
rect 8416 8582 8433 8599
rect 7495 8582 7512 8599
rect 7935 8582 7952 8599
rect 7935 8582 7952 8599
rect 8055 8582 8072 8599
rect 7575 8582 7592 8599
rect 8095 8582 8112 8599
rect 7495 8582 7512 8599
rect 8255 8582 8272 8599
rect 8215 8582 8232 8599
rect 7735 8582 7752 8599
rect 8175 8582 8192 8599
rect 8416 8582 8433 8599
rect 8135 8582 8152 8599
rect 8015 8582 8032 8599
rect 8335 8582 8352 8599
rect 7375 8582 7392 8599
rect 7455 8582 7472 8599
rect 7255 8582 7272 8599
rect 7775 8582 7792 8599
rect 7735 8582 7752 8599
rect 7335 8582 7352 8599
rect 7895 8582 7912 8599
rect 7615 8582 7632 8599
rect 8295 8582 8312 8599
rect 7295 8582 7312 8599
rect 7815 8582 7832 8599
rect 8175 8582 8192 8599
rect 7455 8582 7472 8599
rect 7415 8582 7432 8599
rect 7855 8582 7872 8599
rect 7855 8582 7872 8599
rect 7375 8582 7392 8599
rect 8255 8582 8272 8599
rect 8376 8582 8393 8599
rect 7895 8582 7912 8599
rect 7335 8582 7352 8599
rect 8215 8582 8232 8599
rect 7295 8582 7312 8599
rect 8376 8582 8393 8599
rect 7535 8582 7552 8599
rect 7415 8582 7432 8599
rect 7695 8582 7712 8599
rect 6055 8582 6072 8599
rect 6055 8582 6072 8599
rect 6255 8582 6272 8599
rect 7055 8582 7072 8599
rect 7175 8582 7192 8599
rect 7095 8582 7112 8599
rect 6215 8582 6232 8599
rect 6495 8582 6512 8599
rect 6375 8582 6392 8599
rect 6175 8582 6192 8599
rect 6735 8582 6752 8599
rect 6415 8582 6432 8599
rect 6935 8582 6952 8599
rect 6775 8582 6792 8599
rect 6655 8582 6672 8599
rect 6255 8582 6272 8599
rect 6215 8582 6232 8599
rect 6935 8582 6952 8599
rect 6655 8582 6672 8599
rect 6815 8582 6832 8599
rect 6135 8582 6152 8599
rect 6455 8582 6472 8599
rect 6855 8582 6872 8599
rect 6455 8582 6472 8599
rect 7135 8582 7152 8599
rect 6135 8582 6152 8599
rect 6415 8582 6432 8599
rect 7015 8582 7032 8599
rect 6575 8582 6592 8599
rect 6095 8582 6112 8599
rect 6895 8582 6912 8599
rect 6535 8582 6552 8599
rect 7055 8582 7072 8599
rect 6095 8582 6112 8599
rect 6295 8582 6312 8599
rect 6535 8582 6552 8599
rect 6735 8582 6752 8599
rect 6575 8582 6592 8599
rect 6335 8582 6352 8599
rect 6975 8582 6992 8599
rect 6695 8582 6712 8599
rect 7175 8582 7192 8599
rect 6375 8582 6392 8599
rect 6615 8582 6632 8599
rect 7215 8582 7232 8599
rect 6295 8582 6312 8599
rect 6975 8582 6992 8599
rect 6815 8582 6832 8599
rect 6335 8582 6352 8599
rect 7135 8582 7152 8599
rect 6615 8582 6632 8599
rect 6695 8582 6712 8599
rect 6175 8582 6192 8599
rect 7095 8582 7112 8599
rect 7015 8582 7032 8599
rect 6495 8582 6512 8599
rect 6855 8582 6872 8599
rect 7215 8582 7232 8599
rect 6775 8582 6792 8599
rect 6895 8582 6912 8599
rect 5575 8582 5592 8599
rect 5695 8582 5712 8599
rect 5095 8582 5112 8599
rect 5295 8582 5312 8599
rect 5655 8582 5672 8599
rect 5415 8582 5432 8599
rect 5615 8582 5632 8599
rect 4935 8582 4952 8599
rect 5975 8582 5992 8599
rect 4895 8582 4912 8599
rect 5895 8582 5912 8599
rect 5735 8582 5752 8599
rect 5175 8582 5192 8599
rect 5935 8582 5952 8599
rect 5615 8582 5632 8599
rect 5575 8582 5592 8599
rect 5535 8582 5552 8599
rect 5855 8582 5872 8599
rect 5775 8582 5792 8599
rect 5055 8582 5072 8599
rect 5495 8582 5512 8599
rect 5455 8582 5472 8599
rect 5415 8582 5432 8599
rect 5935 8582 5952 8599
rect 4895 8582 4912 8599
rect 5775 8582 5792 8599
rect 5135 8582 5152 8599
rect 5255 8582 5272 8599
rect 5135 8582 5152 8599
rect 6015 8582 6032 8599
rect 5215 8582 5232 8599
rect 5335 8582 5352 8599
rect 5055 8582 5072 8599
rect 5455 8582 5472 8599
rect 5015 8582 5032 8599
rect 4975 8582 4992 8599
rect 4935 8582 4952 8599
rect 5535 8582 5552 8599
rect 5175 8582 5192 8599
rect 5255 8582 5272 8599
rect 5295 8582 5312 8599
rect 5495 8582 5512 8599
rect 5015 8582 5032 8599
rect 5815 8582 5832 8599
rect 6015 8582 6032 8599
rect 5815 8582 5832 8599
rect 5335 8582 5352 8599
rect 5975 8582 5992 8599
rect 5695 8582 5712 8599
rect 5375 8582 5392 8599
rect 5895 8582 5912 8599
rect 5855 8582 5872 8599
rect 5375 8582 5392 8599
rect 5095 8582 5112 8599
rect 5655 8582 5672 8599
rect 5735 8582 5752 8599
rect 5215 8582 5232 8599
rect 4975 8582 4992 8599
rect 3895 8582 3912 8599
rect 4735 8582 4752 8599
rect 4575 8582 4592 8599
rect 4695 8582 4712 8599
rect 4095 8582 4112 8599
rect 4655 8582 4672 8599
rect 4495 8582 4512 8599
rect 4815 8582 4832 8599
rect 3695 8582 3712 8599
rect 4815 8582 4832 8599
rect 3935 8582 3952 8599
rect 4295 8582 4312 8599
rect 4535 8582 4552 8599
rect 4855 8582 4872 8599
rect 3975 8582 3992 8599
rect 4615 8582 4632 8599
rect 4055 8582 4072 8599
rect 4175 8582 4192 8599
rect 4255 8582 4272 8599
rect 3855 8582 3872 8599
rect 4375 8582 4392 8599
rect 4735 8582 4752 8599
rect 3975 8582 3992 8599
rect 4775 8582 4792 8599
rect 3815 8582 3832 8599
rect 4335 8582 4352 8599
rect 4215 8582 4232 8599
rect 4455 8582 4472 8599
rect 4175 8582 4192 8599
rect 4215 8582 4232 8599
rect 3895 8582 3912 8599
rect 4335 8582 4352 8599
rect 4135 8582 4152 8599
rect 4295 8582 4312 8599
rect 4615 8582 4632 8599
rect 3735 8582 3752 8599
rect 3815 8582 3832 8599
rect 3775 8582 3792 8599
rect 4415 8582 4432 8599
rect 3775 8582 3792 8599
rect 4535 8582 4552 8599
rect 4855 8582 4872 8599
rect 3935 8582 3952 8599
rect 3735 8582 3752 8599
rect 4775 8582 4792 8599
rect 4455 8582 4472 8599
rect 4495 8582 4512 8599
rect 4375 8582 4392 8599
rect 4255 8582 4272 8599
rect 4135 8582 4152 8599
rect 4415 8582 4432 8599
rect 4015 8582 4032 8599
rect 3855 8582 3872 8599
rect 4095 8582 4112 8599
rect 4055 8582 4072 8599
rect 4695 8582 4712 8599
rect 4015 8582 4032 8599
rect 4575 8582 4592 8599
rect 3695 8582 3712 8599
rect 4655 8582 4672 8599
rect 3015 8582 3032 8599
rect 2655 8582 2672 8599
rect 3615 8582 3632 8599
rect 2735 8582 2752 8599
rect 2615 8582 2632 8599
rect 2975 8582 2992 8599
rect 2935 8582 2952 8599
rect 3175 8582 3192 8599
rect 3335 8582 3352 8599
rect 3215 8582 3232 8599
rect 3335 8582 3352 8599
rect 3455 8582 3472 8599
rect 2815 8582 2832 8599
rect 3375 8582 3392 8599
rect 3295 8582 3312 8599
rect 2775 8582 2792 8599
rect 2975 8582 2992 8599
rect 2535 8582 2552 8599
rect 3535 8582 3552 8599
rect 3135 8582 3152 8599
rect 2935 8582 2952 8599
rect 3175 8582 3192 8599
rect 2495 8582 2512 8599
rect 3615 8582 3632 8599
rect 3215 8582 3232 8599
rect 2855 8582 2872 8599
rect 3575 8582 3592 8599
rect 2855 8582 2872 8599
rect 3015 8582 3032 8599
rect 2895 8582 2912 8599
rect 3095 8582 3112 8599
rect 2895 8582 2912 8599
rect 2735 8582 2752 8599
rect 2655 8582 2672 8599
rect 3575 8582 3592 8599
rect 2575 8582 2592 8599
rect 2575 8582 2592 8599
rect 3655 8582 3672 8599
rect 2695 8582 2712 8599
rect 2495 8582 2512 8599
rect 2615 8582 2632 8599
rect 3495 8582 3512 8599
rect 3495 8582 3512 8599
rect 3455 8582 3472 8599
rect 3255 8582 3272 8599
rect 2535 8582 2552 8599
rect 2775 8582 2792 8599
rect 3535 8582 3552 8599
rect 3655 8582 3672 8599
rect 2815 8582 2832 8599
rect 3295 8582 3312 8599
rect 3415 8582 3432 8599
rect 3055 8582 3072 8599
rect 2695 8582 2712 8599
rect 3055 8582 3072 8599
rect 3095 8582 3112 8599
rect 3415 8582 3432 8599
rect 3135 8582 3152 8599
rect 3375 8582 3392 8599
rect 3255 8582 3272 8599
rect 1895 8582 1912 8599
rect 2215 8582 2232 8599
rect 2415 8582 2432 8599
rect 2095 8582 2112 8599
rect 2415 8582 2432 8599
rect 2015 8582 2032 8599
rect 2135 8582 2152 8599
rect 1935 8582 1952 8599
rect 2255 8582 2272 8599
rect 2215 8582 2232 8599
rect 316 8582 333 8599
rect 2175 8582 2192 8599
rect 2375 8582 2392 8599
rect 596 8582 613 8599
rect 476 8582 493 8599
rect 196 8582 213 8599
rect 956 8582 973 8599
rect 1036 8582 1053 8599
rect 2055 8582 2072 8599
rect 836 8582 853 8599
rect 2295 8582 2312 8599
rect 996 8582 1013 8599
rect 556 8582 573 8599
rect 1076 8582 1093 8599
rect 236 8582 253 8599
rect 2255 8582 2272 8599
rect 636 8582 653 8599
rect 276 8582 293 8599
rect 2335 8582 2352 8599
rect 676 8582 693 8599
rect 916 8582 933 8599
rect 1116 8582 1133 8599
rect 356 8582 373 8599
rect 1975 8582 1992 8599
rect 716 8582 733 8599
rect 1935 8582 1952 8599
rect 1895 8582 1912 8599
rect 2015 8582 2032 8599
rect 2135 8582 2152 8599
rect 756 8582 773 8599
rect 436 8582 453 8599
rect 1975 8582 1992 8599
rect 796 8582 813 8599
rect 2095 8582 2112 8599
rect 156 8582 173 8599
rect 2455 8582 2472 8599
rect 1156 8582 1173 8599
rect 2175 8582 2192 8599
rect 116 8582 133 8599
rect 2055 8582 2072 8599
rect 2455 8582 2472 8599
rect 396 8582 413 8599
rect 516 8582 533 8599
rect 2295 8582 2312 8599
rect 876 8582 893 8599
rect 2335 8582 2352 8599
rect 2375 8582 2392 8599
rect 6055 4652 6072 4669
rect 6055 4652 6072 4669
rect 6055 4652 6072 4669
rect 6055 4652 6072 4669
rect 6655 4652 6672 4669
rect 6655 4652 6672 4669
rect 6655 4652 6672 4669
rect 6655 4652 6672 4669
rect 7015 4652 7032 4669
rect 6735 4652 6752 4669
rect 6895 4652 6912 4669
rect 6975 4652 6992 4669
rect 6815 4652 6832 4669
rect 7055 4652 7072 4669
rect 6975 4652 6992 4669
rect 6975 4652 6992 4669
rect 7015 4652 7032 4669
rect 6735 4652 6752 4669
rect 7175 4652 7192 4669
rect 6775 4652 6792 4669
rect 6935 4652 6952 4669
rect 7215 4652 7232 4669
rect 6855 4652 6872 4669
rect 7055 4652 7072 4669
rect 7095 4652 7112 4669
rect 6855 4652 6872 4669
rect 7175 4652 7192 4669
rect 7215 4652 7232 4669
rect 6895 4652 6912 4669
rect 6695 4652 6712 4669
rect 6855 4652 6872 4669
rect 7055 4652 7072 4669
rect 6815 4652 6832 4669
rect 7215 4652 7232 4669
rect 6735 4652 6752 4669
rect 6935 4652 6952 4669
rect 7095 4652 7112 4669
rect 7175 4652 7192 4669
rect 6935 4652 6952 4669
rect 6775 4652 6792 4669
rect 6855 4652 6872 4669
rect 7135 4652 7152 4669
rect 6815 4652 6832 4669
rect 6775 4652 6792 4669
rect 6895 4652 6912 4669
rect 7015 4652 7032 4669
rect 6895 4652 6912 4669
rect 7135 4652 7152 4669
rect 7055 4652 7072 4669
rect 6695 4652 6712 4669
rect 6735 4652 6752 4669
rect 7015 4652 7032 4669
rect 6975 4652 6992 4669
rect 6815 4652 6832 4669
rect 7135 4652 7152 4669
rect 6695 4652 6712 4669
rect 7095 4652 7112 4669
rect 6935 4652 6952 4669
rect 7215 4652 7232 4669
rect 6775 4652 6792 4669
rect 7095 4652 7112 4669
rect 6695 4652 6712 4669
rect 7175 4652 7192 4669
rect 7135 4652 7152 4669
rect 6295 4652 6312 4669
rect 6375 4652 6392 4669
rect 6535 4652 6552 4669
rect 6495 4652 6512 4669
rect 6255 4652 6272 4669
rect 6415 4652 6432 4669
rect 6175 4652 6192 4669
rect 6135 4652 6152 4669
rect 6095 4652 6112 4669
rect 6255 4652 6272 4669
rect 6615 4652 6632 4669
rect 6175 4652 6192 4669
rect 6455 4652 6472 4669
rect 6135 4652 6152 4669
rect 6095 4652 6112 4669
rect 6295 4652 6312 4669
rect 6495 4652 6512 4669
rect 6215 4652 6232 4669
rect 6575 4652 6592 4669
rect 6535 4652 6552 4669
rect 6335 4652 6352 4669
rect 6575 4652 6592 4669
rect 6335 4652 6352 4669
rect 6455 4652 6472 4669
rect 6215 4652 6232 4669
rect 6415 4652 6432 4669
rect 6615 4652 6632 4669
rect 6255 4652 6272 4669
rect 6415 4652 6432 4669
rect 6455 4652 6472 4669
rect 6175 4652 6192 4669
rect 6455 4652 6472 4669
rect 6135 4652 6152 4669
rect 6095 4652 6112 4669
rect 6295 4652 6312 4669
rect 6335 4652 6352 4669
rect 6335 4652 6352 4669
rect 6175 4652 6192 4669
rect 6495 4652 6512 4669
rect 6375 4652 6392 4669
rect 6375 4652 6392 4669
rect 6215 4652 6232 4669
rect 6615 4652 6632 4669
rect 6135 4652 6152 4669
rect 6415 4652 6432 4669
rect 6575 4652 6592 4669
rect 6535 4652 6552 4669
rect 6095 4652 6112 4669
rect 6535 4652 6552 4669
rect 6575 4652 6592 4669
rect 6375 4652 6392 4669
rect 6615 4652 6632 4669
rect 6295 4652 6312 4669
rect 6495 4652 6512 4669
rect 6255 4652 6272 4669
rect 6215 4652 6232 4669
rect 5455 4652 5472 4669
rect 5455 4652 5472 4669
rect 5455 4652 5472 4669
rect 5455 4652 5472 4669
rect 5655 4652 5672 4669
rect 5655 4652 5672 4669
rect 5815 4652 5832 4669
rect 5975 4652 5992 4669
rect 5735 4652 5752 4669
rect 5975 4652 5992 4669
rect 5535 4652 5552 4669
rect 5775 4652 5792 4669
rect 6015 4652 6032 4669
rect 5815 4652 5832 4669
rect 5855 4652 5872 4669
rect 5695 4652 5712 4669
rect 5735 4652 5752 4669
rect 5895 4652 5912 4669
rect 5615 4652 5632 4669
rect 5775 4652 5792 4669
rect 5615 4652 5632 4669
rect 5495 4652 5512 4669
rect 5615 4652 5632 4669
rect 6015 4652 6032 4669
rect 5535 4652 5552 4669
rect 5495 4652 5512 4669
rect 5815 4652 5832 4669
rect 5935 4652 5952 4669
rect 5655 4652 5672 4669
rect 5575 4652 5592 4669
rect 5895 4652 5912 4669
rect 5655 4652 5672 4669
rect 5615 4652 5632 4669
rect 5575 4652 5592 4669
rect 5575 4652 5592 4669
rect 5735 4652 5752 4669
rect 5935 4652 5952 4669
rect 5575 4652 5592 4669
rect 5855 4652 5872 4669
rect 5895 4652 5912 4669
rect 5695 4652 5712 4669
rect 5935 4652 5952 4669
rect 5775 4652 5792 4669
rect 5855 4652 5872 4669
rect 6015 4652 6032 4669
rect 5975 4652 5992 4669
rect 5815 4652 5832 4669
rect 5855 4652 5872 4669
rect 5535 4652 5552 4669
rect 5775 4652 5792 4669
rect 5695 4652 5712 4669
rect 5495 4652 5512 4669
rect 6015 4652 6032 4669
rect 5975 4652 5992 4669
rect 5695 4652 5712 4669
rect 5895 4652 5912 4669
rect 5935 4652 5952 4669
rect 5495 4652 5512 4669
rect 5735 4652 5752 4669
rect 5535 4652 5552 4669
rect 5415 4652 5432 4669
rect 5375 4652 5392 4669
rect 4935 4652 4952 4669
rect 5415 4652 5432 4669
rect 5335 4652 5352 4669
rect 4895 4652 4912 4669
rect 5295 4652 5312 4669
rect 5255 4652 5272 4669
rect 4895 4652 4912 4669
rect 5215 4652 5232 4669
rect 5175 4652 5192 4669
rect 5295 4652 5312 4669
rect 5135 4652 5152 4669
rect 5255 4652 5272 4669
rect 5215 4652 5232 4669
rect 5375 4652 5392 4669
rect 5175 4652 5192 4669
rect 5135 4652 5152 4669
rect 5055 4652 5072 4669
rect 5055 4652 5072 4669
rect 5335 4652 5352 4669
rect 5095 4652 5112 4669
rect 5015 4652 5032 4669
rect 5095 4652 5112 4669
rect 4935 4652 4952 4669
rect 4975 4652 4992 4669
rect 5215 4652 5232 4669
rect 5255 4652 5272 4669
rect 5175 4652 5192 4669
rect 5335 4652 5352 4669
rect 5295 4652 5312 4669
rect 5135 4652 5152 4669
rect 4975 4652 4992 4669
rect 5415 4652 5432 4669
rect 5415 4652 5432 4669
rect 4895 4652 4912 4669
rect 5135 4652 5152 4669
rect 5015 4652 5032 4669
rect 5375 4652 5392 4669
rect 5095 4652 5112 4669
rect 4935 4652 4952 4669
rect 4895 4652 4912 4669
rect 5055 4652 5072 4669
rect 4975 4652 4992 4669
rect 5255 4652 5272 4669
rect 5215 4652 5232 4669
rect 5055 4652 5072 4669
rect 5015 4652 5032 4669
rect 4935 4652 4952 4669
rect 5175 4652 5192 4669
rect 5295 4652 5312 4669
rect 5015 4652 5032 4669
rect 5335 4652 5352 4669
rect 5375 4652 5392 4669
rect 5095 4652 5112 4669
rect 4975 4652 4992 4669
rect 9216 4652 9233 4669
rect 9056 4652 9073 4669
rect 9136 4652 9153 4669
rect 9376 4652 9393 4669
rect 9296 4652 9313 4669
rect 9176 4652 9193 4669
rect 9176 4652 9193 4669
rect 9136 4652 9153 4669
rect 9096 4652 9113 4669
rect 9376 4652 9393 4669
rect 9416 4652 9433 4669
rect 9056 4652 9073 4669
rect 9336 4652 9353 4669
rect 9376 4652 9393 4669
rect 9416 4652 9433 4669
rect 9096 4652 9113 4669
rect 9336 4652 9353 4669
rect 9256 4652 9273 4669
rect 9056 4652 9073 4669
rect 9296 4652 9313 4669
rect 9296 4652 9313 4669
rect 9336 4652 9353 4669
rect 9416 4652 9433 4669
rect 9096 4652 9113 4669
rect 9616 4652 9633 4669
rect 9256 4652 9273 4669
rect 9576 4652 9593 4669
rect 9216 4652 9233 4669
rect 9536 4652 9553 4669
rect 9216 4652 9233 4669
rect 9376 4652 9393 4669
rect 9496 4652 9513 4669
rect 9176 4652 9193 4669
rect 9176 4652 9193 4669
rect 9136 4652 9153 4669
rect 9096 4652 9113 4669
rect 9416 4652 9433 4669
rect 9056 4652 9073 4669
rect 9456 4652 9473 4669
rect 9296 4652 9313 4669
rect 9616 4652 9633 4669
rect 9576 4652 9593 4669
rect 9616 4652 9633 4669
rect 9576 4652 9593 4669
rect 9536 4652 9553 4669
rect 9496 4652 9513 4669
rect 9456 4652 9473 4669
rect 9616 4652 9633 4669
rect 9576 4652 9593 4669
rect 9536 4652 9553 4669
rect 9496 4652 9513 4669
rect 9456 4652 9473 4669
rect 9536 4652 9553 4669
rect 9496 4652 9513 4669
rect 9456 4652 9473 4669
rect 9136 4652 9153 4669
rect 9256 4652 9273 4669
rect 9336 4652 9353 4669
rect 9216 4652 9233 4669
rect 9256 4652 9273 4669
rect 8616 4652 8633 4669
rect 8616 4652 8633 4669
rect 8896 4652 8913 4669
rect 8856 4652 8873 4669
rect 8896 4652 8913 4669
rect 8816 4652 8833 4669
rect 8776 4652 8793 4669
rect 8856 4652 8873 4669
rect 8736 4652 8753 4669
rect 8696 4652 8713 4669
rect 8816 4652 8833 4669
rect 8656 4652 8673 4669
rect 8456 4652 8473 4669
rect 8776 4652 8793 4669
rect 8736 4652 8753 4669
rect 9016 4652 9033 4669
rect 8696 4652 8713 4669
rect 8656 4652 8673 4669
rect 8976 4652 8993 4669
rect 8576 4652 8593 4669
rect 8936 4652 8953 4669
rect 8496 4652 8513 4669
rect 9016 4652 9033 4669
rect 8976 4652 8993 4669
rect 8936 4652 8953 4669
rect 8536 4652 8553 4669
rect 8536 4652 8553 4669
rect 8496 4652 8513 4669
rect 8576 4652 8593 4669
rect 8456 4652 8473 4669
rect 8616 4652 8633 4669
rect 8616 4652 8633 4669
rect 8896 4652 8913 4669
rect 8856 4652 8873 4669
rect 8896 4652 8913 4669
rect 8816 4652 8833 4669
rect 8776 4652 8793 4669
rect 8856 4652 8873 4669
rect 8736 4652 8753 4669
rect 8696 4652 8713 4669
rect 8816 4652 8833 4669
rect 8656 4652 8673 4669
rect 8776 4652 8793 4669
rect 8736 4652 8753 4669
rect 9016 4652 9033 4669
rect 8696 4652 8713 4669
rect 8656 4652 8673 4669
rect 8976 4652 8993 4669
rect 8936 4652 8953 4669
rect 9016 4652 9033 4669
rect 8976 4652 8993 4669
rect 8936 4652 8953 4669
rect 8536 4652 8553 4669
rect 8536 4652 8553 4669
rect 8496 4652 8513 4669
rect 8576 4652 8593 4669
rect 8456 4652 8473 4669
rect 8496 4652 8513 4669
rect 8456 4652 8473 4669
rect 8576 4652 8593 4669
rect 7935 4652 7952 4669
rect 7975 4652 7992 4669
rect 8055 4652 8072 4669
rect 8255 4652 8272 4669
rect 7895 4652 7912 4669
rect 8416 4652 8433 4669
rect 8015 4652 8032 4669
rect 8135 4652 8152 4669
rect 7975 4652 7992 4669
rect 8015 4652 8032 4669
rect 8295 4652 8312 4669
rect 7935 4652 7952 4669
rect 8215 4652 8232 4669
rect 7935 4652 7952 4669
rect 7855 4652 7872 4669
rect 8095 4652 8112 4669
rect 8376 4652 8393 4669
rect 8255 4652 8272 4669
rect 8175 4652 8192 4669
rect 8416 4652 8433 4669
rect 8015 4652 8032 4669
rect 8335 4652 8352 4669
rect 8416 4652 8433 4669
rect 8055 4652 8072 4669
rect 8135 4652 8152 4669
rect 8215 4652 8232 4669
rect 7895 4652 7912 4669
rect 8335 4652 8352 4669
rect 8335 4652 8352 4669
rect 7895 4652 7912 4669
rect 8055 4652 8072 4669
rect 8175 4652 8192 4669
rect 8295 4652 8312 4669
rect 8295 4652 8312 4669
rect 8255 4652 8272 4669
rect 8376 4652 8393 4669
rect 8135 4652 8152 4669
rect 8255 4652 8272 4669
rect 8215 4652 8232 4669
rect 8175 4652 8192 4669
rect 7895 4652 7912 4669
rect 7855 4652 7872 4669
rect 8175 4652 8192 4669
rect 7855 4652 7872 4669
rect 8376 4652 8393 4669
rect 8135 4652 8152 4669
rect 8095 4652 8112 4669
rect 8095 4652 8112 4669
rect 8416 4652 8433 4669
rect 8376 4652 8393 4669
rect 7855 4652 7872 4669
rect 8055 4652 8072 4669
rect 8015 4652 8032 4669
rect 8215 4652 8232 4669
rect 7975 4652 7992 4669
rect 8095 4652 8112 4669
rect 7975 4652 7992 4669
rect 8295 4652 8312 4669
rect 8335 4652 8352 4669
rect 7935 4652 7952 4669
rect 7815 4652 7832 4669
rect 7815 4652 7832 4669
rect 7655 4652 7672 4669
rect 7695 4652 7712 4669
rect 7575 4652 7592 4669
rect 7255 4652 7272 4669
rect 7735 4652 7752 4669
rect 7255 4652 7272 4669
rect 7815 4652 7832 4669
rect 7615 4652 7632 4669
rect 7655 4652 7672 4669
rect 7695 4652 7712 4669
rect 7535 4652 7552 4669
rect 7255 4652 7272 4669
rect 7775 4652 7792 4669
rect 7495 4652 7512 4669
rect 7575 4652 7592 4669
rect 7495 4652 7512 4669
rect 7735 4652 7752 4669
rect 7375 4652 7392 4669
rect 7255 4652 7272 4669
rect 7775 4652 7792 4669
rect 7335 4652 7352 4669
rect 7615 4652 7632 4669
rect 7295 4652 7312 4669
rect 7415 4652 7432 4669
rect 7375 4652 7392 4669
rect 7535 4652 7552 4669
rect 7335 4652 7352 4669
rect 7775 4652 7792 4669
rect 7495 4652 7512 4669
rect 7295 4652 7312 4669
rect 7495 4652 7512 4669
rect 7735 4652 7752 4669
rect 7375 4652 7392 4669
rect 7535 4652 7552 4669
rect 7335 4652 7352 4669
rect 7415 4652 7432 4669
rect 7295 4652 7312 4669
rect 7415 4652 7432 4669
rect 7375 4652 7392 4669
rect 7335 4652 7352 4669
rect 7295 4652 7312 4669
rect 7535 4652 7552 4669
rect 7415 4652 7432 4669
rect 7455 4652 7472 4669
rect 7455 4652 7472 4669
rect 7815 4652 7832 4669
rect 7695 4652 7712 4669
rect 7455 4652 7472 4669
rect 7775 4652 7792 4669
rect 7735 4652 7752 4669
rect 7655 4652 7672 4669
rect 7695 4652 7712 4669
rect 7655 4652 7672 4669
rect 7615 4652 7632 4669
rect 7615 4652 7632 4669
rect 7455 4652 7472 4669
rect 7575 4652 7592 4669
rect 7575 4652 7592 4669
rect 1895 4652 1912 4669
rect 2135 4652 2152 4669
rect 2095 4652 2112 4669
rect 2175 4652 2192 4669
rect 2055 4652 2072 4669
rect 2215 4652 2232 4669
rect 2015 4652 2032 4669
rect 2095 4652 2112 4669
rect 2215 4652 2232 4669
rect 2055 4652 2072 4669
rect 1975 4652 1992 4669
rect 2295 4652 2312 4669
rect 1935 4652 1952 4669
rect 2015 4652 2032 4669
rect 1895 4652 1912 4669
rect 2255 4652 2272 4669
rect 2455 4652 2472 4669
rect 2455 4652 2472 4669
rect 2415 4652 2432 4669
rect 2135 4652 2152 4669
rect 2375 4652 2392 4669
rect 2175 4652 2192 4669
rect 2415 4652 2432 4669
rect 1975 4652 1992 4669
rect 2335 4652 2352 4669
rect 2335 4652 2352 4669
rect 2295 4652 2312 4669
rect 2375 4652 2392 4669
rect 1935 4652 1952 4669
rect 2255 4652 2272 4669
rect 1895 4652 1912 4669
rect 2455 4652 2472 4669
rect 2335 4652 2352 4669
rect 2415 4652 2432 4669
rect 2335 4652 2352 4669
rect 1895 4652 1912 4669
rect 2295 4652 2312 4669
rect 1975 4652 1992 4669
rect 2135 4652 2152 4669
rect 2255 4652 2272 4669
rect 2055 4652 2072 4669
rect 1975 4652 1992 4669
rect 2415 4652 2432 4669
rect 2215 4652 2232 4669
rect 2015 4652 2032 4669
rect 2135 4652 2152 4669
rect 2095 4652 2112 4669
rect 2295 4652 2312 4669
rect 2255 4652 2272 4669
rect 2055 4652 2072 4669
rect 2015 4652 2032 4669
rect 2175 4652 2192 4669
rect 2455 4652 2472 4669
rect 2175 4652 2192 4669
rect 1935 4652 1952 4669
rect 2095 4652 2112 4669
rect 1935 4652 1952 4669
rect 2215 4652 2232 4669
rect 2375 4652 2392 4669
rect 2375 4652 2392 4669
rect 236 4652 253 4669
rect 316 4652 333 4669
rect 956 4652 973 4669
rect 556 4652 573 4669
rect 276 4652 293 4669
rect 716 4652 733 4669
rect 436 4652 453 4669
rect 1156 4652 1173 4669
rect 516 4652 533 4669
rect 356 4652 373 4669
rect 1116 4652 1133 4669
rect 876 4652 893 4669
rect 996 4652 1013 4669
rect 316 4652 333 4669
rect 356 4652 373 4669
rect 476 4652 493 4669
rect 396 4652 413 4669
rect 116 4652 133 4669
rect 396 4652 413 4669
rect 436 4652 453 4669
rect 476 4652 493 4669
rect 516 4652 533 4669
rect 196 4652 213 4669
rect 556 4652 573 4669
rect 596 4652 613 4669
rect 596 4652 613 4669
rect 636 4652 653 4669
rect 676 4652 693 4669
rect 796 4652 813 4669
rect 1036 4652 1053 4669
rect 156 4652 173 4669
rect 716 4652 733 4669
rect 916 4652 933 4669
rect 756 4652 773 4669
rect 796 4652 813 4669
rect 836 4652 853 4669
rect 876 4652 893 4669
rect 276 4652 293 4669
rect 916 4652 933 4669
rect 956 4652 973 4669
rect 236 4652 253 4669
rect 996 4652 1013 4669
rect 1076 4652 1093 4669
rect 1036 4652 1053 4669
rect 1076 4652 1093 4669
rect 676 4652 693 4669
rect 1116 4652 1133 4669
rect 836 4652 853 4669
rect 1156 4652 1173 4669
rect 116 4652 133 4669
rect 156 4652 173 4669
rect 636 4652 653 4669
rect 756 4652 773 4669
rect 196 4652 213 4669
rect 633 3967 650 3984
rect 4575 4652 4592 4669
rect 4615 4652 4632 4669
rect 4535 4652 4552 4669
rect 4655 4652 4672 4669
rect 4815 4652 4832 4669
rect 4455 4652 4472 4669
rect 4855 4652 4872 4669
rect 4335 4652 4352 4669
rect 4535 4652 4552 4669
rect 4415 4652 4432 4669
rect 4855 4652 4872 4669
rect 4375 4652 4392 4669
rect 4335 4652 4352 4669
rect 4295 4652 4312 4669
rect 4295 4652 4312 4669
rect 4455 4652 4472 4669
rect 4375 4652 4392 4669
rect 4855 4652 4872 4669
rect 4415 4652 4432 4669
rect 4735 4652 4752 4669
rect 4695 4652 4712 4669
rect 4495 4652 4512 4669
rect 4695 4652 4712 4669
rect 4695 4652 4712 4669
rect 4735 4652 4752 4669
rect 4775 4652 4792 4669
rect 4855 4652 4872 4669
rect 4415 4652 4432 4669
rect 4655 4652 4672 4669
rect 4495 4652 4512 4669
rect 4535 4652 4552 4669
rect 4375 4652 4392 4669
rect 4615 4652 4632 4669
rect 4335 4652 4352 4669
rect 4815 4652 4832 4669
rect 4535 4652 4552 4669
rect 4775 4652 4792 4669
rect 4415 4652 4432 4669
rect 4775 4652 4792 4669
rect 4735 4652 4752 4669
rect 4655 4652 4672 4669
rect 4295 4652 4312 4669
rect 4615 4652 4632 4669
rect 4815 4652 4832 4669
rect 4575 4652 4592 4669
rect 4815 4652 4832 4669
rect 4495 4652 4512 4669
rect 4655 4652 4672 4669
rect 4695 4652 4712 4669
rect 4495 4652 4512 4669
rect 4575 4652 4592 4669
rect 4775 4652 4792 4669
rect 4455 4652 4472 4669
rect 4615 4652 4632 4669
rect 4375 4652 4392 4669
rect 4335 4652 4352 4669
rect 4295 4652 4312 4669
rect 4575 4652 4592 4669
rect 4735 4652 4752 4669
rect 4455 4652 4472 4669
rect 3775 4652 3792 4669
rect 3735 4652 3752 4669
rect 3695 4652 3712 4669
rect 4015 4652 4032 4669
rect 3975 4652 3992 4669
rect 3935 4652 3952 4669
rect 3895 4652 3912 4669
rect 3855 4652 3872 4669
rect 3815 4652 3832 4669
rect 4055 4652 4072 4669
rect 4255 4652 4272 4669
rect 4215 4652 4232 4669
rect 4175 4652 4192 4669
rect 4095 4652 4112 4669
rect 4135 4652 4152 4669
rect 3775 4652 3792 4669
rect 4095 4652 4112 4669
rect 4055 4652 4072 4669
rect 4255 4652 4272 4669
rect 4215 4652 4232 4669
rect 4015 4652 4032 4669
rect 4175 4652 4192 4669
rect 4095 4652 4112 4669
rect 3975 4652 3992 4669
rect 4135 4652 4152 4669
rect 3775 4652 3792 4669
rect 3935 4652 3952 4669
rect 4095 4652 4112 4669
rect 3735 4652 3752 4669
rect 4055 4652 4072 4669
rect 3895 4652 3912 4669
rect 3695 4652 3712 4669
rect 3815 4652 3832 4669
rect 4255 4652 4272 4669
rect 4015 4652 4032 4669
rect 3975 4652 3992 4669
rect 3855 4652 3872 4669
rect 4215 4652 4232 4669
rect 3935 4652 3952 4669
rect 4175 4652 4192 4669
rect 3895 4652 3912 4669
rect 3775 4652 3792 4669
rect 4135 4652 4152 4669
rect 3855 4652 3872 4669
rect 3815 4652 3832 4669
rect 3735 4652 3752 4669
rect 3695 4652 3712 4669
rect 3975 4652 3992 4669
rect 4215 4652 4232 4669
rect 3935 4652 3952 4669
rect 4175 4652 4192 4669
rect 3895 4652 3912 4669
rect 4135 4652 4152 4669
rect 3855 4652 3872 4669
rect 3735 4652 3752 4669
rect 4055 4652 4072 4669
rect 3695 4652 3712 4669
rect 4255 4652 4272 4669
rect 4015 4652 4032 4669
rect 3815 4652 3832 4669
rect 3255 4652 3272 4669
rect 3335 4652 3352 4669
rect 3535 4652 3552 4669
rect 3415 4652 3432 4669
rect 3255 4652 3272 4669
rect 3455 4652 3472 4669
rect 3095 4652 3112 4669
rect 3335 4652 3352 4669
rect 3255 4652 3272 4669
rect 3615 4652 3632 4669
rect 3655 4652 3672 4669
rect 3255 4652 3272 4669
rect 3215 4652 3232 4669
rect 3575 4652 3592 4669
rect 3295 4652 3312 4669
rect 3375 4652 3392 4669
rect 3655 4652 3672 4669
rect 3495 4652 3512 4669
rect 3415 4652 3432 4669
rect 3495 4652 3512 4669
rect 3135 4652 3152 4669
rect 3535 4652 3552 4669
rect 3215 4652 3232 4669
rect 3575 4652 3592 4669
rect 3415 4652 3432 4669
rect 3095 4652 3112 4669
rect 3135 4652 3152 4669
rect 3335 4652 3352 4669
rect 3215 4652 3232 4669
rect 3135 4652 3152 4669
rect 3095 4652 3112 4669
rect 3495 4652 3512 4669
rect 3615 4652 3632 4669
rect 3415 4652 3432 4669
rect 3175 4652 3192 4669
rect 3455 4652 3472 4669
rect 3175 4652 3192 4669
rect 3375 4652 3392 4669
rect 3175 4652 3192 4669
rect 3535 4652 3552 4669
rect 3615 4652 3632 4669
rect 3495 4652 3512 4669
rect 3335 4652 3352 4669
rect 3375 4652 3392 4669
rect 3175 4652 3192 4669
rect 3295 4652 3312 4669
rect 3295 4652 3312 4669
rect 3655 4652 3672 4669
rect 3375 4652 3392 4669
rect 3135 4652 3152 4669
rect 3295 4652 3312 4669
rect 3575 4652 3592 4669
rect 3615 4652 3632 4669
rect 3455 4652 3472 4669
rect 3655 4652 3672 4669
rect 3535 4652 3552 4669
rect 3575 4652 3592 4669
rect 3095 4652 3112 4669
rect 3455 4652 3472 4669
rect 3215 4652 3232 4669
rect 2975 4652 2992 4669
rect 2895 4652 2912 4669
rect 2775 4652 2792 4669
rect 2735 4652 2752 4669
rect 3015 4652 3032 4669
rect 3055 4652 3072 4669
rect 2535 4652 2552 4669
rect 2615 4652 2632 4669
rect 2735 4652 2752 4669
rect 2495 4652 2512 4669
rect 2855 4652 2872 4669
rect 2575 4652 2592 4669
rect 2815 4652 2832 4669
rect 2975 4652 2992 4669
rect 2695 4652 2712 4669
rect 2815 4652 2832 4669
rect 2655 4652 2672 4669
rect 2775 4652 2792 4669
rect 2935 4652 2952 4669
rect 2855 4652 2872 4669
rect 2655 4652 2672 4669
rect 2495 4652 2512 4669
rect 2535 4652 2552 4669
rect 3055 4652 3072 4669
rect 2695 4652 2712 4669
rect 2615 4652 2632 4669
rect 2895 4652 2912 4669
rect 2575 4652 2592 4669
rect 3015 4652 3032 4669
rect 2935 4652 2952 4669
rect 3055 4652 3072 4669
rect 2775 4652 2792 4669
rect 2495 4652 2512 4669
rect 2735 4652 2752 4669
rect 2895 4652 2912 4669
rect 2855 4652 2872 4669
rect 3015 4652 3032 4669
rect 2575 4652 2592 4669
rect 2655 4652 2672 4669
rect 2735 4652 2752 4669
rect 2975 4652 2992 4669
rect 2815 4652 2832 4669
rect 2695 4652 2712 4669
rect 2615 4652 2632 4669
rect 2695 4652 2712 4669
rect 2935 4652 2952 4669
rect 2775 4652 2792 4669
rect 2655 4652 2672 4669
rect 2535 4652 2552 4669
rect 3055 4652 3072 4669
rect 2615 4652 2632 4669
rect 2895 4652 2912 4669
rect 3015 4652 3032 4669
rect 2935 4652 2952 4669
rect 2855 4652 2872 4669
rect 2975 4652 2992 4669
rect 2575 4652 2592 4669
rect 2535 4652 2552 4669
rect 2495 4652 2512 4669
rect 2815 4652 2832 4669
rect 2481 2394 2498 2411
rect 4836 3163 4853 3180
rect 4836 3163 4853 3180
rect 4836 3163 4853 3180
rect 4836 3163 4853 3180
rect 4276 3163 4293 3180
rect 4276 3163 4293 3180
rect 4276 3163 4293 3180
rect 4276 3163 4293 3180
rect 4796 3163 4813 3180
rect 4796 3163 4813 3180
rect 4636 3163 4653 3180
rect 4756 3163 4773 3180
rect 4636 3163 4653 3180
rect 4716 3163 4733 3180
rect 4716 3163 4733 3180
rect 4596 3163 4613 3180
rect 4436 3163 4453 3180
rect 4356 3163 4373 3180
rect 4676 3163 4693 3180
rect 4756 3163 4773 3180
rect 4676 3163 4693 3180
rect 4316 3163 4333 3180
rect 4516 3163 4533 3180
rect 4556 3163 4573 3180
rect 4356 3163 4373 3180
rect 4756 3163 4773 3180
rect 4556 3163 4573 3180
rect 4476 3163 4493 3180
rect 4636 3163 4653 3180
rect 4356 3163 4373 3180
rect 4756 3163 4773 3180
rect 4516 3163 4533 3180
rect 4716 3163 4733 3180
rect 4316 3163 4333 3180
rect 4516 3163 4533 3180
rect 4316 3163 4333 3180
rect 4476 3163 4493 3180
rect 4596 3163 4613 3180
rect 4676 3163 4693 3180
rect 4556 3163 4573 3180
rect 4596 3163 4613 3180
rect 4396 3163 4413 3180
rect 4796 3163 4813 3180
rect 4796 3163 4813 3180
rect 4516 3163 4533 3180
rect 4476 3163 4493 3180
rect 4556 3163 4573 3180
rect 4436 3163 4453 3180
rect 4476 3163 4493 3180
rect 4676 3163 4693 3180
rect 4436 3163 4453 3180
rect 4316 3163 4333 3180
rect 4396 3163 4413 3180
rect 4436 3163 4453 3180
rect 4636 3163 4653 3180
rect 4716 3163 4733 3180
rect 4596 3163 4613 3180
rect 4356 3163 4373 3180
rect 4396 3163 4413 3180
rect 4396 3163 4413 3180
rect 3836 3163 3853 3180
rect 3876 3163 3893 3180
rect 3796 3163 3813 3180
rect 4036 3163 4053 3180
rect 4236 3163 4253 3180
rect 3916 3163 3933 3180
rect 3956 3163 3973 3180
rect 4116 3163 4133 3180
rect 3956 3163 3973 3180
rect 3836 3163 3853 3180
rect 3756 3163 3773 3180
rect 4116 3163 4133 3180
rect 4196 3163 4213 3180
rect 3796 3163 3813 3180
rect 3796 3163 3813 3180
rect 3756 3163 3773 3180
rect 4076 3163 4093 3180
rect 3836 3163 3853 3180
rect 4236 3163 4253 3180
rect 4076 3163 4093 3180
rect 4196 3163 4213 3180
rect 4196 3163 4213 3180
rect 3916 3163 3933 3180
rect 4156 3163 4173 3180
rect 3756 3163 3773 3180
rect 4156 3163 4173 3180
rect 4156 3163 4173 3180
rect 4036 3163 4053 3180
rect 4236 3163 4253 3180
rect 4156 3163 4173 3180
rect 4076 3163 4093 3180
rect 4036 3163 4053 3180
rect 3956 3163 3973 3180
rect 3876 3163 3893 3180
rect 4196 3163 4213 3180
rect 3876 3163 3893 3180
rect 3756 3163 3773 3180
rect 4116 3163 4133 3180
rect 3876 3163 3893 3180
rect 4076 3163 4093 3180
rect 3796 3163 3813 3180
rect 4036 3163 4053 3180
rect 3916 3163 3933 3180
rect 3996 3163 4013 3180
rect 4116 3163 4133 3180
rect 3836 3163 3853 3180
rect 3996 3163 4013 3180
rect 3996 3163 4013 3180
rect 3996 3163 4013 3180
rect 3956 3163 3973 3180
rect 4236 3163 4253 3180
rect 3916 3163 3933 3180
rect 3196 3163 3213 3180
rect 3196 3163 3213 3180
rect 3196 3163 3213 3180
rect 3196 3163 3213 3180
rect 3356 3163 3373 3180
rect 3636 3163 3653 3180
rect 3396 3163 3413 3180
rect 3596 3163 3613 3180
rect 3276 3163 3293 3180
rect 3676 3163 3693 3180
rect 3396 3163 3413 3180
rect 3316 3163 3333 3180
rect 3476 3163 3493 3180
rect 3396 3163 3413 3180
rect 3636 3163 3653 3180
rect 3716 3163 3733 3180
rect 3636 3163 3653 3180
rect 3316 3163 3333 3180
rect 3556 3163 3573 3180
rect 3596 3163 3613 3180
rect 3636 3163 3653 3180
rect 3596 3163 3613 3180
rect 3556 3163 3573 3180
rect 3236 3163 3253 3180
rect 3436 3163 3453 3180
rect 3716 3163 3733 3180
rect 3516 3163 3533 3180
rect 3716 3163 3733 3180
rect 3556 3163 3573 3180
rect 3436 3163 3453 3180
rect 3676 3163 3693 3180
rect 3556 3163 3573 3180
rect 3316 3163 3333 3180
rect 3516 3163 3533 3180
rect 3276 3163 3293 3180
rect 3356 3163 3373 3180
rect 3596 3163 3613 3180
rect 3396 3163 3413 3180
rect 3476 3163 3493 3180
rect 3236 3163 3253 3180
rect 3316 3163 3333 3180
rect 3476 3163 3493 3180
rect 3716 3163 3733 3180
rect 3436 3163 3453 3180
rect 3276 3163 3293 3180
rect 3236 3163 3253 3180
rect 3476 3163 3493 3180
rect 3236 3163 3253 3180
rect 3276 3163 3293 3180
rect 3356 3163 3373 3180
rect 3516 3163 3533 3180
rect 3516 3163 3533 3180
rect 3676 3163 3693 3180
rect 3436 3163 3453 3180
rect 3676 3163 3693 3180
rect 3356 3163 3373 3180
rect 3076 3163 3093 3180
rect 3116 3163 3133 3180
rect 2876 3163 2893 3180
rect 2996 3163 3013 3180
rect 3036 3163 3053 3180
rect 3076 3163 3093 3180
rect 3116 3163 3133 3180
rect 3116 3163 3133 3180
rect 2796 3163 2813 3180
rect 2996 3163 3013 3180
rect 2796 3163 2813 3180
rect 2676 3163 2693 3180
rect 2876 3163 2893 3180
rect 3116 3163 3133 3180
rect 2836 3163 2853 3180
rect 2916 3163 2933 3180
rect 3036 3163 3053 3180
rect 3076 3163 3093 3180
rect 2916 3163 2933 3180
rect 2796 3163 2813 3180
rect 2756 3163 2773 3180
rect 2716 3163 2733 3180
rect 3076 3163 3093 3180
rect 2836 3163 2853 3180
rect 3036 3163 3053 3180
rect 2836 3163 2853 3180
rect 2676 3163 2693 3180
rect 2836 3163 2853 3180
rect 2796 3163 2813 3180
rect 2956 3163 2973 3180
rect 2676 3163 2693 3180
rect 2876 3163 2893 3180
rect 2716 3163 2733 3180
rect 2956 3163 2973 3180
rect 2916 3163 2933 3180
rect 2716 3163 2733 3180
rect 2956 3163 2973 3180
rect 2956 3163 2973 3180
rect 3036 3163 3053 3180
rect 3156 3163 3173 3180
rect 2676 3163 2693 3180
rect 2876 3163 2893 3180
rect 2756 3163 2773 3180
rect 2996 3163 3013 3180
rect 2716 3163 2733 3180
rect 2996 3163 3013 3180
rect 3156 3163 3173 3180
rect 3156 3163 3173 3180
rect 2756 3163 2773 3180
rect 2916 3163 2933 3180
rect 3156 3163 3173 3180
rect 2756 3163 2773 3180
rect 2116 3163 2133 3180
rect 2116 3163 2133 3180
rect 2116 3163 2133 3180
rect 2116 3163 2133 3180
rect 2236 3163 2253 3180
rect 2196 3163 2213 3180
rect 2556 3163 2573 3180
rect 2636 3163 2653 3180
rect 2596 3163 2613 3180
rect 2276 3163 2293 3180
rect 2276 3163 2293 3180
rect 2516 3163 2533 3180
rect 2436 3163 2453 3180
rect 2316 3163 2333 3180
rect 2596 3163 2613 3180
rect 2596 3163 2613 3180
rect 2156 3163 2173 3180
rect 2596 3163 2613 3180
rect 2636 3163 2653 3180
rect 2636 3163 2653 3180
rect 2516 3163 2533 3180
rect 2476 3163 2493 3180
rect 2396 3163 2413 3180
rect 2396 3163 2413 3180
rect 2436 3163 2453 3180
rect 2396 3163 2413 3180
rect 2436 3163 2453 3180
rect 2196 3163 2213 3180
rect 2396 3163 2413 3180
rect 2516 3163 2533 3180
rect 2436 3163 2453 3180
rect 2356 3163 2373 3180
rect 2236 3163 2253 3180
rect 2556 3163 2573 3180
rect 2476 3163 2493 3180
rect 2356 3163 2373 3180
rect 2316 3163 2333 3180
rect 2516 3163 2533 3180
rect 2156 3163 2173 3180
rect 2276 3163 2293 3180
rect 2356 3163 2373 3180
rect 2476 3163 2493 3180
rect 2236 3163 2253 3180
rect 2156 3163 2173 3180
rect 2476 3163 2493 3180
rect 2556 3163 2573 3180
rect 2636 3163 2653 3180
rect 2156 3163 2173 3180
rect 2316 3163 2333 3180
rect 2316 3163 2333 3180
rect 2356 3163 2373 3180
rect 2276 3163 2293 3180
rect 2556 3163 2573 3180
rect 2196 3163 2213 3180
rect 2236 3163 2253 3180
rect 2196 3163 2213 3180
rect 1676 3163 1693 3180
rect 1876 3163 1893 3180
rect 1796 3163 1813 3180
rect 2076 3163 2093 3180
rect 1636 3163 1653 3180
rect 1676 3163 1693 3180
rect 1916 3163 1933 3180
rect 1876 3163 1893 3180
rect 1956 3163 1973 3180
rect 1996 3163 2013 3180
rect 1756 3163 1773 3180
rect 1836 3163 1853 3180
rect 1636 3163 1653 3180
rect 1876 3163 1893 3180
rect 2076 3163 2093 3180
rect 1716 3163 1733 3180
rect 1836 3163 1853 3180
rect 1996 3163 2013 3180
rect 1876 3163 1893 3180
rect 1596 3163 1613 3180
rect 1596 3163 1613 3180
rect 1956 3163 1973 3180
rect 1796 3163 1813 3180
rect 2076 3163 2093 3180
rect 1636 3163 1653 3180
rect 1716 3163 1733 3180
rect 1596 3163 1613 3180
rect 1636 3163 1653 3180
rect 1916 3163 1933 3180
rect 2036 3163 2053 3180
rect 1756 3163 1773 3180
rect 2076 3163 2093 3180
rect 2036 3163 2053 3180
rect 1956 3163 1973 3180
rect 1996 3163 2013 3180
rect 1596 3163 1613 3180
rect 1756 3163 1773 3180
rect 1676 3163 1693 3180
rect 1836 3163 1853 3180
rect 1796 3163 1813 3180
rect 1916 3163 1933 3180
rect 2036 3163 2053 3180
rect 1716 3163 1733 3180
rect 1836 3163 1853 3180
rect 1676 3163 1693 3180
rect 1956 3163 1973 3180
rect 1996 3163 2013 3180
rect 1796 3163 1813 3180
rect 2036 3163 2053 3180
rect 1916 3163 1933 3180
rect 1716 3163 1733 3180
rect 1756 3163 1773 3180
rect 1036 3163 1053 3180
rect 1036 3163 1053 3180
rect 1036 3163 1053 3180
rect 1036 3163 1053 3180
rect 1276 3163 1293 3180
rect 1476 3163 1493 3180
rect 1436 3163 1453 3180
rect 1476 3163 1493 3180
rect 1076 3163 1093 3180
rect 1116 3163 1133 3180
rect 1076 3163 1093 3180
rect 1156 3163 1173 3180
rect 1516 3163 1533 3180
rect 1156 3163 1173 3180
rect 1396 3163 1413 3180
rect 1556 3163 1573 3180
rect 1436 3163 1453 3180
rect 1276 3163 1293 3180
rect 1316 3163 1333 3180
rect 1196 3163 1213 3180
rect 1316 3163 1333 3180
rect 1356 3163 1373 3180
rect 1196 3163 1213 3180
rect 1236 3163 1253 3180
rect 1516 3163 1533 3180
rect 1236 3163 1253 3180
rect 1396 3163 1413 3180
rect 1556 3163 1573 3180
rect 1276 3163 1293 3180
rect 1116 3163 1133 3180
rect 1476 3163 1493 3180
rect 1516 3163 1533 3180
rect 1076 3163 1093 3180
rect 1396 3163 1413 3180
rect 1316 3163 1333 3180
rect 1276 3163 1293 3180
rect 1436 3163 1453 3180
rect 1556 3163 1573 3180
rect 1156 3163 1173 3180
rect 1236 3163 1253 3180
rect 1196 3163 1213 3180
rect 1316 3163 1333 3180
rect 1356 3163 1373 3180
rect 1356 3163 1373 3180
rect 1396 3163 1413 3180
rect 1356 3163 1373 3180
rect 1116 3163 1133 3180
rect 1196 3163 1213 3180
rect 1476 3163 1493 3180
rect 1116 3163 1133 3180
rect 1436 3163 1453 3180
rect 1556 3163 1573 3180
rect 1516 3163 1533 3180
rect 1076 3163 1093 3180
rect 1236 3163 1253 3180
rect 1156 3163 1173 3180
rect 516 3163 533 3180
rect 836 3163 853 3180
rect 556 3163 573 3180
rect 836 3163 853 3180
rect 676 3163 693 3180
rect 596 3163 613 3180
rect 836 3163 853 3180
rect 716 3163 733 3180
rect 596 3163 613 3180
rect 556 3163 573 3180
rect 516 3163 533 3180
rect 916 3163 933 3180
rect 716 3163 733 3180
rect 916 3163 933 3180
rect 756 3163 773 3180
rect 756 3163 773 3180
rect 676 3163 693 3180
rect 516 3163 533 3180
rect 796 3163 813 3180
rect 756 3163 773 3180
rect 996 3163 1013 3180
rect 676 3163 693 3180
rect 636 3163 653 3180
rect 796 3163 813 3180
rect 876 3163 893 3180
rect 916 3163 933 3180
rect 876 3163 893 3180
rect 636 3163 653 3180
rect 756 3163 773 3180
rect 796 3163 813 3180
rect 716 3163 733 3180
rect 836 3163 853 3180
rect 996 3163 1013 3180
rect 716 3163 733 3180
rect 596 3163 613 3180
rect 676 3163 693 3180
rect 556 3163 573 3180
rect 516 3163 533 3180
rect 796 3163 813 3180
rect 956 3163 973 3180
rect 996 3163 1013 3180
rect 636 3163 653 3180
rect 916 3163 933 3180
rect 956 3163 973 3180
rect 996 3163 1013 3180
rect 596 3163 613 3180
rect 956 3163 973 3180
rect 876 3163 893 3180
rect 636 3163 653 3180
rect 876 3163 893 3180
rect 956 3163 973 3180
rect 556 3163 573 3180
rect 276 3163 293 3180
rect 476 3163 493 3180
rect 356 3163 373 3180
rect 396 3163 413 3180
rect 276 3163 293 3180
rect 356 3163 373 3180
rect 156 3163 173 3180
rect 236 3163 253 3180
rect 236 3163 253 3180
rect 276 3163 293 3180
rect 156 3163 173 3180
rect 116 3163 133 3180
rect 236 3163 253 3180
rect 396 3163 413 3180
rect 316 3163 333 3180
rect 476 3163 493 3180
rect 116 3163 133 3180
rect 436 3163 453 3180
rect 436 3163 453 3180
rect 236 3163 253 3180
rect 276 3163 293 3180
rect 156 3163 173 3180
rect 356 3163 373 3180
rect 396 3163 413 3180
rect 476 3163 493 3180
rect 436 3163 453 3180
rect 316 3163 333 3180
rect 116 3163 133 3180
rect 476 3163 493 3180
rect 396 3163 413 3180
rect 356 3163 373 3180
rect 156 3163 173 3180
rect 196 3163 213 3180
rect 196 3163 213 3180
rect 196 3163 213 3180
rect 196 3163 213 3180
rect 316 3163 333 3180
rect 436 3163 453 3180
rect 316 3163 333 3180
rect 116 3163 133 3180
rect 2481 2394 2498 2411
rect 1161 2394 1178 2411
rect 1201 2394 1218 2411
rect 841 2394 858 2411
rect 1841 2394 1858 2411
rect 1481 2394 1498 2411
rect 1001 2394 1018 2411
rect 1001 2394 1018 2411
rect 1201 2394 1218 2411
rect 1361 2394 1378 2411
rect 1801 2394 1818 2411
rect 1121 2394 1138 2411
rect 1321 2394 1338 2411
rect 1721 2394 1738 2411
rect 1601 2394 1618 2411
rect 1241 2394 1258 2411
rect 2441 2394 2458 2411
rect 2001 2394 2018 2411
rect 2241 2394 2258 2411
rect 2201 2394 2218 2411
rect 2361 2394 2378 2411
rect 2001 2394 2018 2411
rect 2121 2394 2138 2411
rect 1921 2394 1938 2411
rect 1961 2394 1978 2411
rect 2161 2394 2178 2411
rect 2041 2394 2058 2411
rect 2401 2394 2418 2411
rect 2161 2394 2178 2411
rect 1921 2394 1938 2411
rect 2201 2394 2218 2411
rect 2281 2394 2298 2411
rect 2121 2394 2138 2411
rect 2321 2394 2338 2411
rect 2041 2394 2058 2411
rect 2081 2394 2098 2411
rect 2441 2394 2458 2411
rect 2361 2394 2378 2411
rect 2081 2394 2098 2411
rect 2281 2394 2298 2411
rect 1961 2394 1978 2411
rect 2401 2394 2418 2411
rect 2321 2394 2338 2411
rect 2241 2394 2258 2411
rect 961 2394 978 2411
rect 1681 2394 1698 2411
rect 881 2394 898 2411
rect 1881 2394 1898 2411
rect 1521 2394 1538 2411
rect 1041 2394 1058 2411
rect 1441 2394 1458 2411
rect 1121 2394 1138 2411
rect 1401 2394 1418 2411
rect 1681 2394 1698 2411
rect 1361 2394 1378 2411
rect 1081 2394 1098 2411
rect 841 2394 858 2411
rect 1081 2394 1098 2411
rect 1481 2394 1498 2411
rect 1521 2394 1538 2411
rect 1801 2394 1818 2411
rect 1881 2394 1898 2411
rect 1321 2394 1338 2411
rect 1721 2394 1738 2411
rect 921 2394 938 2411
rect 1441 2394 1458 2411
rect 1841 2394 1858 2411
rect 1761 2394 1778 2411
rect 1281 2394 1298 2411
rect 1641 2394 1658 2411
rect 1161 2394 1178 2411
rect 1561 2394 1578 2411
rect 1241 2394 1258 2411
rect 1601 2394 1618 2411
rect 1761 2394 1778 2411
rect 1401 2394 1418 2411
rect 921 2394 938 2411
rect 961 2394 978 2411
rect 1041 2394 1058 2411
rect 1561 2394 1578 2411
rect 881 2394 898 2411
rect 1281 2394 1298 2411
rect 1641 2394 1658 2411
rect 3681 2394 3698 2411
rect 3681 2394 3698 2411
rect 2921 2394 2938 2411
rect 2801 2394 2818 2411
rect 2761 2394 2778 2411
rect 2521 2394 2538 2411
rect 2601 2394 2618 2411
rect 2561 2394 2578 2411
rect 2641 2394 2658 2411
rect 2881 2394 2898 2411
rect 2961 2394 2978 2411
rect 2681 2394 2698 2411
rect 2601 2394 2618 2411
rect 2961 2394 2978 2411
rect 2681 2394 2698 2411
rect 2921 2394 2938 2411
rect 2521 2394 2538 2411
rect 2841 2394 2858 2411
rect 3561 2394 3578 2411
rect 3041 2394 3058 2411
rect 3121 2394 3138 2411
rect 3361 2394 3378 2411
rect 3081 2394 3098 2411
rect 3241 2394 3258 2411
rect 3561 2394 3578 2411
rect 3441 2394 3458 2411
rect 3481 2394 3498 2411
rect 3001 2394 3018 2411
rect 3641 2394 3658 2411
rect 3481 2394 3498 2411
rect 3401 2394 3418 2411
rect 3161 2394 3178 2411
rect 3321 2394 3338 2411
rect 3521 2394 3538 2411
rect 3081 2394 3098 2411
rect 3641 2394 3658 2411
rect 3521 2394 3538 2411
rect 3601 2394 3618 2411
rect 3201 2394 3218 2411
rect 3441 2394 3458 2411
rect 3001 2394 3018 2411
rect 3121 2394 3138 2411
rect 3601 2394 3618 2411
rect 3281 2394 3298 2411
rect 2641 2394 2658 2411
rect 3201 2394 3218 2411
rect 3401 2394 3418 2411
rect 3281 2394 3298 2411
rect 3041 2394 3058 2411
rect 2801 2394 2818 2411
rect 3241 2394 3258 2411
rect 3321 2394 3338 2411
rect 3361 2394 3378 2411
rect 3161 2394 3178 2411
rect 2721 2394 2738 2411
rect 2761 2394 2778 2411
rect 2561 2394 2578 2411
rect 2881 2394 2898 2411
rect 2841 2394 2858 2411
rect 2721 2394 2738 2411
rect 4521 2394 4538 2411
rect 4041 2394 4058 2411
rect 4601 2394 4618 2411
rect 4201 2394 4218 2411
rect 4481 2394 4498 2411
rect 3801 2394 3818 2411
rect 4601 2394 4618 2411
rect 4281 2394 4298 2411
rect 4721 2394 4738 2411
rect 4401 2394 4418 2411
rect 4081 2394 4098 2411
rect 4801 2394 4818 2411
rect 4161 2394 4178 2411
rect 3961 2394 3978 2411
rect 4241 2394 4258 2411
rect 4321 2394 4338 2411
rect 3921 2394 3938 2411
rect 4161 2394 4178 2411
rect 4121 2394 4138 2411
rect 3881 2394 3898 2411
rect 4201 2394 4218 2411
rect 4281 2394 4298 2411
rect 4361 2394 4378 2411
rect 4401 2394 4418 2411
rect 3761 2394 3778 2411
rect 3921 2394 3938 2411
rect 4561 2394 4578 2411
rect 4841 2394 4858 2411
rect 3761 2394 3778 2411
rect 4721 2394 4738 2411
rect 4481 2394 4498 2411
rect 3841 2394 3858 2411
rect 3721 2394 3738 2411
rect 4841 2394 4858 2411
rect 3841 2394 3858 2411
rect 3881 2394 3898 2411
rect 3721 2394 3738 2411
rect 4001 2394 4018 2411
rect 4041 2394 4058 2411
rect 4681 2394 4698 2411
rect 4641 2394 4658 2411
rect 3801 2394 3818 2411
rect 4521 2394 4538 2411
rect 4761 2394 4778 2411
rect 4361 2394 4378 2411
rect 4441 2394 4458 2411
rect 4641 2394 4658 2411
rect 4081 2394 4098 2411
rect 4801 2394 4818 2411
rect 4441 2394 4458 2411
rect 4681 2394 4698 2411
rect 4321 2394 4338 2411
rect 4121 2394 4138 2411
rect 4761 2394 4778 2411
rect 4241 2394 4258 2411
rect 4561 2394 4578 2411
rect 3961 2394 3978 2411
rect 4001 2394 4018 2411
rect 7276 3163 7293 3180
rect 7316 3163 7333 3180
rect 7276 3163 7293 3180
rect 7316 3163 7333 3180
rect 7356 3163 7373 3180
rect 7116 3163 7133 3180
rect 7236 3163 7253 3180
rect 7036 3163 7053 3180
rect 6996 3163 7013 3180
rect 7236 3163 7253 3180
rect 7476 3163 7493 3180
rect 7196 3163 7213 3180
rect 7196 3163 7213 3180
rect 7076 3163 7093 3180
rect 7116 3163 7133 3180
rect 6996 3163 7013 3180
rect 7076 3163 7093 3180
rect 7356 3163 7373 3180
rect 7276 3163 7293 3180
rect 7356 3163 7373 3180
rect 7156 3163 7173 3180
rect 7236 3163 7253 3180
rect 7476 3163 7493 3180
rect 7036 3163 7053 3180
rect 7036 3163 7053 3180
rect 6436 3163 6453 3180
rect 6436 3163 6453 3180
rect 6436 3163 6453 3180
rect 6436 3163 6453 3180
rect 6476 3163 6493 3180
rect 6516 3163 6533 3180
rect 6516 3163 6533 3180
rect 6636 3163 6653 3180
rect 6476 3163 6493 3180
rect 6596 3163 6613 3180
rect 6556 3163 6573 3180
rect 6636 3163 6653 3180
rect 6556 3163 6573 3180
rect 6596 3163 6613 3180
rect 6476 3163 6493 3180
rect 6636 3163 6653 3180
rect 6596 3163 6613 3180
rect 6556 3163 6573 3180
rect 6516 3163 6533 3180
rect 6476 3163 6493 3180
rect 6676 3163 6693 3180
rect 6676 3163 6693 3180
rect 6676 3163 6693 3180
rect 6676 3163 6693 3180
rect 6796 3163 6813 3180
rect 6756 3163 6773 3180
rect 6716 3163 6733 3180
rect 6956 3163 6973 3180
rect 6916 3163 6933 3180
rect 6876 3163 6893 3180
rect 6836 3163 6853 3180
rect 6796 3163 6813 3180
rect 6756 3163 6773 3180
rect 6716 3163 6733 3180
rect 6956 3163 6973 3180
rect 6916 3163 6933 3180
rect 6876 3163 6893 3180
rect 6836 3163 6853 3180
rect 6716 3163 6733 3180
rect 6956 3163 6973 3180
rect 6916 3163 6933 3180
rect 6876 3163 6893 3180
rect 6836 3163 6853 3180
rect 6796 3163 6813 3180
rect 6756 3163 6773 3180
rect 6716 3163 6733 3180
rect 6916 3163 6933 3180
rect 6956 3163 6973 3180
rect 6836 3163 6853 3180
rect 6636 3163 6653 3180
rect 6796 3163 6813 3180
rect 6756 3163 6773 3180
rect 6596 3163 6613 3180
rect 6556 3163 6573 3180
rect 6876 3163 6893 3180
rect 6516 3163 6533 3180
rect 6236 3163 6253 3180
rect 6236 3163 6253 3180
rect 5956 3163 5973 3180
rect 5916 3163 5933 3180
rect 5956 3163 5973 3180
rect 6036 3163 6053 3180
rect 6156 3163 6173 3180
rect 6356 3163 6373 3180
rect 6396 3163 6413 3180
rect 6276 3163 6293 3180
rect 6156 3163 6173 3180
rect 5916 3163 5933 3180
rect 6036 3163 6053 3180
rect 6156 3163 6173 3180
rect 5996 3163 6013 3180
rect 6316 3163 6333 3180
rect 6196 3163 6213 3180
rect 6396 3163 6413 3180
rect 6396 3163 6413 3180
rect 6356 3163 6373 3180
rect 6116 3163 6133 3180
rect 6316 3163 6333 3180
rect 6356 3163 6373 3180
rect 6356 3163 6373 3180
rect 6076 3163 6093 3180
rect 6036 3163 6053 3180
rect 6076 3163 6093 3180
rect 6196 3163 6213 3180
rect 5956 3163 5973 3180
rect 5996 3163 6013 3180
rect 6316 3163 6333 3180
rect 6076 3163 6093 3180
rect 5996 3163 6013 3180
rect 6076 3163 6093 3180
rect 5956 3163 5973 3180
rect 6196 3163 6213 3180
rect 6276 3163 6293 3180
rect 5916 3163 5933 3180
rect 6316 3163 6333 3180
rect 6116 3163 6133 3180
rect 6236 3163 6253 3180
rect 6156 3163 6173 3180
rect 5996 3163 6013 3180
rect 5916 3163 5933 3180
rect 6236 3163 6253 3180
rect 6116 3163 6133 3180
rect 6036 3163 6053 3180
rect 6276 3163 6293 3180
rect 6276 3163 6293 3180
rect 6396 3163 6413 3180
rect 6196 3163 6213 3180
rect 6116 3163 6133 3180
rect 5356 3163 5373 3180
rect 5356 3163 5373 3180
rect 5356 3163 5373 3180
rect 5356 3163 5373 3180
rect 5396 3163 5413 3180
rect 5756 3163 5773 3180
rect 5796 3163 5813 3180
rect 5436 3163 5453 3180
rect 5796 3163 5813 3180
rect 5476 3163 5493 3180
rect 5756 3163 5773 3180
rect 5516 3163 5533 3180
rect 5636 3163 5653 3180
rect 5436 3163 5453 3180
rect 5756 3163 5773 3180
rect 5596 3163 5613 3180
rect 5716 3163 5733 3180
rect 5556 3163 5573 3180
rect 5876 3163 5893 3180
rect 5396 3163 5413 3180
rect 5476 3163 5493 3180
rect 5436 3163 5453 3180
rect 5556 3163 5573 3180
rect 5716 3163 5733 3180
rect 5796 3163 5813 3180
rect 5876 3163 5893 3180
rect 5396 3163 5413 3180
rect 5716 3163 5733 3180
rect 5836 3163 5853 3180
rect 5676 3163 5693 3180
rect 5796 3163 5813 3180
rect 5676 3163 5693 3180
rect 5676 3163 5693 3180
rect 5716 3163 5733 3180
rect 5636 3163 5653 3180
rect 5556 3163 5573 3180
rect 5876 3163 5893 3180
rect 5596 3163 5613 3180
rect 5516 3163 5533 3180
rect 5396 3163 5413 3180
rect 5516 3163 5533 3180
rect 5756 3163 5773 3180
rect 5636 3163 5653 3180
rect 5676 3163 5693 3180
rect 5596 3163 5613 3180
rect 5596 3163 5613 3180
rect 5836 3163 5853 3180
rect 5836 3163 5853 3180
rect 5476 3163 5493 3180
rect 5556 3163 5573 3180
rect 5636 3163 5653 3180
rect 5836 3163 5853 3180
rect 5476 3163 5493 3180
rect 5876 3163 5893 3180
rect 5436 3163 5453 3180
rect 5516 3163 5533 3180
rect 5076 3163 5093 3180
rect 5316 3163 5333 3180
rect 5236 3163 5253 3180
rect 5076 3163 5093 3180
rect 4956 3163 4973 3180
rect 4956 3163 4973 3180
rect 7241 2394 7258 2411
rect 5116 3163 5133 3180
rect 7241 2394 7258 2411
rect 5036 3163 5053 3180
rect 5196 3163 5213 3180
rect 5156 3163 5173 3180
rect 5156 3163 5173 3180
rect 4916 3163 4933 3180
rect 5196 3163 5213 3180
rect 4876 3163 4893 3180
rect 4996 3163 5013 3180
rect 5196 3163 5213 3180
rect 5316 3163 5333 3180
rect 5196 3163 5213 3180
rect 4916 3163 4933 3180
rect 5116 3163 5133 3180
rect 5036 3163 5053 3180
rect 4876 3163 4893 3180
rect 5156 3163 5173 3180
rect 4916 3163 4933 3180
rect 5316 3163 5333 3180
rect 4996 3163 5013 3180
rect 4876 3163 4893 3180
rect 4956 3163 4973 3180
rect 5316 3163 5333 3180
rect 5036 3163 5053 3180
rect 5076 3163 5093 3180
rect 5276 3163 5293 3180
rect 5276 3163 5293 3180
rect 5236 3163 5253 3180
rect 5156 3163 5173 3180
rect 4876 3163 4893 3180
rect 5236 3163 5253 3180
rect 5276 3163 5293 3180
rect 5076 3163 5093 3180
rect 5116 3163 5133 3180
rect 5036 3163 5053 3180
rect 4916 3163 4933 3180
rect 4956 3163 4973 3180
rect 4996 3163 5013 3180
rect 5116 3163 5133 3180
rect 4996 3163 5013 3180
rect 5236 3163 5253 3180
rect 5276 3163 5293 3180
rect 9236 3163 9253 3180
rect 9236 3163 9253 3180
rect 9396 3163 9413 3180
rect 9436 3163 9453 3180
rect 9156 3163 9173 3180
rect 9596 3163 9613 3180
rect 9316 3163 9333 3180
rect 9476 3163 9493 3180
rect 9516 3163 9533 3180
rect 9356 3163 9373 3180
rect 9276 3163 9293 3180
rect 9276 3163 9293 3180
rect 9396 3163 9413 3180
rect 9476 3163 9493 3180
rect 9316 3163 9333 3180
rect 9436 3163 9453 3180
rect 9596 3163 9613 3180
rect 9476 3163 9493 3180
rect 9356 3163 9373 3180
rect 9556 3163 9573 3180
rect 9156 3163 9173 3180
rect 9156 3163 9173 3180
rect 9316 3163 9333 3180
rect 9276 3163 9293 3180
rect 9556 3163 9573 3180
rect 9596 3163 9613 3180
rect 9356 3163 9373 3180
rect 9436 3163 9453 3180
rect 9356 3163 9373 3180
rect 9196 3163 9213 3180
rect 9276 3163 9293 3180
rect 9396 3163 9413 3180
rect 9156 3163 9173 3180
rect 9436 3163 9453 3180
rect 9476 3163 9493 3180
rect 9396 3163 9413 3180
rect 9516 3163 9533 3180
rect 9236 3163 9253 3180
rect 9236 3163 9253 3180
rect 9556 3163 9573 3180
rect 9316 3163 9333 3180
rect 9596 3163 9613 3180
rect 9516 3163 9533 3180
rect 9196 3163 9213 3180
rect 9196 3163 9213 3180
rect 9196 3163 9213 3180
rect 9516 3163 9533 3180
rect 9556 3163 9573 3180
rect 8596 3163 8613 3180
rect 8596 3163 8613 3180
rect 8596 3163 8613 3180
rect 8596 3163 8613 3180
rect 8956 3163 8973 3180
rect 8956 3163 8973 3180
rect 8876 3163 8893 3180
rect 8716 3163 8733 3180
rect 8756 3163 8773 3180
rect 8916 3163 8933 3180
rect 8796 3163 8813 3180
rect 8956 3163 8973 3180
rect 8876 3163 8893 3180
rect 9116 3163 9133 3180
rect 8756 3163 8773 3180
rect 9076 3163 9093 3180
rect 9036 3163 9053 3180
rect 8956 3163 8973 3180
rect 8676 3163 8693 3180
rect 9076 3163 9093 3180
rect 8756 3163 8773 3180
rect 8796 3163 8813 3180
rect 8836 3163 8853 3180
rect 8636 3163 8653 3180
rect 8716 3163 8733 3180
rect 8716 3163 8733 3180
rect 8876 3163 8893 3180
rect 8836 3163 8853 3180
rect 8636 3163 8653 3180
rect 8916 3163 8933 3180
rect 9036 3163 9053 3180
rect 9036 3163 9053 3180
rect 8676 3163 8693 3180
rect 9116 3163 9133 3180
rect 8836 3163 8853 3180
rect 8996 3163 9013 3180
rect 8796 3163 8813 3180
rect 9036 3163 9053 3180
rect 9116 3163 9133 3180
rect 8636 3163 8653 3180
rect 8716 3163 8733 3180
rect 8916 3163 8933 3180
rect 8836 3163 8853 3180
rect 8996 3163 9013 3180
rect 9116 3163 9133 3180
rect 8676 3163 8693 3180
rect 9076 3163 9093 3180
rect 8996 3163 9013 3180
rect 8676 3163 8693 3180
rect 8916 3163 8933 3180
rect 8756 3163 8773 3180
rect 8796 3163 8813 3180
rect 8636 3163 8653 3180
rect 8996 3163 9013 3180
rect 9076 3163 9093 3180
rect 8876 3163 8893 3180
rect 8316 3163 8333 3180
rect 8196 3163 8213 3180
rect 8116 3163 8133 3180
rect 8196 3163 8213 3180
rect 8076 3163 8093 3180
rect 8396 3163 8413 3180
rect 8156 3163 8173 3180
rect 8276 3163 8293 3180
rect 8196 3163 8213 3180
rect 8556 3163 8573 3180
rect 8316 3163 8333 3180
rect 8316 3163 8333 3180
rect 8276 3163 8293 3180
rect 8516 3163 8533 3180
rect 8356 3163 8373 3180
rect 8476 3163 8493 3180
rect 8236 3163 8253 3180
rect 8396 3163 8413 3180
rect 8436 3163 8453 3180
rect 8076 3163 8093 3180
rect 8156 3163 8173 3180
rect 8116 3163 8133 3180
rect 8116 3163 8133 3180
rect 8076 3163 8093 3180
rect 8396 3163 8413 3180
rect 8236 3163 8253 3180
rect 8516 3163 8533 3180
rect 8556 3163 8573 3180
rect 8556 3163 8573 3180
rect 8276 3163 8293 3180
rect 8276 3163 8293 3180
rect 8476 3163 8493 3180
rect 8556 3163 8573 3180
rect 8156 3163 8173 3180
rect 8396 3163 8413 3180
rect 8316 3163 8333 3180
rect 8116 3163 8133 3180
rect 8236 3163 8253 3180
rect 8236 3163 8253 3180
rect 8516 3163 8533 3180
rect 8476 3163 8493 3180
rect 8436 3163 8453 3180
rect 8476 3163 8493 3180
rect 8156 3163 8173 3180
rect 8356 3163 8373 3180
rect 8436 3163 8453 3180
rect 8196 3163 8213 3180
rect 8436 3163 8453 3180
rect 8516 3163 8533 3180
rect 8356 3163 8373 3180
rect 8076 3163 8093 3180
rect 8356 3163 8373 3180
rect 7516 3163 7533 3180
rect 7516 3163 7533 3180
rect 7516 3163 7533 3180
rect 7516 3163 7533 3180
rect 7636 3163 7653 3180
rect 7916 3163 7933 3180
rect 7676 3163 7693 3180
rect 7716 3163 7733 3180
rect 7956 3163 7973 3180
rect 7596 3163 7613 3180
rect 7876 3163 7893 3180
rect 7596 3163 7613 3180
rect 7876 3163 7893 3180
rect 7756 3163 7773 3180
rect 8036 3163 8053 3180
rect 8036 3163 8053 3180
rect 7916 3163 7933 3180
rect 7956 3163 7973 3180
rect 7956 3163 7973 3180
rect 8036 3163 8053 3180
rect 7836 3163 7853 3180
rect 7716 3163 7733 3180
rect 7996 3163 8013 3180
rect 7836 3163 7853 3180
rect 7716 3163 7733 3180
rect 7756 3163 7773 3180
rect 7876 3163 7893 3180
rect 7596 3163 7613 3180
rect 7556 3163 7573 3180
rect 7716 3163 7733 3180
rect 7796 3163 7813 3180
rect 7556 3163 7573 3180
rect 7676 3163 7693 3180
rect 7556 3163 7573 3180
rect 7796 3163 7813 3180
rect 7796 3163 7813 3180
rect 7876 3163 7893 3180
rect 7996 3163 8013 3180
rect 7836 3163 7853 3180
rect 7756 3163 7773 3180
rect 7916 3163 7933 3180
rect 8036 3163 8053 3180
rect 7956 3163 7973 3180
rect 7676 3163 7693 3180
rect 7636 3163 7653 3180
rect 7676 3163 7693 3180
rect 7796 3163 7813 3180
rect 7996 3163 8013 3180
rect 7836 3163 7853 3180
rect 7636 3163 7653 3180
rect 7556 3163 7573 3180
rect 7996 3163 8013 3180
rect 7916 3163 7933 3180
rect 7596 3163 7613 3180
rect 7636 3163 7653 3180
rect 7756 3163 7773 3180
rect 7396 3163 7413 3180
rect 7156 3163 7173 3180
rect 6996 3163 7013 3180
rect 7076 3163 7093 3180
rect 7356 3163 7373 3180
rect 7196 3163 7213 3180
rect 7236 3163 7253 3180
rect 7076 3163 7093 3180
rect 7396 3163 7413 3180
rect 7436 3163 7453 3180
rect 7276 3163 7293 3180
rect 7316 3163 7333 3180
rect 7316 3163 7333 3180
rect 7116 3163 7133 3180
rect 7116 3163 7133 3180
rect 7156 3163 7173 3180
rect 7396 3163 7413 3180
rect 7156 3163 7173 3180
rect 7436 3163 7453 3180
rect 7476 3163 7493 3180
rect 6996 3163 7013 3180
rect 7036 3163 7053 3180
rect 7396 3163 7413 3180
rect 7436 3163 7453 3180
rect 7196 3163 7213 3180
rect 7476 3163 7493 3180
rect 9276 3163 9293 3180
rect 9556 3163 9573 3180
rect 9356 3163 9373 3180
rect 9476 3163 9493 3180
rect 9316 3163 9333 3180
rect 9596 3163 9613 3180
rect 9196 3163 9213 3180
rect 8996 3163 9013 3180
rect 9516 3163 9533 3180
rect 9516 3163 9533 3180
rect 8996 3163 9013 3180
rect 9196 3163 9213 3180
rect 9076 3163 9093 3180
rect 9276 3163 9293 3180
rect 9236 3163 9253 3180
rect 9196 3163 9213 3180
rect 9556 3163 9573 3180
rect 9156 3163 9173 3180
rect 9036 3163 9053 3180
rect 9196 3163 9213 3180
rect 9396 3163 9413 3180
rect 9356 3163 9373 3180
rect 9396 3163 9413 3180
rect 9116 3163 9133 3180
rect 9156 3163 9173 3180
rect 9556 3163 9573 3180
rect 9516 3163 9533 3180
rect 9276 3163 9293 3180
rect 9596 3163 9613 3180
rect 9556 3163 9573 3180
rect 9436 3163 9453 3180
rect 9436 3163 9453 3180
rect 9276 3163 9293 3180
rect 9036 3163 9053 3180
rect 9156 3163 9173 3180
rect 9476 3163 9493 3180
rect 9316 3163 9333 3180
rect 9396 3163 9413 3180
rect 9156 3163 9173 3180
rect 8956 3163 8973 3180
rect 9036 3163 9053 3180
rect 8956 3163 8973 3180
rect 9476 3163 9493 3180
rect 9356 3163 9373 3180
rect 9396 3163 9413 3180
rect 8996 3163 9013 3180
rect 9596 3163 9613 3180
rect 9316 3163 9333 3180
rect 9116 3163 9133 3180
rect 8956 3163 8973 3180
rect 9516 3163 9533 3180
rect 9436 3163 9453 3180
rect 9116 3163 9133 3180
rect 9316 3163 9333 3180
rect 9436 3163 9453 3180
rect 9236 3163 9253 3180
rect 9596 3163 9613 3180
rect 9076 3163 9093 3180
rect 9076 3163 9093 3180
rect 9036 3163 9053 3180
rect 9236 3163 9253 3180
rect 9116 3163 9133 3180
rect 8956 3163 8973 3180
rect 9476 3163 9493 3180
rect 9236 3163 9253 3180
rect 8996 3163 9013 3180
rect 9076 3163 9093 3180
rect 9356 3163 9373 3180
rect 8796 3163 8813 3180
rect 8596 3163 8613 3180
rect 8476 3163 8493 3180
rect 8876 3163 8893 3180
rect 8316 3163 8333 3180
rect 8156 3163 8173 3180
rect 8596 3163 8613 3180
rect 8916 3163 8933 3180
rect 8316 3163 8333 3180
rect 8036 3163 8053 3180
rect 8156 3163 8173 3180
rect 8596 3163 8613 3180
rect 8836 3163 8853 3180
rect 8036 3163 8053 3180
rect 7996 3163 8013 3180
rect 8276 3163 8293 3180
rect 8356 3163 8373 3180
rect 8316 3163 8333 3180
rect 8396 3163 8413 3180
rect 8516 3163 8533 3180
rect 8436 3163 8453 3180
rect 8276 3163 8293 3180
rect 8836 3163 8853 3180
rect 8196 3163 8213 3180
rect 8356 3163 8373 3180
rect 8196 3163 8213 3180
rect 8036 3163 8053 3180
rect 8876 3163 8893 3180
rect 8796 3163 8813 3180
rect 8316 3163 8333 3180
rect 8476 3163 8493 3180
rect 8716 3163 8733 3180
rect 8436 3163 8453 3180
rect 8916 3163 8933 3180
rect 8836 3163 8853 3180
rect 8236 3163 8253 3180
rect 7996 3163 8013 3180
rect 8756 3163 8773 3180
rect 8516 3163 8533 3180
rect 8116 3163 8133 3180
rect 8396 3163 8413 3180
rect 8916 3163 8933 3180
rect 8116 3163 8133 3180
rect 8356 3163 8373 3180
rect 8876 3163 8893 3180
rect 8436 3163 8453 3180
rect 8796 3163 8813 3180
rect 8676 3163 8693 3180
rect 8636 3163 8653 3180
rect 8076 3163 8093 3180
rect 8916 3163 8933 3180
rect 8076 3163 8093 3180
rect 8196 3163 8213 3180
rect 8156 3163 8173 3180
rect 8636 3163 8653 3180
rect 8876 3163 8893 3180
rect 8556 3163 8573 3180
rect 8676 3163 8693 3180
rect 8116 3163 8133 3180
rect 8356 3163 8373 3180
rect 8236 3163 8253 3180
rect 8076 3163 8093 3180
rect 8116 3163 8133 3180
rect 8476 3163 8493 3180
rect 8756 3163 8773 3180
rect 8716 3163 8733 3180
rect 8796 3163 8813 3180
rect 8076 3163 8093 3180
rect 8236 3163 8253 3180
rect 8276 3163 8293 3180
rect 8396 3163 8413 3180
rect 8836 3163 8853 3180
rect 8396 3163 8413 3180
rect 8516 3163 8533 3180
rect 8636 3163 8653 3180
rect 7996 3163 8013 3180
rect 8156 3163 8173 3180
rect 8636 3163 8653 3180
rect 8236 3163 8253 3180
rect 8476 3163 8493 3180
rect 8556 3163 8573 3180
rect 8276 3163 8293 3180
rect 7996 3163 8013 3180
rect 8676 3163 8693 3180
rect 8676 3163 8693 3180
rect 8516 3163 8533 3180
rect 8716 3163 8733 3180
rect 8196 3163 8213 3180
rect 8436 3163 8453 3180
rect 8596 3163 8613 3180
rect 8716 3163 8733 3180
rect 8756 3163 8773 3180
rect 8756 3163 8773 3180
rect 8556 3163 8573 3180
rect 8556 3163 8573 3180
rect 8036 3163 8053 3180
rect 7436 3163 7453 3180
rect 4921 2394 4938 2411
rect 4881 2394 4898 2411
rect 4881 2394 4898 2411
rect 4961 2394 4978 2411
rect 5041 2394 5058 2411
rect 5121 2394 5138 2411
rect 5121 2394 5138 2411
rect 5081 2394 5098 2411
rect 4961 2394 4978 2411
rect 5081 2394 5098 2411
rect 5001 2394 5018 2411
rect 5841 2394 5858 2411
rect 5641 2394 5658 2411
rect 5401 2394 5418 2411
rect 5241 2394 5258 2411
rect 6001 2394 6018 2411
rect 5521 2394 5538 2411
rect 5681 2394 5698 2411
rect 5921 2394 5938 2411
rect 5881 2394 5898 2411
rect 5761 2394 5778 2411
rect 5561 2394 5578 2411
rect 5601 2394 5618 2411
rect 5801 2394 5818 2411
rect 5481 2394 5498 2411
rect 5401 2394 5418 2411
rect 5361 2394 5378 2411
rect 5521 2394 5538 2411
rect 5961 2394 5978 2411
rect 5321 2394 5338 2411
rect 5761 2394 5778 2411
rect 5321 2394 5338 2411
rect 5961 2394 5978 2411
rect 5721 2394 5738 2411
rect 5201 2394 5218 2411
rect 5561 2394 5578 2411
rect 5441 2394 5458 2411
rect 5841 2394 5858 2411
rect 5641 2394 5658 2411
rect 5161 2394 5178 2411
rect 5481 2394 5498 2411
rect 6041 2394 6058 2411
rect 5441 2394 5458 2411
rect 5241 2394 5258 2411
rect 5721 2394 5738 2411
rect 5281 2394 5298 2411
rect 6041 2394 6058 2411
rect 5281 2394 5298 2411
rect 6001 2394 6018 2411
rect 5601 2394 5618 2411
rect 5681 2394 5698 2411
rect 5361 2394 5378 2411
rect 5161 2394 5178 2411
rect 5921 2394 5938 2411
rect 5881 2394 5898 2411
rect 5801 2394 5818 2411
rect 5201 2394 5218 2411
rect 5041 2394 5058 2411
rect 5001 2394 5018 2411
rect 4921 2394 4938 2411
rect 6881 2394 6898 2411
rect 6761 2394 6778 2411
rect 6961 2394 6978 2411
rect 6681 2394 6698 2411
rect 6321 2394 6338 2411
rect 6281 2394 6298 2411
rect 7041 2394 7058 2411
rect 6241 2394 6258 2411
rect 6441 2394 6458 2411
rect 6121 2394 6138 2411
rect 6401 2394 6418 2411
rect 6401 2394 6418 2411
rect 6081 2394 6098 2411
rect 6481 2394 6498 2411
rect 6161 2394 6178 2411
rect 6161 2394 6178 2411
rect 7001 2394 7018 2411
rect 6081 2394 6098 2411
rect 7161 2394 7178 2411
rect 6841 2394 6858 2411
rect 6121 2394 6138 2411
rect 6481 2394 6498 2411
rect 6721 2394 6738 2411
rect 6641 2394 6658 2411
rect 6721 2394 6738 2411
rect 7121 2394 7138 2411
rect 6361 2394 6378 2411
rect 6201 2394 6218 2411
rect 6641 2394 6658 2411
rect 7201 2394 7218 2411
rect 7081 2394 7098 2411
rect 7161 2394 7178 2411
rect 6601 2394 6618 2411
rect 6881 2394 6898 2411
rect 6201 2394 6218 2411
rect 7121 2394 7138 2411
rect 6321 2394 6338 2411
rect 6281 2394 6298 2411
rect 6521 2394 6538 2411
rect 6241 2394 6258 2411
rect 6361 2394 6378 2411
rect 6561 2394 6578 2411
rect 6801 2394 6818 2411
rect 6441 2394 6458 2411
rect 7081 2394 7098 2411
rect 7041 2394 7058 2411
rect 6601 2394 6618 2411
rect 6801 2394 6818 2411
rect 6561 2394 6578 2411
rect 6841 2394 6858 2411
rect 7001 2394 7018 2411
rect 7201 2394 7218 2411
rect 6961 2394 6978 2411
rect 6921 2394 6938 2411
rect 6681 2394 6698 2411
rect 6921 2394 6938 2411
rect 6521 2394 6538 2411
rect 6761 2394 6778 2411
rect 8441 2394 8458 2411
rect 8441 2394 8458 2411
rect 7881 2394 7898 2411
rect 8081 2394 8098 2411
rect 7401 2394 7418 2411
rect 7681 2394 7698 2411
rect 7841 2394 7858 2411
rect 7641 2394 7658 2411
rect 8241 2394 8258 2411
rect 7761 2394 7778 2411
rect 7281 2394 7298 2411
rect 7441 2394 7458 2411
rect 7441 2394 7458 2411
rect 7281 2394 7298 2411
rect 8401 2394 8418 2411
rect 8401 2394 8418 2411
rect 7361 2394 7378 2411
rect 7601 2394 7618 2411
rect 8321 2394 8338 2411
rect 7321 2394 7338 2411
rect 8361 2394 8378 2411
rect 8041 2394 8058 2411
rect 7881 2394 7898 2411
rect 8281 2394 8298 2411
rect 8201 2394 8218 2411
rect 8001 2394 8018 2411
rect 8241 2394 8258 2411
rect 7921 2394 7938 2411
rect 7721 2394 7738 2411
rect 8281 2394 8298 2411
rect 7761 2394 7778 2411
rect 7681 2394 7698 2411
rect 7961 2394 7978 2411
rect 7801 2394 7818 2411
rect 7641 2394 7658 2411
rect 8201 2394 8218 2411
rect 7601 2394 7618 2411
rect 8161 2394 8178 2411
rect 7721 2394 7738 2411
rect 7401 2394 7418 2411
rect 8121 2394 8138 2411
rect 7561 2394 7578 2411
rect 7361 2394 7378 2411
rect 8121 2394 8138 2411
rect 7921 2394 7938 2411
rect 7321 2394 7338 2411
rect 7841 2394 7858 2411
rect 8081 2394 8098 2411
rect 7521 2394 7538 2411
rect 7561 2394 7578 2411
rect 8041 2394 8058 2411
rect 8161 2394 8178 2411
rect 7521 2394 7538 2411
rect 7801 2394 7818 2411
rect 8361 2394 8378 2411
rect 7481 2394 7498 2411
rect 7481 2394 7498 2411
rect 8001 2394 8018 2411
rect 8321 2394 8338 2411
rect 7961 2394 7978 2411
rect 9041 2394 9058 2411
rect 9601 2394 9618 2411
rect 9481 2394 9498 2411
rect 8641 2394 8658 2411
rect 9441 2394 9458 2411
rect 9401 2394 9418 2411
rect 8601 2394 8618 2411
rect 9361 2394 9378 2411
rect 9321 2394 9338 2411
rect 8881 2394 8898 2411
rect 8601 2394 8618 2411
rect 9001 2394 9018 2411
rect 9281 2394 9298 2411
rect 9241 2394 9258 2411
rect 8961 2394 8978 2411
rect 9201 2394 9218 2411
rect 9161 2394 9178 2411
rect 8921 2394 8938 2411
rect 9121 2394 9138 2411
rect 9081 2394 9098 2411
rect 8881 2394 8898 2411
rect 9041 2394 9058 2411
rect 8841 2394 8858 2411
rect 8561 2394 8578 2411
rect 8521 2394 8538 2411
rect 8801 2394 8818 2411
rect 9441 2394 9458 2411
rect 8521 2394 8538 2411
rect 8841 2394 8858 2411
rect 9401 2394 9418 2411
rect 8481 2394 8498 2411
rect 8481 2394 8498 2411
rect 9481 2394 9498 2411
rect 8561 2394 8578 2411
rect 9521 2394 9538 2411
rect 8761 2394 8778 2411
rect 9561 2394 9578 2411
rect 9001 2394 9018 2411
rect 8721 2394 8738 2411
rect 8921 2394 8938 2411
rect 8961 2394 8978 2411
rect 8681 2394 8698 2411
rect 8641 2394 8658 2411
rect 9561 2394 9578 2411
rect 9361 2394 9378 2411
rect 8801 2394 8818 2411
rect 9321 2394 9338 2411
rect 9281 2394 9298 2411
rect 8761 2394 8778 2411
rect 9601 2394 9618 2411
rect 9241 2394 9258 2411
rect 9201 2394 9218 2411
rect 8721 2394 8738 2411
rect 9161 2394 9178 2411
rect 9121 2394 9138 2411
rect 9521 2394 9538 2411
rect 8681 2394 8698 2411
rect 9081 2394 9098 2411
rect 15576 4652 15593 4669
rect 15576 4652 15593 4669
rect 15576 4652 15593 4669
rect 15576 4652 15593 4669
rect 16176 4652 16193 4669
rect 16176 4652 16193 4669
rect 16176 4652 16193 4669
rect 16176 4652 16193 4669
rect 16616 4652 16633 4669
rect 16616 4652 16633 4669
rect 16216 4652 16233 4669
rect 16576 4652 16593 4669
rect 16456 4652 16473 4669
rect 16536 4652 16553 4669
rect 16656 4652 16673 4669
rect 16496 4652 16513 4669
rect 16456 4652 16473 4669
rect 16456 4652 16473 4669
rect 16696 4652 16713 4669
rect 16416 4652 16433 4669
rect 16536 4652 16553 4669
rect 16496 4652 16513 4669
rect 16376 4652 16393 4669
rect 16456 4652 16473 4669
rect 16696 4652 16713 4669
rect 16416 4652 16433 4669
rect 16656 4652 16673 4669
rect 16576 4652 16593 4669
rect 16416 4652 16433 4669
rect 16376 4652 16393 4669
rect 16336 4652 16353 4669
rect 16536 4652 16553 4669
rect 16336 4652 16353 4669
rect 16296 4652 16313 4669
rect 16496 4652 16513 4669
rect 16736 4652 16753 4669
rect 16256 4652 16273 4669
rect 16696 4652 16713 4669
rect 16656 4652 16673 4669
rect 16616 4652 16633 4669
rect 16616 4652 16633 4669
rect 16216 4652 16233 4669
rect 16576 4652 16593 4669
rect 16296 4652 16313 4669
rect 16736 4652 16753 4669
rect 16256 4652 16273 4669
rect 16216 4652 16233 4669
rect 16376 4652 16393 4669
rect 16336 4652 16353 4669
rect 16256 4652 16273 4669
rect 16536 4652 16553 4669
rect 16216 4652 16233 4669
rect 16336 4652 16353 4669
rect 16296 4652 16313 4669
rect 16696 4652 16713 4669
rect 16416 4652 16433 4669
rect 16576 4652 16593 4669
rect 16256 4652 16273 4669
rect 16296 4652 16313 4669
rect 16736 4652 16753 4669
rect 16496 4652 16513 4669
rect 16376 4652 16393 4669
rect 16736 4652 16753 4669
rect 16656 4652 16673 4669
rect 16056 4652 16073 4669
rect 16016 4652 16033 4669
rect 15976 4652 15993 4669
rect 15936 4652 15953 4669
rect 16056 4652 16073 4669
rect 16096 4652 16113 4669
rect 16096 4652 16113 4669
rect 16136 4652 16153 4669
rect 16136 4652 16153 4669
rect 15696 4652 15713 4669
rect 15816 4652 15833 4669
rect 15896 4652 15913 4669
rect 15776 4652 15793 4669
rect 15736 4652 15753 4669
rect 15656 4652 15673 4669
rect 15696 4652 15713 4669
rect 15816 4652 15833 4669
rect 15656 4652 15673 4669
rect 15856 4652 15873 4669
rect 15856 4652 15873 4669
rect 15736 4652 15753 4669
rect 15896 4652 15913 4669
rect 15776 4652 15793 4669
rect 15616 4652 15633 4669
rect 15616 4652 15633 4669
rect 16016 4652 16033 4669
rect 16136 4652 16153 4669
rect 15696 4652 15713 4669
rect 15816 4652 15833 4669
rect 15896 4652 15913 4669
rect 15776 4652 15793 4669
rect 15736 4652 15753 4669
rect 15656 4652 15673 4669
rect 15696 4652 15713 4669
rect 15816 4652 15833 4669
rect 15656 4652 15673 4669
rect 15856 4652 15873 4669
rect 15856 4652 15873 4669
rect 15736 4652 15753 4669
rect 15896 4652 15913 4669
rect 15776 4652 15793 4669
rect 16016 4652 16033 4669
rect 15976 4652 15993 4669
rect 15616 4652 15633 4669
rect 15936 4652 15953 4669
rect 16056 4652 16073 4669
rect 16016 4652 16033 4669
rect 15976 4652 15993 4669
rect 15936 4652 15953 4669
rect 16056 4652 16073 4669
rect 15616 4652 15633 4669
rect 16096 4652 16113 4669
rect 16096 4652 16113 4669
rect 15976 4652 15993 4669
rect 16136 4652 16153 4669
rect 15936 4652 15953 4669
rect 14976 4652 14993 4669
rect 14976 4652 14993 4669
rect 14976 4652 14993 4669
rect 14976 4652 14993 4669
rect 15016 4652 15033 4669
rect 15016 4652 15033 4669
rect 15056 4652 15073 4669
rect 15136 4652 15153 4669
rect 15176 4652 15193 4669
rect 15416 4652 15433 4669
rect 15376 4652 15393 4669
rect 15416 4652 15433 4669
rect 15496 4652 15513 4669
rect 15136 4652 15153 4669
rect 15096 4652 15113 4669
rect 15296 4652 15313 4669
rect 15216 4652 15233 4669
rect 15256 4652 15273 4669
rect 15376 4652 15393 4669
rect 15096 4652 15113 4669
rect 15296 4652 15313 4669
rect 15096 4652 15113 4669
rect 15496 4652 15513 4669
rect 15216 4652 15233 4669
rect 15536 4652 15553 4669
rect 15496 4652 15513 4669
rect 15056 4652 15073 4669
rect 15056 4652 15073 4669
rect 15336 4652 15353 4669
rect 15496 4652 15513 4669
rect 15176 4652 15193 4669
rect 15536 4652 15553 4669
rect 15456 4652 15473 4669
rect 15456 4652 15473 4669
rect 15016 4652 15033 4669
rect 15016 4652 15033 4669
rect 15336 4652 15353 4669
rect 15136 4652 15153 4669
rect 15336 4652 15353 4669
rect 15176 4652 15193 4669
rect 15216 4652 15233 4669
rect 15416 4652 15433 4669
rect 15256 4652 15273 4669
rect 15416 4652 15433 4669
rect 15456 4652 15473 4669
rect 15216 4652 15233 4669
rect 15456 4652 15473 4669
rect 15136 4652 15153 4669
rect 15176 4652 15193 4669
rect 15256 4652 15273 4669
rect 15536 4652 15553 4669
rect 15376 4652 15393 4669
rect 15296 4652 15313 4669
rect 15096 4652 15113 4669
rect 15536 4652 15553 4669
rect 15256 4652 15273 4669
rect 15376 4652 15393 4669
rect 15296 4652 15313 4669
rect 15336 4652 15353 4669
rect 15056 4652 15073 4669
rect 14896 4652 14913 4669
rect 14896 4652 14913 4669
rect 14856 4652 14873 4669
rect 14656 4652 14673 4669
rect 14616 4652 14633 4669
rect 14576 4652 14593 4669
rect 14536 4652 14553 4669
rect 14496 4652 14513 4669
rect 14456 4652 14473 4669
rect 14416 4652 14433 4669
rect 14816 4652 14833 4669
rect 14776 4652 14793 4669
rect 14736 4652 14753 4669
rect 14696 4652 14713 4669
rect 14656 4652 14673 4669
rect 14616 4652 14633 4669
rect 14576 4652 14593 4669
rect 14536 4652 14553 4669
rect 14496 4652 14513 4669
rect 14456 4652 14473 4669
rect 14416 4652 14433 4669
rect 14816 4652 14833 4669
rect 14776 4652 14793 4669
rect 14736 4652 14753 4669
rect 14696 4652 14713 4669
rect 14496 4652 14513 4669
rect 14616 4652 14633 4669
rect 14456 4652 14473 4669
rect 14936 4652 14953 4669
rect 14416 4652 14433 4669
rect 14816 4652 14833 4669
rect 14576 4652 14593 4669
rect 14776 4652 14793 4669
rect 14736 4652 14753 4669
rect 14856 4652 14873 4669
rect 14696 4652 14713 4669
rect 14536 4652 14553 4669
rect 14496 4652 14513 4669
rect 14936 4652 14953 4669
rect 14456 4652 14473 4669
rect 14416 4652 14433 4669
rect 14856 4652 14873 4669
rect 14816 4652 14833 4669
rect 14776 4652 14793 4669
rect 14736 4652 14753 4669
rect 14696 4652 14713 4669
rect 14656 4652 14673 4669
rect 14856 4652 14873 4669
rect 14616 4652 14633 4669
rect 14936 4652 14953 4669
rect 14656 4652 14673 4669
rect 14576 4652 14593 4669
rect 14896 4652 14913 4669
rect 14536 4652 14553 4669
rect 14896 4652 14913 4669
rect 14936 4652 14953 4669
rect 18616 4652 18633 4669
rect 18616 4652 18633 4669
rect 18976 4652 18993 4669
rect 18936 4652 18953 4669
rect 18896 4652 18913 4669
rect 18856 4652 18873 4669
rect 18816 4652 18833 4669
rect 18776 4652 18793 4669
rect 18736 4652 18753 4669
rect 19136 4652 19153 4669
rect 19096 4652 19113 4669
rect 19056 4652 19073 4669
rect 19016 4652 19033 4669
rect 18976 4652 18993 4669
rect 18936 4652 18953 4669
rect 18896 4652 18913 4669
rect 18856 4652 18873 4669
rect 18816 4652 18833 4669
rect 18776 4652 18793 4669
rect 18736 4652 18753 4669
rect 19136 4652 19153 4669
rect 19096 4652 19113 4669
rect 19056 4652 19073 4669
rect 19016 4652 19033 4669
rect 18696 4652 18713 4669
rect 18656 4652 18673 4669
rect 18696 4652 18713 4669
rect 18656 4652 18673 4669
rect 18736 4652 18753 4669
rect 19136 4652 19153 4669
rect 18576 4652 18593 4669
rect 19096 4652 19113 4669
rect 19056 4652 19073 4669
rect 19016 4652 19033 4669
rect 18976 4652 18993 4669
rect 18576 4652 18593 4669
rect 18936 4652 18953 4669
rect 18896 4652 18913 4669
rect 18856 4652 18873 4669
rect 18816 4652 18833 4669
rect 18776 4652 18793 4669
rect 18576 4652 18593 4669
rect 18736 4652 18753 4669
rect 19136 4652 19153 4669
rect 19096 4652 19113 4669
rect 19056 4652 19073 4669
rect 19016 4652 19033 4669
rect 18696 4652 18713 4669
rect 18656 4652 18673 4669
rect 18696 4652 18713 4669
rect 18656 4652 18673 4669
rect 18976 4652 18993 4669
rect 18936 4652 18953 4669
rect 18576 4652 18593 4669
rect 18896 4652 18913 4669
rect 18856 4652 18873 4669
rect 18816 4652 18833 4669
rect 18616 4652 18633 4669
rect 18616 4652 18633 4669
rect 18776 4652 18793 4669
rect 18336 4652 18353 4669
rect 18536 4652 18553 4669
rect 18256 4652 18273 4669
rect 18496 4652 18513 4669
rect 18216 4652 18233 4669
rect 18176 4652 18193 4669
rect 18136 4652 18153 4669
rect 18096 4652 18113 4669
rect 18456 4652 18473 4669
rect 18416 4652 18433 4669
rect 18376 4652 18393 4669
rect 18536 4652 18553 4669
rect 18496 4652 18513 4669
rect 18456 4652 18473 4669
rect 18416 4652 18433 4669
rect 18376 4652 18393 4669
rect 18336 4652 18353 4669
rect 18296 4652 18313 4669
rect 18256 4652 18273 4669
rect 18216 4652 18233 4669
rect 18176 4652 18193 4669
rect 18136 4652 18153 4669
rect 18096 4652 18113 4669
rect 17976 4652 17993 4669
rect 18016 4652 18033 4669
rect 18056 4652 18073 4669
rect 18016 4652 18033 4669
rect 18056 4652 18073 4669
rect 17976 4652 17993 4669
rect 18016 4652 18033 4669
rect 18056 4652 18073 4669
rect 17976 4652 17993 4669
rect 18296 4652 18313 4669
rect 18336 4652 18353 4669
rect 18536 4652 18553 4669
rect 18256 4652 18273 4669
rect 18496 4652 18513 4669
rect 18216 4652 18233 4669
rect 18176 4652 18193 4669
rect 18136 4652 18153 4669
rect 18096 4652 18113 4669
rect 18456 4652 18473 4669
rect 18416 4652 18433 4669
rect 18376 4652 18393 4669
rect 17976 4652 17993 4669
rect 18016 4652 18033 4669
rect 18056 4652 18073 4669
rect 18536 4652 18553 4669
rect 18496 4652 18513 4669
rect 18456 4652 18473 4669
rect 18416 4652 18433 4669
rect 18376 4652 18393 4669
rect 18336 4652 18353 4669
rect 18296 4652 18313 4669
rect 18256 4652 18273 4669
rect 18216 4652 18233 4669
rect 18176 4652 18193 4669
rect 18136 4652 18153 4669
rect 18096 4652 18113 4669
rect 18296 4652 18313 4669
rect 17936 4652 17953 4669
rect 17616 4652 17633 4669
rect 17576 4652 17593 4669
rect 17376 4652 17393 4669
rect 17616 4652 17633 4669
rect 17456 4652 17473 4669
rect 17776 4652 17793 4669
rect 17776 4652 17793 4669
rect 17536 4652 17553 4669
rect 17536 4652 17553 4669
rect 17936 4652 17953 4669
rect 17416 4652 17433 4669
rect 17496 4652 17513 4669
rect 17496 4652 17513 4669
rect 17376 4652 17393 4669
rect 17656 4652 17673 4669
rect 17736 4652 17753 4669
rect 17896 4652 17913 4669
rect 17936 4652 17953 4669
rect 17416 4652 17433 4669
rect 17856 4652 17873 4669
rect 17536 4652 17553 4669
rect 17616 4652 17633 4669
rect 17856 4652 17873 4669
rect 17536 4652 17553 4669
rect 17576 4652 17593 4669
rect 17816 4652 17833 4669
rect 17816 4652 17833 4669
rect 17776 4652 17793 4669
rect 17376 4652 17393 4669
rect 17736 4652 17753 4669
rect 17456 4652 17473 4669
rect 17696 4652 17713 4669
rect 17656 4652 17673 4669
rect 17656 4652 17673 4669
rect 17896 4652 17913 4669
rect 17936 4652 17953 4669
rect 17896 4652 17913 4669
rect 17416 4652 17433 4669
rect 17496 4652 17513 4669
rect 17376 4652 17393 4669
rect 17696 4652 17713 4669
rect 17456 4652 17473 4669
rect 17856 4652 17873 4669
rect 17456 4652 17473 4669
rect 17616 4652 17633 4669
rect 17736 4652 17753 4669
rect 17856 4652 17873 4669
rect 17896 4652 17913 4669
rect 17696 4652 17713 4669
rect 17416 4652 17433 4669
rect 17576 4652 17593 4669
rect 17816 4652 17833 4669
rect 17816 4652 17833 4669
rect 17776 4652 17793 4669
rect 17576 4652 17593 4669
rect 17736 4652 17753 4669
rect 17496 4652 17513 4669
rect 17696 4652 17713 4669
rect 17656 4652 17673 4669
rect 16856 4652 16873 4669
rect 16816 4652 16833 4669
rect 16776 4652 16793 4669
rect 17216 4652 17233 4669
rect 17256 4652 17273 4669
rect 17256 4652 17273 4669
rect 17016 4652 17033 4669
rect 16976 4652 16993 4669
rect 17336 4652 17353 4669
rect 17296 4652 17313 4669
rect 16936 4652 16953 4669
rect 16896 4652 16913 4669
rect 16856 4652 16873 4669
rect 16976 4652 16993 4669
rect 16816 4652 16833 4669
rect 16936 4652 16953 4669
rect 17176 4652 17193 4669
rect 17176 4652 17193 4669
rect 17056 4652 17073 4669
rect 17136 4652 17153 4669
rect 17216 4652 17233 4669
rect 17096 4652 17113 4669
rect 17016 4652 17033 4669
rect 17056 4652 17073 4669
rect 16896 4652 16913 4669
rect 17336 4652 17353 4669
rect 17296 4652 17313 4669
rect 17136 4652 17153 4669
rect 16776 4652 16793 4669
rect 17096 4652 17113 4669
rect 16856 4652 16873 4669
rect 17216 4652 17233 4669
rect 17256 4652 17273 4669
rect 17256 4652 17273 4669
rect 17016 4652 17033 4669
rect 17056 4652 17073 4669
rect 16936 4652 16953 4669
rect 17336 4652 17353 4669
rect 16896 4652 16913 4669
rect 17296 4652 17313 4669
rect 17136 4652 17153 4669
rect 17096 4652 17113 4669
rect 16856 4652 16873 4669
rect 16976 4652 16993 4669
rect 16816 4652 16833 4669
rect 17336 4652 17353 4669
rect 17296 4652 17313 4669
rect 16816 4652 16833 4669
rect 16776 4652 16793 4669
rect 16976 4652 16993 4669
rect 17176 4652 17193 4669
rect 17176 4652 17193 4669
rect 17056 4652 17073 4669
rect 16936 4652 16953 4669
rect 16896 4652 16913 4669
rect 17136 4652 17153 4669
rect 17216 4652 17233 4669
rect 17096 4652 17113 4669
rect 17016 4652 17033 4669
rect 16776 4652 16793 4669
rect 10816 4652 10833 4669
rect 10816 4652 10833 4669
rect 10816 4652 10833 4669
rect 10816 4652 10833 4669
rect 11416 4652 11433 4669
rect 11416 4652 11433 4669
rect 11416 4652 11433 4669
rect 11416 4652 11433 4669
rect 11776 4652 11793 4669
rect 11816 4652 11833 4669
rect 11656 4652 11673 4669
rect 11776 4652 11793 4669
rect 11456 4652 11473 4669
rect 11776 4652 11793 4669
rect 11576 4652 11593 4669
rect 11896 4652 11913 4669
rect 11976 4652 11993 4669
rect 11696 4652 11713 4669
rect 11456 4652 11473 4669
rect 11976 4652 11993 4669
rect 11616 4652 11633 4669
rect 11656 4652 11673 4669
rect 11656 4652 11673 4669
rect 11456 4652 11473 4669
rect 11536 4652 11553 4669
rect 11936 4652 11953 4669
rect 11536 4652 11553 4669
rect 11936 4652 11953 4669
rect 11736 4652 11753 4669
rect 11896 4652 11913 4669
rect 11616 4652 11633 4669
rect 11536 4652 11553 4669
rect 11536 4652 11553 4669
rect 11616 4652 11633 4669
rect 11856 4652 11873 4669
rect 11896 4652 11913 4669
rect 11736 4652 11753 4669
rect 11696 4652 11713 4669
rect 11856 4652 11873 4669
rect 11816 4652 11833 4669
rect 11976 4652 11993 4669
rect 11736 4652 11753 4669
rect 11496 4652 11513 4669
rect 11656 4652 11673 4669
rect 11856 4652 11873 4669
rect 11576 4652 11593 4669
rect 11616 4652 11633 4669
rect 11496 4652 11513 4669
rect 11576 4652 11593 4669
rect 11736 4652 11753 4669
rect 11976 4652 11993 4669
rect 11936 4652 11953 4669
rect 11816 4652 11833 4669
rect 11576 4652 11593 4669
rect 11776 4652 11793 4669
rect 11936 4652 11953 4669
rect 11896 4652 11913 4669
rect 11856 4652 11873 4669
rect 11816 4652 11833 4669
rect 11696 4652 11713 4669
rect 11696 4652 11713 4669
rect 11496 4652 11513 4669
rect 11496 4652 11513 4669
rect 11456 4652 11473 4669
rect 11336 4652 11353 4669
rect 11376 4652 11393 4669
rect 11296 4652 11313 4669
rect 11176 4652 11193 4669
rect 11176 4652 11193 4669
rect 11216 4652 11233 4669
rect 11136 4652 11153 4669
rect 10856 4652 10873 4669
rect 10856 4652 10873 4669
rect 11096 4652 11113 4669
rect 11096 4652 11113 4669
rect 10936 4652 10953 4669
rect 11056 4652 11073 4669
rect 11256 4652 11273 4669
rect 11256 4652 11273 4669
rect 11216 4652 11233 4669
rect 11056 4652 11073 4669
rect 11056 4652 11073 4669
rect 10976 4652 10993 4669
rect 11176 4652 11193 4669
rect 11336 4652 11353 4669
rect 11216 4652 11233 4669
rect 11136 4652 11153 4669
rect 11376 4652 11393 4669
rect 11256 4652 11273 4669
rect 10856 4652 10873 4669
rect 10976 4652 10993 4669
rect 11096 4652 11113 4669
rect 11016 4652 11033 4669
rect 11096 4652 11113 4669
rect 11256 4652 11273 4669
rect 11176 4652 11193 4669
rect 11336 4652 11353 4669
rect 11016 4652 11033 4669
rect 11296 4652 11313 4669
rect 10896 4652 10913 4669
rect 11376 4652 11393 4669
rect 11136 4652 11153 4669
rect 10976 4652 10993 4669
rect 10896 4652 10913 4669
rect 10936 4652 10953 4669
rect 10856 4652 10873 4669
rect 11336 4652 11353 4669
rect 10936 4652 10953 4669
rect 11296 4652 11313 4669
rect 11056 4652 11073 4669
rect 11216 4652 11233 4669
rect 11016 4652 11033 4669
rect 10896 4652 10913 4669
rect 11136 4652 11153 4669
rect 10896 4652 10913 4669
rect 11016 4652 11033 4669
rect 11296 4652 11313 4669
rect 10976 4652 10993 4669
rect 10936 4652 10953 4669
rect 11376 4652 11393 4669
rect 10216 4652 10233 4669
rect 10216 4652 10233 4669
rect 10216 4652 10233 4669
rect 10216 4652 10233 4669
rect 10776 4652 10793 4669
rect 10376 4652 10393 4669
rect 10776 4652 10793 4669
rect 10336 4652 10353 4669
rect 10656 4652 10673 4669
rect 10456 4652 10473 4669
rect 10776 4652 10793 4669
rect 10296 4652 10313 4669
rect 10416 4652 10433 4669
rect 10616 4652 10633 4669
rect 10376 4652 10393 4669
rect 10536 4652 10553 4669
rect 10576 4652 10593 4669
rect 10496 4652 10513 4669
rect 10576 4652 10593 4669
rect 10456 4652 10473 4669
rect 10736 4652 10753 4669
rect 10256 4652 10273 4669
rect 10616 4652 10633 4669
rect 10576 4652 10593 4669
rect 10696 4652 10713 4669
rect 10496 4652 10513 4669
rect 10736 4652 10753 4669
rect 10736 4652 10753 4669
rect 10576 4652 10593 4669
rect 10656 4652 10673 4669
rect 10336 4652 10353 4669
rect 10696 4652 10713 4669
rect 10736 4652 10753 4669
rect 10536 4652 10553 4669
rect 10696 4652 10713 4669
rect 10296 4652 10313 4669
rect 10496 4652 10513 4669
rect 10656 4652 10673 4669
rect 10256 4652 10273 4669
rect 10336 4652 10353 4669
rect 10296 4652 10313 4669
rect 10256 4652 10273 4669
rect 10656 4652 10673 4669
rect 10616 4652 10633 4669
rect 10456 4652 10473 4669
rect 10416 4652 10433 4669
rect 10696 4652 10713 4669
rect 10496 4652 10513 4669
rect 10456 4652 10473 4669
rect 10616 4652 10633 4669
rect 10416 4652 10433 4669
rect 10536 4652 10553 4669
rect 10376 4652 10393 4669
rect 10776 4652 10793 4669
rect 10336 4652 10353 4669
rect 10296 4652 10313 4669
rect 10256 4652 10273 4669
rect 10416 4652 10433 4669
rect 10376 4652 10393 4669
rect 10536 4652 10553 4669
rect 9856 4652 9873 4669
rect 9696 4652 9713 4669
rect 10136 4652 10153 4669
rect 10096 4652 10113 4669
rect 9656 4652 9673 4669
rect 9816 4652 9833 4669
rect 9936 4652 9953 4669
rect 9776 4652 9793 4669
rect 9736 4652 9753 4669
rect 9896 4652 9913 4669
rect 9936 4652 9953 4669
rect 9896 4652 9913 4669
rect 9856 4652 9873 4669
rect 9816 4652 9833 4669
rect 9776 4652 9793 4669
rect 9736 4652 9753 4669
rect 9696 4652 9713 4669
rect 9656 4652 9673 4669
rect 9856 4652 9873 4669
rect 9896 4652 9913 4669
rect 9816 4652 9833 4669
rect 10136 4652 10153 4669
rect 9776 4652 9793 4669
rect 10096 4652 10113 4669
rect 9736 4652 9753 4669
rect 9856 4652 9873 4669
rect 9696 4652 9713 4669
rect 9656 4652 9673 4669
rect 10096 4652 10113 4669
rect 9936 4652 9953 4669
rect 9976 4652 9993 4669
rect 10136 4652 10153 4669
rect 9816 4652 9833 4669
rect 10056 4652 10073 4669
rect 10176 4652 10193 4669
rect 10016 4652 10033 4669
rect 9776 4652 9793 4669
rect 10056 4652 10073 4669
rect 9736 4652 9753 4669
rect 9976 4652 9993 4669
rect 10056 4652 10073 4669
rect 10016 4652 10033 4669
rect 9936 4652 9953 4669
rect 10016 4652 10033 4669
rect 9896 4652 9913 4669
rect 9696 4652 9713 4669
rect 9656 4652 9673 4669
rect 10176 4652 10193 4669
rect 10056 4652 10073 4669
rect 10176 4652 10193 4669
rect 10136 4652 10153 4669
rect 10096 4652 10113 4669
rect 9976 4652 9993 4669
rect 10016 4652 10033 4669
rect 10176 4652 10193 4669
rect 9976 4652 9993 4669
rect 13856 4652 13873 4669
rect 13816 4652 13833 4669
rect 14176 4652 14193 4669
rect 13896 4652 13913 4669
rect 13856 4652 13873 4669
rect 13816 4652 13833 4669
rect 13936 4652 13953 4669
rect 14136 4652 14153 4669
rect 14096 4652 14113 4669
rect 14056 4652 14073 4669
rect 14256 4652 14273 4669
rect 14296 4652 14313 4669
rect 14296 4652 14313 4669
rect 14376 4652 14393 4669
rect 14336 4652 14353 4669
rect 14376 4652 14393 4669
rect 14336 4652 14353 4669
rect 13976 4652 13993 4669
rect 14016 4652 14033 4669
rect 14256 4652 14273 4669
rect 14216 4652 14233 4669
rect 14216 4652 14233 4669
rect 14296 4652 14313 4669
rect 14296 4652 14313 4669
rect 14376 4652 14393 4669
rect 14336 4652 14353 4669
rect 14376 4652 14393 4669
rect 14336 4652 14353 4669
rect 13976 4652 13993 4669
rect 14016 4652 14033 4669
rect 14256 4652 14273 4669
rect 14216 4652 14233 4669
rect 13936 4652 13953 4669
rect 14176 4652 14193 4669
rect 13896 4652 13913 4669
rect 13856 4652 13873 4669
rect 13816 4652 13833 4669
rect 14176 4652 14193 4669
rect 14136 4652 14153 4669
rect 14096 4652 14113 4669
rect 14056 4652 14073 4669
rect 14256 4652 14273 4669
rect 14216 4652 14233 4669
rect 14176 4652 14193 4669
rect 14136 4652 14153 4669
rect 14096 4652 14113 4669
rect 14056 4652 14073 4669
rect 14016 4652 14033 4669
rect 13976 4652 13993 4669
rect 13936 4652 13953 4669
rect 13896 4652 13913 4669
rect 13856 4652 13873 4669
rect 13816 4652 13833 4669
rect 14136 4652 14153 4669
rect 14096 4652 14113 4669
rect 14056 4652 14073 4669
rect 14016 4652 14033 4669
rect 13976 4652 13993 4669
rect 13936 4652 13953 4669
rect 13896 4652 13913 4669
rect 13696 4652 13713 4669
rect 13256 4652 13273 4669
rect 13496 4652 13513 4669
rect 13496 4652 13513 4669
rect 13456 4652 13473 4669
rect 13416 4652 13433 4669
rect 13736 4652 13753 4669
rect 13376 4652 13393 4669
rect 13336 4652 13353 4669
rect 13616 4652 13633 4669
rect 13296 4652 13313 4669
rect 13256 4652 13273 4669
rect 13456 4652 13473 4669
rect 13216 4652 13233 4669
rect 13216 4652 13233 4669
rect 13696 4652 13713 4669
rect 13736 4652 13753 4669
rect 13416 4652 13433 4669
rect 13656 4652 13673 4669
rect 13576 4652 13593 4669
rect 13376 4652 13393 4669
rect 13776 4652 13793 4669
rect 13776 4652 13793 4669
rect 13656 4652 13673 4669
rect 13336 4652 13353 4669
rect 13576 4652 13593 4669
rect 13536 4652 13553 4669
rect 13296 4652 13313 4669
rect 13536 4652 13553 4669
rect 13696 4652 13713 4669
rect 13256 4652 13273 4669
rect 13496 4652 13513 4669
rect 13496 4652 13513 4669
rect 13456 4652 13473 4669
rect 13416 4652 13433 4669
rect 13736 4652 13753 4669
rect 13376 4652 13393 4669
rect 13336 4652 13353 4669
rect 13616 4652 13633 4669
rect 13296 4652 13313 4669
rect 13256 4652 13273 4669
rect 13456 4652 13473 4669
rect 13216 4652 13233 4669
rect 13216 4652 13233 4669
rect 13696 4652 13713 4669
rect 13736 4652 13753 4669
rect 13416 4652 13433 4669
rect 13656 4652 13673 4669
rect 13576 4652 13593 4669
rect 13376 4652 13393 4669
rect 13616 4652 13633 4669
rect 13616 4652 13633 4669
rect 13776 4652 13793 4669
rect 13776 4652 13793 4669
rect 13656 4652 13673 4669
rect 13336 4652 13353 4669
rect 13576 4652 13593 4669
rect 13536 4652 13553 4669
rect 13296 4652 13313 4669
rect 13536 4652 13553 4669
rect 12936 4652 12953 4669
rect 12776 4652 12793 4669
rect 12616 4652 12633 4669
rect 12616 4652 12633 4669
rect 12776 4652 12793 4669
rect 12816 4652 12833 4669
rect 12656 4652 12673 4669
rect 12656 4652 12673 4669
rect 12896 4652 12913 4669
rect 12696 4652 12713 4669
rect 12936 4652 12953 4669
rect 13176 4652 13193 4669
rect 12696 4652 12713 4669
rect 13136 4652 13153 4669
rect 13056 4652 13073 4669
rect 13096 4652 13113 4669
rect 13096 4652 13113 4669
rect 13016 4652 13033 4669
rect 13176 4652 13193 4669
rect 12616 4652 12633 4669
rect 13056 4652 13073 4669
rect 13016 4652 13033 4669
rect 13136 4652 13153 4669
rect 12976 4652 12993 4669
rect 12976 4652 12993 4669
rect 12776 4652 12793 4669
rect 12736 4652 12753 4669
rect 13176 4652 13193 4669
rect 12896 4652 12913 4669
rect 12856 4652 12873 4669
rect 12816 4652 12833 4669
rect 13136 4652 13153 4669
rect 13096 4652 13113 4669
rect 13176 4652 13193 4669
rect 13096 4652 13113 4669
rect 12856 4652 12873 4669
rect 12856 4652 12873 4669
rect 13056 4652 13073 4669
rect 12736 4652 12753 4669
rect 12816 4652 12833 4669
rect 13056 4652 13073 4669
rect 12656 4652 12673 4669
rect 13016 4652 13033 4669
rect 12616 4652 12633 4669
rect 12896 4652 12913 4669
rect 12776 4652 12793 4669
rect 12696 4652 12713 4669
rect 12736 4652 12753 4669
rect 13136 4652 13153 4669
rect 12976 4652 12993 4669
rect 13016 4652 13033 4669
rect 12896 4652 12913 4669
rect 12936 4652 12953 4669
rect 12936 4652 12953 4669
rect 12856 4652 12873 4669
rect 12976 4652 12993 4669
rect 12736 4652 12753 4669
rect 12816 4652 12833 4669
rect 12656 4652 12673 4669
rect 12696 4652 12713 4669
rect 12456 4652 12473 4669
rect 12136 4652 12153 4669
rect 12376 4652 12393 4669
rect 12416 4652 12433 4669
rect 12056 4652 12073 4669
rect 12016 4652 12033 4669
rect 12536 4652 12553 4669
rect 12216 4652 12233 4669
rect 12016 4652 12033 4669
rect 12496 4652 12513 4669
rect 12056 4652 12073 4669
rect 12016 4652 12033 4669
rect 12536 4652 12553 4669
rect 12216 4652 12233 4669
rect 12416 4652 12433 4669
rect 12376 4652 12393 4669
rect 12016 4652 12033 4669
rect 12496 4652 12513 4669
rect 12336 4652 12353 4669
rect 12576 4652 12593 4669
rect 12296 4652 12313 4669
rect 12096 4652 12113 4669
rect 12456 4652 12473 4669
rect 12256 4652 12273 4669
rect 12296 4652 12313 4669
rect 12536 4652 12553 4669
rect 12176 4652 12193 4669
rect 12576 4652 12593 4669
rect 12096 4652 12113 4669
rect 12256 4652 12273 4669
rect 12496 4652 12513 4669
rect 12576 4652 12593 4669
rect 12456 4652 12473 4669
rect 12536 4652 12553 4669
rect 12496 4652 12513 4669
rect 12176 4652 12193 4669
rect 12456 4652 12473 4669
rect 12416 4652 12433 4669
rect 12136 4652 12153 4669
rect 12416 4652 12433 4669
rect 12056 4652 12073 4669
rect 12376 4652 12393 4669
rect 12336 4652 12353 4669
rect 12296 4652 12313 4669
rect 12296 4652 12313 4669
rect 12256 4652 12273 4669
rect 12136 4652 12153 4669
rect 12216 4652 12233 4669
rect 12176 4652 12193 4669
rect 12136 4652 12153 4669
rect 12376 4652 12393 4669
rect 12096 4652 12113 4669
rect 12216 4652 12233 4669
rect 12096 4652 12113 4669
rect 12256 4652 12273 4669
rect 12576 4652 12593 4669
rect 12056 4652 12073 4669
rect 12336 4652 12353 4669
rect 12176 4652 12193 4669
rect 12336 4652 12353 4669
rect 10796 3163 10813 3180
rect 11116 3163 11133 3180
rect 11076 3163 11093 3180
rect 11036 3163 11053 3180
rect 10996 3163 11013 3180
rect 10956 3163 10973 3180
rect 10916 3163 10933 3180
rect 10876 3163 10893 3180
rect 11116 3163 11133 3180
rect 11076 3163 11093 3180
rect 11036 3163 11053 3180
rect 10796 3163 10813 3180
rect 11076 3163 11093 3180
rect 10956 3163 10973 3180
rect 11276 3163 11293 3180
rect 11276 3163 11293 3180
rect 11156 3163 11173 3180
rect 11156 3163 11173 3180
rect 10916 3163 10933 3180
rect 10876 3163 10893 3180
rect 10996 3163 11013 3180
rect 11196 3163 11213 3180
rect 11116 3163 11133 3180
rect 11036 3163 11053 3180
rect 10956 3163 10973 3180
rect 10876 3163 10893 3180
rect 10996 3163 11013 3180
rect 11236 3163 11253 3180
rect 11236 3163 11253 3180
rect 10916 3163 10933 3180
rect 10916 3163 10933 3180
rect 10796 3163 10813 3180
rect 11236 3163 11253 3180
rect 10876 3163 10893 3180
rect 11156 3163 11173 3180
rect 10676 3163 10693 3180
rect 10236 3163 10253 3180
rect 10276 3163 10293 3180
rect 10476 3163 10493 3180
rect 10436 3163 10453 3180
rect 10316 3163 10333 3180
rect 10556 3163 10573 3180
rect 10396 3163 10413 3180
rect 10716 3163 10733 3180
rect 10716 3163 10733 3180
rect 10516 3163 10533 3180
rect 10716 3163 10733 3180
rect 10476 3163 10493 3180
rect 10356 3163 10373 3180
rect 10556 3163 10573 3180
rect 10316 3163 10333 3180
rect 10436 3163 10453 3180
rect 10396 3163 10413 3180
rect 10436 3163 10453 3180
rect 10356 3163 10373 3180
rect 10236 3163 10253 3180
rect 10596 3163 10613 3180
rect 10676 3163 10693 3180
rect 10396 3163 10413 3180
rect 10276 3163 10293 3180
rect 10276 3163 10293 3180
rect 10636 3163 10653 3180
rect 10396 3163 10413 3180
rect 10556 3163 10573 3180
rect 10516 3163 10533 3180
rect 10636 3163 10653 3180
rect 10676 3163 10693 3180
rect 10236 3163 10253 3180
rect 10516 3163 10533 3180
rect 10676 3163 10693 3180
rect 10716 3163 10733 3180
rect 10596 3163 10613 3180
rect 10516 3163 10533 3180
rect 10636 3163 10653 3180
rect 10276 3163 10293 3180
rect 10316 3163 10333 3180
rect 10476 3163 10493 3180
rect 10436 3163 10453 3180
rect 10636 3163 10653 3180
rect 10476 3163 10493 3180
rect 10316 3163 10333 3180
rect 10356 3163 10373 3180
rect 10596 3163 10613 3180
rect 10356 3163 10373 3180
rect 10596 3163 10613 3180
rect 10556 3163 10573 3180
rect 10236 3163 10253 3180
rect 9676 3163 9693 3180
rect 9676 3163 9693 3180
rect 9676 3163 9693 3180
rect 9676 3163 9693 3180
rect 10116 3163 10133 3180
rect 9916 3163 9933 3180
rect 9836 3163 9853 3180
rect 9876 3163 9893 3180
rect 9836 3163 9853 3180
rect 9716 3163 9733 3180
rect 9956 3163 9973 3180
rect 9796 3163 9813 3180
rect 9996 3163 10013 3180
rect 9916 3163 9933 3180
rect 9796 3163 9813 3180
rect 10076 3163 10093 3180
rect 10196 3163 10213 3180
rect 9956 3163 9973 3180
rect 10196 3163 10213 3180
rect 9956 3163 9973 3180
rect 10156 3163 10173 3180
rect 9996 3163 10013 3180
rect 9796 3163 9813 3180
rect 9916 3163 9933 3180
rect 9916 3163 9933 3180
rect 9876 3163 9893 3180
rect 10076 3163 10093 3180
rect 9756 3163 9773 3180
rect 9836 3163 9853 3180
rect 10116 3163 10133 3180
rect 9756 3163 9773 3180
rect 9796 3163 9813 3180
rect 10036 3163 10053 3180
rect 9876 3163 9893 3180
rect 10036 3163 10053 3180
rect 10196 3163 10213 3180
rect 9716 3163 9733 3180
rect 9716 3163 9733 3180
rect 9996 3163 10013 3180
rect 9876 3163 9893 3180
rect 10196 3163 10213 3180
rect 9756 3163 9773 3180
rect 9756 3163 9773 3180
rect 10156 3163 10173 3180
rect 10156 3163 10173 3180
rect 10116 3163 10133 3180
rect 10036 3163 10053 3180
rect 10036 3163 10053 3180
rect 10076 3163 10093 3180
rect 9716 3163 9733 3180
rect 9956 3163 9973 3180
rect 9836 3163 9853 3180
rect 10156 3163 10173 3180
rect 10076 3163 10093 3180
rect 9996 3163 10013 3180
rect 10116 3163 10133 3180
rect 9636 3163 9653 3180
rect 9636 3163 9653 3180
rect 9636 3163 9653 3180
rect 9636 3163 9653 3180
rect 14277 3163 14294 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 14357 3163 14374 3180
rect 13997 3163 14014 3180
rect 14277 3163 14294 3180
rect 14357 3163 14374 3180
rect 14317 3163 14334 3180
rect 14357 3163 14374 3180
rect 14277 3163 14294 3180
rect 14317 3163 14334 3180
rect 14237 3163 14254 3180
rect 14277 3163 14294 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14357 3163 14374 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14317 3163 14334 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14317 3163 14334 3180
rect 13837 3163 13854 3180
rect 13957 3163 13974 3180
rect 13917 3163 13934 3180
rect 13877 3163 13894 3180
rect 13837 3163 13854 3180
rect 13917 3163 13934 3180
rect 13917 3163 13934 3180
rect 13517 3163 13534 3180
rect 13597 3163 13614 3180
rect 13597 3163 13614 3180
rect 13877 3163 13894 3180
rect 13677 3163 13694 3180
rect 13837 3163 13854 3180
rect 13837 3163 13854 3180
rect 13557 3163 13574 3180
rect 13957 3163 13974 3180
rect 13877 3163 13894 3180
rect 13957 3163 13974 3180
rect 13637 3163 13654 3180
rect 13957 3163 13974 3180
rect 13917 3163 13934 3180
rect 13757 3163 13774 3180
rect 13877 3163 13894 3180
rect 13477 3163 13494 3180
rect 13797 3163 13814 3180
rect 13717 3163 13734 3180
rect 13797 3163 13814 3180
rect 13797 3163 13814 3180
rect 13757 3163 13774 3180
rect 13757 3163 13774 3180
rect 13717 3163 13734 3180
rect 13677 3163 13694 3180
rect 13637 3163 13654 3180
rect 13677 3163 13694 3180
rect 13597 3163 13614 3180
rect 13557 3163 13574 3180
rect 13517 3163 13534 3180
rect 13477 3163 13494 3180
rect 13557 3163 13574 3180
rect 13717 3163 13734 3180
rect 13637 3163 13654 3180
rect 13677 3163 13694 3180
rect 13597 3163 13614 3180
rect 13717 3163 13734 3180
rect 13637 3163 13654 3180
rect 13517 3163 13534 3180
rect 13557 3163 13574 3180
rect 13477 3163 13494 3180
rect 13757 3163 13774 3180
rect 13517 3163 13534 3180
rect 13797 3163 13814 3180
rect 13477 3163 13494 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 13237 3163 13254 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13397 3163 13414 3180
rect 13037 3163 13054 3180
rect 13397 3163 13414 3180
rect 13197 3163 13214 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13357 3163 13374 3180
rect 13117 3163 13134 3180
rect 13437 3163 13454 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13037 3163 13054 3180
rect 13277 3163 13294 3180
rect 12997 3163 13014 3180
rect 13277 3163 13294 3180
rect 12957 3163 12974 3180
rect 13237 3163 13254 3180
rect 13197 3163 13214 3180
rect 13277 3163 13294 3180
rect 12957 3163 12974 3180
rect 13237 3163 13254 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13437 3163 13454 3180
rect 12997 3163 13014 3180
rect 13277 3163 13294 3180
rect 12997 3163 13014 3180
rect 13437 3163 13454 3180
rect 13197 3163 13214 3180
rect 13117 3163 13134 3180
rect 13117 3163 13134 3180
rect 13037 3163 13054 3180
rect 13037 3163 13054 3180
rect 13117 3163 13134 3180
rect 12957 3163 12974 3180
rect 13197 3163 13214 3180
rect 13077 3163 13094 3180
rect 13157 3163 13174 3180
rect 12997 3163 13014 3180
rect 13397 3163 13414 3180
rect 13357 3163 13374 3180
rect 13357 3163 13374 3180
rect 13357 3163 13374 3180
rect 13237 3163 13254 3180
rect 13437 3163 13454 3180
rect 12957 3163 12974 3180
rect 13397 3163 13414 3180
rect 12637 3163 12654 3180
rect 12677 3163 12694 3180
rect 12437 3163 12454 3180
rect 12517 3163 12534 3180
rect 12757 3163 12774 3180
rect 12637 3163 12654 3180
rect 12437 3163 12454 3180
rect 12757 3163 12774 3180
rect 12637 3163 12654 3180
rect 12517 3163 12534 3180
rect 12637 3163 12654 3180
rect 12797 3163 12814 3180
rect 12597 3163 12614 3180
rect 12477 3163 12494 3180
rect 12837 3163 12854 3180
rect 12797 3163 12814 3180
rect 12397 3163 12414 3180
rect 12597 3163 12614 3180
rect 12717 3163 12734 3180
rect 12877 3163 12894 3180
rect 12597 3163 12614 3180
rect 12877 3163 12894 3180
rect 12877 3163 12894 3180
rect 12757 3163 12774 3180
rect 12717 3163 12734 3180
rect 12557 3163 12574 3180
rect 12717 3163 12734 3180
rect 12477 3163 12494 3180
rect 12837 3163 12854 3180
rect 12477 3163 12494 3180
rect 12397 3163 12414 3180
rect 12397 3163 12414 3180
rect 12717 3163 12734 3180
rect 12557 3163 12574 3180
rect 12877 3163 12894 3180
rect 12677 3163 12694 3180
rect 12837 3163 12854 3180
rect 12797 3163 12814 3180
rect 12557 3163 12574 3180
rect 12477 3163 12494 3180
rect 12837 3163 12854 3180
rect 12757 3163 12774 3180
rect 12677 3163 12694 3180
rect 12437 3163 12454 3180
rect 12557 3163 12574 3180
rect 12397 3163 12414 3180
rect 12677 3163 12694 3180
rect 12797 3163 12814 3180
rect 12597 3163 12614 3180
rect 12517 3163 12534 3180
rect 12517 3163 12534 3180
rect 12437 3163 12454 3180
rect 11837 3163 11854 3180
rect 11837 3163 11854 3180
rect 11837 3163 11854 3180
rect 11837 3163 11854 3180
rect 12197 3163 12214 3180
rect 12277 3163 12294 3180
rect 12117 3163 12134 3180
rect 12237 3163 12254 3180
rect 11917 3163 11934 3180
rect 12037 3163 12054 3180
rect 11877 3163 11894 3180
rect 12357 3163 12374 3180
rect 12157 3163 12174 3180
rect 12357 3163 12374 3180
rect 12317 3163 12334 3180
rect 11957 3163 11974 3180
rect 12237 3163 12254 3180
rect 12317 3163 12334 3180
rect 11997 3163 12014 3180
rect 12237 3163 12254 3180
rect 12277 3163 12294 3180
rect 12197 3163 12214 3180
rect 11997 3163 12014 3180
rect 12117 3163 12134 3180
rect 11877 3163 11894 3180
rect 11877 3163 11894 3180
rect 12037 3163 12054 3180
rect 12197 3163 12214 3180
rect 12157 3163 12174 3180
rect 12077 3163 12094 3180
rect 12117 3163 12134 3180
rect 12077 3163 12094 3180
rect 12037 3163 12054 3180
rect 12197 3163 12214 3180
rect 11997 3163 12014 3180
rect 11957 3163 11974 3180
rect 12357 3163 12374 3180
rect 12317 3163 12334 3180
rect 12277 3163 12294 3180
rect 12317 3163 12334 3180
rect 12237 3163 12254 3180
rect 12077 3163 12094 3180
rect 11957 3163 11974 3180
rect 12357 3163 12374 3180
rect 12157 3163 12174 3180
rect 11997 3163 12014 3180
rect 11917 3163 11934 3180
rect 12037 3163 12054 3180
rect 12157 3163 12174 3180
rect 12117 3163 12134 3180
rect 11917 3163 11934 3180
rect 11957 3163 11974 3180
rect 12277 3163 12294 3180
rect 11917 3163 11934 3180
rect 12077 3163 12094 3180
rect 11877 3163 11894 3180
rect 11317 3163 11334 3180
rect 11397 3163 11414 3180
rect 11397 3163 11414 3180
rect 11637 3163 11654 3180
rect 11397 3163 11414 3180
rect 11717 3163 11734 3180
rect 11557 3163 11574 3180
rect 11637 3163 11654 3180
rect 11597 3163 11614 3180
rect 11477 3163 11494 3180
rect 11637 3163 11654 3180
rect 11757 3163 11774 3180
rect 11797 3163 11814 3180
rect 11557 3163 11574 3180
rect 11357 3163 11374 3180
rect 11437 3163 11454 3180
rect 11677 3163 11694 3180
rect 11397 3163 11414 3180
rect 11717 3163 11734 3180
rect 11517 3163 11534 3180
rect 11637 3163 11654 3180
rect 11357 3163 11374 3180
rect 11557 3163 11574 3180
rect 11677 3163 11694 3180
rect 11317 3163 11334 3180
rect 11797 3163 11814 3180
rect 11477 3163 11494 3180
rect 11437 3163 11454 3180
rect 11517 3163 11534 3180
rect 11437 3163 11454 3180
rect 11757 3163 11774 3180
rect 11437 3163 11454 3180
rect 11797 3163 11814 3180
rect 11477 3163 11494 3180
rect 11517 3163 11534 3180
rect 11317 3163 11334 3180
rect 11677 3163 11694 3180
rect 11757 3163 11774 3180
rect 11717 3163 11734 3180
rect 11597 3163 11614 3180
rect 11317 3163 11334 3180
rect 11357 3163 11374 3180
rect 11717 3163 11734 3180
rect 11797 3163 11814 3180
rect 11357 3163 11374 3180
rect 11517 3163 11534 3180
rect 11557 3163 11574 3180
rect 11597 3163 11614 3180
rect 11477 3163 11494 3180
rect 11597 3163 11614 3180
rect 11677 3163 11694 3180
rect 11757 3163 11774 3180
rect 10756 3163 10773 3180
rect 10756 3163 10773 3180
rect 10756 3163 10773 3180
rect 10756 3163 10773 3180
rect 11196 3163 11213 3180
rect 10836 3163 10853 3180
rect 10836 3163 10853 3180
rect 11036 3163 11053 3180
rect 10796 3163 10813 3180
rect 10836 3163 10853 3180
rect 11196 3163 11213 3180
rect 10836 3163 10853 3180
rect 11116 3163 11133 3180
rect 10996 3163 11013 3180
rect 11076 3163 11093 3180
rect 10956 3163 10973 3180
rect 11276 3163 11293 3180
rect 11236 3163 11253 3180
rect 11196 3163 11213 3180
rect 11276 3163 11293 3180
rect 11797 3163 11814 3180
rect 11797 3163 11814 3180
rect 11797 3163 11814 3180
rect 11797 3163 11814 3180
rect 14357 3163 14374 3180
rect 14317 3163 14334 3180
rect 14357 3163 14374 3180
rect 14277 3163 14294 3180
rect 14317 3163 14334 3180
rect 14237 3163 14254 3180
rect 14277 3163 14294 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14357 3163 14374 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14317 3163 14334 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14317 3163 14334 3180
rect 13837 3163 13854 3180
rect 13957 3163 13974 3180
rect 13917 3163 13934 3180
rect 13877 3163 13894 3180
rect 13837 3163 13854 3180
rect 13917 3163 13934 3180
rect 13917 3163 13934 3180
rect 13877 3163 13894 3180
rect 13837 3163 13854 3180
rect 13837 3163 13854 3180
rect 13957 3163 13974 3180
rect 13877 3163 13894 3180
rect 13957 3163 13974 3180
rect 13957 3163 13974 3180
rect 13917 3163 13934 3180
rect 13757 3163 13774 3180
rect 13877 3163 13894 3180
rect 13797 3163 13814 3180
rect 13717 3163 13734 3180
rect 13797 3163 13814 3180
rect 13797 3163 13814 3180
rect 13757 3163 13774 3180
rect 13757 3163 13774 3180
rect 13717 3163 13734 3180
rect 13717 3163 13734 3180
rect 13717 3163 13734 3180
rect 13757 3163 13774 3180
rect 13797 3163 13814 3180
rect 14277 3163 14294 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 13997 3163 14014 3180
rect 14237 3163 14254 3180
rect 14197 3163 14214 3180
rect 14157 3163 14174 3180
rect 14117 3163 14134 3180
rect 14077 3163 14094 3180
rect 14037 3163 14054 3180
rect 14357 3163 14374 3180
rect 13997 3163 14014 3180
rect 14277 3163 14294 3180
rect 12757 3163 12774 3180
rect 12757 3163 12774 3180
rect 12757 3163 12774 3180
rect 12757 3163 12774 3180
rect 12837 3163 12854 3180
rect 12837 3163 12854 3180
rect 12797 3163 12814 3180
rect 12797 3163 12814 3180
rect 13517 3163 13534 3180
rect 13597 3163 13614 3180
rect 13597 3163 13614 3180
rect 13677 3163 13694 3180
rect 13557 3163 13574 3180
rect 13637 3163 13654 3180
rect 12877 3163 12894 3180
rect 13477 3163 13494 3180
rect 13677 3163 13694 3180
rect 13637 3163 13654 3180
rect 13677 3163 13694 3180
rect 13597 3163 13614 3180
rect 13557 3163 13574 3180
rect 13517 3163 13534 3180
rect 13477 3163 13494 3180
rect 13557 3163 13574 3180
rect 13637 3163 13654 3180
rect 13677 3163 13694 3180
rect 13597 3163 13614 3180
rect 13637 3163 13654 3180
rect 13517 3163 13534 3180
rect 13557 3163 13574 3180
rect 13477 3163 13494 3180
rect 13517 3163 13534 3180
rect 13477 3163 13494 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 12917 3163 12934 3180
rect 13237 3163 13254 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13397 3163 13414 3180
rect 13037 3163 13054 3180
rect 13397 3163 13414 3180
rect 13197 3163 13214 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13357 3163 13374 3180
rect 13117 3163 13134 3180
rect 13437 3163 13454 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13037 3163 13054 3180
rect 13277 3163 13294 3180
rect 12997 3163 13014 3180
rect 13277 3163 13294 3180
rect 12957 3163 12974 3180
rect 13237 3163 13254 3180
rect 13197 3163 13214 3180
rect 13277 3163 13294 3180
rect 12957 3163 12974 3180
rect 13237 3163 13254 3180
rect 13077 3163 13094 3180
rect 13317 3163 13334 3180
rect 13157 3163 13174 3180
rect 13437 3163 13454 3180
rect 12997 3163 13014 3180
rect 13277 3163 13294 3180
rect 12997 3163 13014 3180
rect 13437 3163 13454 3180
rect 13197 3163 13214 3180
rect 13117 3163 13134 3180
rect 13117 3163 13134 3180
rect 13037 3163 13054 3180
rect 13037 3163 13054 3180
rect 12837 3163 12854 3180
rect 13117 3163 13134 3180
rect 12957 3163 12974 3180
rect 13197 3163 13214 3180
rect 13077 3163 13094 3180
rect 13157 3163 13174 3180
rect 12997 3163 13014 3180
rect 13397 3163 13414 3180
rect 13357 3163 13374 3180
rect 12797 3163 12814 3180
rect 13357 3163 13374 3180
rect 13357 3163 13374 3180
rect 13237 3163 13254 3180
rect 13437 3163 13454 3180
rect 12877 3163 12894 3180
rect 12957 3163 12974 3180
rect 13397 3163 13414 3180
rect 12877 3163 12894 3180
rect 12877 3163 12894 3180
rect 12797 3163 12814 3180
rect 12837 3163 12854 3180
rect 12197 3163 12214 3180
rect 12557 3163 12574 3180
rect 12477 3163 12494 3180
rect 11997 3163 12014 3180
rect 12437 3163 12454 3180
rect 11997 3163 12014 3180
rect 12237 3163 12254 3180
rect 12437 3163 12454 3180
rect 11957 3163 11974 3180
rect 11957 3163 11974 3180
rect 12597 3163 12614 3180
rect 12357 3163 12374 3180
rect 11837 3163 11854 3180
rect 12277 3163 12294 3180
rect 12317 3163 12334 3180
rect 12557 3163 12574 3180
rect 12277 3163 12294 3180
rect 11837 3163 11854 3180
rect 12197 3163 12214 3180
rect 12317 3163 12334 3180
rect 12557 3163 12574 3180
rect 12237 3163 12254 3180
rect 11837 3163 11854 3180
rect 12077 3163 12094 3180
rect 12677 3163 12694 3180
rect 11957 3163 11974 3180
rect 12397 3163 12414 3180
rect 11997 3163 12014 3180
rect 12397 3163 12414 3180
rect 12317 3163 12334 3180
rect 12117 3163 12134 3180
rect 12237 3163 12254 3180
rect 12197 3163 12214 3180
rect 11877 3163 11894 3180
rect 11997 3163 12014 3180
rect 12677 3163 12694 3180
rect 11837 3163 11854 3180
rect 11877 3163 11894 3180
rect 11917 3163 11934 3180
rect 12397 3163 12414 3180
rect 12277 3163 12294 3180
rect 12037 3163 12054 3180
rect 12037 3163 12054 3180
rect 12357 3163 12374 3180
rect 12717 3163 12734 3180
rect 12677 3163 12694 3180
rect 12157 3163 12174 3180
rect 12197 3163 12214 3180
rect 12117 3163 12134 3180
rect 12397 3163 12414 3180
rect 12117 3163 12134 3180
rect 12157 3163 12174 3180
rect 12717 3163 12734 3180
rect 12597 3163 12614 3180
rect 11917 3163 11934 3180
rect 12157 3163 12174 3180
rect 12237 3163 12254 3180
rect 12077 3163 12094 3180
rect 11957 3163 11974 3180
rect 12717 3163 12734 3180
rect 12117 3163 12134 3180
rect 12517 3163 12534 3180
rect 12277 3163 12294 3180
rect 12077 3163 12094 3180
rect 11917 3163 11934 3180
rect 12637 3163 12654 3180
rect 11917 3163 11934 3180
rect 12677 3163 12694 3180
rect 12557 3163 12574 3180
rect 12437 3163 12454 3180
rect 12077 3163 12094 3180
rect 12517 3163 12534 3180
rect 12037 3163 12054 3180
rect 12717 3163 12734 3180
rect 11877 3163 11894 3180
rect 12637 3163 12654 3180
rect 12477 3163 12494 3180
rect 12437 3163 12454 3180
rect 11877 3163 11894 3180
rect 12037 3163 12054 3180
rect 12477 3163 12494 3180
rect 12637 3163 12654 3180
rect 12357 3163 12374 3180
rect 12517 3163 12534 3180
rect 12597 3163 12614 3180
rect 12637 3163 12654 3180
rect 12157 3163 12174 3180
rect 12317 3163 12334 3180
rect 12517 3163 12534 3180
rect 12597 3163 12614 3180
rect 12357 3163 12374 3180
rect 12477 3163 12494 3180
rect 10836 3163 10853 3180
rect 10836 3163 10853 3180
rect 10836 3163 10853 3180
rect 10836 3163 10853 3180
rect 11757 3163 11774 3180
rect 11717 3163 11734 3180
rect 11597 3163 11614 3180
rect 11317 3163 11334 3180
rect 11357 3163 11374 3180
rect 11717 3163 11734 3180
rect 11357 3163 11374 3180
rect 11517 3163 11534 3180
rect 11557 3163 11574 3180
rect 11597 3163 11614 3180
rect 11477 3163 11494 3180
rect 11597 3163 11614 3180
rect 11677 3163 11694 3180
rect 11757 3163 11774 3180
rect 11196 3163 11213 3180
rect 11477 3163 11494 3180
rect 11517 3163 11534 3180
rect 11036 3163 11053 3180
rect 11317 3163 11334 3180
rect 11196 3163 11213 3180
rect 11677 3163 11694 3180
rect 11116 3163 11133 3180
rect 10996 3163 11013 3180
rect 11076 3163 11093 3180
rect 10956 3163 10973 3180
rect 11276 3163 11293 3180
rect 11236 3163 11253 3180
rect 11196 3163 11213 3180
rect 11276 3163 11293 3180
rect 11156 3163 11173 3180
rect 11116 3163 11133 3180
rect 11076 3163 11093 3180
rect 11036 3163 11053 3180
rect 10996 3163 11013 3180
rect 10956 3163 10973 3180
rect 10916 3163 10933 3180
rect 10876 3163 10893 3180
rect 11116 3163 11133 3180
rect 11076 3163 11093 3180
rect 11036 3163 11053 3180
rect 11076 3163 11093 3180
rect 10956 3163 10973 3180
rect 11276 3163 11293 3180
rect 11276 3163 11293 3180
rect 11156 3163 11173 3180
rect 11156 3163 11173 3180
rect 10916 3163 10933 3180
rect 10876 3163 10893 3180
rect 11317 3163 11334 3180
rect 10996 3163 11013 3180
rect 11196 3163 11213 3180
rect 11116 3163 11133 3180
rect 11397 3163 11414 3180
rect 11036 3163 11053 3180
rect 10956 3163 10973 3180
rect 10876 3163 10893 3180
rect 11397 3163 11414 3180
rect 10996 3163 11013 3180
rect 11236 3163 11253 3180
rect 11236 3163 11253 3180
rect 11637 3163 11654 3180
rect 10916 3163 10933 3180
rect 10916 3163 10933 3180
rect 11397 3163 11414 3180
rect 11236 3163 11253 3180
rect 10876 3163 10893 3180
rect 11156 3163 11173 3180
rect 11717 3163 11734 3180
rect 11557 3163 11574 3180
rect 11637 3163 11654 3180
rect 11597 3163 11614 3180
rect 11477 3163 11494 3180
rect 11637 3163 11654 3180
rect 11757 3163 11774 3180
rect 11557 3163 11574 3180
rect 11357 3163 11374 3180
rect 11437 3163 11454 3180
rect 11677 3163 11694 3180
rect 11397 3163 11414 3180
rect 11717 3163 11734 3180
rect 11517 3163 11534 3180
rect 11637 3163 11654 3180
rect 11357 3163 11374 3180
rect 11557 3163 11574 3180
rect 11677 3163 11694 3180
rect 11317 3163 11334 3180
rect 11477 3163 11494 3180
rect 11437 3163 11454 3180
rect 11517 3163 11534 3180
rect 11437 3163 11454 3180
rect 11757 3163 11774 3180
rect 11437 3163 11454 3180
rect 10196 3163 10213 3180
rect 9916 3163 9933 3180
rect 10756 3163 10773 3180
rect 10676 3163 10693 3180
rect 10236 3163 10253 3180
rect 9956 3163 9973 3180
rect 10276 3163 10293 3180
rect 9996 3163 10013 3180
rect 10476 3163 10493 3180
rect 10436 3163 10453 3180
rect 10116 3163 10133 3180
rect 10316 3163 10333 3180
rect 9956 3163 9973 3180
rect 10556 3163 10573 3180
rect 10396 3163 10413 3180
rect 10716 3163 10733 3180
rect 10116 3163 10133 3180
rect 10716 3163 10733 3180
rect 10516 3163 10533 3180
rect 10156 3163 10173 3180
rect 10716 3163 10733 3180
rect 10756 3163 10773 3180
rect 10476 3163 10493 3180
rect 10356 3163 10373 3180
rect 10556 3163 10573 3180
rect 10756 3163 10773 3180
rect 10316 3163 10333 3180
rect 10436 3163 10453 3180
rect 10396 3163 10413 3180
rect 10196 3163 10213 3180
rect 10436 3163 10453 3180
rect 10356 3163 10373 3180
rect 9916 3163 9933 3180
rect 10236 3163 10253 3180
rect 10116 3163 10133 3180
rect 10596 3163 10613 3180
rect 10676 3163 10693 3180
rect 10396 3163 10413 3180
rect 10796 3163 10813 3180
rect 10276 3163 10293 3180
rect 10076 3163 10093 3180
rect 10276 3163 10293 3180
rect 10156 3163 10173 3180
rect 10636 3163 10653 3180
rect 9956 3163 9973 3180
rect 10396 3163 10413 3180
rect 10156 3163 10173 3180
rect 10556 3163 10573 3180
rect 10036 3163 10053 3180
rect 10516 3163 10533 3180
rect 10076 3163 10093 3180
rect 10636 3163 10653 3180
rect 10116 3163 10133 3180
rect 10676 3163 10693 3180
rect 10236 3163 10253 3180
rect 10196 3163 10213 3180
rect 10516 3163 10533 3180
rect 10796 3163 10813 3180
rect 10676 3163 10693 3180
rect 10036 3163 10053 3180
rect 10716 3163 10733 3180
rect 9916 3163 9933 3180
rect 10596 3163 10613 3180
rect 10196 3163 10213 3180
rect 10516 3163 10533 3180
rect 9916 3163 9933 3180
rect 10636 3163 10653 3180
rect 9996 3163 10013 3180
rect 10276 3163 10293 3180
rect 9996 3163 10013 3180
rect 10036 3163 10053 3180
rect 10316 3163 10333 3180
rect 10476 3163 10493 3180
rect 10076 3163 10093 3180
rect 10436 3163 10453 3180
rect 10036 3163 10053 3180
rect 9996 3163 10013 3180
rect 10636 3163 10653 3180
rect 10476 3163 10493 3180
rect 10796 3163 10813 3180
rect 10316 3163 10333 3180
rect 10156 3163 10173 3180
rect 10356 3163 10373 3180
rect 10596 3163 10613 3180
rect 10796 3163 10813 3180
rect 10356 3163 10373 3180
rect 10076 3163 10093 3180
rect 10596 3163 10613 3180
rect 10556 3163 10573 3180
rect 10756 3163 10773 3180
rect 10236 3163 10253 3180
rect 9956 3163 9973 3180
rect 12001 2394 12018 2411
rect 12001 2394 12018 2411
rect 9876 3163 9893 3180
rect 9836 3163 9853 3180
rect 9636 3163 9653 3180
rect 9836 3163 9853 3180
rect 9876 3163 9893 3180
rect 9636 3163 9653 3180
rect 9636 3163 9653 3180
rect 9676 3163 9693 3180
rect 9716 3163 9733 3180
rect 9676 3163 9693 3180
rect 9756 3163 9773 3180
rect 9836 3163 9853 3180
rect 9636 3163 9653 3180
rect 9716 3163 9733 3180
rect 9756 3163 9773 3180
rect 9756 3163 9773 3180
rect 9796 3163 9813 3180
rect 9796 3163 9813 3180
rect 9716 3163 9733 3180
rect 9756 3163 9773 3180
rect 9796 3163 9813 3180
rect 9716 3163 9733 3180
rect 9876 3163 9893 3180
rect 9836 3163 9853 3180
rect 9796 3163 9813 3180
rect 9876 3163 9893 3180
rect 9676 3163 9693 3180
rect 9676 3163 9693 3180
rect 11156 3163 11173 3180
rect 10041 2394 10058 2411
rect 10721 2394 10738 2411
rect 10601 2394 10618 2411
rect 9801 2394 9818 2411
rect 9881 2394 9898 2411
rect 10521 2394 10538 2411
rect 10721 2394 10738 2411
rect 10201 2394 10218 2411
rect 10201 2394 10218 2411
rect 9681 2394 9698 2411
rect 9641 2394 9658 2411
rect 10441 2394 10458 2411
rect 10281 2394 10298 2411
rect 10241 2394 10258 2411
rect 10561 2394 10578 2411
rect 10121 2394 10138 2411
rect 10641 2394 10658 2411
rect 9641 2394 9658 2411
rect 10001 2394 10018 2411
rect 10281 2394 10298 2411
rect 9681 2394 9698 2411
rect 9841 2394 9858 2411
rect 10681 2394 10698 2411
rect 10081 2394 10098 2411
rect 10761 2394 10778 2411
rect 10601 2394 10618 2411
rect 9841 2394 9858 2411
rect 9801 2394 9818 2411
rect 10801 2394 10818 2411
rect 10761 2394 10778 2411
rect 10161 2394 10178 2411
rect 9721 2394 9738 2411
rect 10481 2394 10498 2411
rect 10321 2394 10338 2411
rect 9761 2394 9778 2411
rect 10081 2394 10098 2411
rect 10001 2394 10018 2411
rect 10481 2394 10498 2411
rect 10441 2394 10458 2411
rect 9721 2394 9738 2411
rect 10041 2394 10058 2411
rect 9921 2394 9938 2411
rect 9961 2394 9978 2411
rect 10241 2394 10258 2411
rect 10361 2394 10378 2411
rect 9961 2394 9978 2411
rect 9761 2394 9778 2411
rect 9881 2394 9898 2411
rect 10401 2394 10418 2411
rect 10361 2394 10378 2411
rect 10121 2394 10138 2411
rect 10521 2394 10538 2411
rect 9921 2394 9938 2411
rect 10401 2394 10418 2411
rect 10801 2394 10818 2411
rect 10561 2394 10578 2411
rect 10681 2394 10698 2411
rect 10321 2394 10338 2411
rect 10161 2394 10178 2411
rect 10641 2394 10658 2411
rect 11881 2394 11898 2411
rect 11601 2394 11618 2411
rect 11961 2394 11978 2411
rect 11041 2394 11058 2411
rect 11161 2394 11178 2411
rect 11561 2394 11578 2411
rect 11081 2394 11098 2411
rect 11001 2394 11018 2411
rect 11321 2394 11338 2411
rect 11041 2394 11058 2411
rect 11881 2394 11898 2411
rect 11721 2394 11738 2411
rect 11841 2394 11858 2411
rect 11841 2394 11858 2411
rect 11921 2394 11938 2411
rect 11801 2394 11818 2411
rect 11961 2394 11978 2411
rect 11201 2394 11218 2411
rect 11761 2394 11778 2411
rect 10961 2394 10978 2411
rect 11801 2394 11818 2411
rect 11641 2394 11658 2411
rect 11641 2394 11658 2411
rect 11721 2394 11738 2411
rect 11481 2394 11498 2411
rect 11161 2394 11178 2411
rect 10921 2394 10938 2411
rect 11681 2394 11698 2411
rect 11601 2394 11618 2411
rect 11681 2394 11698 2411
rect 10961 2394 10978 2411
rect 11761 2394 11778 2411
rect 11441 2394 11458 2411
rect 11561 2394 11578 2411
rect 11281 2394 11298 2411
rect 11521 2394 11538 2411
rect 10841 2394 10858 2411
rect 11401 2394 11418 2411
rect 11481 2394 11498 2411
rect 10921 2394 10938 2411
rect 11441 2394 11458 2411
rect 11121 2394 11138 2411
rect 11001 2394 11018 2411
rect 11401 2394 11418 2411
rect 11361 2394 11378 2411
rect 10881 2394 10898 2411
rect 11361 2394 11378 2411
rect 11521 2394 11538 2411
rect 11321 2394 11338 2411
rect 11281 2394 11298 2411
rect 11241 2394 11258 2411
rect 11921 2394 11938 2411
rect 11241 2394 11258 2411
rect 10841 2394 10858 2411
rect 11201 2394 11218 2411
rect 11081 2394 11098 2411
rect 10881 2394 10898 2411
rect 11121 2394 11138 2411
rect 13201 2394 13218 2411
rect 13201 2394 13218 2411
rect 12321 2394 12338 2411
rect 12241 2394 12258 2411
rect 12201 2394 12218 2411
rect 12081 2394 12098 2411
rect 12281 2394 12298 2411
rect 12281 2394 12298 2411
rect 12041 2394 12058 2411
rect 12041 2394 12058 2411
rect 12321 2394 12338 2411
rect 12521 2394 12538 2411
rect 12561 2394 12578 2411
rect 12161 2394 12178 2411
rect 12161 2394 12178 2411
rect 12081 2394 12098 2411
rect 12121 2394 12138 2411
rect 12401 2394 12418 2411
rect 12601 2394 12618 2411
rect 13121 2394 13138 2411
rect 13081 2394 13098 2411
rect 13041 2394 13058 2411
rect 13001 2394 13018 2411
rect 12961 2394 12978 2411
rect 12921 2394 12938 2411
rect 12881 2394 12898 2411
rect 12841 2394 12858 2411
rect 12801 2394 12818 2411
rect 12761 2394 12778 2411
rect 12721 2394 12738 2411
rect 12401 2394 12418 2411
rect 13161 2394 13178 2411
rect 13121 2394 13138 2411
rect 13081 2394 13098 2411
rect 13041 2394 13058 2411
rect 13001 2394 13018 2411
rect 12961 2394 12978 2411
rect 12921 2394 12938 2411
rect 12881 2394 12898 2411
rect 12841 2394 12858 2411
rect 12801 2394 12818 2411
rect 12761 2394 12778 2411
rect 12721 2394 12738 2411
rect 12681 2394 12698 2411
rect 13161 2394 13178 2411
rect 12361 2394 12378 2411
rect 12481 2394 12498 2411
rect 12681 2394 12698 2411
rect 12641 2394 12658 2411
rect 12601 2394 12618 2411
rect 12561 2394 12578 2411
rect 12521 2394 12538 2411
rect 12481 2394 12498 2411
rect 12241 2394 12258 2411
rect 12441 2394 12458 2411
rect 12441 2394 12458 2411
rect 12121 2394 12138 2411
rect 12641 2394 12658 2411
rect 12201 2394 12218 2411
rect 12361 2394 12378 2411
rect 14242 2394 14259 2411
rect 13802 2394 13819 2411
rect 14202 2394 14219 2411
rect 14322 2394 14339 2411
rect 14002 2394 14019 2411
rect 14242 2394 14259 2411
rect 13962 2394 13979 2411
rect 13842 2394 13859 2411
rect 13761 2394 13778 2411
rect 13641 2394 13658 2411
rect 14202 2394 14219 2411
rect 13721 2394 13738 2411
rect 14162 2394 14179 2411
rect 13601 2394 13618 2411
rect 13882 2394 13899 2411
rect 13561 2394 13578 2411
rect 13521 2394 13538 2411
rect 13481 2394 13498 2411
rect 13441 2394 13458 2411
rect 14042 2394 14059 2411
rect 14082 2394 14099 2411
rect 13401 2394 13418 2411
rect 13361 2394 13378 2411
rect 13321 2394 13338 2411
rect 14362 2394 14379 2411
rect 13842 2394 13859 2411
rect 13882 2394 13899 2411
rect 14002 2394 14019 2411
rect 13802 2394 13819 2411
rect 14362 2394 14379 2411
rect 14122 2394 14139 2411
rect 14322 2394 14339 2411
rect 13922 2394 13939 2411
rect 14282 2394 14299 2411
rect 13962 2394 13979 2411
rect 14122 2394 14139 2411
rect 13922 2394 13939 2411
rect 14082 2394 14099 2411
rect 14042 2394 14059 2411
rect 13641 2394 13658 2411
rect 13601 2394 13618 2411
rect 14162 2394 14179 2411
rect 13681 2394 13698 2411
rect 13561 2394 13578 2411
rect 13521 2394 13538 2411
rect 14282 2394 14299 2411
rect 13721 2394 13738 2411
rect 13681 2394 13698 2411
rect 13281 2394 13298 2411
rect 13241 2394 13258 2411
rect 13481 2394 13498 2411
rect 13441 2394 13458 2411
rect 13401 2394 13418 2411
rect 13361 2394 13378 2411
rect 13321 2394 13338 2411
rect 13761 2394 13778 2411
rect 13281 2394 13298 2411
rect 13241 2394 13258 2411
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 15077 3163 15094 3180
rect 15117 3163 15134 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 14717 3163 14734 3180
rect 14997 3163 15014 3180
rect 14797 3163 14814 3180
rect 14997 3163 15014 3180
rect 14677 3163 14694 3180
rect 14957 3163 14974 3180
rect 14877 3163 14894 3180
rect 14997 3163 15014 3180
rect 14917 3163 14934 3180
rect 14917 3163 14934 3180
rect 14957 3163 14974 3180
rect 14917 3163 14934 3180
rect 14877 3163 14894 3180
rect 14877 3163 14894 3180
rect 14837 3163 14854 3180
rect 14837 3163 14854 3180
rect 14837 3163 14854 3180
rect 15037 3163 15054 3180
rect 14797 3163 14814 3180
rect 14797 3163 14814 3180
rect 14917 3163 14934 3180
rect 14757 3163 14774 3180
rect 14757 3163 14774 3180
rect 14757 3163 14774 3180
rect 15037 3163 15054 3180
rect 14717 3163 14734 3180
rect 14717 3163 14734 3180
rect 14877 3163 14894 3180
rect 15037 3163 15054 3180
rect 14677 3163 14694 3180
rect 14677 3163 14694 3180
rect 15037 3163 15054 3180
rect 14957 3163 14974 3180
rect 14837 3163 14854 3180
rect 14677 3163 14694 3180
rect 14797 3163 14814 3180
rect 14717 3163 14734 3180
rect 14997 3163 15014 3180
rect 14957 3163 14974 3180
rect 14757 3163 14774 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 15077 3163 15094 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 15077 3163 15094 3180
rect 15077 3163 15094 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15077 3163 15094 3180
rect 14397 3163 14414 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 14557 3163 14574 3180
rect 14397 3163 14414 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 14477 3163 14494 3180
rect 14437 3163 14454 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 14517 3163 14534 3180
rect 14477 3163 14494 3180
rect 14437 3163 14454 3180
rect 15077 3163 15094 3180
rect 15077 3163 15094 3180
rect 15517 3163 15534 3180
rect 14517 3163 14534 3180
rect 15477 3163 15494 3180
rect 14477 3163 14494 3180
rect 14517 3163 14534 3180
rect 14477 3163 14494 3180
rect 14597 3163 14614 3180
rect 14437 3163 14454 3180
rect 14517 3163 14534 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15077 3163 15094 3180
rect 15117 3163 15134 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15597 3163 15614 3180
rect 15557 3163 15574 3180
rect 15517 3163 15534 3180
rect 15477 3163 15494 3180
rect 15437 3163 15454 3180
rect 15397 3163 15414 3180
rect 15357 3163 15374 3180
rect 15317 3163 15334 3180
rect 15277 3163 15294 3180
rect 15237 3163 15254 3180
rect 15197 3163 15214 3180
rect 15157 3163 15174 3180
rect 15117 3163 15134 3180
rect 14717 3163 14734 3180
rect 14637 3163 14654 3180
rect 14637 3163 14654 3180
rect 14637 3163 14654 3180
rect 14597 3163 14614 3180
rect 14557 3163 14574 3180
rect 14637 3163 14654 3180
rect 14557 3163 14574 3180
rect 14557 3163 14574 3180
rect 14597 3163 14614 3180
rect 14597 3163 14614 3180
rect 14997 3163 15014 3180
rect 14797 3163 14814 3180
rect 14437 3163 14454 3180
rect 14997 3163 15014 3180
rect 14677 3163 14694 3180
rect 14957 3163 14974 3180
rect 14877 3163 14894 3180
rect 14997 3163 15014 3180
rect 14557 3163 14574 3180
rect 14917 3163 14934 3180
rect 14917 3163 14934 3180
rect 14957 3163 14974 3180
rect 14917 3163 14934 3180
rect 14877 3163 14894 3180
rect 14397 3163 14414 3180
rect 14877 3163 14894 3180
rect 14597 3163 14614 3180
rect 14837 3163 14854 3180
rect 14837 3163 14854 3180
rect 14397 3163 14414 3180
rect 14837 3163 14854 3180
rect 14557 3163 14574 3180
rect 15037 3163 15054 3180
rect 14797 3163 14814 3180
rect 14797 3163 14814 3180
rect 14917 3163 14934 3180
rect 14757 3163 14774 3180
rect 14757 3163 14774 3180
rect 14757 3163 14774 3180
rect 14637 3163 14654 3180
rect 15037 3163 15054 3180
rect 14717 3163 14734 3180
rect 14717 3163 14734 3180
rect 14877 3163 14894 3180
rect 15037 3163 15054 3180
rect 14677 3163 14694 3180
rect 14677 3163 14694 3180
rect 15037 3163 15054 3180
rect 14637 3163 14654 3180
rect 14957 3163 14974 3180
rect 14837 3163 14854 3180
rect 14597 3163 14614 3180
rect 14557 3163 14574 3180
rect 14677 3163 14694 3180
rect 14797 3163 14814 3180
rect 14717 3163 14734 3180
rect 14637 3163 14654 3180
rect 14597 3163 14614 3180
rect 14557 3163 14574 3180
rect 14637 3163 14654 3180
rect 14997 3163 15014 3180
rect 14957 3163 14974 3180
rect 14757 3163 14774 3180
rect 14597 3163 14614 3180
rect 16762 2394 16779 2411
rect 16762 2394 16779 2411
rect 14437 3163 14454 3180
rect 14397 3163 14414 3180
rect 14397 3163 14414 3180
rect 14397 3163 14414 3180
rect 14397 3163 14414 3180
rect 14477 3163 14494 3180
rect 14437 3163 14454 3180
rect 14517 3163 14534 3180
rect 14477 3163 14494 3180
rect 14437 3163 14454 3180
rect 14517 3163 14534 3180
rect 14477 3163 14494 3180
rect 14517 3163 14534 3180
rect 14477 3163 14494 3180
rect 14437 3163 14454 3180
rect 14517 3163 14534 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 17757 3163 17774 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 16637 3163 16654 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17197 3163 17214 3180
rect 17477 3163 17494 3180
rect 17717 3163 17734 3180
rect 17717 3163 17734 3180
rect 17517 3163 17534 3180
rect 17637 3163 17654 3180
rect 17477 3163 17494 3180
rect 17677 3163 17694 3180
rect 17637 3163 17654 3180
rect 17597 3163 17614 3180
rect 17597 3163 17614 3180
rect 17557 3163 17574 3180
rect 17517 3163 17534 3180
rect 17597 3163 17614 3180
rect 17557 3163 17574 3180
rect 17637 3163 17654 3180
rect 17477 3163 17494 3180
rect 17597 3163 17614 3180
rect 17517 3163 17534 3180
rect 17517 3163 17534 3180
rect 17477 3163 17494 3180
rect 17717 3163 17734 3180
rect 17677 3163 17694 3180
rect 17677 3163 17694 3180
rect 17677 3163 17694 3180
rect 17557 3163 17574 3180
rect 17557 3163 17574 3180
rect 17637 3163 17654 3180
rect 17477 3163 17494 3180
rect 17717 3163 17734 3180
rect 17717 3163 17734 3180
rect 17557 3163 17574 3180
rect 17717 3163 17734 3180
rect 17517 3163 17534 3180
rect 17637 3163 17654 3180
rect 17477 3163 17494 3180
rect 17677 3163 17694 3180
rect 17637 3163 17654 3180
rect 17597 3163 17614 3180
rect 17597 3163 17614 3180
rect 17557 3163 17574 3180
rect 17517 3163 17534 3180
rect 17597 3163 17614 3180
rect 17557 3163 17574 3180
rect 17637 3163 17654 3180
rect 17477 3163 17494 3180
rect 17597 3163 17614 3180
rect 17517 3163 17534 3180
rect 17517 3163 17534 3180
rect 17477 3163 17494 3180
rect 17717 3163 17734 3180
rect 17677 3163 17694 3180
rect 17677 3163 17694 3180
rect 17677 3163 17694 3180
rect 17557 3163 17574 3180
rect 17717 3163 17734 3180
rect 17637 3163 17654 3180
rect 17357 3163 17374 3180
rect 17237 3163 17254 3180
rect 17357 3163 17374 3180
rect 17437 3163 17454 3180
rect 17437 3163 17454 3180
rect 17357 3163 17374 3180
rect 17357 3163 17374 3180
rect 17437 3163 17454 3180
rect 17277 3163 17294 3180
rect 17437 3163 17454 3180
rect 17397 3163 17414 3180
rect 17437 3163 17454 3180
rect 17357 3163 17374 3180
rect 17397 3163 17414 3180
rect 17317 3163 17334 3180
rect 17277 3163 17294 3180
rect 17277 3163 17294 3180
rect 17317 3163 17334 3180
rect 17317 3163 17334 3180
rect 17397 3163 17414 3180
rect 17277 3163 17294 3180
rect 17237 3163 17254 3180
rect 17397 3163 17414 3180
rect 17237 3163 17254 3180
rect 17237 3163 17254 3180
rect 17317 3163 17334 3180
rect 17237 3163 17254 3180
rect 17317 3163 17334 3180
rect 17397 3163 17414 3180
rect 17437 3163 17454 3180
rect 17437 3163 17454 3180
rect 17357 3163 17374 3180
rect 17357 3163 17374 3180
rect 17437 3163 17454 3180
rect 17277 3163 17294 3180
rect 17237 3163 17254 3180
rect 17397 3163 17414 3180
rect 17277 3163 17294 3180
rect 17317 3163 17334 3180
rect 17317 3163 17334 3180
rect 17397 3163 17414 3180
rect 17237 3163 17254 3180
rect 17357 3163 17374 3180
rect 17277 3163 17294 3180
rect 17277 3163 17294 3180
rect 17237 3163 17254 3180
rect 17397 3163 17414 3180
rect 17317 3163 17334 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 16917 3163 16934 3180
rect 17117 3163 17134 3180
rect 17037 3163 17054 3180
rect 17117 3163 17134 3180
rect 17117 3163 17134 3180
rect 16997 3163 17014 3180
rect 17037 3163 17054 3180
rect 17077 3163 17094 3180
rect 17077 3163 17094 3180
rect 16957 3163 16974 3180
rect 16997 3163 17014 3180
rect 16957 3163 16974 3180
rect 17077 3163 17094 3180
rect 17157 3163 17174 3180
rect 17077 3163 17094 3180
rect 17037 3163 17054 3180
rect 17077 3163 17094 3180
rect 17157 3163 17174 3180
rect 17157 3163 17174 3180
rect 17157 3163 17174 3180
rect 17117 3163 17134 3180
rect 17157 3163 17174 3180
rect 16997 3163 17014 3180
rect 17117 3163 17134 3180
rect 16997 3163 17014 3180
rect 17117 3163 17134 3180
rect 16957 3163 16974 3180
rect 17077 3163 17094 3180
rect 17117 3163 17134 3180
rect 17037 3163 17054 3180
rect 16957 3163 16974 3180
rect 17157 3163 17174 3180
rect 17037 3163 17054 3180
rect 16957 3163 16974 3180
rect 17037 3163 17054 3180
rect 16997 3163 17014 3180
rect 16997 3163 17014 3180
rect 16997 3163 17014 3180
rect 17157 3163 17174 3180
rect 17077 3163 17094 3180
rect 16957 3163 16974 3180
rect 17077 3163 17094 3180
rect 17037 3163 17054 3180
rect 16957 3163 16974 3180
rect 17037 3163 17054 3180
rect 16997 3163 17014 3180
rect 16957 3163 16974 3180
rect 17117 3163 17134 3180
rect 17157 3163 17174 3180
rect 16877 3163 16894 3180
rect 16677 3163 16694 3180
rect 16757 3163 16774 3180
rect 16677 3163 16694 3180
rect 16797 3163 16814 3180
rect 16837 3163 16854 3180
rect 16877 3163 16894 3180
rect 16877 3163 16894 3180
rect 16757 3163 16774 3180
rect 16877 3163 16894 3180
rect 16877 3163 16894 3180
rect 16837 3163 16854 3180
rect 16797 3163 16814 3180
rect 16837 3163 16854 3180
rect 16877 3163 16894 3180
rect 16717 3163 16734 3180
rect 16837 3163 16854 3180
rect 16837 3163 16854 3180
rect 16717 3163 16734 3180
rect 16797 3163 16814 3180
rect 16757 3163 16774 3180
rect 16757 3163 16774 3180
rect 16677 3163 16694 3180
rect 16677 3163 16694 3180
rect 16757 3163 16774 3180
rect 16797 3163 16814 3180
rect 16677 3163 16694 3180
rect 16677 3163 16694 3180
rect 16877 3163 16894 3180
rect 16757 3163 16774 3180
rect 16837 3163 16854 3180
rect 16717 3163 16734 3180
rect 16837 3163 16854 3180
rect 16877 3163 16894 3180
rect 16717 3163 16734 3180
rect 16757 3163 16774 3180
rect 16717 3163 16734 3180
rect 16677 3163 16694 3180
rect 16797 3163 16814 3180
rect 16717 3163 16734 3180
rect 16797 3163 16814 3180
rect 16837 3163 16854 3180
rect 16797 3163 16814 3180
rect 16757 3163 16774 3180
rect 16717 3163 16734 3180
rect 16677 3163 16694 3180
rect 16717 3163 16734 3180
rect 16797 3163 16814 3180
rect 16597 3163 16614 3180
rect 16437 3163 16454 3180
rect 16517 3163 16534 3180
rect 16557 3163 16574 3180
rect 16397 3163 16414 3180
rect 16557 3163 16574 3180
rect 16477 3163 16494 3180
rect 16397 3163 16414 3180
rect 16597 3163 16614 3180
rect 16397 3163 16414 3180
rect 16597 3163 16614 3180
rect 16477 3163 16494 3180
rect 16517 3163 16534 3180
rect 16517 3163 16534 3180
rect 16557 3163 16574 3180
rect 16397 3163 16414 3180
rect 16597 3163 16614 3180
rect 16437 3163 16454 3180
rect 16477 3163 16494 3180
rect 16437 3163 16454 3180
rect 16517 3163 16534 3180
rect 16437 3163 16454 3180
rect 16437 3163 16454 3180
rect 16557 3163 16574 3180
rect 16557 3163 16574 3180
rect 16517 3163 16534 3180
rect 16437 3163 16454 3180
rect 16397 3163 16414 3180
rect 16597 3163 16614 3180
rect 16557 3163 16574 3180
rect 16597 3163 16614 3180
rect 16517 3163 16534 3180
rect 16397 3163 16414 3180
rect 16597 3163 16614 3180
rect 16477 3163 16494 3180
rect 16477 3163 16494 3180
rect 16517 3163 16534 3180
rect 16437 3163 16454 3180
rect 16557 3163 16574 3180
rect 16477 3163 16494 3180
rect 16437 3163 16454 3180
rect 16477 3163 16494 3180
rect 16597 3163 16614 3180
rect 16397 3163 16414 3180
rect 16477 3163 16494 3180
rect 16557 3163 16574 3180
rect 16517 3163 16534 3180
rect 16397 3163 16414 3180
rect 16317 3163 16334 3180
rect 16197 3163 16214 3180
rect 16357 3163 16374 3180
rect 16277 3163 16294 3180
rect 16277 3163 16294 3180
rect 16117 3163 16134 3180
rect 16157 3163 16174 3180
rect 16237 3163 16254 3180
rect 16157 3163 16174 3180
rect 16117 3163 16134 3180
rect 16197 3163 16214 3180
rect 16197 3163 16214 3180
rect 16317 3163 16334 3180
rect 16277 3163 16294 3180
rect 16237 3163 16254 3180
rect 16157 3163 16174 3180
rect 16157 3163 16174 3180
rect 16197 3163 16214 3180
rect 16157 3163 16174 3180
rect 16357 3163 16374 3180
rect 16237 3163 16254 3180
rect 16237 3163 16254 3180
rect 16317 3163 16334 3180
rect 16157 3163 16174 3180
rect 16357 3163 16374 3180
rect 16237 3163 16254 3180
rect 16357 3163 16374 3180
rect 16317 3163 16334 3180
rect 16277 3163 16294 3180
rect 16317 3163 16334 3180
rect 16117 3163 16134 3180
rect 16317 3163 16334 3180
rect 16357 3163 16374 3180
rect 16117 3163 16134 3180
rect 16117 3163 16134 3180
rect 16317 3163 16334 3180
rect 16117 3163 16134 3180
rect 16157 3163 16174 3180
rect 16237 3163 16254 3180
rect 16157 3163 16174 3180
rect 16197 3163 16214 3180
rect 16117 3163 16134 3180
rect 16277 3163 16294 3180
rect 16277 3163 16294 3180
rect 16357 3163 16374 3180
rect 16197 3163 16214 3180
rect 16357 3163 16374 3180
rect 16277 3163 16294 3180
rect 16197 3163 16214 3180
rect 16237 3163 16254 3180
rect 16237 3163 16254 3180
rect 16357 3163 16374 3180
rect 16117 3163 16134 3180
rect 16197 3163 16214 3180
rect 16317 3163 16334 3180
rect 16277 3163 16294 3180
rect 16037 3163 16054 3180
rect 15997 3163 16014 3180
rect 15957 3163 15974 3180
rect 15997 3163 16014 3180
rect 15877 3163 15894 3180
rect 15837 3163 15854 3180
rect 15877 3163 15894 3180
rect 15877 3163 15894 3180
rect 15837 3163 15854 3180
rect 15957 3163 15974 3180
rect 16077 3163 16094 3180
rect 15837 3163 15854 3180
rect 15917 3163 15934 3180
rect 15917 3163 15934 3180
rect 16037 3163 16054 3180
rect 15877 3163 15894 3180
rect 15957 3163 15974 3180
rect 15997 3163 16014 3180
rect 16037 3163 16054 3180
rect 16077 3163 16094 3180
rect 15957 3163 15974 3180
rect 16077 3163 16094 3180
rect 15837 3163 15854 3180
rect 15997 3163 16014 3180
rect 16077 3163 16094 3180
rect 15877 3163 15894 3180
rect 16037 3163 16054 3180
rect 15877 3163 15894 3180
rect 15917 3163 15934 3180
rect 15837 3163 15854 3180
rect 15917 3163 15934 3180
rect 15997 3163 16014 3180
rect 15837 3163 15854 3180
rect 15957 3163 15974 3180
rect 16077 3163 16094 3180
rect 15877 3163 15894 3180
rect 15837 3163 15854 3180
rect 15997 3163 16014 3180
rect 15957 3163 15974 3180
rect 15917 3163 15934 3180
rect 15877 3163 15894 3180
rect 16037 3163 16054 3180
rect 15917 3163 15934 3180
rect 16037 3163 16054 3180
rect 15997 3163 16014 3180
rect 15957 3163 15974 3180
rect 16077 3163 16094 3180
rect 16037 3163 16054 3180
rect 15917 3163 15934 3180
rect 15997 3163 16014 3180
rect 15837 3163 15854 3180
rect 16077 3163 16094 3180
rect 16077 3163 16094 3180
rect 15917 3163 15934 3180
rect 16037 3163 16054 3180
rect 15957 3163 15974 3180
rect 15757 3163 15774 3180
rect 15557 3163 15574 3180
rect 15637 3163 15654 3180
rect 15557 3163 15574 3180
rect 15717 3163 15734 3180
rect 15797 3163 15814 3180
rect 15677 3163 15694 3180
rect 15757 3163 15774 3180
rect 15717 3163 15734 3180
rect 15797 3163 15814 3180
rect 15557 3163 15574 3180
rect 15557 3163 15574 3180
rect 15637 3163 15654 3180
rect 15597 3163 15614 3180
rect 15757 3163 15774 3180
rect 15557 3163 15574 3180
rect 15797 3163 15814 3180
rect 15797 3163 15814 3180
rect 15677 3163 15694 3180
rect 15637 3163 15654 3180
rect 15597 3163 15614 3180
rect 15757 3163 15774 3180
rect 15797 3163 15814 3180
rect 15717 3163 15734 3180
rect 15677 3163 15694 3180
rect 15717 3163 15734 3180
rect 15677 3163 15694 3180
rect 15597 3163 15614 3180
rect 15597 3163 15614 3180
rect 15797 3163 15814 3180
rect 15717 3163 15734 3180
rect 15757 3163 15774 3180
rect 15757 3163 15774 3180
rect 15677 3163 15694 3180
rect 15717 3163 15734 3180
rect 15637 3163 15654 3180
rect 15757 3163 15774 3180
rect 15677 3163 15694 3180
rect 15717 3163 15734 3180
rect 15557 3163 15574 3180
rect 15797 3163 15814 3180
rect 15597 3163 15614 3180
rect 15637 3163 15654 3180
rect 15557 3163 15574 3180
rect 15597 3163 15614 3180
rect 15637 3163 15654 3180
rect 15797 3163 15814 3180
rect 15637 3163 15654 3180
rect 15677 3163 15694 3180
rect 15557 3163 15574 3180
rect 15637 3163 15654 3180
rect 15597 3163 15614 3180
rect 15597 3163 15614 3180
rect 15717 3163 15734 3180
rect 15757 3163 15774 3180
rect 15677 3163 15694 3180
rect 15317 3163 15334 3180
rect 14522 2394 14539 2411
rect 15082 2394 15099 2411
rect 14882 2394 14899 2411
rect 15402 2394 15419 2411
rect 15522 2394 15539 2411
rect 15042 2394 15059 2411
rect 14922 2394 14939 2411
rect 15562 2394 15579 2411
rect 15002 2394 15019 2411
rect 14882 2394 14899 2411
rect 15162 2394 15179 2411
rect 15362 2394 15379 2411
rect 14962 2394 14979 2411
rect 14962 2394 14979 2411
rect 15442 2394 15459 2411
rect 15122 2394 15139 2411
rect 14922 2394 14939 2411
rect 15322 2394 15339 2411
rect 15562 2394 15579 2411
rect 15522 2394 15539 2411
rect 15482 2394 15499 2411
rect 15442 2394 15459 2411
rect 15402 2394 15419 2411
rect 15362 2394 15379 2411
rect 15322 2394 15339 2411
rect 15242 2394 15259 2411
rect 15282 2394 15299 2411
rect 15282 2394 15299 2411
rect 15202 2394 15219 2411
rect 15162 2394 15179 2411
rect 15242 2394 15259 2411
rect 15122 2394 15139 2411
rect 15482 2394 15499 2411
rect 15082 2394 15099 2411
rect 15202 2394 15219 2411
rect 15042 2394 15059 2411
rect 15002 2394 15019 2411
rect 14482 2394 14499 2411
rect 14482 2394 14499 2411
rect 14442 2394 14459 2411
rect 14402 2394 14419 2411
rect 14682 2394 14699 2411
rect 14842 2394 14859 2411
rect 14802 2394 14819 2411
rect 14442 2394 14459 2411
rect 14762 2394 14779 2411
rect 14402 2394 14419 2411
rect 14642 2394 14659 2411
rect 14842 2394 14859 2411
rect 14602 2394 14619 2411
rect 14802 2394 14819 2411
rect 14762 2394 14779 2411
rect 14562 2394 14579 2411
rect 14722 2394 14739 2411
rect 14682 2394 14699 2411
rect 14642 2394 14659 2411
rect 14722 2394 14739 2411
rect 14602 2394 14619 2411
rect 14522 2394 14539 2411
rect 14562 2394 14579 2411
rect 16402 2394 16419 2411
rect 15882 2394 15899 2411
rect 15762 2394 15779 2411
rect 15922 2394 15939 2411
rect 15842 2394 15859 2411
rect 15882 2394 15899 2411
rect 15922 2394 15939 2411
rect 16682 2394 16699 2411
rect 15682 2394 15699 2411
rect 16242 2394 16259 2411
rect 16362 2394 16379 2411
rect 16202 2394 16219 2411
rect 16322 2394 16339 2411
rect 16642 2394 16659 2411
rect 16362 2394 16379 2411
rect 15722 2394 15739 2411
rect 16322 2394 16339 2411
rect 16602 2394 16619 2411
rect 16282 2394 16299 2411
rect 15682 2394 15699 2411
rect 16282 2394 16299 2411
rect 15642 2394 15659 2411
rect 16562 2394 16579 2411
rect 16522 2394 16539 2411
rect 15602 2394 15619 2411
rect 16242 2394 16259 2411
rect 16482 2394 16499 2411
rect 15642 2394 15659 2411
rect 16202 2394 16219 2411
rect 16162 2394 16179 2411
rect 15722 2394 15739 2411
rect 16402 2394 16419 2411
rect 16442 2394 16459 2411
rect 16162 2394 16179 2411
rect 16722 2394 16739 2411
rect 16682 2394 16699 2411
rect 16642 2394 16659 2411
rect 16602 2394 16619 2411
rect 16562 2394 16579 2411
rect 16522 2394 16539 2411
rect 15802 2394 15819 2411
rect 16482 2394 16499 2411
rect 16122 2394 16139 2411
rect 15602 2394 15619 2411
rect 16082 2394 16099 2411
rect 16042 2394 16059 2411
rect 16002 2394 16019 2411
rect 15802 2394 15819 2411
rect 15962 2394 15979 2411
rect 16082 2394 16099 2411
rect 15762 2394 15779 2411
rect 16042 2394 16059 2411
rect 16002 2394 16019 2411
rect 16442 2394 16459 2411
rect 16122 2394 16139 2411
rect 16722 2394 16739 2411
rect 15962 2394 15979 2411
rect 15842 2394 15859 2411
rect 17362 2394 17379 2411
rect 17322 2394 17339 2411
rect 17282 2394 17299 2411
rect 17242 2394 17259 2411
rect 16882 2394 16899 2411
rect 16842 2394 16859 2411
rect 18082 2394 18099 2411
rect 18042 2394 18059 2411
rect 17002 2394 17019 2411
rect 17002 2394 17019 2411
rect 16962 2394 16979 2411
rect 18002 2394 18019 2411
rect 17962 2394 17979 2411
rect 16802 2394 16819 2411
rect 17922 2394 17939 2411
rect 16962 2394 16979 2411
rect 17882 2394 17899 2411
rect 16842 2394 16859 2411
rect 16922 2394 16939 2411
rect 17842 2394 17859 2411
rect 17802 2394 17819 2411
rect 16922 2394 16939 2411
rect 17202 2394 17219 2411
rect 17762 2394 17779 2411
rect 17722 2394 17739 2411
rect 17682 2394 17699 2411
rect 17642 2394 17659 2411
rect 17602 2394 17619 2411
rect 16802 2394 16819 2411
rect 17562 2394 17579 2411
rect 17162 2394 17179 2411
rect 16882 2394 16899 2411
rect 18082 2394 18099 2411
rect 17122 2394 17139 2411
rect 17082 2394 17099 2411
rect 17042 2394 17059 2411
rect 18042 2394 18059 2411
rect 17122 2394 17139 2411
rect 18002 2394 18019 2411
rect 17082 2394 17099 2411
rect 17042 2394 17059 2411
rect 17482 2394 17499 2411
rect 17442 2394 17459 2411
rect 17522 2394 17539 2411
rect 17962 2394 17979 2411
rect 17522 2394 17539 2411
rect 17922 2394 17939 2411
rect 17882 2394 17899 2411
rect 17842 2394 17859 2411
rect 17802 2394 17819 2411
rect 17762 2394 17779 2411
rect 17722 2394 17739 2411
rect 17682 2394 17699 2411
rect 17642 2394 17659 2411
rect 17602 2394 17619 2411
rect 17562 2394 17579 2411
rect 17402 2394 17419 2411
rect 17362 2394 17379 2411
rect 17322 2394 17339 2411
rect 17282 2394 17299 2411
rect 17242 2394 17259 2411
rect 17202 2394 17219 2411
rect 17162 2394 17179 2411
rect 17482 2394 17499 2411
rect 17442 2394 17459 2411
rect 17402 2394 17419 2411
rect -9412 2394 -9395 2411
rect -9412 2394 -9395 2411
rect -325 8582 -308 8599
rect -285 8582 -268 8599
rect -245 8582 -228 8599
rect -205 8582 -188 8599
rect -165 8582 -148 8599
rect -125 8582 -108 8599
rect -85 8582 -68 8599
rect -45 8582 -28 8599
rect -5 8582 13 8599
rect 36 8582 53 8599
rect 76 8582 93 8599
rect -1685 8582 -1668 8599
rect -1725 8582 -1708 8599
rect -1765 8582 -1748 8599
rect -1805 8582 -1788 8599
rect -1845 8582 -1828 8599
rect -1885 8582 -1868 8599
rect -1925 8582 -1908 8599
rect -1965 8582 -1948 8599
rect -2005 8582 -1988 8599
rect -2045 8582 -2028 8599
rect -2085 8582 -2068 8599
rect -2125 8582 -2108 8599
rect -2165 8582 -2148 8599
rect -2205 8582 -2188 8599
rect -965 8582 -948 8599
rect -1685 8582 -1668 8599
rect -1725 8582 -1708 8599
rect -1765 8582 -1748 8599
rect -1805 8582 -1788 8599
rect -1845 8582 -1828 8599
rect -1885 8582 -1868 8599
rect -1925 8582 -1908 8599
rect -1965 8582 -1948 8599
rect -2005 8582 -1988 8599
rect -2045 8582 -2028 8599
rect -2085 8582 -2068 8599
rect -2125 8582 -2108 8599
rect -2165 8582 -2148 8599
rect -2205 8582 -2188 8599
rect -925 8582 -908 8599
rect -2245 8582 -2228 8599
rect -2245 8582 -2228 8599
rect -885 8582 -868 8599
rect -845 8582 -828 8599
rect -805 8582 -788 8599
rect -765 8582 -748 8599
rect -725 8582 -708 8599
rect -685 8582 -668 8599
rect -645 8582 -628 8599
rect -605 8582 -588 8599
rect -565 8582 -548 8599
rect -525 8582 -508 8599
rect -485 8582 -468 8599
rect -445 8582 -428 8599
rect -405 8582 -388 8599
rect -365 8582 -348 8599
rect -2485 8582 -2468 8599
rect -2725 8582 -2708 8599
rect -2565 8582 -2548 8599
rect -2285 8582 -2268 8599
rect -3285 8582 -3268 8599
rect -2765 8582 -2748 8599
rect -2805 8582 -2788 8599
rect -2765 8582 -2748 8599
rect -3085 8582 -3068 8599
rect -2805 8582 -2788 8599
rect -2525 8582 -2508 8599
rect -3325 8582 -3308 8599
rect -3405 8582 -3388 8599
rect -3325 8582 -3308 8599
rect -2525 8582 -2508 8599
rect -2325 8582 -2308 8599
rect -2365 8582 -2348 8599
rect -2965 8582 -2948 8599
rect -3125 8582 -3108 8599
rect -2565 8582 -2548 8599
rect -2645 8582 -2628 8599
rect -3445 8582 -3428 8599
rect -2605 8582 -2588 8599
rect -3285 8582 -3268 8599
rect -2405 8582 -2388 8599
rect -2365 8582 -2348 8599
rect -2685 8582 -2668 8599
rect -2845 8582 -2828 8599
rect -3165 8582 -3148 8599
rect -2845 8582 -2828 8599
rect -2605 8582 -2588 8599
rect -3365 8582 -3348 8599
rect -2885 8582 -2868 8599
rect -2925 8582 -2908 8599
rect -3445 8582 -3428 8599
rect -2405 8582 -2388 8599
rect -2285 8582 -2268 8599
rect -3405 8582 -3388 8599
rect -3005 8582 -2988 8599
rect -2325 8582 -2308 8599
rect -2885 8582 -2868 8599
rect -2445 8582 -2428 8599
rect -2685 8582 -2668 8599
rect -2725 8582 -2708 8599
rect -2925 8582 -2908 8599
rect -3205 8582 -3188 8599
rect -3365 8582 -3348 8599
rect -2645 8582 -2628 8599
rect -2965 8582 -2948 8599
rect -3005 8582 -2988 8599
rect -3045 8582 -3028 8599
rect -3085 8582 -3068 8599
rect -2445 8582 -2428 8599
rect -3125 8582 -3108 8599
rect -3165 8582 -3148 8599
rect -3205 8582 -3188 8599
rect -3245 8582 -3228 8599
rect -3045 8582 -3028 8599
rect -2485 8582 -2468 8599
rect -3245 8582 -3228 8599
rect -4485 8582 -4468 8599
rect -4405 8582 -4388 8599
rect -3765 8582 -3748 8599
rect -4285 8582 -4268 8599
rect -4325 8582 -4308 8599
rect -3565 8582 -3548 8599
rect -4565 8582 -4548 8599
rect -3685 8582 -3668 8599
rect -3605 8582 -3588 8599
rect -3765 8582 -3748 8599
rect -3885 8582 -3868 8599
rect -4205 8582 -4188 8599
rect -3885 8582 -3868 8599
rect -4245 8582 -4228 8599
rect -3605 8582 -3588 8599
rect -3805 8582 -3788 8599
rect -3485 8582 -3468 8599
rect -4485 8582 -4468 8599
rect -3645 8582 -3628 8599
rect -4125 8582 -4108 8599
rect -3485 8582 -3468 8599
rect -3965 8582 -3948 8599
rect -3805 8582 -3788 8599
rect -3725 8582 -3708 8599
rect -4445 8582 -4428 8599
rect -4165 8582 -4148 8599
rect -3645 8582 -3628 8599
rect -4445 8582 -4428 8599
rect -4365 8582 -4348 8599
rect -4605 8582 -4588 8599
rect -4405 8582 -4388 8599
rect -3965 8582 -3948 8599
rect -4045 8582 -4028 8599
rect -4005 8582 -3988 8599
rect -3845 8582 -3828 8599
rect -4285 8582 -4268 8599
rect -4605 8582 -4588 8599
rect -4325 8582 -4308 8599
rect -3845 8582 -3828 8599
rect -4645 8582 -4628 8599
rect -3565 8582 -3548 8599
rect -4085 8582 -4068 8599
rect -4525 8582 -4508 8599
rect -4365 8582 -4348 8599
rect -4245 8582 -4228 8599
rect -3525 8582 -3508 8599
rect -4165 8582 -4148 8599
rect -4645 8582 -4628 8599
rect -3525 8582 -3508 8599
rect -4525 8582 -4508 8599
rect -3685 8582 -3668 8599
rect -4085 8582 -4068 8599
rect -4005 8582 -3988 8599
rect -4205 8582 -4188 8599
rect -3925 8582 -3908 8599
rect -3725 8582 -3708 8599
rect -4125 8582 -4108 8599
rect -4565 8582 -4548 8599
rect -4045 8582 -4028 8599
rect -3925 8582 -3908 8599
rect -5845 8582 -5828 8599
rect -5845 8582 -5828 8599
rect -4925 8582 -4908 8599
rect -5445 8582 -5428 8599
rect -5365 8582 -5348 8599
rect -5165 8582 -5148 8599
rect -5165 8582 -5148 8599
rect -4965 8582 -4948 8599
rect -5445 8582 -5428 8599
rect -5485 8582 -5468 8599
rect -5245 8582 -5228 8599
rect -5005 8582 -4988 8599
rect -5525 8582 -5508 8599
rect -4765 8582 -4748 8599
rect -4805 8582 -4788 8599
rect -5765 8582 -5748 8599
rect -5525 8582 -5508 8599
rect -5565 8582 -5548 8599
rect -5125 8582 -5108 8599
rect -5565 8582 -5548 8599
rect -5605 8582 -5588 8599
rect -4885 8582 -4868 8599
rect -5045 8582 -5028 8599
rect -5685 8582 -5668 8599
rect -5085 8582 -5068 8599
rect -5805 8582 -5788 8599
rect -5605 8582 -5588 8599
rect -5645 8582 -5628 8599
rect -5205 8582 -5188 8599
rect -5685 8582 -5668 8599
rect -4845 8582 -4828 8599
rect -4925 8582 -4908 8599
rect -5725 8582 -5708 8599
rect -4685 8582 -4668 8599
rect -5205 8582 -5188 8599
rect -5765 8582 -5748 8599
rect -4685 8582 -4668 8599
rect -5405 8582 -5388 8599
rect -4965 8582 -4948 8599
rect -4845 8582 -4828 8599
rect -5285 8582 -5268 8599
rect -5805 8582 -5788 8599
rect -5325 8582 -5308 8599
rect -4765 8582 -4748 8599
rect -4805 8582 -4788 8599
rect -5005 8582 -4988 8599
rect -4885 8582 -4868 8599
rect -5125 8582 -5108 8599
rect -5645 8582 -5628 8599
rect -5365 8582 -5348 8599
rect -5085 8582 -5068 8599
rect -5045 8582 -5028 8599
rect -4725 8582 -4708 8599
rect -5325 8582 -5308 8599
rect -5725 8582 -5708 8599
rect -4725 8582 -4708 8599
rect -5245 8582 -5228 8599
rect -5485 8582 -5468 8599
rect -5405 8582 -5388 8599
rect -5285 8582 -5268 8599
rect -6446 8582 -6429 8599
rect -6926 8582 -6909 8599
rect -6766 8582 -6749 8599
rect -6246 8582 -6229 8599
rect -5965 8582 -5948 8599
rect -6046 8582 -6029 8599
rect -6886 8582 -6869 8599
rect -6486 8582 -6469 8599
rect -6446 8582 -6429 8599
rect -6806 8582 -6789 8599
rect -6046 8582 -6029 8599
rect -5885 8582 -5868 8599
rect -6326 8582 -6309 8599
rect -6526 8582 -6509 8599
rect -6686 8582 -6669 8599
rect -6646 8582 -6629 8599
rect -6126 8582 -6109 8599
rect -6766 8582 -6749 8599
rect -6246 8582 -6229 8599
rect -6566 8582 -6549 8599
rect -6326 8582 -6309 8599
rect -5925 8582 -5908 8599
rect -6806 8582 -6789 8599
rect -6006 8582 -5989 8599
rect -6366 8582 -6349 8599
rect -7006 8582 -6989 8599
rect -6566 8582 -6549 8599
rect -6486 8582 -6469 8599
rect -6086 8582 -6069 8599
rect -6846 8582 -6829 8599
rect -6006 8582 -5989 8599
rect -5965 8582 -5948 8599
rect -6966 8582 -6949 8599
rect -6366 8582 -6349 8599
rect -6286 8582 -6269 8599
rect -6166 8582 -6149 8599
rect -6846 8582 -6829 8599
rect -6966 8582 -6949 8599
rect -6526 8582 -6509 8599
rect -6206 8582 -6189 8599
rect -6606 8582 -6589 8599
rect -6726 8582 -6709 8599
rect -7006 8582 -6989 8599
rect -6926 8582 -6909 8599
rect -6126 8582 -6109 8599
rect -6726 8582 -6709 8599
rect -5885 8582 -5868 8599
rect -5925 8582 -5908 8599
rect -6646 8582 -6629 8599
rect -6406 8582 -6389 8599
rect -6286 8582 -6269 8599
rect -6206 8582 -6189 8599
rect -6606 8582 -6589 8599
rect -6406 8582 -6389 8599
rect -6686 8582 -6669 8599
rect -6086 8582 -6069 8599
rect -6886 8582 -6869 8599
rect -6166 8582 -6149 8599
rect -7366 8582 -7349 8599
rect -7766 8582 -7749 8599
rect -7086 8582 -7069 8599
rect -8126 8582 -8109 8599
rect -7086 8582 -7069 8599
rect -7806 8582 -7789 8599
rect -7966 8582 -7949 8599
rect -7886 8582 -7869 8599
rect -7726 8582 -7709 8599
rect -7286 8582 -7269 8599
rect -7566 8582 -7549 8599
rect -7806 8582 -7789 8599
rect -7326 8582 -7309 8599
rect -7206 8582 -7189 8599
rect -8126 8582 -8109 8599
rect -8166 8582 -8149 8599
rect -7646 8582 -7629 8599
rect -7686 8582 -7669 8599
rect -7126 8582 -7109 8599
rect -7646 8582 -7629 8599
rect -8166 8582 -8149 8599
rect -7446 8582 -7429 8599
rect -8006 8582 -7989 8599
rect -7486 8582 -7469 8599
rect -7046 8582 -7029 8599
rect -7166 8582 -7149 8599
rect -7966 8582 -7949 8599
rect -7446 8582 -7429 8599
rect -8086 8582 -8069 8599
rect -8006 8582 -7989 8599
rect -7046 8582 -7029 8599
rect -7326 8582 -7309 8599
rect -7406 8582 -7389 8599
rect -8206 8582 -8189 8599
rect -7526 8582 -7509 8599
rect -7166 8582 -7149 8599
rect -7606 8582 -7589 8599
rect -7766 8582 -7749 8599
rect -7486 8582 -7469 8599
rect -8206 8582 -8189 8599
rect -7246 8582 -7229 8599
rect -8046 8582 -8029 8599
rect -7686 8582 -7669 8599
rect -7206 8582 -7189 8599
rect -7886 8582 -7869 8599
rect -7726 8582 -7709 8599
rect -7526 8582 -7509 8599
rect -7366 8582 -7349 8599
rect -7846 8582 -7829 8599
rect -7926 8582 -7909 8599
rect -7406 8582 -7389 8599
rect -7846 8582 -7829 8599
rect -7246 8582 -7229 8599
rect -7566 8582 -7549 8599
rect -7606 8582 -7589 8599
rect -8046 8582 -8029 8599
rect -7126 8582 -7109 8599
rect -8086 8582 -8069 8599
rect -7926 8582 -7909 8599
rect -7286 8582 -7269 8599
rect -8886 8582 -8869 8599
rect -8606 8582 -8589 8599
rect -8926 8582 -8909 8599
rect -9166 8582 -9149 8599
rect -8246 8582 -8229 8599
rect -8286 8582 -8269 8599
rect -8446 8582 -8429 8599
rect -8686 8582 -8669 8599
rect -8286 8582 -8269 8599
rect -8606 8582 -8589 8599
rect -8566 8582 -8549 8599
rect -8406 8582 -8389 8599
rect -9366 8582 -9349 8599
rect -8926 8582 -8909 8599
rect -8486 8582 -8469 8599
rect -8846 8582 -8829 8599
rect -9286 8582 -9269 8599
rect -8806 8582 -8789 8599
rect -8526 8582 -8509 8599
rect -8966 8582 -8949 8599
rect -8766 8582 -8749 8599
rect -9366 8582 -9349 8599
rect -9086 8582 -9069 8599
rect -8246 8582 -8229 8599
rect -8486 8582 -8469 8599
rect -9326 8582 -9309 8599
rect -8886 8582 -8869 8599
rect -8526 8582 -8509 8599
rect -9326 8582 -9309 8599
rect -9006 8582 -8989 8599
rect -9206 8582 -9189 8599
rect -9166 8582 -9149 8599
rect -8646 8582 -8629 8599
rect -8846 8582 -8829 8599
rect -9206 8582 -9189 8599
rect -8366 8582 -8349 8599
rect -9246 8582 -9229 8599
rect -8326 8582 -8309 8599
rect -9286 8582 -9269 8599
rect -8726 8582 -8709 8599
rect -9126 8582 -9109 8599
rect -9246 8582 -9229 8599
rect -8686 8582 -8669 8599
rect -9406 8582 -9389 8599
rect -8966 8582 -8949 8599
rect -9406 8582 -9389 8599
rect -9046 8582 -9029 8599
rect -8446 8582 -8429 8599
rect -8326 8582 -8309 8599
rect -8646 8582 -8629 8599
rect -9046 8582 -9029 8599
rect -8366 8582 -8349 8599
rect -8766 8582 -8749 8599
rect -9126 8582 -9109 8599
rect -8566 8582 -8549 8599
rect -8406 8582 -8389 8599
rect -9006 8582 -8989 8599
rect -9086 8582 -9069 8599
rect -8726 8582 -8709 8599
rect -8806 8582 -8789 8599
rect -10606 8582 -10589 8599
rect -10606 8582 -10589 8599
rect -10406 8582 -10389 8599
rect -10086 8582 -10069 8599
rect -10446 8582 -10429 8599
rect -10366 8582 -10349 8599
rect -10406 8582 -10389 8599
rect -10486 8582 -10469 8599
rect -9646 8582 -9629 8599
rect -10126 8582 -10109 8599
rect -9686 8582 -9669 8599
rect -10246 8582 -10229 8599
rect -9726 8582 -9709 8599
rect -10446 8582 -10429 8599
rect -10526 8582 -10509 8599
rect -9806 8582 -9789 8599
rect -9486 8582 -9469 8599
rect -9886 8582 -9869 8599
rect -10246 8582 -10229 8599
rect -10046 8582 -10029 8599
rect -9606 8582 -9589 8599
rect -10126 8582 -10109 8599
rect -10566 8582 -10549 8599
rect -10006 8582 -9989 8599
rect -9526 8582 -9509 8599
rect -9446 8582 -9429 8599
rect -9446 8582 -9429 8599
rect -10286 8582 -10269 8599
rect -10086 8582 -10069 8599
rect -9526 8582 -9509 8599
rect -10046 8582 -10029 8599
rect -9726 8582 -9709 8599
rect -10006 8582 -9989 8599
rect -9846 8582 -9829 8599
rect -10366 8582 -10349 8599
rect -10206 8582 -10189 8599
rect -10166 8582 -10149 8599
rect -9886 8582 -9869 8599
rect -9806 8582 -9789 8599
rect -9966 8582 -9949 8599
rect -9486 8582 -9469 8599
rect -9686 8582 -9669 8599
rect -10486 8582 -10469 8599
rect -9766 8582 -9749 8599
rect -9966 8582 -9949 8599
rect -10526 8582 -10509 8599
rect -9926 8582 -9909 8599
rect -9566 8582 -9549 8599
rect -10326 8582 -10309 8599
rect -9566 8582 -9549 8599
rect -9646 8582 -9629 8599
rect -10206 8582 -10189 8599
rect -10566 8582 -10549 8599
rect -9846 8582 -9829 8599
rect -9766 8582 -9749 8599
rect -10166 8582 -10149 8599
rect -10286 8582 -10269 8599
rect -9926 8582 -9909 8599
rect -9606 8582 -9589 8599
rect -10326 8582 -10309 8599
rect -11606 8582 -11589 8599
rect -11166 8582 -11149 8599
rect -10686 8582 -10669 8599
rect -10806 8582 -10789 8599
rect -11366 8582 -11349 8599
rect -11646 8582 -11629 8599
rect -10886 8582 -10869 8599
rect -11126 8582 -11109 8599
rect -11006 8582 -10989 8599
rect -10726 8582 -10709 8599
rect -11086 8582 -11069 8599
rect -11406 8582 -11389 8599
rect -11526 8582 -11509 8599
rect -11486 8582 -11469 8599
rect -11686 8582 -11669 8599
rect -11326 8582 -11309 8599
rect -11126 8582 -11109 8599
rect -11406 8582 -11389 8599
rect -11086 8582 -11069 8599
rect -10926 8582 -10909 8599
rect -11286 8582 -11269 8599
rect -11686 8582 -11669 8599
rect -11566 8582 -11549 8599
rect -11166 8582 -11149 8599
rect -10766 8582 -10749 8599
rect -11646 8582 -11629 8599
rect -10966 8582 -10949 8599
rect -11246 8582 -11229 8599
rect -11446 8582 -11429 8599
rect -11766 8582 -11749 8599
rect -10766 8582 -10749 8599
rect -11046 8582 -11029 8599
rect -11486 8582 -11469 8599
rect -11566 8582 -11549 8599
rect -11446 8582 -11429 8599
rect -11726 8582 -11709 8599
rect -11246 8582 -11229 8599
rect -11606 8582 -11589 8599
rect -11366 8582 -11349 8599
rect -11046 8582 -11029 8599
rect -10846 8582 -10829 8599
rect -10926 8582 -10909 8599
rect -11326 8582 -11309 8599
rect -10646 8582 -10629 8599
rect -10646 8582 -10629 8599
rect -10806 8582 -10789 8599
rect -11766 8582 -11749 8599
rect -11006 8582 -10989 8599
rect -11206 8582 -11189 8599
rect -11206 8582 -11189 8599
rect -10846 8582 -10829 8599
rect -11726 8582 -11709 8599
rect -10886 8582 -10869 8599
rect -11286 8582 -11269 8599
rect -10686 8582 -10669 8599
rect -11526 8582 -11509 8599
rect -10966 8582 -10949 8599
rect -10726 8582 -10709 8599
rect -12566 8582 -12549 8599
rect -12046 8582 -12029 8599
rect -12126 8582 -12109 8599
rect -12286 8582 -12269 8599
rect -12886 8582 -12869 8599
rect -12806 8582 -12789 8599
rect -12686 8582 -12669 8599
rect -11926 8582 -11909 8599
rect -12406 8582 -12389 8599
rect -12606 8582 -12589 8599
rect -12366 8582 -12349 8599
rect -12526 8582 -12509 8599
rect -12006 8582 -11989 8599
rect -12966 8582 -12949 8599
rect -12446 8582 -12429 8599
rect -11966 8582 -11949 8599
rect -12206 8582 -12189 8599
rect -12766 8582 -12749 8599
rect -12926 8582 -12909 8599
rect -12646 8582 -12629 8599
rect -12726 8582 -12709 8599
rect -11846 8582 -11829 8599
rect -11886 8582 -11869 8599
rect -12966 8582 -12949 8599
rect -11846 8582 -11829 8599
rect -11966 8582 -11949 8599
rect -12326 8582 -12309 8599
rect -12606 8582 -12589 8599
rect -12686 8582 -12669 8599
rect -12086 8582 -12069 8599
rect -12726 8582 -12709 8599
rect -12166 8582 -12149 8599
rect -12886 8582 -12869 8599
rect -12206 8582 -12189 8599
rect -11886 8582 -11869 8599
rect -12006 8582 -11989 8599
rect -12766 8582 -12749 8599
rect -12246 8582 -12229 8599
rect -12926 8582 -12909 8599
rect -12246 8582 -12229 8599
rect -12086 8582 -12069 8599
rect -12806 8582 -12789 8599
rect -12406 8582 -12389 8599
rect -12366 8582 -12349 8599
rect -12486 8582 -12469 8599
rect -12446 8582 -12429 8599
rect -12846 8582 -12829 8599
rect -12486 8582 -12469 8599
rect -11926 8582 -11909 8599
rect -12286 8582 -12269 8599
rect -12846 8582 -12829 8599
rect -12126 8582 -12109 8599
rect -11806 8582 -11789 8599
rect -12326 8582 -12309 8599
rect -12046 8582 -12029 8599
rect -11806 8582 -11789 8599
rect -12566 8582 -12549 8599
rect -12646 8582 -12629 8599
rect -12526 8582 -12509 8599
rect -12166 8582 -12149 8599
rect -13166 8582 -13149 8599
rect -13406 8582 -13389 8599
rect -13686 8582 -13669 8599
rect -13966 8582 -13949 8599
rect -13966 8582 -13949 8599
rect -13486 8582 -13469 8599
rect -14006 8582 -13989 8599
rect -14126 8582 -14109 8599
rect -14006 8582 -13989 8599
rect -13486 8582 -13469 8599
rect -13886 8582 -13869 8599
rect -13606 8582 -13589 8599
rect -13566 8582 -13549 8599
rect -14046 8582 -14029 8599
rect -13046 8582 -13029 8599
rect -13286 8582 -13269 8599
rect -13606 8582 -13589 8599
rect -13206 8582 -13189 8599
rect -13646 8582 -13629 8599
rect -13526 8582 -13509 8599
rect -13926 8582 -13909 8599
rect -13006 8582 -12989 8599
rect -13766 8582 -13749 8599
rect -13846 8582 -13829 8599
rect -13566 8582 -13549 8599
rect -13726 8582 -13709 8599
rect -13086 8582 -13069 8599
rect -14166 8582 -14149 8599
rect -13206 8582 -13189 8599
rect -13326 8582 -13309 8599
rect -13086 8582 -13069 8599
rect -13726 8582 -13709 8599
rect -13686 8582 -13669 8599
rect -13366 8582 -13349 8599
rect -13126 8582 -13109 8599
rect -13046 8582 -13029 8599
rect -13286 8582 -13269 8599
rect -13406 8582 -13389 8599
rect -13246 8582 -13229 8599
rect -14086 8582 -14069 8599
rect -13446 8582 -13429 8599
rect -13366 8582 -13349 8599
rect -14086 8582 -14069 8599
rect -14126 8582 -14109 8599
rect -14166 8582 -14149 8599
rect -13766 8582 -13749 8599
rect -13846 8582 -13829 8599
rect -13446 8582 -13429 8599
rect -13166 8582 -13149 8599
rect -13326 8582 -13309 8599
rect -13886 8582 -13869 8599
rect -13806 8582 -13789 8599
rect -13006 8582 -12989 8599
rect -13646 8582 -13629 8599
rect -13526 8582 -13509 8599
rect -13926 8582 -13909 8599
rect -14046 8582 -14029 8599
rect -13126 8582 -13109 8599
rect -13806 8582 -13789 8599
rect -13246 8582 -13229 8599
rect -15366 8582 -15349 8599
rect -15366 8582 -15349 8599
rect -14966 8582 -14949 8599
rect -14606 8582 -14589 8599
rect -15166 8582 -15149 8599
rect -15126 8582 -15109 8599
rect -15206 8582 -15189 8599
rect -14686 8582 -14669 8599
rect -15046 8582 -15029 8599
rect -14526 8582 -14509 8599
rect -15086 8582 -15069 8599
rect -14406 8582 -14389 8599
rect -14926 8582 -14909 8599
rect -14766 8582 -14749 8599
rect -14566 8582 -14549 8599
rect -14366 8582 -14349 8599
rect -15326 8582 -15309 8599
rect -14246 8582 -14229 8599
rect -15006 8582 -14989 8599
rect -15326 8582 -15309 8599
rect -14526 8582 -14509 8599
rect -14326 8582 -14309 8599
rect -14646 8582 -14629 8599
rect -15246 8582 -15229 8599
rect -14726 8582 -14709 8599
rect -14646 8582 -14629 8599
rect -14486 8582 -14469 8599
rect -15286 8582 -15269 8599
rect -14726 8582 -14709 8599
rect -14846 8582 -14829 8599
rect -14286 8582 -14269 8599
rect -15246 8582 -15229 8599
rect -14606 8582 -14589 8599
rect -14686 8582 -14669 8599
rect -15006 8582 -14989 8599
rect -14206 8582 -14189 8599
rect -14286 8582 -14269 8599
rect -15046 8582 -15029 8599
rect -14886 8582 -14869 8599
rect -14926 8582 -14909 8599
rect -15166 8582 -15149 8599
rect -15286 8582 -15269 8599
rect -14566 8582 -14549 8599
rect -14966 8582 -14949 8599
rect -14366 8582 -14349 8599
rect -15086 8582 -15069 8599
rect -14806 8582 -14789 8599
rect -14206 8582 -14189 8599
rect -14406 8582 -14389 8599
rect -14446 8582 -14429 8599
rect -14766 8582 -14749 8599
rect -14326 8582 -14309 8599
rect -14806 8582 -14789 8599
rect -14846 8582 -14829 8599
rect -14486 8582 -14469 8599
rect -14446 8582 -14429 8599
rect -14886 8582 -14869 8599
rect -14246 8582 -14229 8599
rect -15206 8582 -15189 8599
rect -15126 8582 -15109 8599
rect -15726 8582 -15709 8599
rect -15846 8582 -15829 8599
rect -16246 8582 -16229 8599
rect -16006 8582 -15989 8599
rect -15846 8582 -15829 8599
rect -15766 8582 -15749 8599
rect -15766 8582 -15749 8599
rect -16126 8582 -16109 8599
rect -16526 8582 -16509 8599
rect -16006 8582 -15989 8599
rect -16326 8582 -16309 8599
rect -15526 8582 -15509 8599
rect -16046 8582 -16029 8599
rect -16046 8582 -16029 8599
rect -15646 8582 -15629 8599
rect -15646 8582 -15629 8599
rect -15566 8582 -15549 8599
rect -15406 8582 -15389 8599
rect -15686 8582 -15669 8599
rect -16486 8582 -16469 8599
rect -16366 8582 -16349 8599
rect -15486 8582 -15469 8599
rect -15406 8582 -15389 8599
rect -15686 8582 -15669 8599
rect -15886 8582 -15869 8599
rect -15886 8582 -15869 8599
rect -15926 8582 -15909 8599
rect -16286 8582 -16269 8599
rect -16446 8582 -16429 8599
rect -15606 8582 -15589 8599
rect -15526 8582 -15509 8599
rect -16486 8582 -16469 8599
rect -15726 8582 -15709 8599
rect -16206 8582 -16189 8599
rect -16206 8582 -16189 8599
rect -15966 8582 -15949 8599
rect -15446 8582 -15429 8599
rect -15446 8582 -15429 8599
rect -16086 8582 -16069 8599
rect -16166 8582 -16149 8599
rect -16366 8582 -16349 8599
rect -16286 8582 -16269 8599
rect -16086 8582 -16069 8599
rect -16166 8582 -16149 8599
rect -15966 8582 -15949 8599
rect -16446 8582 -16429 8599
rect -16326 8582 -16309 8599
rect -16406 8582 -16389 8599
rect -16126 8582 -16109 8599
rect -15806 8582 -15789 8599
rect -15606 8582 -15589 8599
rect -16406 8582 -16389 8599
rect -16526 8582 -16509 8599
rect -15566 8582 -15549 8599
rect -16246 8582 -16229 8599
rect -15806 8582 -15789 8599
rect -15926 8582 -15909 8599
rect -15486 8582 -15469 8599
rect -17206 8582 -17189 8599
rect -17246 8582 -17229 8599
rect -16846 8582 -16829 8599
rect -17566 8582 -17549 8599
rect -16606 8582 -16589 8599
rect -16686 8582 -16669 8599
rect -17406 8582 -17389 8599
rect -16766 8582 -16749 8599
rect -17446 8582 -17429 8599
rect -17046 8582 -17029 8599
rect -16966 8582 -16949 8599
rect -16806 8582 -16789 8599
rect -17126 8582 -17109 8599
rect -16926 8582 -16909 8599
rect -17686 8582 -17669 8599
rect -17726 8582 -17709 8599
rect -17606 8582 -17589 8599
rect -16886 8582 -16869 8599
rect -17486 8582 -17469 8599
rect -16726 8582 -16709 8599
rect -17286 8582 -17269 8599
rect -16886 8582 -16869 8599
rect -17366 8582 -17349 8599
rect -17486 8582 -17469 8599
rect -17726 8582 -17709 8599
rect -16966 8582 -16949 8599
rect -16646 8582 -16629 8599
rect -17286 8582 -17269 8599
rect -17526 8582 -17509 8599
rect -17566 8582 -17549 8599
rect -17686 8582 -17669 8599
rect -17206 8582 -17189 8599
rect -16646 8582 -16629 8599
rect -17326 8582 -17309 8599
rect -17406 8582 -17389 8599
rect -17006 8582 -16989 8599
rect -17246 8582 -17229 8599
rect -16846 8582 -16829 8599
rect -16926 8582 -16909 8599
rect -17046 8582 -17029 8599
rect -17526 8582 -17509 8599
rect -17606 8582 -17589 8599
rect -16686 8582 -16669 8599
rect -17086 8582 -17069 8599
rect -17086 8582 -17069 8599
rect -17646 8582 -17629 8599
rect -16606 8582 -16589 8599
rect -17646 8582 -17629 8599
rect -16566 8582 -16549 8599
rect -16766 8582 -16749 8599
rect -17366 8582 -17349 8599
rect -17166 8582 -17149 8599
rect -16806 8582 -16789 8599
rect -17446 8582 -17429 8599
rect -17166 8582 -17149 8599
rect -17006 8582 -16989 8599
rect -16566 8582 -16549 8599
rect -17126 8582 -17109 8599
rect -16726 8582 -16709 8599
rect -17326 8582 -17309 8599
rect -18166 8582 -18149 8599
rect -18086 8582 -18069 8599
rect -18606 8582 -18589 8599
rect -18006 8582 -17989 8599
rect -18006 8582 -17989 8599
rect -18486 8582 -18469 8599
rect -18446 8582 -18429 8599
rect -17926 8582 -17909 8599
rect -18246 8582 -18229 8599
rect -18926 8582 -18909 8599
rect -18846 8582 -18829 8599
rect -18046 8582 -18029 8599
rect -18806 8582 -18789 8599
rect -18246 8582 -18229 8599
rect -17926 8582 -17909 8599
rect -18326 8582 -18309 8599
rect -18406 8582 -18389 8599
rect -18686 8582 -18669 8599
rect -18566 8582 -18549 8599
rect -18086 8582 -18069 8599
rect -17806 8582 -17789 8599
rect -18686 8582 -18669 8599
rect -18766 8582 -18749 8599
rect -18046 8582 -18029 8599
rect -17886 8582 -17869 8599
rect -18326 8582 -18309 8599
rect -18206 8582 -18189 8599
rect -18126 8582 -18109 8599
rect -18286 8582 -18269 8599
rect -18526 8582 -18509 8599
rect -18366 8582 -18349 8599
rect -18526 8582 -18509 8599
rect -18446 8582 -18429 8599
rect -18766 8582 -18749 8599
rect -17966 8582 -17949 8599
rect -18646 8582 -18629 8599
rect -17846 8582 -17829 8599
rect -18126 8582 -18109 8599
rect -18646 8582 -18629 8599
rect -18926 8582 -18909 8599
rect -18486 8582 -18469 8599
rect -18286 8582 -18269 8599
rect -18206 8582 -18189 8599
rect -18366 8582 -18349 8599
rect -17766 8582 -17749 8599
rect -18886 8582 -18869 8599
rect -18726 8582 -18709 8599
rect -17886 8582 -17869 8599
rect -18566 8582 -18549 8599
rect -18406 8582 -18389 8599
rect -18726 8582 -18709 8599
rect -18806 8582 -18789 8599
rect -17766 8582 -17749 8599
rect -17806 8582 -17789 8599
rect -18166 8582 -18149 8599
rect -18846 8582 -18829 8599
rect -18886 8582 -18869 8599
rect -17966 8582 -17949 8599
rect -18606 8582 -18589 8599
rect -17846 8582 -17829 8599
rect -14173 2394 -14156 2411
rect -14173 2394 -14156 2411
rect -11966 4652 -11949 4669
rect -11926 4652 -11909 4669
rect -12006 4652 -11989 4669
rect -12046 4652 -12029 4669
rect -11966 4652 -11949 4669
rect -12086 4652 -12069 4669
rect -12126 4652 -12109 4669
rect -12006 4652 -11989 4669
rect -12166 4652 -12149 4669
rect -12046 4652 -12029 4669
rect -12086 4652 -12069 4669
rect -11806 4652 -11789 4669
rect -12126 4652 -12109 4669
rect -12166 4652 -12149 4669
rect -12206 4652 -12189 4669
rect -11846 4652 -11829 4669
rect -12246 4652 -12229 4669
rect -12286 4652 -12269 4669
rect -12326 4652 -12309 4669
rect -11886 4652 -11869 4669
rect -12366 4652 -12349 4669
rect -12006 4652 -11989 4669
rect -12206 4652 -12189 4669
rect -12206 4652 -12189 4669
rect -12246 4652 -12229 4669
rect -12286 4652 -12269 4669
rect -12326 4652 -12309 4669
rect -11806 4652 -11789 4669
rect -12366 4652 -12349 4669
rect -11966 4652 -11949 4669
rect -11846 4652 -11829 4669
rect -11846 4652 -11829 4669
rect -11886 4652 -11869 4669
rect -11886 4652 -11869 4669
rect -12166 4652 -12149 4669
rect -12006 4652 -11989 4669
rect -11846 4652 -11829 4669
rect -12206 4652 -12189 4669
rect -11966 4652 -11949 4669
rect -12326 4652 -12309 4669
rect -12246 4652 -12229 4669
rect -12086 4652 -12069 4669
rect -12126 4652 -12109 4669
rect -12286 4652 -12269 4669
rect -11886 4652 -11869 4669
rect -12046 4652 -12029 4669
rect -12246 4652 -12229 4669
rect -12086 4652 -12069 4669
rect -11806 4652 -11789 4669
rect -12366 4652 -12349 4669
rect -12166 4652 -12149 4669
rect -12126 4652 -12109 4669
rect -11926 4652 -11909 4669
rect -12046 4652 -12029 4669
rect -12326 4652 -12309 4669
rect -11806 4652 -11789 4669
rect -12286 4652 -12269 4669
rect -11926 4652 -11909 4669
rect -12366 4652 -12349 4669
rect -11926 4652 -11909 4669
rect -12486 4652 -12469 4669
rect -12726 4652 -12709 4669
rect -12606 4652 -12589 4669
rect -12926 4652 -12909 4669
rect -12486 4652 -12469 4669
rect -12646 4652 -12629 4669
rect -12526 4652 -12509 4669
rect -12566 4652 -12549 4669
rect -12686 4652 -12669 4669
rect -12406 4652 -12389 4669
rect -12606 4652 -12589 4669
rect -12526 4652 -12509 4669
rect -12966 4652 -12949 4669
rect -12446 4652 -12429 4669
rect -12766 4652 -12749 4669
rect -12926 4652 -12909 4669
rect -12646 4652 -12629 4669
rect -12966 4652 -12949 4669
rect -12686 4652 -12669 4669
rect -12726 4652 -12709 4669
rect -12886 4652 -12869 4669
rect -12766 4652 -12749 4669
rect -12806 4652 -12789 4669
rect -12446 4652 -12429 4669
rect -12846 4652 -12829 4669
rect -12846 4652 -12829 4669
rect -12566 4652 -12549 4669
rect -12886 4652 -12869 4669
rect -12406 4652 -12389 4669
rect -12406 4652 -12389 4669
rect -12446 4652 -12429 4669
rect -12406 4652 -12389 4669
rect -12446 4652 -12429 4669
rect -12726 4652 -12709 4669
rect -12526 4652 -12509 4669
rect -12886 4652 -12869 4669
rect -12566 4652 -12549 4669
rect -12806 4652 -12789 4669
rect -12606 4652 -12589 4669
rect -12926 4652 -12909 4669
rect -12486 4652 -12469 4669
rect -12646 4652 -12629 4669
rect -12526 4652 -12509 4669
rect -12566 4652 -12549 4669
rect -12686 4652 -12669 4669
rect -12606 4652 -12589 4669
rect -12646 4652 -12629 4669
rect -12966 4652 -12949 4669
rect -12686 4652 -12669 4669
rect -12726 4652 -12709 4669
rect -12766 4652 -12749 4669
rect -12806 4652 -12789 4669
rect -12846 4652 -12829 4669
rect -12846 4652 -12829 4669
rect -12886 4652 -12869 4669
rect -12926 4652 -12909 4669
rect -12486 4652 -12469 4669
rect -12966 4652 -12949 4669
rect -12766 4652 -12749 4669
rect -12806 4652 -12789 4669
rect -13126 4652 -13109 4669
rect -13246 4652 -13229 4669
rect -13566 4652 -13549 4669
rect -13286 4652 -13269 4669
rect -13406 4652 -13389 4669
rect -13006 4652 -12989 4669
rect -13166 4652 -13149 4669
rect -13326 4652 -13309 4669
rect -13446 4652 -13429 4669
rect -13126 4652 -13109 4669
rect -13046 4652 -13029 4669
rect -13206 4652 -13189 4669
rect -13246 4652 -13229 4669
rect -13366 4652 -13349 4669
rect -13526 4652 -13509 4669
rect -13326 4652 -13309 4669
rect -13246 4652 -13229 4669
rect -13486 4652 -13469 4669
rect -13006 4652 -12989 4669
rect -13486 4652 -13469 4669
rect -13446 4652 -13429 4669
rect -13006 4652 -12989 4669
rect -13286 4652 -13269 4669
rect -13006 4652 -12989 4669
rect -13086 4652 -13069 4669
rect -13046 4652 -13029 4669
rect -13326 4652 -13309 4669
rect -13566 4652 -13549 4669
rect -13406 4652 -13389 4669
rect -13126 4652 -13109 4669
rect -13526 4652 -13509 4669
rect -13166 4652 -13149 4669
rect -13086 4652 -13069 4669
rect -13126 4652 -13109 4669
rect -13166 4652 -13149 4669
rect -13206 4652 -13189 4669
rect -13206 4652 -13189 4669
rect -13246 4652 -13229 4669
rect -13286 4652 -13269 4669
rect -13286 4652 -13269 4669
rect -13046 4652 -13029 4669
rect -13166 4652 -13149 4669
rect -13566 4652 -13549 4669
rect -13326 4652 -13309 4669
rect -13566 4652 -13549 4669
rect -13086 4652 -13069 4669
rect -13086 4652 -13069 4669
rect -13446 4652 -13429 4669
rect -13486 4652 -13469 4669
rect -13526 4652 -13509 4669
rect -13406 4652 -13389 4669
rect -13446 4652 -13429 4669
rect -13486 4652 -13469 4669
rect -13526 4652 -13509 4669
rect -13406 4652 -13389 4669
rect -13366 4652 -13349 4669
rect -13366 4652 -13349 4669
rect -13046 4652 -13029 4669
rect -13366 4652 -13349 4669
rect -13206 4652 -13189 4669
rect -14086 4652 -14069 4669
rect -13606 4652 -13589 4669
rect -14126 4652 -14109 4669
rect -13806 4652 -13789 4669
rect -14046 4652 -14029 4669
rect -13686 4652 -13669 4669
rect -13966 4652 -13949 4669
rect -14166 4652 -14149 4669
rect -14126 4652 -14109 4669
rect -13886 4652 -13869 4669
rect -13966 4652 -13949 4669
rect -13646 4652 -13629 4669
rect -14086 4652 -14069 4669
rect -13766 4652 -13749 4669
rect -13606 4652 -13589 4669
rect -13766 4652 -13749 4669
rect -13846 4652 -13829 4669
rect -13686 4652 -13669 4669
rect -13926 4652 -13909 4669
rect -13646 4652 -13629 4669
rect -14006 4652 -13989 4669
rect -13886 4652 -13869 4669
rect -13726 4652 -13709 4669
rect -14006 4652 -13989 4669
rect -13926 4652 -13909 4669
rect -14166 4652 -14149 4669
rect -13806 4652 -13789 4669
rect -13726 4652 -13709 4669
rect -14046 4652 -14029 4669
rect -13766 4652 -13749 4669
rect -13646 4652 -13629 4669
rect -14126 4652 -14109 4669
rect -14006 4652 -13989 4669
rect -13686 4652 -13669 4669
rect -13806 4652 -13789 4669
rect -13766 4652 -13749 4669
rect -14086 4652 -14069 4669
rect -14166 4652 -14149 4669
rect -14126 4652 -14109 4669
rect -13646 4652 -13629 4669
rect -13846 4652 -13829 4669
rect -14166 4652 -14149 4669
rect -13846 4652 -13829 4669
rect -13886 4652 -13869 4669
rect -13886 4652 -13869 4669
rect -13686 4652 -13669 4669
rect -13726 4652 -13709 4669
rect -13926 4652 -13909 4669
rect -13806 4652 -13789 4669
rect -13606 4652 -13589 4669
rect -13966 4652 -13949 4669
rect -13966 4652 -13949 4669
rect -13926 4652 -13909 4669
rect -14006 4652 -13989 4669
rect -13606 4652 -13589 4669
rect -13726 4652 -13709 4669
rect -14046 4652 -14029 4669
rect -14046 4652 -14029 4669
rect -14086 4652 -14069 4669
rect -13846 4652 -13829 4669
rect -10606 4652 -10589 4669
rect -10606 4652 -10589 4669
rect -10606 4652 -10589 4669
rect -10606 4652 -10589 4669
rect -10006 4652 -9989 4669
rect -10006 4652 -9989 4669
rect -10006 4652 -9989 4669
rect -10006 4652 -9989 4669
rect -9526 4652 -9509 4669
rect -9606 4652 -9589 4669
rect -9846 4652 -9829 4669
rect -9886 4652 -9869 4669
rect -9686 4652 -9669 4669
rect -9726 4652 -9709 4669
rect -9966 4652 -9949 4669
rect -9806 4652 -9789 4669
rect -9886 4652 -9869 4669
rect -9726 4652 -9709 4669
rect -9606 4652 -9589 4669
rect -9726 4652 -9709 4669
rect -9526 4652 -9509 4669
rect -9446 4652 -9429 4669
rect -9606 4652 -9589 4669
rect -9566 4652 -9549 4669
rect -9846 4652 -9829 4669
rect -9766 4652 -9749 4669
rect -9886 4652 -9869 4669
rect -9966 4652 -9949 4669
rect -9566 4652 -9549 4669
rect -9966 4652 -9949 4669
rect -9646 4652 -9629 4669
rect -9646 4652 -9629 4669
rect -9446 4652 -9429 4669
rect -9806 4652 -9789 4669
rect -9926 4652 -9909 4669
rect -9686 4652 -9669 4669
rect -9486 4652 -9469 4669
rect -9806 4652 -9789 4669
rect -9646 4652 -9629 4669
rect -9526 4652 -9509 4669
rect -9926 4652 -9909 4669
rect -9606 4652 -9589 4669
rect -9686 4652 -9669 4669
rect -9446 4652 -9429 4669
rect -9726 4652 -9709 4669
rect -9686 4652 -9669 4669
rect -9766 4652 -9749 4669
rect -9846 4652 -9829 4669
rect -9446 4652 -9429 4669
rect -9886 4652 -9869 4669
rect -9646 4652 -9629 4669
rect -9486 4652 -9469 4669
rect -9806 4652 -9789 4669
rect -9486 4652 -9469 4669
rect -9926 4652 -9909 4669
rect -9486 4652 -9469 4669
rect -9966 4652 -9949 4669
rect -9766 4652 -9749 4669
rect -9526 4652 -9509 4669
rect -9566 4652 -9549 4669
rect -9846 4652 -9829 4669
rect -9766 4652 -9749 4669
rect -9566 4652 -9549 4669
rect -9926 4652 -9909 4669
rect -10046 4652 -10029 4669
rect -10246 4652 -10229 4669
rect -10086 4652 -10069 4669
rect -10126 4652 -10109 4669
rect -10286 4652 -10269 4669
rect -10486 4652 -10469 4669
rect -10526 4652 -10509 4669
rect -10566 4652 -10549 4669
rect -10126 4652 -10109 4669
rect -10326 4652 -10309 4669
rect -10366 4652 -10349 4669
rect -10406 4652 -10389 4669
rect -10446 4652 -10429 4669
rect -10486 4652 -10469 4669
rect -10526 4652 -10509 4669
rect -10566 4652 -10549 4669
rect -10046 4652 -10029 4669
rect -10326 4652 -10309 4669
rect -10366 4652 -10349 4669
rect -10406 4652 -10389 4669
rect -10446 4652 -10429 4669
rect -10566 4652 -10549 4669
rect -10086 4652 -10069 4669
rect -10206 4652 -10189 4669
rect -10166 4652 -10149 4669
rect -10326 4652 -10309 4669
rect -10086 4652 -10069 4669
rect -10366 4652 -10349 4669
rect -10406 4652 -10389 4669
rect -10126 4652 -10109 4669
rect -10446 4652 -10429 4669
rect -10246 4652 -10229 4669
rect -10286 4652 -10269 4669
rect -10286 4652 -10269 4669
rect -10046 4652 -10029 4669
rect -10206 4652 -10189 4669
rect -10486 4652 -10469 4669
rect -10526 4652 -10509 4669
rect -10206 4652 -10189 4669
rect -10566 4652 -10549 4669
rect -10166 4652 -10149 4669
rect -10286 4652 -10269 4669
rect -10366 4652 -10349 4669
rect -10126 4652 -10109 4669
rect -10326 4652 -10309 4669
rect -10446 4652 -10429 4669
rect -10486 4652 -10469 4669
rect -10246 4652 -10229 4669
rect -10526 4652 -10509 4669
rect -10046 4652 -10029 4669
rect -10166 4652 -10149 4669
rect -10206 4652 -10189 4669
rect -10246 4652 -10229 4669
rect -10086 4652 -10069 4669
rect -10406 4652 -10389 4669
rect -10166 4652 -10149 4669
rect -11206 4652 -11189 4669
rect -11206 4652 -11189 4669
rect -11206 4652 -11189 4669
rect -11206 4652 -11189 4669
rect -10846 4652 -10829 4669
rect -11166 4652 -11149 4669
rect -11006 4652 -10989 4669
rect -10686 4652 -10669 4669
rect -10726 4652 -10709 4669
rect -10766 4652 -10749 4669
rect -10726 4652 -10709 4669
rect -10646 4652 -10629 4669
rect -11046 4652 -11029 4669
rect -10686 4652 -10669 4669
rect -10886 4652 -10869 4669
rect -10646 4652 -10629 4669
rect -10926 4652 -10909 4669
rect -10806 4652 -10789 4669
rect -11126 4652 -11109 4669
rect -11086 4652 -11069 4669
rect -10886 4652 -10869 4669
rect -11086 4652 -11069 4669
rect -10966 4652 -10949 4669
rect -11166 4652 -11149 4669
rect -11086 4652 -11069 4669
rect -10766 4652 -10749 4669
rect -10766 4652 -10749 4669
rect -11126 4652 -11109 4669
rect -10646 4652 -10629 4669
rect -10806 4652 -10789 4669
rect -11006 4652 -10989 4669
rect -11126 4652 -11109 4669
rect -10686 4652 -10669 4669
rect -10846 4652 -10829 4669
rect -10966 4652 -10949 4669
rect -10646 4652 -10629 4669
rect -10726 4652 -10709 4669
rect -10886 4652 -10869 4669
rect -10926 4652 -10909 4669
rect -11166 4652 -11149 4669
rect -10966 4652 -10949 4669
rect -10926 4652 -10909 4669
rect -10926 4652 -10909 4669
rect -11086 4652 -11069 4669
rect -10686 4652 -10669 4669
rect -10966 4652 -10949 4669
rect -10806 4652 -10789 4669
rect -11006 4652 -10989 4669
rect -10846 4652 -10829 4669
rect -10846 4652 -10829 4669
rect -11126 4652 -11109 4669
rect -10726 4652 -10709 4669
rect -11046 4652 -11029 4669
rect -11006 4652 -10989 4669
rect -10886 4652 -10869 4669
rect -10766 4652 -10749 4669
rect -11166 4652 -11149 4669
rect -11046 4652 -11029 4669
rect -10806 4652 -10789 4669
rect -11046 4652 -11029 4669
rect -11726 4652 -11709 4669
rect -11406 4652 -11389 4669
rect -11766 4652 -11749 4669
rect -11606 4652 -11589 4669
rect -11526 4652 -11509 4669
rect -11246 4652 -11229 4669
rect -11286 4652 -11269 4669
rect -11326 4652 -11309 4669
rect -11366 4652 -11349 4669
rect -11686 4652 -11669 4669
rect -11446 4652 -11429 4669
rect -11246 4652 -11229 4669
rect -11446 4652 -11429 4669
rect -11646 4652 -11629 4669
rect -11526 4652 -11509 4669
rect -11246 4652 -11229 4669
rect -11286 4652 -11269 4669
rect -11486 4652 -11469 4669
rect -11286 4652 -11269 4669
rect -11246 4652 -11229 4669
rect -11566 4652 -11549 4669
rect -11326 4652 -11309 4669
rect -11646 4652 -11629 4669
rect -11366 4652 -11349 4669
rect -11566 4652 -11549 4669
rect -11606 4652 -11589 4669
rect -11326 4652 -11309 4669
rect -11406 4652 -11389 4669
rect -11766 4652 -11749 4669
rect -11726 4652 -11709 4669
rect -11766 4652 -11749 4669
rect -11526 4652 -11509 4669
rect -11606 4652 -11589 4669
rect -11686 4652 -11669 4669
rect -11686 4652 -11669 4669
rect -11446 4652 -11429 4669
rect -11446 4652 -11429 4669
rect -11366 4652 -11349 4669
rect -11726 4652 -11709 4669
rect -11406 4652 -11389 4669
rect -11646 4652 -11629 4669
rect -11486 4652 -11469 4669
rect -11646 4652 -11629 4669
rect -11406 4652 -11389 4669
rect -11726 4652 -11709 4669
rect -11486 4652 -11469 4669
rect -11566 4652 -11549 4669
rect -11766 4652 -11749 4669
rect -11526 4652 -11509 4669
rect -11286 4652 -11269 4669
rect -11486 4652 -11469 4669
rect -11326 4652 -11309 4669
rect -11366 4652 -11349 4669
rect -11566 4652 -11549 4669
rect -11606 4652 -11589 4669
rect -11686 4652 -11669 4669
rect -16646 4652 -16629 4669
rect -16686 4652 -16669 4669
rect -16726 4652 -16709 4669
rect -16766 4652 -16749 4669
rect -16566 4652 -16549 4669
rect -16606 4652 -16589 4669
rect -16646 4652 -16629 4669
rect -16686 4652 -16669 4669
rect -16726 4652 -16709 4669
rect -16766 4652 -16749 4669
rect -16566 4652 -16549 4669
rect -17126 4652 -17109 4669
rect -16646 4652 -16629 4669
rect -16566 4652 -16549 4669
rect -16766 4652 -16749 4669
rect -16606 4652 -16589 4669
rect -16926 4652 -16909 4669
rect -17006 4652 -16989 4669
rect -16686 4652 -16669 4669
rect -16846 4652 -16829 4669
rect -17086 4652 -17069 4669
rect -16766 4652 -16749 4669
rect -16566 4652 -16549 4669
rect -16886 4652 -16869 4669
rect -16846 4652 -16829 4669
rect -16726 4652 -16709 4669
rect -16886 4652 -16869 4669
rect -16966 4652 -16949 4669
rect -17046 4652 -17029 4669
rect -16806 4652 -16789 4669
rect -16646 4652 -16629 4669
rect -17046 4652 -17029 4669
rect -17046 4652 -17029 4669
rect -17086 4652 -17069 4669
rect -17126 4652 -17109 4669
rect -16806 4652 -16789 4669
rect -17006 4652 -16989 4669
rect -16806 4652 -16789 4669
rect -16846 4652 -16829 4669
rect -16886 4652 -16869 4669
rect -16926 4652 -16909 4669
rect -16966 4652 -16949 4669
rect -17006 4652 -16989 4669
rect -17046 4652 -17029 4669
rect -17086 4652 -17069 4669
rect -17126 4652 -17109 4669
rect -16606 4652 -16589 4669
rect -16726 4652 -16709 4669
rect -16806 4652 -16789 4669
rect -16846 4652 -16829 4669
rect -16886 4652 -16869 4669
rect -16926 4652 -16909 4669
rect -16926 4652 -16909 4669
rect -17086 4652 -17069 4669
rect -16966 4652 -16949 4669
rect -16686 4652 -16669 4669
rect -17006 4652 -16989 4669
rect -17126 4652 -17109 4669
rect -16966 4652 -16949 4669
rect -16606 4652 -16589 4669
rect -17486 4652 -17469 4669
rect -17686 4652 -17669 4669
rect -17166 4652 -17149 4669
rect -17726 4652 -17709 4669
rect -17566 4652 -17549 4669
rect -17486 4652 -17469 4669
rect -17406 4652 -17389 4669
rect -17286 4652 -17269 4669
rect -17446 4652 -17429 4669
rect -17446 4652 -17429 4669
rect -17606 4652 -17589 4669
rect -17566 4652 -17549 4669
rect -17646 4652 -17629 4669
rect -17326 4652 -17309 4669
rect -17726 4652 -17709 4669
rect -17526 4652 -17509 4669
rect -17246 4652 -17229 4669
rect -17326 4652 -17309 4669
rect -17166 4652 -17149 4669
rect -17286 4652 -17269 4669
rect -17526 4652 -17509 4669
rect -17646 4652 -17629 4669
rect -17206 4652 -17189 4669
rect -17406 4652 -17389 4669
rect -17606 4652 -17589 4669
rect -17366 4652 -17349 4669
rect -17206 4652 -17189 4669
rect -17366 4652 -17349 4669
rect -17246 4652 -17229 4669
rect -17246 4652 -17229 4669
rect -17526 4652 -17509 4669
rect -17286 4652 -17269 4669
rect -17566 4652 -17549 4669
rect -17246 4652 -17229 4669
rect -17286 4652 -17269 4669
rect -17326 4652 -17309 4669
rect -17366 4652 -17349 4669
rect -17406 4652 -17389 4669
rect -17446 4652 -17429 4669
rect -17486 4652 -17469 4669
rect -17526 4652 -17509 4669
rect -17566 4652 -17549 4669
rect -17606 4652 -17589 4669
rect -17646 4652 -17629 4669
rect -17686 4652 -17669 4669
rect -17726 4652 -17709 4669
rect -17326 4652 -17309 4669
rect -17606 4652 -17589 4669
rect -17366 4652 -17349 4669
rect -17646 4652 -17629 4669
rect -17166 4652 -17149 4669
rect -17206 4652 -17189 4669
rect -17166 4652 -17149 4669
rect -17206 4652 -17189 4669
rect -17406 4652 -17389 4669
rect -17686 4652 -17669 4669
rect -17446 4652 -17429 4669
rect -17726 4652 -17709 4669
rect -17486 4652 -17469 4669
rect -17686 4652 -17669 4669
rect -17766 4652 -17749 4669
rect -17766 4652 -17749 4669
rect -17806 4652 -17789 4669
rect -17846 4652 -17829 4669
rect -18046 4652 -18029 4669
rect -17806 4652 -17789 4669
rect -17926 4652 -17909 4669
rect -17846 4652 -17829 4669
rect -17886 4652 -17869 4669
rect -18086 4652 -18069 4669
rect -18126 4652 -18109 4669
rect -18326 4652 -18309 4669
rect -18126 4652 -18109 4669
rect -17766 4652 -17749 4669
rect -18166 4652 -18149 4669
rect -18126 4652 -18109 4669
rect -18206 4652 -18189 4669
rect -18166 4652 -18149 4669
rect -17886 4652 -17869 4669
rect -18286 4652 -18269 4669
rect -18246 4652 -18229 4669
rect -17966 4652 -17949 4669
rect -18286 4652 -18269 4669
rect -17806 4652 -17789 4669
rect -18006 4652 -17989 4669
rect -18246 4652 -18229 4669
rect -18326 4652 -18309 4669
rect -17926 4652 -17909 4669
rect -18206 4652 -18189 4669
rect -18166 4652 -18149 4669
rect -17806 4652 -17789 4669
rect -17926 4652 -17909 4669
rect -18246 4652 -18229 4669
rect -17886 4652 -17869 4669
rect -18086 4652 -18069 4669
rect -18006 4652 -17989 4669
rect -18326 4652 -18309 4669
rect -18126 4652 -18109 4669
rect -17966 4652 -17949 4669
rect -18046 4652 -18029 4669
rect -17926 4652 -17909 4669
rect -17886 4652 -17869 4669
rect -18206 4652 -18189 4669
rect -17966 4652 -17949 4669
rect -18046 4652 -18029 4669
rect -18246 4652 -18229 4669
rect -18006 4652 -17989 4669
rect -18286 4652 -18269 4669
rect -17966 4652 -17949 4669
rect -17766 4652 -17749 4669
rect -18286 4652 -18269 4669
rect -18166 4652 -18149 4669
rect -18046 4652 -18029 4669
rect -18006 4652 -17989 4669
rect -18086 4652 -18069 4669
rect -17846 4652 -17829 4669
rect -18326 4652 -18309 4669
rect -18206 4652 -18189 4669
rect -18086 4652 -18069 4669
rect -17846 4652 -17829 4669
rect -18846 4652 -18829 4669
rect -18766 4652 -18749 4669
rect -18566 4652 -18549 4669
rect -18686 4652 -18669 4669
rect -18646 4652 -18629 4669
rect -18406 4652 -18389 4669
rect -18886 4652 -18869 4669
rect -18806 4652 -18789 4669
rect -18606 4652 -18589 4669
rect -18446 4652 -18429 4669
rect -18366 4652 -18349 4669
rect -18606 4652 -18589 4669
rect -18406 4652 -18389 4669
rect -18726 4652 -18709 4669
rect -18486 4652 -18469 4669
rect -18486 4652 -18469 4669
rect -18846 4652 -18829 4669
rect -18646 4652 -18629 4669
rect -18526 4652 -18509 4669
rect -18926 4652 -18909 4669
rect -18806 4652 -18789 4669
rect -18446 4652 -18429 4669
rect -18926 4652 -18909 4669
rect -18886 4652 -18869 4669
rect -18766 4652 -18749 4669
rect -18686 4652 -18669 4669
rect -18526 4652 -18509 4669
rect -18566 4652 -18549 4669
rect -18726 4652 -18709 4669
rect -18766 4652 -18749 4669
rect -18806 4652 -18789 4669
rect -18366 4652 -18349 4669
rect -18846 4652 -18829 4669
rect -18886 4652 -18869 4669
rect -18926 4652 -18909 4669
rect -18686 4652 -18669 4669
rect -18726 4652 -18709 4669
rect -18766 4652 -18749 4669
rect -18806 4652 -18789 4669
rect -18846 4652 -18829 4669
rect -18886 4652 -18869 4669
rect -18926 4652 -18909 4669
rect -18366 4652 -18349 4669
rect -18406 4652 -18389 4669
rect -18446 4652 -18429 4669
rect -18406 4652 -18389 4669
rect -18486 4652 -18469 4669
rect -18526 4652 -18509 4669
rect -18446 4652 -18429 4669
rect -18566 4652 -18549 4669
rect -18606 4652 -18589 4669
rect -18486 4652 -18469 4669
rect -18646 4652 -18629 4669
rect -18526 4652 -18509 4669
rect -18566 4652 -18549 4669
rect -18606 4652 -18589 4669
rect -18646 4652 -18629 4669
rect -18686 4652 -18669 4669
rect -18726 4652 -18709 4669
rect -18366 4652 -18349 4669
rect -15366 4652 -15349 4669
rect -15366 4652 -15349 4669
rect -15366 4652 -15349 4669
rect -15366 4652 -15349 4669
rect -14766 4652 -14749 4669
rect -14766 4652 -14749 4669
rect -14766 4652 -14749 4669
rect -14766 4652 -14749 4669
rect -14646 4652 -14629 4669
rect -14246 4652 -14229 4669
rect -14286 4652 -14269 4669
rect -14446 4652 -14429 4669
rect -14726 4652 -14709 4669
rect -14606 4652 -14589 4669
rect -14686 4652 -14669 4669
rect -14726 4652 -14709 4669
rect -14326 4652 -14309 4669
rect -14206 4652 -14189 4669
rect -14366 4652 -14349 4669
rect -14486 4652 -14469 4669
rect -14486 4652 -14469 4669
rect -14566 4652 -14549 4669
rect -14686 4652 -14669 4669
rect -14566 4652 -14549 4669
rect -14246 4652 -14229 4669
rect -14486 4652 -14469 4669
rect -14406 4652 -14389 4669
rect -14286 4652 -14269 4669
rect -14366 4652 -14349 4669
rect -14526 4652 -14509 4669
rect -14326 4652 -14309 4669
rect -14286 4652 -14269 4669
rect -14646 4652 -14629 4669
rect -14726 4652 -14709 4669
rect -14446 4652 -14429 4669
rect -14606 4652 -14589 4669
rect -14646 4652 -14629 4669
rect -14646 4652 -14629 4669
rect -14486 4652 -14469 4669
rect -14366 4652 -14349 4669
rect -14526 4652 -14509 4669
rect -14686 4652 -14669 4669
rect -14406 4652 -14389 4669
rect -14566 4652 -14549 4669
rect -14326 4652 -14309 4669
rect -14246 4652 -14229 4669
rect -14286 4652 -14269 4669
rect -14406 4652 -14389 4669
rect -14446 4652 -14429 4669
rect -14606 4652 -14589 4669
rect -14206 4652 -14189 4669
rect -14526 4652 -14509 4669
rect -14446 4652 -14429 4669
rect -14326 4652 -14309 4669
rect -14566 4652 -14549 4669
rect -14406 4652 -14389 4669
rect -14206 4652 -14189 4669
rect -14366 4652 -14349 4669
rect -14526 4652 -14509 4669
rect -14246 4652 -14229 4669
rect -14606 4652 -14589 4669
rect -14686 4652 -14669 4669
rect -14206 4652 -14189 4669
rect -14726 4652 -14709 4669
rect -15166 4652 -15149 4669
rect -15206 4652 -15189 4669
rect -15246 4652 -15229 4669
rect -15286 4652 -15269 4669
rect -15326 4652 -15309 4669
rect -14846 4652 -14829 4669
rect -15166 4652 -15149 4669
rect -15206 4652 -15189 4669
rect -14886 4652 -14869 4669
rect -14926 4652 -14909 4669
rect -14966 4652 -14949 4669
rect -15006 4652 -14989 4669
rect -15046 4652 -15029 4669
rect -15006 4652 -14989 4669
rect -14806 4652 -14789 4669
rect -14846 4652 -14829 4669
rect -14886 4652 -14869 4669
rect -14926 4652 -14909 4669
rect -14966 4652 -14949 4669
rect -15006 4652 -14989 4669
rect -15046 4652 -15029 4669
rect -15086 4652 -15069 4669
rect -15246 4652 -15229 4669
rect -14806 4652 -14789 4669
rect -15286 4652 -15269 4669
rect -14846 4652 -14829 4669
rect -15326 4652 -15309 4669
rect -15326 4652 -15309 4669
rect -15046 4652 -15029 4669
rect -15166 4652 -15149 4669
rect -15006 4652 -14989 4669
rect -15126 4652 -15109 4669
rect -15286 4652 -15269 4669
rect -15126 4652 -15109 4669
rect -14806 4652 -14789 4669
rect -15206 4652 -15189 4669
rect -15086 4652 -15069 4669
rect -15326 4652 -15309 4669
rect -14846 4652 -14829 4669
rect -15086 4652 -15069 4669
rect -15126 4652 -15109 4669
rect -15246 4652 -15229 4669
rect -14886 4652 -14869 4669
rect -14886 4652 -14869 4669
rect -15166 4652 -15149 4669
rect -14926 4652 -14909 4669
rect -14806 4652 -14789 4669
rect -15206 4652 -15189 4669
rect -14966 4652 -14949 4669
rect -15046 4652 -15029 4669
rect -14926 4652 -14909 4669
rect -15286 4652 -15269 4669
rect -15246 4652 -15229 4669
rect -15086 4652 -15069 4669
rect -14966 4652 -14949 4669
rect -15126 4652 -15109 4669
rect -15966 4652 -15949 4669
rect -15966 4652 -15949 4669
rect -15966 4652 -15949 4669
rect -15966 4652 -15949 4669
rect -15806 4652 -15789 4669
rect -15766 4652 -15749 4669
rect -15686 4652 -15669 4669
rect -15726 4652 -15709 4669
rect -15406 4652 -15389 4669
rect -15846 4652 -15829 4669
rect -15446 4652 -15429 4669
rect -15766 4652 -15749 4669
rect -15526 4652 -15509 4669
rect -15486 4652 -15469 4669
rect -15526 4652 -15509 4669
rect -15606 4652 -15589 4669
rect -15926 4652 -15909 4669
rect -15446 4652 -15429 4669
rect -15526 4652 -15509 4669
rect -15526 4652 -15509 4669
rect -15406 4652 -15389 4669
rect -15566 4652 -15549 4669
rect -15486 4652 -15469 4669
rect -15606 4652 -15589 4669
rect -15646 4652 -15629 4669
rect -15686 4652 -15669 4669
rect -15926 4652 -15909 4669
rect -15726 4652 -15709 4669
rect -15886 4652 -15869 4669
rect -15566 4652 -15549 4669
rect -15446 4652 -15429 4669
rect -15806 4652 -15789 4669
rect -15766 4652 -15749 4669
rect -15566 4652 -15549 4669
rect -15846 4652 -15829 4669
rect -15606 4652 -15589 4669
rect -15726 4652 -15709 4669
rect -15646 4652 -15629 4669
rect -15766 4652 -15749 4669
rect -15806 4652 -15789 4669
rect -15406 4652 -15389 4669
rect -15886 4652 -15869 4669
rect -15846 4652 -15829 4669
rect -15446 4652 -15429 4669
rect -15846 4652 -15829 4669
rect -15726 4652 -15709 4669
rect -15566 4652 -15549 4669
rect -15926 4652 -15909 4669
rect -15486 4652 -15469 4669
rect -15686 4652 -15669 4669
rect -15806 4652 -15789 4669
rect -15406 4652 -15389 4669
rect -15606 4652 -15589 4669
rect -15886 4652 -15869 4669
rect -15646 4652 -15629 4669
rect -15486 4652 -15469 4669
rect -15886 4652 -15869 4669
rect -15686 4652 -15669 4669
rect -15926 4652 -15909 4669
rect -15646 4652 -15629 4669
rect -16166 4652 -16149 4669
rect -16006 4652 -15989 4669
rect -16526 4652 -16509 4669
rect -16046 4652 -16029 4669
rect -16006 4652 -15989 4669
rect -16086 4652 -16069 4669
rect -16366 4652 -16349 4669
rect -16126 4652 -16109 4669
rect -16166 4652 -16149 4669
rect -16206 4652 -16189 4669
rect -16006 4652 -15989 4669
rect -16246 4652 -16229 4669
rect -16286 4652 -16269 4669
rect -16246 4652 -16229 4669
rect -16326 4652 -16309 4669
rect -16366 4652 -16349 4669
rect -16526 4652 -16509 4669
rect -16086 4652 -16069 4669
rect -16126 4652 -16109 4669
rect -16326 4652 -16309 4669
rect -16406 4652 -16389 4669
rect -16206 4652 -16189 4669
rect -16206 4652 -16189 4669
rect -16486 4652 -16469 4669
rect -16486 4652 -16469 4669
rect -16006 4652 -15989 4669
rect -16446 4652 -16429 4669
rect -16286 4652 -16269 4669
rect -16166 4652 -16149 4669
rect -16246 4652 -16229 4669
rect -16046 4652 -16029 4669
rect -16166 4652 -16149 4669
rect -16446 4652 -16429 4669
rect -16286 4652 -16269 4669
rect -16366 4652 -16349 4669
rect -16406 4652 -16389 4669
rect -16526 4652 -16509 4669
rect -16446 4652 -16429 4669
rect -16286 4652 -16269 4669
rect -16326 4652 -16309 4669
rect -16406 4652 -16389 4669
rect -16326 4652 -16309 4669
rect -16486 4652 -16469 4669
rect -16206 4652 -16189 4669
rect -16126 4652 -16109 4669
rect -16046 4652 -16029 4669
rect -16086 4652 -16069 4669
rect -16366 4652 -16349 4669
rect -16046 4652 -16029 4669
rect -16246 4652 -16229 4669
rect -16086 4652 -16069 4669
rect -16406 4652 -16389 4669
rect -16126 4652 -16109 4669
rect -16446 4652 -16429 4669
rect -16486 4652 -16469 4669
rect -16526 4652 -16509 4669
rect -18846 3163 -18829 3180
rect -18486 3163 -18469 3180
rect -18686 3163 -18669 3180
rect -18726 3163 -18709 3180
rect -18446 3163 -18429 3180
rect -18446 3163 -18429 3180
rect -18886 3163 -18869 3180
rect -18566 3163 -18549 3180
rect -18486 3163 -18469 3180
rect -18886 3163 -18869 3180
rect -18886 3163 -18869 3180
rect -18606 3163 -18589 3180
rect -18766 3163 -18749 3180
rect -18686 3163 -18669 3180
rect -18566 3163 -18549 3180
rect -18486 3163 -18469 3180
rect -18646 3163 -18629 3180
rect -18606 3163 -18589 3180
rect -18406 3163 -18389 3180
rect -18926 3163 -18909 3180
rect -18926 3163 -18909 3180
rect -18406 3163 -18389 3180
rect -18686 3163 -18669 3180
rect -18726 3163 -18709 3180
rect -18446 3163 -18429 3180
rect -18606 3163 -18589 3180
rect -18726 3163 -18709 3180
rect -18406 3163 -18389 3180
rect -18806 3163 -18789 3180
rect -18566 3163 -18549 3180
rect -18806 3163 -18789 3180
rect -18526 3163 -18509 3180
rect -18846 3163 -18829 3180
rect -18446 3163 -18429 3180
rect -18766 3163 -18749 3180
rect -18646 3163 -18629 3180
rect -18846 3163 -18829 3180
rect -18926 3163 -18909 3180
rect -18686 3163 -18669 3180
rect -18646 3163 -18629 3180
rect -18926 3163 -18909 3180
rect -18886 3163 -18869 3180
rect -18766 3163 -18749 3180
rect -18486 3163 -18469 3180
rect -18766 3163 -18749 3180
rect -18726 3163 -18709 3180
rect -18526 3163 -18509 3180
rect -18526 3163 -18509 3180
rect -18846 3163 -18829 3180
rect -18526 3163 -18509 3180
rect -18566 3163 -18549 3180
rect -18646 3163 -18629 3180
rect -18406 3163 -18389 3180
rect -18606 3163 -18589 3180
rect -18806 3163 -18789 3180
rect -18806 3163 -18789 3180
rect -14366 3163 -14349 3180
rect -14526 3163 -14509 3180
rect -14206 3163 -14189 3180
rect -14326 3163 -14309 3180
rect -14286 3163 -14269 3180
rect -14326 3163 -14309 3180
rect -14246 3163 -14229 3180
rect -14486 3163 -14469 3180
rect -14286 3163 -14269 3180
rect -14566 3163 -14549 3180
rect -14566 3163 -14549 3180
rect -14406 3163 -14389 3180
rect -14286 3163 -14269 3180
rect -14406 3163 -14389 3180
rect -14366 3163 -14349 3180
rect -14246 3163 -14229 3180
rect -14446 3163 -14429 3180
rect -14446 3163 -14429 3180
rect -14326 3163 -14309 3180
rect -14486 3163 -14469 3180
rect -14606 3163 -14589 3180
rect -14206 3163 -14189 3180
rect -14246 3163 -14229 3180
rect -14486 3163 -14469 3180
rect -14206 3163 -14189 3180
rect -14606 3163 -14589 3180
rect -14526 3163 -14509 3180
rect -14406 3163 -14389 3180
rect -14606 3163 -14589 3180
rect -14486 3163 -14469 3180
rect -14566 3163 -14549 3180
rect -14606 3163 -14589 3180
rect -14366 3163 -14349 3180
rect -14446 3163 -14429 3180
rect -14246 3163 -14229 3180
rect -14206 3163 -14189 3180
rect -14526 3163 -14509 3180
rect -14526 3163 -14509 3180
rect -14286 3163 -14269 3180
rect -14446 3163 -14429 3180
rect -14366 3163 -14349 3180
rect -14406 3163 -14389 3180
rect -14566 3163 -14549 3180
rect -14326 3163 -14309 3180
rect -15166 3163 -15149 3180
rect -15166 3163 -15149 3180
rect -15166 3163 -15149 3180
rect -15166 3163 -15149 3180
rect -15126 3163 -15109 3180
rect -14806 3163 -14789 3180
rect -15086 3163 -15069 3180
rect -14846 3163 -14829 3180
rect -15086 3163 -15069 3180
rect -14766 3163 -14749 3180
rect -15126 3163 -15109 3180
rect -14766 3163 -14749 3180
rect -14886 3163 -14869 3180
rect -14886 3163 -14869 3180
rect -14766 3163 -14749 3180
rect -15046 3163 -15029 3180
rect -14926 3163 -14909 3180
rect -14766 3163 -14749 3180
rect -14806 3163 -14789 3180
rect -15126 3163 -15109 3180
rect -14966 3163 -14949 3180
rect -15006 3163 -14989 3180
rect -15046 3163 -15029 3180
rect -14926 3163 -14909 3180
rect -15086 3163 -15069 3180
rect -14966 3163 -14949 3180
rect -14726 3163 -14709 3180
rect -14646 3163 -14629 3180
rect -14846 3163 -14829 3180
rect -15126 3163 -15109 3180
rect -14726 3163 -14709 3180
rect -14686 3163 -14669 3180
rect -14886 3163 -14869 3180
rect -14726 3163 -14709 3180
rect -14926 3163 -14909 3180
rect -14966 3163 -14949 3180
rect -15006 3163 -14989 3180
rect -15046 3163 -15029 3180
rect -15006 3163 -14989 3180
rect -14686 3163 -14669 3180
rect -14806 3163 -14789 3180
rect -14846 3163 -14829 3180
rect -14886 3163 -14869 3180
rect -14926 3163 -14909 3180
rect -14966 3163 -14949 3180
rect -15006 3163 -14989 3180
rect -15046 3163 -15029 3180
rect -14646 3163 -14629 3180
rect -14726 3163 -14709 3180
rect -15086 3163 -15069 3180
rect -14646 3163 -14629 3180
rect -14806 3163 -14789 3180
rect -14646 3163 -14629 3180
rect -14686 3163 -14669 3180
rect -14846 3163 -14829 3180
rect -14686 3163 -14669 3180
rect -15286 3163 -15269 3180
rect -15606 3163 -15589 3180
rect -15406 3163 -15389 3180
rect -15326 3163 -15309 3180
rect -15686 3163 -15669 3180
rect -15246 3163 -15229 3180
rect -15286 3163 -15269 3180
rect -15566 3163 -15549 3180
rect -15366 3163 -15349 3180
rect -15206 3163 -15189 3180
rect -15406 3163 -15389 3180
rect -15446 3163 -15429 3180
rect -15566 3163 -15549 3180
rect -15686 3163 -15669 3180
rect -15326 3163 -15309 3180
rect -15566 3163 -15549 3180
rect -15206 3163 -15189 3180
rect -15686 3163 -15669 3180
rect -15486 3163 -15469 3180
rect -15446 3163 -15429 3180
rect -15486 3163 -15469 3180
rect -15566 3163 -15549 3180
rect -15366 3163 -15349 3180
rect -15366 3163 -15349 3180
rect -15486 3163 -15469 3180
rect -15646 3163 -15629 3180
rect -15606 3163 -15589 3180
rect -15406 3163 -15389 3180
rect -15206 3163 -15189 3180
rect -15606 3163 -15589 3180
rect -15606 3163 -15589 3180
rect -15526 3163 -15509 3180
rect -15646 3163 -15629 3180
rect -15326 3163 -15309 3180
rect -15526 3163 -15509 3180
rect -15646 3163 -15629 3180
rect -15446 3163 -15429 3180
rect -15526 3163 -15509 3180
rect -15206 3163 -15189 3180
rect -15406 3163 -15389 3180
rect -15286 3163 -15269 3180
rect -15246 3163 -15229 3180
rect -15646 3163 -15629 3180
rect -15686 3163 -15669 3180
rect -15246 3163 -15229 3180
rect -15246 3163 -15229 3180
rect -15286 3163 -15269 3180
rect -15446 3163 -15429 3180
rect -15486 3163 -15469 3180
rect -15526 3163 -15509 3180
rect -15366 3163 -15349 3180
rect -15326 3163 -15309 3180
rect -16246 3163 -16229 3180
rect -16246 3163 -16229 3180
rect -16246 3163 -16229 3180
rect -16246 3163 -16229 3180
rect -15806 3163 -15789 3180
rect -16126 3163 -16109 3180
rect -15806 3163 -15789 3180
rect -15926 3163 -15909 3180
rect -16126 3163 -16109 3180
rect -16206 3163 -16189 3180
rect -16006 3163 -15989 3180
rect -15766 3163 -15749 3180
rect -15886 3163 -15869 3180
rect -16046 3163 -16029 3180
rect -15926 3163 -15909 3180
rect -15726 3163 -15709 3180
rect -15966 3163 -15949 3180
rect -15846 3163 -15829 3180
rect -16166 3163 -16149 3180
rect -15726 3163 -15709 3180
rect -15966 3163 -15949 3180
rect -16086 3163 -16069 3180
rect -16046 3163 -16029 3180
rect -16166 3163 -16149 3180
rect -16206 3163 -16189 3180
rect -15726 3163 -15709 3180
rect -16086 3163 -16069 3180
rect -15926 3163 -15909 3180
rect -16166 3163 -16149 3180
rect -15846 3163 -15829 3180
rect -15766 3163 -15749 3180
rect -16126 3163 -16109 3180
rect -16006 3163 -15989 3180
rect -16086 3163 -16069 3180
rect -15806 3163 -15789 3180
rect -15966 3163 -15949 3180
rect -16086 3163 -16069 3180
rect -15726 3163 -15709 3180
rect -16006 3163 -15989 3180
rect -16126 3163 -16109 3180
rect -16206 3163 -16189 3180
rect -15806 3163 -15789 3180
rect -15886 3163 -15869 3180
rect -15926 3163 -15909 3180
rect -15766 3163 -15749 3180
rect -15846 3163 -15829 3180
rect -15886 3163 -15869 3180
rect -16166 3163 -16149 3180
rect -16046 3163 -16029 3180
rect -16006 3163 -15989 3180
rect -16206 3163 -16189 3180
rect -15766 3163 -15749 3180
rect -15846 3163 -15829 3180
rect -15966 3163 -15949 3180
rect -16046 3163 -16029 3180
rect -15886 3163 -15869 3180
rect -16406 3163 -16389 3180
rect -16446 3163 -16429 3180
rect -16766 3163 -16749 3180
rect -16526 3163 -16509 3180
rect -16486 3163 -16469 3180
rect -16486 3163 -16469 3180
rect -16566 3163 -16549 3180
rect -16286 3163 -16269 3180
rect -16326 3163 -16309 3180
rect -16726 3163 -16709 3180
rect -16286 3163 -16269 3180
rect -16406 3163 -16389 3180
rect -16326 3163 -16309 3180
rect -16646 3163 -16629 3180
rect -16366 3163 -16349 3180
rect -16526 3163 -16509 3180
rect -16646 3163 -16629 3180
rect -16606 3163 -16589 3180
rect -16766 3163 -16749 3180
rect -16566 3163 -16549 3180
rect -16366 3163 -16349 3180
rect -16606 3163 -16589 3180
rect -16366 3163 -16349 3180
rect -16566 3163 -16549 3180
rect -16766 3163 -16749 3180
rect -16326 3163 -16309 3180
rect -16446 3163 -16429 3180
rect -16606 3163 -16589 3180
rect -16726 3163 -16709 3180
rect -16366 3163 -16349 3180
rect -16606 3163 -16589 3180
rect -16526 3163 -16509 3180
rect -16486 3163 -16469 3180
rect -16406 3163 -16389 3180
rect -16526 3163 -16509 3180
rect -16446 3163 -16429 3180
rect -16686 3163 -16669 3180
rect -16486 3163 -16469 3180
rect -16646 3163 -16629 3180
rect -16286 3163 -16269 3180
rect -16646 3163 -16629 3180
rect -16726 3163 -16709 3180
rect -16326 3163 -16309 3180
rect -16766 3163 -16749 3180
rect -16686 3163 -16669 3180
rect -16446 3163 -16429 3180
rect -16286 3163 -16269 3180
rect -16406 3163 -16389 3180
rect -16566 3163 -16549 3180
rect -16686 3163 -16669 3180
rect -16726 3163 -16709 3180
rect -16686 3163 -16669 3180
rect -16806 3163 -16789 3180
rect -17166 3163 -17149 3180
rect -17206 3163 -17189 3180
rect -17126 3163 -17109 3180
rect -17046 3163 -17029 3180
rect -16846 3163 -16829 3180
rect -17246 3163 -17229 3180
rect -16926 3163 -16909 3180
rect -17166 3163 -17149 3180
rect -17046 3163 -17029 3180
rect -16846 3163 -16829 3180
rect -17086 3163 -17069 3180
rect -17286 3163 -17269 3180
rect -17006 3163 -16989 3180
rect -17286 3163 -17269 3180
rect -16886 3163 -16869 3180
rect -17046 3163 -17029 3180
rect -17206 3163 -17189 3180
rect -17006 3163 -16989 3180
rect -16966 3163 -16949 3180
rect -17286 3163 -17269 3180
rect -16886 3163 -16869 3180
rect -17246 3163 -17229 3180
rect -16886 3163 -16869 3180
rect -17206 3163 -17189 3180
rect -16806 3163 -16789 3180
rect -17086 3163 -17069 3180
rect -17126 3163 -17109 3180
rect -16966 3163 -16949 3180
rect -17126 3163 -17109 3180
rect -16926 3163 -16909 3180
rect -16846 3163 -16829 3180
rect -17286 3163 -17269 3180
rect -17006 3163 -16989 3180
rect -16886 3163 -16869 3180
rect -16966 3163 -16949 3180
rect -17126 3163 -17109 3180
rect -16806 3163 -16789 3180
rect -16926 3163 -16909 3180
rect -17006 3163 -16989 3180
rect -16966 3163 -16949 3180
rect -17046 3163 -17029 3180
rect -17086 3163 -17069 3180
rect -17246 3163 -17229 3180
rect -17166 3163 -17149 3180
rect -16846 3163 -16829 3180
rect -17086 3163 -17069 3180
rect -16806 3163 -16789 3180
rect -16926 3163 -16909 3180
rect -17206 3163 -17189 3180
rect -17166 3163 -17149 3180
rect -17246 3163 -17229 3180
rect -17566 3163 -17549 3180
rect -17846 3163 -17829 3180
rect -17446 3163 -17429 3180
rect -17766 3163 -17749 3180
rect -17686 3163 -17669 3180
rect -17606 3163 -17589 3180
rect -17686 3163 -17669 3180
rect -17726 3163 -17709 3180
rect -17486 3163 -17469 3180
rect -17406 3163 -17389 3180
rect -17486 3163 -17469 3180
rect -17566 3163 -17549 3180
rect -17486 3163 -17469 3180
rect -17526 3163 -17509 3180
rect -17646 3163 -17629 3180
rect -17326 3163 -17309 3180
rect -17726 3163 -17709 3180
rect -17806 3163 -17789 3180
rect -17766 3163 -17749 3180
rect -17526 3163 -17509 3180
rect -17526 3163 -17509 3180
rect -17566 3163 -17549 3180
rect -17606 3163 -17589 3180
rect -17766 3163 -17749 3180
rect -17326 3163 -17309 3180
rect -17846 3163 -17829 3180
rect -17686 3163 -17669 3180
rect -17366 3163 -17349 3180
rect -17486 3163 -17469 3180
rect -17846 3163 -17829 3180
rect -17766 3163 -17749 3180
rect -17726 3163 -17709 3180
rect -17366 3163 -17349 3180
rect -17566 3163 -17549 3180
rect -17406 3163 -17389 3180
rect -17526 3163 -17509 3180
rect -17646 3163 -17629 3180
rect -17446 3163 -17429 3180
rect -17686 3163 -17669 3180
rect -17326 3163 -17309 3180
rect -17406 3163 -17389 3180
rect -17446 3163 -17429 3180
rect -17606 3163 -17589 3180
rect -17606 3163 -17589 3180
rect -17806 3163 -17789 3180
rect -17406 3163 -17389 3180
rect -17806 3163 -17789 3180
rect -17726 3163 -17709 3180
rect -17326 3163 -17309 3180
rect -17646 3163 -17629 3180
rect -17366 3163 -17349 3180
rect -17646 3163 -17629 3180
rect -17446 3163 -17429 3180
rect -17806 3163 -17789 3180
rect -17366 3163 -17349 3180
rect -17846 3163 -17829 3180
rect -18166 3163 -18149 3180
rect -17926 3163 -17909 3180
rect -17966 3163 -17949 3180
rect -18006 3163 -17989 3180
rect -17886 3163 -17869 3180
rect -18206 3163 -18189 3180
rect -17926 3163 -17909 3180
rect -18046 3163 -18029 3180
rect -18326 3163 -18309 3180
rect -18286 3163 -18269 3180
rect -18286 3163 -18269 3180
rect -18366 3163 -18349 3180
rect -18166 3163 -18149 3180
rect -18006 3163 -17989 3180
rect -18126 3163 -18109 3180
rect -18046 3163 -18029 3180
rect -18366 3163 -18349 3180
rect -17926 3163 -17909 3180
rect -18046 3163 -18029 3180
rect -18246 3163 -18229 3180
rect -18246 3163 -18229 3180
rect -17926 3163 -17909 3180
rect -18366 3163 -18349 3180
rect -18126 3163 -18109 3180
rect -18126 3163 -18109 3180
rect -17966 3163 -17949 3180
rect -18326 3163 -18309 3180
rect -18206 3163 -18189 3180
rect -18246 3163 -18229 3180
rect -18086 3163 -18069 3180
rect -17966 3163 -17949 3180
rect -18246 3163 -18229 3180
rect -17966 3163 -17949 3180
rect -18326 3163 -18309 3180
rect -18326 3163 -18309 3180
rect -17886 3163 -17869 3180
rect -18046 3163 -18029 3180
rect -18126 3163 -18109 3180
rect -18206 3163 -18189 3180
rect -18286 3163 -18269 3180
rect -17886 3163 -17869 3180
rect -18206 3163 -18189 3180
rect -18166 3163 -18149 3180
rect -18086 3163 -18069 3180
rect -18286 3163 -18269 3180
rect -17886 3163 -17869 3180
rect -18006 3163 -17989 3180
rect -18006 3163 -17989 3180
rect -18366 3163 -18349 3180
rect -18086 3163 -18069 3180
rect -18086 3163 -18069 3180
rect -18166 3163 -18149 3180
rect -17373 2394 -17356 2411
rect -16653 2394 -16636 2411
rect -16613 2394 -16596 2411
rect -17213 2394 -17196 2411
rect -17253 2394 -17236 2411
rect -16813 2394 -16796 2411
rect -17413 2394 -17396 2411
rect -16853 2394 -16836 2411
rect -17453 2394 -17436 2411
rect -16853 2394 -16836 2411
rect -17133 2394 -17116 2411
rect -17413 2394 -17396 2411
rect -17453 2394 -17436 2411
rect -17293 2394 -17276 2411
rect -16573 2394 -16556 2411
rect -16893 2394 -16876 2411
rect -17293 2394 -17276 2411
rect -16573 2394 -16556 2411
rect -16693 2394 -16676 2411
rect -17253 2394 -17236 2411
rect -16693 2394 -16676 2411
rect -16933 2394 -16916 2411
rect -17173 2394 -17156 2411
rect -16773 2394 -16756 2411
rect -17053 2394 -17036 2411
rect -16973 2394 -16956 2411
rect -17333 2394 -17316 2411
rect -17173 2394 -17156 2411
rect -16933 2394 -16916 2411
rect -17013 2394 -16996 2411
rect -17333 2394 -17316 2411
rect -17213 2394 -17196 2411
rect -17013 2394 -16996 2411
rect -16893 2394 -16876 2411
rect -17133 2394 -17116 2411
rect -17093 2394 -17076 2411
rect -17053 2394 -17036 2411
rect -16773 2394 -16756 2411
rect -16613 2394 -16596 2411
rect -16813 2394 -16796 2411
rect -16973 2394 -16956 2411
rect -16653 2394 -16636 2411
rect -17373 2394 -17356 2411
rect -16733 2394 -16716 2411
rect -17093 2394 -17076 2411
rect -16733 2394 -16716 2411
rect -15373 2394 -15356 2411
rect -15373 2394 -15356 2411
rect -16053 2394 -16036 2411
rect -15493 2394 -15476 2411
rect -15693 2394 -15676 2411
rect -16373 2394 -16356 2411
rect -15453 2394 -15436 2411
rect -15973 2394 -15956 2411
rect -15853 2394 -15836 2411
rect -16093 2394 -16076 2411
rect -15893 2394 -15876 2411
rect -15533 2394 -15516 2411
rect -16133 2394 -16116 2411
rect -15733 2394 -15716 2411
rect -16253 2394 -16236 2411
rect -15773 2394 -15756 2411
rect -15893 2394 -15876 2411
rect -16133 2394 -16116 2411
rect -15573 2394 -15556 2411
rect -16293 2394 -16276 2411
rect -15493 2394 -15476 2411
rect -16173 2394 -16156 2411
rect -16333 2394 -16316 2411
rect -15933 2394 -15916 2411
rect -16173 2394 -16156 2411
rect -15573 2394 -15556 2411
rect -15853 2394 -15836 2411
rect -16373 2394 -16356 2411
rect -16093 2394 -16076 2411
rect -15413 2394 -15396 2411
rect -15613 2394 -15596 2411
rect -15613 2394 -15596 2411
rect -16013 2394 -15996 2411
rect -16213 2394 -16196 2411
rect -15653 2394 -15636 2411
rect -15413 2394 -15396 2411
rect -15813 2394 -15796 2411
rect -15693 2394 -15676 2411
rect -15973 2394 -15956 2411
rect -15813 2394 -15796 2411
rect -15453 2394 -15436 2411
rect -15733 2394 -15716 2411
rect -16253 2394 -16236 2411
rect -15533 2394 -15516 2411
rect -15773 2394 -15756 2411
rect -16013 2394 -15996 2411
rect -15933 2394 -15916 2411
rect -16213 2394 -16196 2411
rect -16293 2394 -16276 2411
rect -15653 2394 -15636 2411
rect -16053 2394 -16036 2411
rect -16533 2394 -16516 2411
rect -16493 2394 -16476 2411
rect -16413 2394 -16396 2411
rect -16533 2394 -16516 2411
rect -16413 2394 -16396 2411
rect -16453 2394 -16436 2411
rect -16453 2394 -16436 2411
rect -16493 2394 -16476 2411
rect -16333 2394 -16316 2411
rect -14693 2394 -14676 2411
rect -15173 2394 -15156 2411
rect -14373 2394 -14356 2411
rect -14213 2394 -14196 2411
rect -14213 2394 -14196 2411
rect -14893 2394 -14876 2411
rect -15293 2394 -15276 2411
rect -14733 2394 -14716 2411
rect -14253 2394 -14236 2411
rect -14373 2394 -14356 2411
rect -14573 2394 -14556 2411
rect -15173 2394 -15156 2411
rect -14413 2394 -14396 2411
rect -15213 2394 -15196 2411
rect -14493 2394 -14476 2411
rect -14333 2394 -14316 2411
rect -14333 2394 -14316 2411
rect -14853 2394 -14836 2411
rect -15333 2394 -15316 2411
rect -15013 2394 -14996 2411
rect -15253 2394 -15236 2411
rect -14933 2394 -14916 2411
rect -14813 2394 -14796 2411
rect -14733 2394 -14716 2411
rect -14493 2394 -14476 2411
rect -14653 2394 -14636 2411
rect -15253 2394 -15236 2411
rect -14453 2394 -14436 2411
rect -14933 2394 -14916 2411
rect -15333 2394 -15316 2411
rect -15293 2394 -15276 2411
rect -14533 2394 -14516 2411
rect -14813 2394 -14796 2411
rect -14893 2394 -14876 2411
rect -15013 2394 -14996 2411
rect -15053 2394 -15036 2411
rect -15053 2394 -15036 2411
rect -14773 2394 -14756 2411
rect -14613 2394 -14596 2411
rect -14973 2394 -14956 2411
rect -14573 2394 -14556 2411
rect -14853 2394 -14836 2411
rect -14653 2394 -14636 2411
rect -14693 2394 -14676 2411
rect -14293 2394 -14276 2411
rect -15093 2394 -15076 2411
rect -15133 2394 -15116 2411
rect -15093 2394 -15076 2411
rect -14253 2394 -14236 2411
rect -14413 2394 -14396 2411
rect -14973 2394 -14956 2411
rect -14293 2394 -14276 2411
rect -15133 2394 -15116 2411
rect -14773 2394 -14756 2411
rect -14533 2394 -14516 2411
rect -14613 2394 -14596 2411
rect -14453 2394 -14436 2411
rect -15213 2394 -15196 2411
rect -10605 3163 -10588 3180
rect -10605 3163 -10588 3180
rect -10605 3163 -10588 3180
rect -10605 3163 -10588 3180
rect -10485 3163 -10468 3180
rect -10525 3163 -10508 3180
rect -10565 3163 -10548 3180
rect -10325 3163 -10308 3180
rect -10365 3163 -10348 3180
rect -10405 3163 -10388 3180
rect -10445 3163 -10428 3180
rect -10485 3163 -10468 3180
rect -10525 3163 -10508 3180
rect -10565 3163 -10548 3180
rect -10325 3163 -10308 3180
rect -10365 3163 -10348 3180
rect -10405 3163 -10388 3180
rect -10445 3163 -10428 3180
rect -10565 3163 -10548 3180
rect -10325 3163 -10308 3180
rect -10365 3163 -10348 3180
rect -10405 3163 -10388 3180
rect -10445 3163 -10428 3180
rect -10485 3163 -10468 3180
rect -10525 3163 -10508 3180
rect -10565 3163 -10548 3180
rect -10365 3163 -10348 3180
rect -10325 3163 -10308 3180
rect -10445 3163 -10428 3180
rect -10645 3163 -10628 3180
rect -10485 3163 -10468 3180
rect -10525 3163 -10508 3180
rect -10685 3163 -10668 3180
rect -10725 3163 -10708 3180
rect -10405 3163 -10388 3180
rect -10765 3163 -10748 3180
rect -11045 3163 -11028 3180
rect -11045 3163 -11028 3180
rect -11325 3163 -11308 3180
rect -11365 3163 -11348 3180
rect -11325 3163 -11308 3180
rect -11245 3163 -11228 3180
rect -11125 3163 -11108 3180
rect -10925 3163 -10908 3180
rect -10885 3163 -10868 3180
rect -11005 3163 -10988 3180
rect -11125 3163 -11108 3180
rect -11365 3163 -11348 3180
rect -11245 3163 -11228 3180
rect -11125 3163 -11108 3180
rect -11285 3163 -11268 3180
rect -10965 3163 -10948 3180
rect -11085 3163 -11068 3180
rect -10885 3163 -10868 3180
rect -10885 3163 -10868 3180
rect -10925 3163 -10908 3180
rect -11165 3163 -11148 3180
rect -10965 3163 -10948 3180
rect -10925 3163 -10908 3180
rect -10925 3163 -10908 3180
rect -11205 3163 -11188 3180
rect -11245 3163 -11228 3180
rect -11205 3163 -11188 3180
rect -11085 3163 -11068 3180
rect -11325 3163 -11308 3180
rect -11285 3163 -11268 3180
rect -10965 3163 -10948 3180
rect -11205 3163 -11188 3180
rect -11285 3163 -11268 3180
rect -11205 3163 -11188 3180
rect -11325 3163 -11308 3180
rect -11085 3163 -11068 3180
rect -11005 3163 -10988 3180
rect -11365 3163 -11348 3180
rect -10965 3163 -10948 3180
rect -11165 3163 -11148 3180
rect -11045 3163 -11028 3180
rect -11125 3163 -11108 3180
rect -11285 3163 -11268 3180
rect -11365 3163 -11348 3180
rect -11045 3163 -11028 3180
rect -11165 3163 -11148 3180
rect -11245 3163 -11228 3180
rect -11005 3163 -10988 3180
rect -11005 3163 -10988 3180
rect -10885 3163 -10868 3180
rect -11085 3163 -11068 3180
rect -11165 3163 -11148 3180
rect -11925 3163 -11908 3180
rect -11925 3163 -11908 3180
rect -11925 3163 -11908 3180
rect -11925 3163 -11908 3180
rect -11765 3163 -11748 3180
rect -11525 3163 -11508 3180
rect -11605 3163 -11588 3180
rect -11685 3163 -11668 3180
rect -11685 3163 -11668 3180
rect -11445 3163 -11428 3180
rect -11445 3163 -11428 3180
rect -11805 3163 -11788 3180
rect -11725 3163 -11708 3180
rect -11445 3163 -11428 3180
rect -11805 3163 -11788 3180
rect -11405 3163 -11388 3180
rect -11845 3163 -11828 3180
rect -11765 3163 -11748 3180
rect -11645 3163 -11628 3180
rect -11845 3163 -11828 3180
rect -11485 3163 -11468 3180
rect -11485 3163 -11468 3180
rect -11525 3163 -11508 3180
rect -11645 3163 -11628 3180
rect -11405 3163 -11388 3180
rect -11805 3163 -11788 3180
rect -11845 3163 -11828 3180
rect -11725 3163 -11708 3180
rect -11885 3163 -11868 3180
rect -11485 3163 -11468 3180
rect -11885 3163 -11868 3180
rect -11605 3163 -11588 3180
rect -11565 3163 -11548 3180
rect -11445 3163 -11428 3180
rect -11765 3163 -11748 3180
rect -11525 3163 -11508 3180
rect -11885 3163 -11868 3180
rect -11485 3163 -11468 3180
rect -11565 3163 -11548 3180
rect -11645 3163 -11628 3180
rect -11685 3163 -11668 3180
rect -11565 3163 -11548 3180
rect -11605 3163 -11588 3180
rect -11805 3163 -11788 3180
rect -11885 3163 -11868 3180
rect -11725 3163 -11708 3180
rect -11645 3163 -11628 3180
rect -11725 3163 -11708 3180
rect -11565 3163 -11548 3180
rect -11605 3163 -11588 3180
rect -11405 3163 -11388 3180
rect -11525 3163 -11508 3180
rect -11765 3163 -11748 3180
rect -11685 3163 -11668 3180
rect -11845 3163 -11828 3180
rect -11405 3163 -11388 3180
rect -12125 3163 -12108 3180
rect -12125 3163 -12108 3180
rect -12125 3163 -12108 3180
rect -12325 3163 -12308 3180
rect -12285 3163 -12268 3180
rect -12285 3163 -12268 3180
rect -12045 3163 -12028 3180
rect -12245 3163 -12228 3180
rect -12245 3163 -12228 3180
rect -12045 3163 -12028 3180
rect -12445 3163 -12428 3180
rect -12365 3163 -12348 3180
rect -12365 3163 -12348 3180
rect -12125 3163 -12108 3180
rect -12245 3163 -12228 3180
rect -12245 3163 -12228 3180
rect -12325 3163 -12308 3180
rect -12405 3163 -12388 3180
rect -12325 3163 -12308 3180
rect -12405 3163 -12388 3180
rect -12085 3163 -12068 3180
rect -12205 3163 -12188 3180
rect -12445 3163 -12428 3180
rect -12085 3163 -12068 3180
rect -12405 3163 -12388 3180
rect -12405 3163 -12388 3180
rect -12165 3163 -12148 3180
rect -12045 3163 -12028 3180
rect -12445 3163 -12428 3180
rect -12085 3163 -12068 3180
rect -12365 3163 -12348 3180
rect -11965 3163 -11948 3180
rect -12005 3163 -11988 3180
rect -12005 3163 -11988 3180
rect -12285 3163 -12268 3180
rect -11965 3163 -11948 3180
rect -12005 3163 -11988 3180
rect -12285 3163 -12268 3180
rect -12165 3163 -12148 3180
rect -12165 3163 -12148 3180
rect -12205 3163 -12188 3180
rect -12445 3163 -12428 3180
rect -12365 3163 -12348 3180
rect -11965 3163 -11948 3180
rect -12005 3163 -11988 3180
rect -12045 3163 -12028 3180
rect -12165 3163 -12148 3180
rect -12085 3163 -12068 3180
rect -11965 3163 -11948 3180
rect -12205 3163 -12188 3180
rect -12205 3163 -12188 3180
rect -12325 3163 -12308 3180
rect -13006 3163 -12989 3180
rect -13006 3163 -12989 3180
rect -13006 3163 -12989 3180
rect -13006 3163 -12989 3180
rect -12766 3163 -12749 3180
rect -12806 3163 -12789 3180
rect -12486 3163 -12469 3180
rect -12726 3163 -12709 3180
rect -12966 3163 -12949 3180
rect -12686 3163 -12669 3180
rect -12606 3163 -12589 3180
rect -12926 3163 -12909 3180
rect -12486 3163 -12469 3180
rect -12646 3163 -12629 3180
rect -12526 3163 -12509 3180
rect -12566 3163 -12549 3180
rect -12686 3163 -12669 3180
rect -12606 3163 -12589 3180
rect -12526 3163 -12509 3180
rect -12966 3163 -12949 3180
rect -12766 3163 -12749 3180
rect -12926 3163 -12909 3180
rect -12726 3163 -12709 3180
rect -12646 3163 -12629 3180
rect -12766 3163 -12749 3180
rect -12966 3163 -12949 3180
rect -12966 3163 -12949 3180
rect -12686 3163 -12669 3180
rect -12726 3163 -12709 3180
rect -12886 3163 -12869 3180
rect -12766 3163 -12749 3180
rect -12806 3163 -12789 3180
rect -12846 3163 -12829 3180
rect -12846 3163 -12829 3180
rect -12846 3163 -12829 3180
rect -12566 3163 -12549 3180
rect -12886 3163 -12869 3180
rect -12886 3163 -12869 3180
rect -12846 3163 -12829 3180
rect -12486 3163 -12469 3180
rect -12806 3163 -12789 3180
rect -12726 3163 -12709 3180
rect -12526 3163 -12509 3180
rect -12886 3163 -12869 3180
rect -12566 3163 -12549 3180
rect -12806 3163 -12789 3180
rect -12606 3163 -12589 3180
rect -12926 3163 -12909 3180
rect -12486 3163 -12469 3180
rect -12646 3163 -12629 3180
rect -12926 3163 -12909 3180
rect -12526 3163 -12509 3180
rect -12566 3163 -12549 3180
rect -12686 3163 -12669 3180
rect -12606 3163 -12589 3180
rect -12646 3163 -12629 3180
rect -13286 3163 -13269 3180
rect -13086 3163 -13069 3180
rect -13486 3163 -13469 3180
rect -13046 3163 -13029 3180
rect -13206 3163 -13189 3180
rect -13046 3163 -13029 3180
rect -13166 3163 -13149 3180
rect -13046 3163 -13029 3180
rect -13166 3163 -13149 3180
rect -13526 3163 -13509 3180
rect -13126 3163 -13109 3180
rect -13126 3163 -13109 3180
rect -13246 3163 -13229 3180
rect -13326 3163 -13309 3180
rect -13166 3163 -13149 3180
rect -13406 3163 -13389 3180
rect -13086 3163 -13069 3180
rect -13326 3163 -13309 3180
rect -13086 3163 -13069 3180
rect -13446 3163 -13429 3180
rect -13486 3163 -13469 3180
rect -13326 3163 -13309 3180
rect -13486 3163 -13469 3180
rect -13206 3163 -13189 3180
rect -13126 3163 -13109 3180
rect -13206 3163 -13189 3180
rect -13526 3163 -13509 3180
rect -13406 3163 -13389 3180
rect -13286 3163 -13269 3180
rect -13446 3163 -13429 3180
rect -13246 3163 -13229 3180
rect -13326 3163 -13309 3180
rect -13526 3163 -13509 3180
rect -13486 3163 -13469 3180
rect -13446 3163 -13429 3180
rect -13086 3163 -13069 3180
rect -13526 3163 -13509 3180
rect -13246 3163 -13229 3180
rect -13246 3163 -13229 3180
rect -13406 3163 -13389 3180
rect -13206 3163 -13189 3180
rect -13286 3163 -13269 3180
rect -13166 3163 -13149 3180
rect -13286 3163 -13269 3180
rect -13366 3163 -13349 3180
rect -13126 3163 -13109 3180
rect -13366 3163 -13349 3180
rect -13366 3163 -13349 3180
rect -13406 3163 -13389 3180
rect -13446 3163 -13429 3180
rect -13046 3163 -13029 3180
rect -13366 3163 -13349 3180
rect -14086 3163 -14069 3180
rect -14086 3163 -14069 3180
rect -14086 3163 -14069 3180
rect -14086 3163 -14069 3180
rect -13726 3163 -13709 3180
rect -13566 3163 -13549 3180
rect -13766 3163 -13749 3180
rect -13966 3163 -13949 3180
rect -13926 3163 -13909 3180
rect -13646 3163 -13629 3180
rect -13566 3163 -13549 3180
rect -13686 3163 -13669 3180
rect -13966 3163 -13949 3180
rect -13646 3163 -13629 3180
rect -13646 3163 -13629 3180
rect -13646 3163 -13629 3180
rect -13566 3163 -13549 3180
rect -13846 3163 -13829 3180
rect -13966 3163 -13949 3180
rect -13686 3163 -13669 3180
rect -14046 3163 -14029 3180
rect -14006 3163 -13989 3180
rect -13806 3163 -13789 3180
rect -13766 3163 -13749 3180
rect -13846 3163 -13829 3180
rect -13846 3163 -13829 3180
rect -13926 3163 -13909 3180
rect -13926 3163 -13909 3180
rect -13886 3163 -13869 3180
rect -14006 3163 -13989 3180
rect -13606 3163 -13589 3180
rect -13886 3163 -13869 3180
rect -13806 3163 -13789 3180
rect -13886 3163 -13869 3180
rect -13566 3163 -13549 3180
rect -13966 3163 -13949 3180
rect -13686 3163 -13669 3180
rect -13686 3163 -13669 3180
rect -13726 3163 -13709 3180
rect -14046 3163 -14029 3180
rect -13766 3163 -13749 3180
rect -13726 3163 -13709 3180
rect -13606 3163 -13589 3180
rect -13726 3163 -13709 3180
rect -14006 3163 -13989 3180
rect -13926 3163 -13909 3180
rect -13886 3163 -13869 3180
rect -13806 3163 -13789 3180
rect -13806 3163 -13789 3180
rect -13846 3163 -13829 3180
rect -14046 3163 -14029 3180
rect -14046 3163 -14029 3180
rect -14006 3163 -13989 3180
rect -13766 3163 -13749 3180
rect -13606 3163 -13589 3180
rect -13606 3163 -13589 3180
rect -9765 3163 -9748 3180
rect -9765 3163 -9748 3180
rect -9765 3163 -9748 3180
rect -14126 3163 -14109 3180
rect -9765 3163 -9748 3180
rect -14126 3163 -14109 3180
rect -9685 3163 -9668 3180
rect -9605 3163 -9588 3180
rect -9725 3163 -9708 3180
rect -9565 3163 -9548 3180
rect -9485 3163 -9468 3180
rect -9605 3163 -9588 3180
rect -14166 3163 -14149 3180
rect -9645 3163 -9628 3180
rect -9485 3163 -9468 3180
rect -9525 3163 -9508 3180
rect -9565 3163 -9548 3180
rect -9445 3163 -9428 3180
rect -9565 3163 -9548 3180
rect -9525 3163 -9508 3180
rect -9485 3163 -9468 3180
rect -9565 3163 -9548 3180
rect -9445 3163 -9428 3180
rect -9485 3163 -9468 3180
rect -9645 3163 -9628 3180
rect -9605 3163 -9588 3180
rect -9445 3163 -9428 3180
rect -9725 3163 -9708 3180
rect -9725 3163 -9708 3180
rect -9445 3163 -9428 3180
rect -9685 3163 -9668 3180
rect -14166 3163 -14149 3180
rect -9725 3163 -9708 3180
rect -9645 3163 -9628 3180
rect -9645 3163 -9628 3180
rect -14166 3163 -14149 3180
rect -9525 3163 -9508 3180
rect -9525 3163 -9508 3180
rect -9605 3163 -9588 3180
rect -9685 3163 -9668 3180
rect -9685 3163 -9668 3180
rect -10285 3163 -10268 3180
rect -9845 3163 -9828 3180
rect -14126 3163 -14109 3180
rect -10285 3163 -10268 3180
rect -14166 3163 -14149 3180
rect -10005 3163 -9988 3180
rect -10005 3163 -9988 3180
rect -10005 3163 -9988 3180
rect -14126 3163 -14109 3180
rect -10005 3163 -9988 3180
rect -10045 3163 -10028 3180
rect -9965 3163 -9948 3180
rect -10125 3163 -10108 3180
rect -9965 3163 -9948 3180
rect -9805 3163 -9788 3180
rect -10285 3163 -10268 3180
rect -10125 3163 -10108 3180
rect -9885 3163 -9868 3180
rect -10045 3163 -10028 3180
rect -10205 3163 -10188 3180
rect -9925 3163 -9908 3180
rect -9925 3163 -9908 3180
rect -10245 3163 -10228 3180
rect -10085 3163 -10068 3180
rect -9925 3163 -9908 3180
rect -10245 3163 -10228 3180
rect -10165 3163 -10148 3180
rect -9965 3163 -9948 3180
rect -9885 3163 -9868 3180
rect -9805 3163 -9788 3180
rect -10125 3163 -10108 3180
rect -10085 3163 -10068 3180
rect -10045 3163 -10028 3180
rect -10085 3163 -10068 3180
rect -10245 3163 -10228 3180
rect -10285 3163 -10268 3180
rect -10165 3163 -10148 3180
rect -10205 3163 -10188 3180
rect -9805 3163 -9788 3180
rect -9925 3163 -9908 3180
rect -10205 3163 -10188 3180
rect -10205 3163 -10188 3180
rect -9885 3163 -9868 3180
rect -9845 3163 -9828 3180
rect -10245 3163 -10228 3180
rect -10125 3163 -10108 3180
rect -10045 3163 -10028 3180
rect -9885 3163 -9868 3180
rect -10085 3163 -10068 3180
rect -9805 3163 -9788 3180
rect -9845 3163 -9828 3180
rect -10165 3163 -10148 3180
rect -9965 3163 -9948 3180
rect -10165 3163 -10148 3180
rect -9845 3163 -9828 3180
rect -10845 3163 -10828 3180
rect -10845 3163 -10828 3180
rect -10845 3163 -10828 3180
rect -10845 3163 -10828 3180
rect -10805 3163 -10788 3180
rect -10765 3163 -10748 3180
rect -10765 3163 -10748 3180
rect -10645 3163 -10628 3180
rect -10805 3163 -10788 3180
rect -10685 3163 -10668 3180
rect -10725 3163 -10708 3180
rect -10645 3163 -10628 3180
rect -10725 3163 -10708 3180
rect -10685 3163 -10668 3180
rect -10805 3163 -10788 3180
rect -10645 3163 -10628 3180
rect -10685 3163 -10668 3180
rect -10725 3163 -10708 3180
rect -10765 3163 -10748 3180
rect -10805 3163 -10788 3180
rect -13053 2394 -13036 2411
rect -13013 2394 -12996 2411
rect -13733 2394 -13716 2411
rect -13573 2394 -13556 2411
rect -14093 2394 -14076 2411
rect -13173 2394 -13156 2411
rect -13973 2394 -13956 2411
rect -13213 2394 -13196 2411
rect -14013 2394 -13996 2411
rect -13253 2394 -13236 2411
rect -13293 2394 -13276 2411
rect -13413 2394 -13396 2411
rect -13773 2394 -13756 2411
rect -14133 2394 -14116 2411
rect -14053 2394 -14036 2411
rect -13613 2394 -13596 2411
rect -13333 2394 -13316 2411
rect -13453 2394 -13436 2411
rect -13813 2394 -13796 2411
rect -13373 2394 -13356 2411
rect -13893 2394 -13876 2411
rect -14093 2394 -14076 2411
rect -13493 2394 -13476 2411
rect -14133 2394 -14116 2411
rect -13533 2394 -13516 2411
rect -13653 2394 -13636 2411
rect -14013 2394 -13996 2411
rect -13853 2394 -13836 2411
rect -13573 2394 -13556 2411
rect -13933 2394 -13916 2411
rect -13173 2394 -13156 2411
rect -13933 2394 -13916 2411
rect -13213 2394 -13196 2411
rect -13613 2394 -13596 2411
rect -13253 2394 -13236 2411
rect -13653 2394 -13636 2411
rect -13293 2394 -13276 2411
rect -13693 2394 -13676 2411
rect -13333 2394 -13316 2411
rect -13693 2394 -13676 2411
rect -14053 2394 -14036 2411
rect -13893 2394 -13876 2411
rect -13373 2394 -13356 2411
rect -13733 2394 -13716 2411
rect -13853 2394 -13836 2411
rect -13413 2394 -13396 2411
rect -13773 2394 -13756 2411
rect -13973 2394 -13956 2411
rect -13453 2394 -13436 2411
rect -13813 2394 -13796 2411
rect -13493 2394 -13476 2411
rect -13533 2394 -13516 2411
rect -13053 2394 -13036 2411
rect -13093 2394 -13076 2411
rect -13013 2394 -12996 2411
rect -13133 2394 -13116 2411
rect -13093 2394 -13076 2411
rect -13133 2394 -13116 2411
rect -12453 2394 -12436 2411
rect -12493 2394 -12476 2411
rect -12253 2394 -12236 2411
rect -12893 2394 -12876 2411
rect -12213 2394 -12196 2411
rect -12253 2394 -12236 2411
rect -12773 2394 -12756 2411
rect -12293 2394 -12276 2411
rect -12613 2394 -12596 2411
rect -12933 2394 -12916 2411
rect -12373 2394 -12356 2411
rect -11813 2394 -11796 2411
rect -11813 2394 -11796 2411
rect -11853 2394 -11836 2411
rect -11973 2394 -11956 2411
rect -12013 2394 -11996 2411
rect -12053 2394 -12036 2411
rect -11853 2394 -11836 2411
rect -11933 2394 -11916 2411
rect -11973 2394 -11956 2411
rect -12013 2394 -11996 2411
rect -12053 2394 -12036 2411
rect -11933 2394 -11916 2411
rect -11893 2394 -11876 2411
rect -11893 2394 -11876 2411
rect -12693 2394 -12676 2411
rect -12333 2394 -12316 2411
rect -12613 2394 -12596 2411
rect -12693 2394 -12676 2411
rect -12653 2394 -12636 2411
rect -12573 2394 -12556 2411
rect -12093 2394 -12076 2411
rect -12653 2394 -12636 2411
rect -12493 2394 -12476 2411
rect -12773 2394 -12756 2411
rect -12413 2394 -12396 2411
rect -12533 2394 -12516 2411
rect -12813 2394 -12796 2411
rect -12933 2394 -12916 2411
rect -12533 2394 -12516 2411
rect -12333 2394 -12316 2411
rect -12973 2394 -12956 2411
rect -12853 2394 -12836 2411
rect -12813 2394 -12796 2411
rect -12853 2394 -12836 2411
rect -12973 2394 -12956 2411
rect -12133 2394 -12116 2411
rect -12173 2394 -12156 2411
rect -12573 2394 -12556 2411
rect -12413 2394 -12396 2411
rect -12093 2394 -12076 2411
rect -12453 2394 -12436 2411
rect -12893 2394 -12876 2411
rect -12293 2394 -12276 2411
rect -12173 2394 -12156 2411
rect -12373 2394 -12356 2411
rect -12133 2394 -12116 2411
rect -12213 2394 -12196 2411
rect -12733 2394 -12716 2411
rect -12733 2394 -12716 2411
rect -10612 2394 -10595 2411
rect -10612 2394 -10595 2411
rect -10652 2394 -10635 2411
rect -10652 2394 -10635 2411
rect -10692 2394 -10675 2411
rect -10732 2394 -10715 2411
rect -10772 2394 -10755 2411
rect -10812 2394 -10795 2411
rect -10852 2394 -10835 2411
rect -11613 2394 -11596 2411
rect -11653 2394 -11636 2411
rect -11693 2394 -11676 2411
rect -11253 2394 -11236 2411
rect -11733 2394 -11716 2411
rect -11773 2394 -11756 2411
rect -11053 2394 -11036 2411
rect -11573 2394 -11556 2411
rect -11413 2394 -11396 2411
rect -11093 2394 -11076 2411
rect -11613 2394 -11596 2411
rect -11533 2394 -11516 2411
rect -11333 2394 -11316 2411
rect -11013 2394 -10996 2411
rect -11293 2394 -11276 2411
rect -11133 2394 -11116 2411
rect -11453 2394 -11436 2411
rect -11013 2394 -10996 2411
rect -11573 2394 -11556 2411
rect -11653 2394 -11636 2411
rect -11173 2394 -11156 2411
rect -11053 2394 -11036 2411
rect -11093 2394 -11076 2411
rect -11213 2394 -11196 2411
rect -11133 2394 -11116 2411
rect -11693 2394 -11676 2411
rect -11173 2394 -11156 2411
rect -11493 2394 -11476 2411
rect -11213 2394 -11196 2411
rect -11253 2394 -11236 2411
rect -11493 2394 -11476 2411
rect -11733 2394 -11716 2411
rect -11453 2394 -11436 2411
rect -11293 2394 -11276 2411
rect -11333 2394 -11316 2411
rect -11373 2394 -11356 2411
rect -11373 2394 -11356 2411
rect -11773 2394 -11756 2411
rect -11413 2394 -11396 2411
rect -11533 2394 -11516 2411
rect -10892 2394 -10875 2411
rect -10932 2394 -10915 2411
rect -10972 2394 -10955 2411
rect -10732 2394 -10715 2411
rect -10772 2394 -10755 2411
rect -10812 2394 -10795 2411
rect -10852 2394 -10835 2411
rect -10892 2394 -10875 2411
rect -10932 2394 -10915 2411
rect -10972 2394 -10955 2411
rect -10692 2394 -10675 2411
rect -9972 2394 -9955 2411
rect -10252 2394 -10235 2411
rect -10412 2394 -10395 2411
rect -9532 2394 -9515 2411
rect -10012 2394 -9995 2411
rect -10092 2394 -10075 2411
rect -10292 2394 -10275 2411
rect -10052 2394 -10035 2411
rect -10572 2394 -10555 2411
rect -10012 2394 -9995 2411
rect -10532 2394 -10515 2411
rect -9492 2394 -9475 2411
rect -10332 2394 -10315 2411
rect -10572 2394 -10555 2411
rect -9572 2394 -9555 2411
rect -10092 2394 -10075 2411
rect -10532 2394 -10515 2411
rect -10132 2394 -10115 2411
rect -10492 2394 -10475 2411
rect -9612 2394 -9595 2411
rect -9652 2394 -9635 2411
rect -9692 2394 -9675 2411
rect -9732 2394 -9715 2411
rect -9452 2394 -9435 2411
rect -9732 2394 -9715 2411
rect -9492 2394 -9475 2411
rect -9772 2394 -9755 2411
rect -9812 2394 -9795 2411
rect -9852 2394 -9835 2411
rect -9892 2394 -9875 2411
rect -9532 2394 -9515 2411
rect -9572 2394 -9555 2411
rect -9612 2394 -9595 2411
rect -9772 2394 -9755 2411
rect -10172 2394 -10155 2411
rect -9812 2394 -9795 2411
rect -10172 2394 -10155 2411
rect -9852 2394 -9835 2411
rect -10212 2394 -10195 2411
rect -10372 2394 -10355 2411
rect -10252 2394 -10235 2411
rect -9892 2394 -9875 2411
rect -9932 2394 -9915 2411
rect -9652 2394 -9635 2411
rect -10292 2394 -10275 2411
rect -9452 2394 -9435 2411
rect -10332 2394 -10315 2411
rect -10212 2394 -10195 2411
rect -9692 2394 -9675 2411
rect -10452 2394 -10435 2411
rect -10052 2394 -10035 2411
rect -9972 2394 -9955 2411
rect -10492 2394 -10475 2411
rect -10372 2394 -10355 2411
rect -10452 2394 -10435 2411
rect -10132 2394 -10115 2411
rect -10412 2394 -10395 2411
rect -9932 2394 -9915 2411
rect -4652 2394 -4635 2411
rect -4652 2394 -4635 2411
rect -2365 4652 -2348 4669
rect -2405 4652 -2388 4669
rect -2445 4652 -2428 4669
rect -2485 4652 -2468 4669
rect -2725 4652 -2708 4669
rect -2805 4652 -2788 4669
rect -2525 4652 -2508 4669
rect -2565 4652 -2548 4669
rect -2605 4652 -2588 4669
rect -2845 4652 -2828 4669
rect -2365 4652 -2348 4669
rect -2405 4652 -2388 4669
rect -2445 4652 -2428 4669
rect -2485 4652 -2468 4669
rect -2525 4652 -2508 4669
rect -2565 4652 -2548 4669
rect -2605 4652 -2588 4669
rect -2325 4652 -2308 4669
rect -2285 4652 -2268 4669
rect -2285 4652 -2268 4669
rect -2325 4652 -2308 4669
rect -2285 4652 -2268 4669
rect -2365 4652 -2348 4669
rect -2325 4652 -2308 4669
rect -2405 4652 -2388 4669
rect -2685 4652 -2668 4669
rect -2445 4652 -2428 4669
rect -2725 4652 -2708 4669
rect -2485 4652 -2468 4669
rect -2365 4652 -2348 4669
rect -2525 4652 -2508 4669
rect -2645 4652 -2628 4669
rect -2565 4652 -2548 4669
rect -2405 4652 -2388 4669
rect -2605 4652 -2588 4669
rect -2845 4652 -2828 4669
rect -2645 4652 -2628 4669
rect -2445 4652 -2428 4669
rect -2685 4652 -2668 4669
rect -2725 4652 -2708 4669
rect -2765 4652 -2748 4669
rect -2805 4652 -2788 4669
rect -2845 4652 -2828 4669
rect -2605 4652 -2588 4669
rect -2485 4652 -2468 4669
rect -2565 4652 -2548 4669
rect -2765 4652 -2748 4669
rect -2645 4652 -2628 4669
rect -2685 4652 -2668 4669
rect -2725 4652 -2708 4669
rect -2765 4652 -2748 4669
rect -2805 4652 -2788 4669
rect -2845 4652 -2828 4669
rect -2765 4652 -2748 4669
rect -2645 4652 -2628 4669
rect -2285 4652 -2268 4669
rect -2325 4652 -2308 4669
rect -2525 4652 -2508 4669
rect -2685 4652 -2668 4669
rect -2805 4652 -2788 4669
rect -2925 4652 -2908 4669
rect -3405 4652 -3388 4669
rect -3005 4652 -2988 4669
rect -2885 4652 -2868 4669
rect -2925 4652 -2908 4669
rect -3365 4652 -3348 4669
rect -2965 4652 -2948 4669
rect -3005 4652 -2988 4669
rect -3045 4652 -3028 4669
rect -3085 4652 -3068 4669
rect -3125 4652 -3108 4669
rect -3165 4652 -3148 4669
rect -3205 4652 -3188 4669
rect -3245 4652 -3228 4669
rect -3285 4652 -3268 4669
rect -3325 4652 -3308 4669
rect -3365 4652 -3348 4669
rect -3405 4652 -3388 4669
rect -3445 4652 -3428 4669
rect -2965 4652 -2948 4669
rect -3045 4652 -3028 4669
rect -3085 4652 -3068 4669
rect -3125 4652 -3108 4669
rect -3445 4652 -3428 4669
rect -3165 4652 -3148 4669
rect -3205 4652 -3188 4669
rect -3245 4652 -3228 4669
rect -3285 4652 -3268 4669
rect -2965 4652 -2948 4669
rect -3005 4652 -2988 4669
rect -3045 4652 -3028 4669
rect -3085 4652 -3068 4669
rect -3125 4652 -3108 4669
rect -3165 4652 -3148 4669
rect -3205 4652 -3188 4669
rect -3245 4652 -3228 4669
rect -3285 4652 -3268 4669
rect -3325 4652 -3308 4669
rect -3365 4652 -3348 4669
rect -3405 4652 -3388 4669
rect -3445 4652 -3428 4669
rect -3045 4652 -3028 4669
rect -3085 4652 -3068 4669
rect -3125 4652 -3108 4669
rect -3165 4652 -3148 4669
rect -3205 4652 -3188 4669
rect -3245 4652 -3228 4669
rect -3285 4652 -3268 4669
rect -3325 4652 -3308 4669
rect -3365 4652 -3348 4669
rect -3405 4652 -3388 4669
rect -3445 4652 -3428 4669
rect -2885 4652 -2868 4669
rect -2925 4652 -2908 4669
rect -2965 4652 -2948 4669
rect -3005 4652 -2988 4669
rect -2885 4652 -2868 4669
rect -2925 4652 -2908 4669
rect -3325 4652 -3308 4669
rect -2885 4652 -2868 4669
rect -3925 4652 -3908 4669
rect -3485 4652 -3468 4669
rect -3925 4652 -3908 4669
rect -3925 4652 -3908 4669
rect -4045 4652 -4028 4669
rect -3565 4652 -3548 4669
rect -3485 4652 -3468 4669
rect -3485 4652 -3468 4669
rect -3525 4652 -3508 4669
rect -3845 4652 -3828 4669
rect -3525 4652 -3508 4669
rect -3565 4652 -3548 4669
rect -4045 4652 -4028 4669
rect -3605 4652 -3588 4669
rect -3645 4652 -3628 4669
rect -3885 4652 -3868 4669
rect -3605 4652 -3588 4669
rect -3685 4652 -3668 4669
rect -3725 4652 -3708 4669
rect -3765 4652 -3748 4669
rect -3885 4652 -3868 4669
rect -3805 4652 -3788 4669
rect -3965 4652 -3948 4669
rect -3925 4652 -3908 4669
rect -3845 4652 -3828 4669
rect -3965 4652 -3948 4669
rect -4005 4652 -3988 4669
rect -4005 4652 -3988 4669
rect -3725 4652 -3708 4669
rect -4045 4652 -4028 4669
rect -4005 4652 -3988 4669
rect -3565 4652 -3548 4669
rect -3645 4652 -3628 4669
rect -4045 4652 -4028 4669
rect -3605 4652 -3588 4669
rect -3685 4652 -3668 4669
rect -3565 4652 -3548 4669
rect -3645 4652 -3628 4669
rect -3765 4652 -3748 4669
rect -3965 4652 -3948 4669
rect -3725 4652 -3708 4669
rect -3805 4652 -3788 4669
rect -3845 4652 -3828 4669
rect -4005 4652 -3988 4669
rect -3525 4652 -3508 4669
rect -3765 4652 -3748 4669
rect -3485 4652 -3468 4669
rect -3805 4652 -3788 4669
rect -3845 4652 -3828 4669
rect -3525 4652 -3508 4669
rect -3685 4652 -3668 4669
rect -3605 4652 -3588 4669
rect -3885 4652 -3868 4669
rect -3725 4652 -3708 4669
rect -3645 4652 -3628 4669
rect -3805 4652 -3788 4669
rect -3765 4652 -3748 4669
rect -3965 4652 -3948 4669
rect -3685 4652 -3668 4669
rect -3885 4652 -3868 4669
rect -4085 4652 -4068 4669
rect -4605 4652 -4588 4669
rect -4525 4652 -4508 4669
rect -4645 4652 -4628 4669
rect -4285 4652 -4268 4669
rect -4565 4652 -4548 4669
rect -4165 4652 -4148 4669
rect -4605 4652 -4588 4669
rect -4325 4652 -4308 4669
rect -4645 4652 -4628 4669
rect -4365 4652 -4348 4669
rect -4205 4652 -4188 4669
rect -4405 4652 -4388 4669
rect -4125 4652 -4108 4669
rect -4445 4652 -4428 4669
rect -4245 4652 -4228 4669
rect -4085 4652 -4068 4669
rect -4125 4652 -4108 4669
rect -4165 4652 -4148 4669
rect -4205 4652 -4188 4669
rect -4245 4652 -4228 4669
rect -4285 4652 -4268 4669
rect -4325 4652 -4308 4669
rect -4365 4652 -4348 4669
rect -4405 4652 -4388 4669
rect -4445 4652 -4428 4669
rect -4525 4652 -4508 4669
rect -4485 4652 -4468 4669
rect -4485 4652 -4468 4669
rect -4605 4652 -4588 4669
rect -4645 4652 -4628 4669
rect -4525 4652 -4508 4669
rect -4325 4652 -4308 4669
rect -4205 4652 -4188 4669
rect -4645 4652 -4628 4669
rect -4125 4652 -4108 4669
rect -4285 4652 -4268 4669
rect -4365 4652 -4348 4669
rect -4445 4652 -4428 4669
rect -4085 4652 -4068 4669
rect -4165 4652 -4148 4669
rect -4405 4652 -4388 4669
rect -4565 4652 -4548 4669
rect -4365 4652 -4348 4669
rect -4245 4652 -4228 4669
rect -4565 4652 -4548 4669
rect -4245 4652 -4228 4669
rect -4445 4652 -4428 4669
rect -4165 4652 -4148 4669
rect -4605 4652 -4588 4669
rect -4325 4652 -4308 4669
rect -4525 4652 -4508 4669
rect -4085 4652 -4068 4669
rect -4205 4652 -4188 4669
rect -4125 4652 -4108 4669
rect -4485 4652 -4468 4669
rect -4285 4652 -4268 4669
rect -4485 4652 -4468 4669
rect -4405 4652 -4388 4669
rect -4565 4652 -4548 4669
rect -885 4652 -868 4669
rect -845 4652 -828 4669
rect -805 4652 -788 4669
rect -765 4652 -748 4669
rect -725 4652 -708 4669
rect -685 4652 -668 4669
rect -645 4652 -628 4669
rect -605 4652 -588 4669
rect -565 4652 -548 4669
rect -525 4652 -508 4669
rect -485 4652 -468 4669
rect -885 4652 -868 4669
rect -965 4652 -948 4669
rect -845 4652 -828 4669
rect -805 4652 -788 4669
rect -765 4652 -748 4669
rect -725 4652 -708 4669
rect -685 4652 -668 4669
rect -645 4652 -628 4669
rect -605 4652 -588 4669
rect -565 4652 -548 4669
rect -525 4652 -508 4669
rect -485 4652 -468 4669
rect -445 4652 -428 4669
rect -405 4652 -388 4669
rect -365 4652 -348 4669
rect -325 4652 -308 4669
rect -285 4652 -268 4669
rect -245 4652 -228 4669
rect -205 4652 -188 4669
rect -165 4652 -148 4669
rect -125 4652 -108 4669
rect -85 4652 -68 4669
rect -45 4652 -28 4669
rect -5 4652 13 4669
rect 36 4652 53 4669
rect 76 4652 93 4669
rect -965 4652 -948 4669
rect -925 4652 -908 4669
rect -445 4652 -428 4669
rect -405 4652 -388 4669
rect -365 4652 -348 4669
rect -325 4652 -308 4669
rect -285 4652 -268 4669
rect -245 4652 -228 4669
rect -205 4652 -188 4669
rect -165 4652 -148 4669
rect -125 4652 -108 4669
rect -85 4652 -68 4669
rect -45 4652 -28 4669
rect -5 4652 13 4669
rect 36 4652 53 4669
rect 76 4652 93 4669
rect -925 4652 -908 4669
rect -2005 4652 -1988 4669
rect -2045 4652 -2028 4669
rect -2085 4652 -2068 4669
rect -2125 4652 -2108 4669
rect -2165 4652 -2148 4669
rect -2205 4652 -2188 4669
rect -2245 4652 -2228 4669
rect -1685 4652 -1668 4669
rect -1725 4652 -1708 4669
rect -1765 4652 -1748 4669
rect -1805 4652 -1788 4669
rect -1845 4652 -1828 4669
rect -1885 4652 -1868 4669
rect -1925 4652 -1908 4669
rect -1965 4652 -1948 4669
rect -2005 4652 -1988 4669
rect -2045 4652 -2028 4669
rect -2085 4652 -2068 4669
rect -2125 4652 -2108 4669
rect -2165 4652 -2148 4669
rect -2205 4652 -2188 4669
rect -2205 4652 -2188 4669
rect -1765 4652 -1748 4669
rect -1805 4652 -1788 4669
rect -1845 4652 -1828 4669
rect -1885 4652 -1868 4669
rect -1925 4652 -1908 4669
rect -1965 4652 -1948 4669
rect -2005 4652 -1988 4669
rect -2045 4652 -2028 4669
rect -2085 4652 -2068 4669
rect -2125 4652 -2108 4669
rect -2205 4652 -2188 4669
rect -2165 4652 -2148 4669
rect -2245 4652 -2228 4669
rect -1685 4652 -1668 4669
rect -1725 4652 -1708 4669
rect -2245 4652 -2228 4669
rect -2245 4652 -2228 4669
rect -1685 4652 -1668 4669
rect -1725 4652 -1708 4669
rect -1765 4652 -1748 4669
rect -1805 4652 -1788 4669
rect -1845 4652 -1828 4669
rect -1885 4652 -1868 4669
rect -1925 4652 -1908 4669
rect -1685 4652 -1668 4669
rect -1725 4652 -1708 4669
rect -1765 4652 -1748 4669
rect -1805 4652 -1788 4669
rect -1845 4652 -1828 4669
rect -1885 4652 -1868 4669
rect -1925 4652 -1908 4669
rect -1965 4652 -1948 4669
rect -2005 4652 -1988 4669
rect -2045 4652 -2028 4669
rect -2085 4652 -2068 4669
rect -2125 4652 -2108 4669
rect -2165 4652 -2148 4669
rect -1965 4652 -1948 4669
rect -7206 4652 -7189 4669
rect -7606 4652 -7589 4669
rect -7406 4652 -7389 4669
rect -7126 4652 -7109 4669
rect -7446 4652 -7429 4669
rect -7446 4652 -7429 4669
rect -7486 4652 -7469 4669
rect -7166 4652 -7149 4669
rect -7446 4652 -7429 4669
rect -7486 4652 -7469 4669
rect -7046 4652 -7029 4669
rect -7326 4652 -7309 4669
rect -7406 4652 -7389 4669
rect -7526 4652 -7509 4669
rect -7526 4652 -7509 4669
rect -7486 4652 -7469 4669
rect -7246 4652 -7229 4669
rect -7566 4652 -7549 4669
rect -7406 4652 -7389 4669
rect -7526 4652 -7509 4669
rect -7526 4652 -7509 4669
rect -7606 4652 -7589 4669
rect -7246 4652 -7229 4669
rect -7566 4652 -7549 4669
rect -7606 4652 -7589 4669
rect -7126 4652 -7109 4669
rect -7286 4652 -7269 4669
rect -7606 4652 -7589 4669
rect -7566 4652 -7549 4669
rect -7246 4652 -7229 4669
rect -7166 4652 -7149 4669
rect -7366 4652 -7349 4669
rect -7446 4652 -7429 4669
rect -7046 4652 -7029 4669
rect -7406 4652 -7389 4669
rect -7566 4652 -7549 4669
rect -7326 4652 -7309 4669
rect -7286 4652 -7269 4669
rect -7366 4652 -7349 4669
rect -7206 4652 -7189 4669
rect -7086 4652 -7069 4669
rect -7326 4652 -7309 4669
rect -7086 4652 -7069 4669
rect -7126 4652 -7109 4669
rect -7286 4652 -7269 4669
rect -7486 4652 -7469 4669
rect -7366 4652 -7349 4669
rect -7366 4652 -7349 4669
rect -7046 4652 -7029 4669
rect -7206 4652 -7189 4669
rect -7166 4652 -7149 4669
rect -7246 4652 -7229 4669
rect -7086 4652 -7069 4669
rect -7046 4652 -7029 4669
rect -7286 4652 -7269 4669
rect -7086 4652 -7069 4669
rect -7126 4652 -7109 4669
rect -7166 4652 -7149 4669
rect -7206 4652 -7189 4669
rect -7326 4652 -7309 4669
rect -8206 4652 -8189 4669
rect -8126 4652 -8109 4669
rect -8126 4652 -8109 4669
rect -8046 4652 -8029 4669
rect -7646 4652 -7629 4669
rect -8086 4652 -8069 4669
rect -7686 4652 -7669 4669
rect -8086 4652 -8069 4669
rect -8166 4652 -8149 4669
rect -7726 4652 -7709 4669
rect -8006 4652 -7989 4669
rect -7766 4652 -7749 4669
rect -7806 4652 -7789 4669
rect -8206 4652 -8189 4669
rect -7646 4652 -7629 4669
rect -8006 4652 -7989 4669
rect -7966 4652 -7949 4669
rect -7686 4652 -7669 4669
rect -7726 4652 -7709 4669
rect -7766 4652 -7749 4669
rect -7846 4652 -7829 4669
rect -7806 4652 -7789 4669
rect -8046 4652 -8029 4669
rect -7846 4652 -7829 4669
rect -7886 4652 -7869 4669
rect -7886 4652 -7869 4669
rect -7926 4652 -7909 4669
rect -7926 4652 -7909 4669
rect -7966 4652 -7949 4669
rect -8046 4652 -8029 4669
rect -7926 4652 -7909 4669
rect -7766 4652 -7749 4669
rect -7966 4652 -7949 4669
rect -7806 4652 -7789 4669
rect -7646 4652 -7629 4669
rect -7686 4652 -7669 4669
rect -7646 4652 -7629 4669
rect -7966 4652 -7949 4669
rect -8086 4652 -8069 4669
rect -7766 4652 -7749 4669
rect -8206 4652 -8189 4669
rect -8046 4652 -8029 4669
rect -7686 4652 -7669 4669
rect -7886 4652 -7869 4669
rect -7926 4652 -7909 4669
rect -8166 4652 -8149 4669
rect -8086 4652 -8069 4669
rect -7846 4652 -7829 4669
rect -7726 4652 -7709 4669
rect -8166 4652 -8149 4669
rect -7846 4652 -7829 4669
rect -7726 4652 -7709 4669
rect -7886 4652 -7869 4669
rect -8206 4652 -8189 4669
rect -7806 4652 -7789 4669
rect -8126 4652 -8109 4669
rect -8006 4652 -7989 4669
rect -8006 4652 -7989 4669
rect -8126 4652 -8109 4669
rect -8166 4652 -8149 4669
rect -8406 4652 -8389 4669
rect -8366 4652 -8349 4669
rect -8286 4652 -8269 4669
rect -8406 4652 -8389 4669
rect -8486 4652 -8469 4669
rect -8526 4652 -8509 4669
rect -8446 4652 -8429 4669
rect -8606 4652 -8589 4669
rect -8486 4652 -8469 4669
rect -8526 4652 -8509 4669
rect -8246 4652 -8229 4669
rect -8526 4652 -8509 4669
rect -8446 4652 -8429 4669
rect -8566 4652 -8549 4669
rect -8686 4652 -8669 4669
rect -8766 4652 -8749 4669
rect -8606 4652 -8589 4669
rect -8766 4652 -8749 4669
rect -8646 4652 -8629 4669
rect -8726 4652 -8709 4669
rect -8806 4652 -8789 4669
rect -8686 4652 -8669 4669
rect -8446 4652 -8429 4669
rect -8726 4652 -8709 4669
rect -8286 4652 -8269 4669
rect -8606 4652 -8589 4669
rect -8766 4652 -8749 4669
rect -8646 4652 -8629 4669
rect -8806 4652 -8789 4669
rect -8406 4652 -8389 4669
rect -8726 4652 -8709 4669
rect -8806 4652 -8789 4669
rect -8326 4652 -8309 4669
rect -8406 4652 -8389 4669
rect -8526 4652 -8509 4669
rect -8366 4652 -8349 4669
rect -8326 4652 -8309 4669
rect -8246 4652 -8229 4669
rect -8446 4652 -8429 4669
rect -8246 4652 -8229 4669
rect -8566 4652 -8549 4669
rect -8566 4652 -8549 4669
rect -8486 4652 -8469 4669
rect -8646 4652 -8629 4669
rect -8286 4652 -8269 4669
rect -8606 4652 -8589 4669
rect -8566 4652 -8549 4669
rect -8686 4652 -8669 4669
rect -8806 4652 -8789 4669
rect -8326 4652 -8309 4669
rect -8766 4652 -8749 4669
rect -8486 4652 -8469 4669
rect -8726 4652 -8709 4669
rect -8246 4652 -8229 4669
rect -8366 4652 -8349 4669
rect -8366 4652 -8349 4669
rect -8286 4652 -8269 4669
rect -8686 4652 -8669 4669
rect -8326 4652 -8309 4669
rect -8646 4652 -8629 4669
rect -9166 4652 -9149 4669
rect -8846 4652 -8829 4669
rect -9366 4652 -9349 4669
rect -8846 4652 -8829 4669
rect -9246 4652 -9229 4669
rect -8886 4652 -8869 4669
rect -8886 4652 -8869 4669
rect -8926 4652 -8909 4669
rect -9086 4652 -9069 4669
rect -8966 4652 -8949 4669
rect -9326 4652 -9309 4669
rect -9006 4652 -8989 4669
rect -8846 4652 -8829 4669
rect -8886 4652 -8869 4669
rect -8966 4652 -8949 4669
rect -9406 4652 -9389 4669
rect -9326 4652 -9309 4669
rect -9166 4652 -9149 4669
rect -8926 4652 -8909 4669
rect -9046 4652 -9029 4669
rect -8966 4652 -8949 4669
rect -9086 4652 -9069 4669
rect -9006 4652 -8989 4669
rect -9206 4652 -9189 4669
rect -8966 4652 -8949 4669
rect -9126 4652 -9109 4669
rect -9406 4652 -9389 4669
rect -9366 4652 -9349 4669
rect -9046 4652 -9029 4669
rect -8886 4652 -8869 4669
rect -8846 4652 -8829 4669
rect -9006 4652 -8989 4669
rect -9286 4652 -9269 4669
rect -9246 4652 -9229 4669
rect -9246 4652 -9229 4669
rect -9126 4652 -9109 4669
rect -9366 4652 -9349 4669
rect -9166 4652 -9149 4669
rect -9366 4652 -9349 4669
rect -9406 4652 -9389 4669
rect -9206 4652 -9189 4669
rect -9286 4652 -9269 4669
rect -9286 4652 -9269 4669
rect -9406 4652 -9389 4669
rect -9086 4652 -9069 4669
rect -9126 4652 -9109 4669
rect -9326 4652 -9309 4669
rect -9166 4652 -9149 4669
rect -9206 4652 -9189 4669
rect -9086 4652 -9069 4669
rect -9326 4652 -9309 4669
rect -9046 4652 -9029 4669
rect -9046 4652 -9029 4669
rect -9006 4652 -8989 4669
rect -9126 4652 -9109 4669
rect -9206 4652 -9189 4669
rect -8926 4652 -8909 4669
rect -9246 4652 -9229 4669
rect -9286 4652 -9269 4669
rect -8926 4652 -8909 4669
rect -5845 4652 -5828 4669
rect -5845 4652 -5828 4669
rect -5845 4652 -5828 4669
rect -5845 4652 -5828 4669
rect -5245 4652 -5228 4669
rect -5245 4652 -5228 4669
rect -5245 4652 -5228 4669
rect -5245 4652 -5228 4669
rect -4845 4652 -4828 4669
rect -4765 4652 -4748 4669
rect -4885 4652 -4868 4669
rect -5125 4652 -5108 4669
rect -4805 4652 -4788 4669
rect -4885 4652 -4868 4669
rect -4805 4652 -4788 4669
rect -4765 4652 -4748 4669
rect -4845 4652 -4828 4669
rect -4845 4652 -4828 4669
rect -5085 4652 -5068 4669
rect -4685 4652 -4668 4669
rect -4885 4652 -4868 4669
rect -4685 4652 -4668 4669
rect -4925 4652 -4908 4669
rect -4965 4652 -4948 4669
rect -5005 4652 -4988 4669
rect -5045 4652 -5028 4669
rect -4885 4652 -4868 4669
rect -5085 4652 -5068 4669
rect -5125 4652 -5108 4669
rect -4725 4652 -4708 4669
rect -5165 4652 -5148 4669
rect -5205 4652 -5188 4669
rect -5085 4652 -5068 4669
rect -4925 4652 -4908 4669
rect -4725 4652 -4708 4669
rect -4965 4652 -4948 4669
rect -4725 4652 -4708 4669
rect -4965 4652 -4948 4669
rect -5045 4652 -5028 4669
rect -4925 4652 -4908 4669
rect -4805 4652 -4788 4669
rect -5125 4652 -5108 4669
rect -5165 4652 -5148 4669
rect -4765 4652 -4748 4669
rect -5005 4652 -4988 4669
rect -4765 4652 -4748 4669
rect -5005 4652 -4988 4669
rect -4685 4652 -4668 4669
rect -5205 4652 -5188 4669
rect -5165 4652 -5148 4669
rect -4925 4652 -4908 4669
rect -4965 4652 -4948 4669
rect -4805 4652 -4788 4669
rect -5005 4652 -4988 4669
rect -5045 4652 -5028 4669
rect -5085 4652 -5068 4669
rect -5125 4652 -5108 4669
rect -5045 4652 -5028 4669
rect -5165 4652 -5148 4669
rect -5205 4652 -5188 4669
rect -5205 4652 -5188 4669
rect -4845 4652 -4828 4669
rect -4685 4652 -4668 4669
rect -4725 4652 -4708 4669
rect -5765 4652 -5748 4669
rect -5805 4652 -5788 4669
rect -5725 4652 -5708 4669
rect -5645 4652 -5628 4669
rect -5285 4652 -5268 4669
rect -5725 4652 -5708 4669
rect -5685 4652 -5668 4669
rect -5285 4652 -5268 4669
rect -5325 4652 -5308 4669
rect -5365 4652 -5348 4669
rect -5405 4652 -5388 4669
rect -5445 4652 -5428 4669
rect -5485 4652 -5468 4669
rect -5525 4652 -5508 4669
rect -5565 4652 -5548 4669
rect -5605 4652 -5588 4669
rect -5645 4652 -5628 4669
rect -5685 4652 -5668 4669
rect -5285 4652 -5268 4669
rect -5765 4652 -5748 4669
rect -5325 4652 -5308 4669
rect -5365 4652 -5348 4669
rect -5805 4652 -5788 4669
rect -5405 4652 -5388 4669
rect -5445 4652 -5428 4669
rect -5485 4652 -5468 4669
rect -5405 4652 -5388 4669
rect -5525 4652 -5508 4669
rect -5285 4652 -5268 4669
rect -5565 4652 -5548 4669
rect -5325 4652 -5308 4669
rect -5365 4652 -5348 4669
rect -5605 4652 -5588 4669
rect -5325 4652 -5308 4669
rect -5405 4652 -5388 4669
rect -5645 4652 -5628 4669
rect -5365 4652 -5348 4669
rect -5445 4652 -5428 4669
rect -5645 4652 -5628 4669
rect -5685 4652 -5668 4669
rect -5725 4652 -5708 4669
rect -5765 4652 -5748 4669
rect -5805 4652 -5788 4669
rect -5805 4652 -5788 4669
rect -5485 4652 -5468 4669
rect -5445 4652 -5428 4669
rect -5485 4652 -5468 4669
rect -5525 4652 -5508 4669
rect -5525 4652 -5508 4669
rect -5565 4652 -5548 4669
rect -5565 4652 -5548 4669
rect -5605 4652 -5588 4669
rect -5685 4652 -5668 4669
rect -5605 4652 -5588 4669
rect -5765 4652 -5748 4669
rect -5725 4652 -5708 4669
rect -6446 4652 -6429 4669
rect -6446 4652 -6429 4669
rect -6446 4652 -6429 4669
rect -6446 4652 -6429 4669
rect -6086 4652 -6069 4669
rect -6086 4652 -6069 4669
rect -6246 4652 -6229 4669
rect -5885 4652 -5868 4669
rect -5885 4652 -5868 4669
rect -5925 4652 -5908 4669
rect -5965 4652 -5948 4669
rect -5925 4652 -5908 4669
rect -6006 4652 -5989 4669
rect -6086 4652 -6069 4669
rect -6126 4652 -6109 4669
rect -6166 4652 -6149 4669
rect -6286 4652 -6269 4669
rect -5885 4652 -5868 4669
rect -6206 4652 -6189 4669
rect -6326 4652 -6309 4669
rect -6006 4652 -5989 4669
rect -6046 4652 -6029 4669
rect -6086 4652 -6069 4669
rect -6006 4652 -5989 4669
rect -6126 4652 -6109 4669
rect -6166 4652 -6149 4669
rect -6206 4652 -6189 4669
rect -6246 4652 -6229 4669
rect -6286 4652 -6269 4669
rect -6326 4652 -6309 4669
rect -6366 4652 -6349 4669
rect -6406 4652 -6389 4669
rect -6166 4652 -6149 4669
rect -6206 4652 -6189 4669
rect -6246 4652 -6229 4669
rect -6206 4652 -6189 4669
rect -6326 4652 -6309 4669
rect -5925 4652 -5908 4669
rect -6006 4652 -5989 4669
rect -6126 4652 -6109 4669
rect -6126 4652 -6109 4669
rect -6366 4652 -6349 4669
rect -6406 4652 -6389 4669
rect -6286 4652 -6269 4669
rect -5965 4652 -5948 4669
rect -6166 4652 -6149 4669
rect -6246 4652 -6229 4669
rect -6326 4652 -6309 4669
rect -5965 4652 -5948 4669
rect -6286 4652 -6269 4669
rect -6046 4652 -6029 4669
rect -6046 4652 -6029 4669
rect -6366 4652 -6349 4669
rect -6366 4652 -6349 4669
rect -5885 4652 -5868 4669
rect -6046 4652 -6029 4669
rect -6406 4652 -6389 4669
rect -5965 4652 -5948 4669
rect -5925 4652 -5908 4669
rect -6406 4652 -6389 4669
rect -7006 4652 -6989 4669
rect -6526 4652 -6509 4669
rect -7006 4652 -6989 4669
rect -6886 4652 -6869 4669
rect -6886 4652 -6869 4669
rect -6486 4652 -6469 4669
rect -6806 4652 -6789 4669
rect -6526 4652 -6509 4669
rect -6766 4652 -6749 4669
rect -6566 4652 -6549 4669
rect -6566 4652 -6549 4669
rect -6486 4652 -6469 4669
rect -6966 4652 -6949 4669
rect -6606 4652 -6589 4669
rect -6926 4652 -6909 4669
rect -6646 4652 -6629 4669
rect -6606 4652 -6589 4669
rect -6926 4652 -6909 4669
rect -6486 4652 -6469 4669
rect -6926 4652 -6909 4669
rect -6966 4652 -6949 4669
rect -6766 4652 -6749 4669
rect -6806 4652 -6789 4669
rect -6846 4652 -6829 4669
rect -6886 4652 -6869 4669
rect -6926 4652 -6909 4669
rect -6966 4652 -6949 4669
rect -7006 4652 -6989 4669
rect -6646 4652 -6629 4669
rect -6486 4652 -6469 4669
rect -6526 4652 -6509 4669
rect -6566 4652 -6549 4669
rect -6606 4652 -6589 4669
rect -6646 4652 -6629 4669
rect -6686 4652 -6669 4669
rect -6526 4652 -6509 4669
rect -6566 4652 -6549 4669
rect -6686 4652 -6669 4669
rect -6726 4652 -6709 4669
rect -6606 4652 -6589 4669
rect -6766 4652 -6749 4669
rect -6686 4652 -6669 4669
rect -6806 4652 -6789 4669
rect -6846 4652 -6829 4669
rect -6966 4652 -6949 4669
rect -6846 4652 -6829 4669
rect -6726 4652 -6709 4669
rect -6686 4652 -6669 4669
rect -6886 4652 -6869 4669
rect -6726 4652 -6709 4669
rect -7006 4652 -6989 4669
rect -6726 4652 -6709 4669
rect -6766 4652 -6749 4669
rect -6806 4652 -6789 4669
rect -6846 4652 -6829 4669
rect -6646 4652 -6629 4669
rect -8485 3163 -8468 3180
rect -8445 3163 -8428 3180
rect -8645 3163 -8628 3180
rect -8565 3163 -8548 3180
rect -8565 3163 -8548 3180
rect -8405 3163 -8388 3180
rect -8445 3163 -8428 3180
rect -8645 3163 -8628 3180
rect -8365 3163 -8348 3180
rect -8245 3163 -8228 3180
rect -8245 3163 -8228 3180
rect -8605 3163 -8588 3180
rect -8165 3163 -8148 3180
rect -8445 3163 -8428 3180
rect -8285 3163 -8268 3180
rect -8485 3163 -8468 3180
rect -8245 3163 -8228 3180
rect -8165 3163 -8148 3180
rect -8645 3163 -8628 3180
rect -8565 3163 -8548 3180
rect -8365 3163 -8348 3180
rect -9165 3163 -9148 3180
rect -9085 3163 -9068 3180
rect -9205 3163 -9188 3180
rect -9125 3163 -9108 3180
rect -9005 3163 -8988 3180
rect -8725 3163 -8708 3180
rect -9005 3163 -8988 3180
rect -8925 3163 -8908 3180
rect -8805 3163 -8788 3180
rect -8885 3163 -8868 3180
rect -8845 3163 -8828 3180
rect -9125 3163 -9108 3180
rect -9165 3163 -9148 3180
rect -8885 3163 -8868 3180
rect -8765 3163 -8748 3180
rect -8725 3163 -8708 3180
rect -9005 3163 -8988 3180
rect -8805 3163 -8788 3180
rect -8725 3163 -8708 3180
rect -8885 3163 -8868 3180
rect -8965 3163 -8948 3180
rect -9045 3163 -9028 3180
rect -8765 3163 -8748 3180
rect -8845 3163 -8828 3180
rect -8805 3163 -8788 3180
rect -8925 3163 -8908 3180
rect -8845 3163 -8828 3180
rect -8845 3163 -8828 3180
rect -8925 3163 -8908 3180
rect -8925 3163 -8908 3180
rect -9045 3163 -9028 3180
rect -9045 3163 -9028 3180
rect -8805 3163 -8788 3180
rect -8965 3163 -8948 3180
rect -8765 3163 -8748 3180
rect -9085 3163 -9068 3180
rect -9125 3163 -9108 3180
rect -9005 3163 -8988 3180
rect -9165 3163 -9148 3180
rect -9205 3163 -9188 3180
rect -9205 3163 -9188 3180
rect -9165 3163 -9148 3180
rect -9085 3163 -9068 3180
rect -8965 3163 -8948 3180
rect -9085 3163 -9068 3180
rect -8765 3163 -8748 3180
rect -9125 3163 -9108 3180
rect -8965 3163 -8948 3180
rect -9045 3163 -9028 3180
rect -8725 3163 -8708 3180
rect -8885 3163 -8868 3180
rect -9205 3163 -9188 3180
rect -9245 3163 -9228 3180
rect -9365 3163 -9348 3180
rect -9285 3163 -9268 3180
rect -9325 3163 -9308 3180
rect -9365 3163 -9348 3180
rect -9285 3163 -9268 3180
rect -9405 3163 -9388 3180
rect -9405 3163 -9388 3180
rect -9285 3163 -9268 3180
rect -9245 3163 -9228 3180
rect -9325 3163 -9308 3180
rect -9325 3163 -9308 3180
rect -9365 3163 -9348 3180
rect -9405 3163 -9388 3180
rect -9245 3163 -9228 3180
rect -9405 3163 -9388 3180
rect -9365 3163 -9348 3180
rect -9285 3163 -9268 3180
rect -9325 3163 -9308 3180
rect -9245 3163 -9228 3180
rect -4885 3163 -4868 3180
rect -4725 3163 -4708 3180
rect -4725 3163 -4708 3180
rect -4725 3163 -4708 3180
rect -4845 3163 -4828 3180
rect -4725 3163 -4708 3180
rect -4765 3163 -4748 3180
rect -4805 3163 -4788 3180
rect -4885 3163 -4868 3180
rect -4765 3163 -4748 3180
rect -4765 3163 -4748 3180
rect -4805 3163 -4788 3180
rect -4685 3163 -4668 3180
rect -4805 3163 -4788 3180
rect -4885 3163 -4868 3180
rect -4805 3163 -4788 3180
rect -4845 3163 -4828 3180
rect -4685 3163 -4668 3180
rect -4765 3163 -4748 3180
rect -4845 3163 -4828 3180
rect -4845 3163 -4828 3180
rect -4685 3163 -4668 3180
rect -4885 3163 -4868 3180
rect -4685 3163 -4668 3180
rect -5445 3163 -5428 3180
rect -5445 3163 -5428 3180
rect -5445 3163 -5428 3180
rect -5445 3163 -5428 3180
rect -5405 3163 -5388 3180
rect -5085 3163 -5068 3180
rect -5125 3163 -5108 3180
rect -5165 3163 -5148 3180
rect -5205 3163 -5188 3180
rect -5085 3163 -5068 3180
rect -5285 3163 -5268 3180
rect -4925 3163 -4908 3180
rect -4965 3163 -4948 3180
rect -4965 3163 -4948 3180
rect -5045 3163 -5028 3180
rect -5325 3163 -5308 3180
rect -4925 3163 -4908 3180
rect -5285 3163 -5268 3180
rect -5365 3163 -5348 3180
rect -5125 3163 -5108 3180
rect -5165 3163 -5148 3180
rect -5325 3163 -5308 3180
rect -5005 3163 -4988 3180
rect -5405 3163 -5388 3180
rect -5125 3163 -5108 3180
rect -5005 3163 -4988 3180
rect -5285 3163 -5268 3180
rect -5325 3163 -5308 3180
rect -5245 3163 -5228 3180
rect -5205 3163 -5188 3180
rect -5165 3163 -5148 3180
rect -4925 3163 -4908 3180
rect -4965 3163 -4948 3180
rect -5245 3163 -5228 3180
rect -5005 3163 -4988 3180
rect -5365 3163 -5348 3180
rect -5045 3163 -5028 3180
rect -5085 3163 -5068 3180
rect -5365 3163 -5348 3180
rect -5125 3163 -5108 3180
rect -4965 3163 -4948 3180
rect -5045 3163 -5028 3180
rect -5285 3163 -5268 3180
rect -5165 3163 -5148 3180
rect -5205 3163 -5188 3180
rect -5325 3163 -5308 3180
rect -5205 3163 -5188 3180
rect -5245 3163 -5228 3180
rect -5365 3163 -5348 3180
rect -5405 3163 -5388 3180
rect -5085 3163 -5068 3180
rect -5405 3163 -5388 3180
rect -5005 3163 -4988 3180
rect -5045 3163 -5028 3180
rect -5245 3163 -5228 3180
rect -4925 3163 -4908 3180
rect -5645 3163 -5628 3180
rect -5845 3163 -5828 3180
rect -5925 3163 -5908 3180
rect -5805 3163 -5788 3180
rect -5845 3163 -5828 3180
rect -5525 3163 -5508 3180
rect -5565 3163 -5548 3180
rect -5885 3163 -5868 3180
rect -5685 3163 -5668 3180
rect -5485 3163 -5468 3180
rect -5605 3163 -5588 3180
rect -5645 3163 -5628 3180
rect -5965 3163 -5948 3180
rect -5765 3163 -5748 3180
rect -5485 3163 -5468 3180
rect -5605 3163 -5588 3180
rect -5965 3163 -5948 3180
rect -5925 3163 -5908 3180
rect -5685 3163 -5668 3180
rect -5685 3163 -5668 3180
rect -5525 3163 -5508 3180
rect -5845 3163 -5828 3180
rect -5645 3163 -5628 3180
rect -5805 3163 -5788 3180
rect -5565 3163 -5548 3180
rect -5685 3163 -5668 3180
rect -5885 3163 -5868 3180
rect -5725 3163 -5708 3180
rect -5605 3163 -5588 3180
rect -5765 3163 -5748 3180
rect -5765 3163 -5748 3180
rect -5965 3163 -5948 3180
rect -5725 3163 -5708 3180
rect -5805 3163 -5788 3180
rect -5525 3163 -5508 3180
rect -5925 3163 -5908 3180
rect -5885 3163 -5868 3180
rect -5765 3163 -5748 3180
rect -5725 3163 -5708 3180
rect -5485 3163 -5468 3180
rect -5845 3163 -5828 3180
rect -5525 3163 -5508 3180
rect -5805 3163 -5788 3180
rect -5965 3163 -5948 3180
rect -5565 3163 -5548 3180
rect -5925 3163 -5908 3180
rect -5485 3163 -5468 3180
rect -5725 3163 -5708 3180
rect -5605 3163 -5588 3180
rect -5885 3163 -5868 3180
rect -5645 3163 -5628 3180
rect -5565 3163 -5548 3180
rect -6525 3163 -6508 3180
rect -6525 3163 -6508 3180
rect -6525 3163 -6508 3180
rect -6525 3163 -6508 3180
rect -6165 3163 -6148 3180
rect -6285 3163 -6268 3180
rect -6205 3163 -6188 3180
rect -6325 3163 -6308 3180
rect -6005 3163 -5988 3180
rect -6045 3163 -6028 3180
rect -6085 3163 -6068 3180
rect -6005 3163 -5988 3180
rect -6125 3163 -6108 3180
rect -6165 3163 -6148 3180
rect -6205 3163 -6188 3180
rect -6245 3163 -6228 3180
rect -6285 3163 -6268 3180
rect -6325 3163 -6308 3180
rect -6365 3163 -6348 3180
rect -6405 3163 -6388 3180
rect -6165 3163 -6148 3180
rect -6205 3163 -6188 3180
rect -6245 3163 -6228 3180
rect -6485 3163 -6468 3180
rect -6205 3163 -6188 3180
rect -6325 3163 -6308 3180
rect -6005 3163 -5988 3180
rect -6005 3163 -5988 3180
rect -6125 3163 -6108 3180
rect -6125 3163 -6108 3180
rect -6365 3163 -6348 3180
rect -6405 3163 -6388 3180
rect -6285 3163 -6268 3180
rect -6085 3163 -6068 3180
rect -6165 3163 -6148 3180
rect -6245 3163 -6228 3180
rect -6325 3163 -6308 3180
rect -6285 3163 -6268 3180
rect -6045 3163 -6028 3180
rect -6045 3163 -6028 3180
rect -6365 3163 -6348 3180
rect -6365 3163 -6348 3180
rect -6485 3163 -6468 3180
rect -6045 3163 -6028 3180
rect -6405 3163 -6388 3180
rect -6125 3163 -6108 3180
rect -6405 3163 -6388 3180
rect -6085 3163 -6068 3180
rect -6445 3163 -6428 3180
rect -6445 3163 -6428 3180
rect -6445 3163 -6428 3180
rect -6085 3163 -6068 3180
rect -6445 3163 -6428 3180
rect -6245 3163 -6228 3180
rect -6485 3163 -6468 3180
rect -6485 3163 -6468 3180
rect -6685 3163 -6668 3180
rect -7045 3163 -7028 3180
rect -6965 3163 -6948 3180
rect -6565 3163 -6548 3180
rect -6565 3163 -6548 3180
rect -6965 3163 -6948 3180
rect -6845 3163 -6828 3180
rect -6605 3163 -6588 3180
rect -7005 3163 -6988 3180
rect -6765 3163 -6748 3180
rect -7045 3163 -7028 3180
rect -6765 3163 -6748 3180
rect -6965 3163 -6948 3180
rect -6645 3163 -6628 3180
rect -6605 3163 -6588 3180
rect -6925 3163 -6908 3180
rect -6645 3163 -6628 3180
rect -6685 3163 -6668 3180
rect -6805 3163 -6788 3180
rect -6885 3163 -6868 3180
rect -6925 3163 -6908 3180
rect -6925 3163 -6908 3180
rect -6725 3163 -6708 3180
rect -7045 3163 -7028 3180
rect -7005 3163 -6988 3180
rect -6725 3163 -6708 3180
rect -6565 3163 -6548 3180
rect -6765 3163 -6748 3180
rect -6805 3163 -6788 3180
rect -6925 3163 -6908 3180
rect -6845 3163 -6828 3180
rect -7045 3163 -7028 3180
rect -6685 3163 -6668 3180
rect -6885 3163 -6868 3180
rect -6645 3163 -6628 3180
rect -6725 3163 -6708 3180
rect -6605 3163 -6588 3180
rect -6765 3163 -6748 3180
rect -6685 3163 -6668 3180
rect -6645 3163 -6628 3180
rect -6805 3163 -6788 3180
rect -6845 3163 -6828 3180
rect -6965 3163 -6948 3180
rect -6845 3163 -6828 3180
rect -6725 3163 -6708 3180
rect -7005 3163 -6988 3180
rect -6605 3163 -6588 3180
rect -6805 3163 -6788 3180
rect -7005 3163 -6988 3180
rect -6885 3163 -6868 3180
rect -6885 3163 -6868 3180
rect -6565 3163 -6548 3180
rect -7605 3163 -7588 3180
rect -7605 3163 -7588 3180
rect -7605 3163 -7588 3180
rect -7605 3163 -7588 3180
rect -7165 3163 -7148 3180
rect -7445 3163 -7428 3180
rect -7485 3163 -7468 3180
rect -7325 3163 -7308 3180
rect -7405 3163 -7388 3180
rect -7525 3163 -7508 3180
rect -7525 3163 -7508 3180
rect -7485 3163 -7468 3180
rect -7245 3163 -7228 3180
rect -7565 3163 -7548 3180
rect -7405 3163 -7388 3180
rect -7525 3163 -7508 3180
rect -7525 3163 -7508 3180
rect -7125 3163 -7108 3180
rect -7245 3163 -7228 3180
rect -7565 3163 -7548 3180
rect -7445 3163 -7428 3180
rect -7125 3163 -7108 3180
rect -7285 3163 -7268 3180
rect -7445 3163 -7428 3180
rect -7565 3163 -7548 3180
rect -7245 3163 -7228 3180
rect -7165 3163 -7148 3180
rect -7365 3163 -7348 3180
rect -7445 3163 -7428 3180
rect -7405 3163 -7388 3180
rect -7565 3163 -7548 3180
rect -7325 3163 -7308 3180
rect -7285 3163 -7268 3180
rect -7365 3163 -7348 3180
rect -7205 3163 -7188 3180
rect -7085 3163 -7068 3180
rect -7325 3163 -7308 3180
rect -7085 3163 -7068 3180
rect -7125 3163 -7108 3180
rect -7285 3163 -7268 3180
rect -7485 3163 -7468 3180
rect -7365 3163 -7348 3180
rect -7365 3163 -7348 3180
rect -7205 3163 -7188 3180
rect -7165 3163 -7148 3180
rect -7245 3163 -7228 3180
rect -7085 3163 -7068 3180
rect -7285 3163 -7268 3180
rect -7085 3163 -7068 3180
rect -7125 3163 -7108 3180
rect -7165 3163 -7148 3180
rect -7205 3163 -7188 3180
rect -7325 3163 -7308 3180
rect -7205 3163 -7188 3180
rect -7485 3163 -7468 3180
rect -7405 3163 -7388 3180
rect -7765 3163 -7748 3180
rect -7645 3163 -7628 3180
rect -7845 3163 -7828 3180
rect -7965 3163 -7948 3180
rect -8045 3163 -8028 3180
rect -8005 3163 -7988 3180
rect -7685 3163 -7668 3180
rect -7725 3163 -7708 3180
rect -8125 3163 -8108 3180
rect -7805 3163 -7788 3180
rect -7925 3163 -7908 3180
rect -7885 3163 -7868 3180
rect -7685 3163 -7668 3180
rect -7925 3163 -7908 3180
rect -8085 3163 -8068 3180
rect -8085 3163 -8068 3180
rect -7725 3163 -7708 3180
rect -8045 3163 -8028 3180
rect -7845 3163 -7828 3180
rect -7965 3163 -7948 3180
rect -7725 3163 -7708 3180
rect -7805 3163 -7788 3180
rect -7765 3163 -7748 3180
rect -7845 3163 -7828 3180
rect -8125 3163 -8108 3180
rect -7845 3163 -7828 3180
rect -7885 3163 -7868 3180
rect -8045 3163 -8028 3180
rect -8085 3163 -8068 3180
rect -7725 3163 -7708 3180
rect -7645 3163 -7628 3180
rect -7885 3163 -7868 3180
rect -7685 3163 -7668 3180
rect -7805 3163 -7788 3180
rect -8005 3163 -7988 3180
rect -7885 3163 -7868 3180
rect -7965 3163 -7948 3180
rect -7805 3163 -7788 3180
rect -7925 3163 -7908 3180
rect -8125 3163 -8108 3180
rect -8005 3163 -7988 3180
rect -7685 3163 -7668 3180
rect -7925 3163 -7908 3180
rect -8005 3163 -7988 3180
rect -8125 3163 -8108 3180
rect -7645 3163 -7628 3180
rect -8045 3163 -8028 3180
rect -7965 3163 -7948 3180
rect -7765 3163 -7748 3180
rect -8085 3163 -8068 3180
rect -7645 3163 -7628 3180
rect -7765 3163 -7748 3180
rect -8685 3163 -8668 3180
rect -8685 3163 -8668 3180
rect -8685 3163 -8668 3180
rect -8685 3163 -8668 3180
rect -8205 3163 -8188 3180
rect -8285 3163 -8268 3180
rect -8605 3163 -8588 3180
rect -8365 3163 -8348 3180
rect -8525 3163 -8508 3180
rect -8485 3163 -8468 3180
rect -8645 3163 -8628 3180
rect -8285 3163 -8268 3180
rect -8205 3163 -8188 3180
rect -8405 3163 -8388 3180
rect -8445 3163 -8428 3180
rect -8285 3163 -8268 3180
rect -8165 3163 -8148 3180
rect -8605 3163 -8588 3180
rect -8325 3163 -8308 3180
rect -8325 3163 -8308 3180
rect -8405 3163 -8388 3180
rect -8565 3163 -8548 3180
rect -8525 3163 -8508 3180
rect -8365 3163 -8348 3180
rect -8485 3163 -8468 3180
rect -8325 3163 -8308 3180
rect -8405 3163 -8388 3180
rect -8165 3163 -8148 3180
rect -8525 3163 -8508 3180
rect -8205 3163 -8188 3180
rect -8245 3163 -8228 3180
rect -8325 3163 -8308 3180
rect -8605 3163 -8588 3180
rect -8205 3163 -8188 3180
rect -8525 3163 -8508 3180
rect -9292 2394 -9275 2411
rect -8492 2394 -8475 2411
rect -9332 2394 -9315 2411
rect -9372 2394 -9355 2411
rect -8772 2394 -8755 2411
rect -8572 2394 -8555 2411
rect -8812 2394 -8795 2411
rect -9372 2394 -9355 2411
rect -9012 2394 -8995 2411
rect -9052 2394 -9035 2411
rect -9092 2394 -9075 2411
rect -9132 2394 -9115 2411
rect -9172 2394 -9155 2411
rect -9212 2394 -9195 2411
rect -9252 2394 -9235 2411
rect -8852 2394 -8835 2411
rect -8892 2394 -8875 2411
rect -8932 2394 -8915 2411
rect -8972 2394 -8955 2411
rect -9012 2394 -8995 2411
rect -9052 2394 -9035 2411
rect -9092 2394 -9075 2411
rect -9132 2394 -9115 2411
rect -9172 2394 -9155 2411
rect -9212 2394 -9195 2411
rect -9252 2394 -9235 2411
rect -8852 2394 -8835 2411
rect -8892 2394 -8875 2411
rect -8772 2394 -8755 2411
rect -8972 2394 -8955 2411
rect -8372 2394 -8355 2411
rect -8692 2394 -8675 2411
rect -8652 2394 -8635 2411
rect -8652 2394 -8635 2411
rect -8412 2394 -8395 2411
rect -8252 2394 -8235 2411
rect -8292 2394 -8275 2411
rect -9292 2394 -9275 2411
rect -8332 2394 -8315 2411
rect -8252 2394 -8235 2411
rect -9332 2394 -9315 2411
rect -8732 2394 -8715 2411
rect -8532 2394 -8515 2411
rect -8532 2394 -8515 2411
rect -8732 2394 -8715 2411
rect -8332 2394 -8315 2411
rect -8492 2394 -8475 2411
rect -8292 2394 -8275 2411
rect -8692 2394 -8675 2411
rect -8612 2394 -8595 2411
rect -8452 2394 -8435 2411
rect -8372 2394 -8355 2411
rect -8452 2394 -8435 2411
rect -8932 2394 -8915 2411
rect -8412 2394 -8395 2411
rect -8812 2394 -8795 2411
rect -8572 2394 -8555 2411
rect -8612 2394 -8595 2411
rect -7612 2394 -7595 2411
rect -7772 2394 -7755 2411
rect -7852 2394 -7835 2411
rect -7732 2394 -7715 2411
rect -7092 2394 -7075 2411
rect -7972 2394 -7955 2411
rect -8052 2394 -8035 2411
rect -8172 2394 -8155 2411
rect -8052 2394 -8035 2411
rect -7772 2394 -7755 2411
rect -7492 2394 -7475 2411
rect -7852 2394 -7835 2411
rect -7932 2394 -7915 2411
rect -8172 2394 -8155 2411
rect -7332 2394 -7315 2411
rect -7652 2394 -7635 2411
rect -7572 2394 -7555 2411
rect -8012 2394 -7995 2411
rect -7692 2394 -7675 2411
rect -7572 2394 -7555 2411
rect -7132 2394 -7115 2411
rect -7372 2394 -7355 2411
rect -7732 2394 -7715 2411
rect -7652 2394 -7635 2411
rect -7972 2394 -7955 2411
rect -8012 2394 -7995 2411
rect -7332 2394 -7315 2411
rect -7612 2394 -7595 2411
rect -8132 2394 -8115 2411
rect -7452 2394 -7435 2411
rect -7372 2394 -7355 2411
rect -7172 2394 -7155 2411
rect -7292 2394 -7275 2411
rect -7412 2394 -7395 2411
rect -7052 2394 -7035 2411
rect -7532 2394 -7515 2411
rect -7052 2394 -7035 2411
rect -7452 2394 -7435 2411
rect -7092 2394 -7075 2411
rect -7212 2394 -7195 2411
rect -7412 2394 -7395 2411
rect -7252 2394 -7235 2411
rect -7132 2394 -7115 2411
rect -7692 2394 -7675 2411
rect -7172 2394 -7155 2411
rect -7492 2394 -7475 2411
rect -7212 2394 -7195 2411
rect -7292 2394 -7275 2411
rect -7252 2394 -7235 2411
rect -7532 2394 -7515 2411
rect -8092 2394 -8075 2411
rect -8212 2394 -8195 2411
rect -8092 2394 -8075 2411
rect -7892 2394 -7875 2411
rect -7892 2394 -7875 2411
rect -8212 2394 -8195 2411
rect -7812 2394 -7795 2411
rect -7812 2394 -7795 2411
rect -8132 2394 -8115 2411
rect -7932 2394 -7915 2411
rect -5852 2394 -5835 2411
rect -5852 2394 -5835 2411
rect -6852 2394 -6835 2411
rect -6892 2394 -6875 2411
rect -6932 2394 -6915 2411
rect -6932 2394 -6915 2411
rect -6772 2394 -6755 2411
rect -6972 2394 -6955 2411
rect -7012 2394 -6995 2411
rect -6692 2394 -6675 2411
rect -6732 2394 -6715 2411
rect -6972 2394 -6955 2411
rect -6372 2394 -6355 2411
rect -6132 2394 -6115 2411
rect -6412 2394 -6395 2411
rect -6332 2394 -6315 2411
rect -5892 2394 -5875 2411
rect -5892 2394 -5875 2411
rect -6412 2394 -6395 2411
rect -6572 2394 -6555 2411
rect -6292 2394 -6275 2411
rect -6292 2394 -6275 2411
rect -6372 2394 -6355 2411
rect -5932 2394 -5915 2411
rect -6452 2394 -6435 2411
rect -6052 2394 -6035 2411
rect -6092 2394 -6075 2411
rect -6452 2394 -6435 2411
rect -6332 2394 -6315 2411
rect -6172 2394 -6155 2411
rect -6492 2394 -6475 2411
rect -6772 2394 -6755 2411
rect -6892 2394 -6875 2411
rect -6532 2394 -6515 2411
rect -6132 2394 -6115 2411
rect -6492 2394 -6475 2411
rect -6652 2394 -6635 2411
rect -6652 2394 -6635 2411
rect -6572 2394 -6555 2411
rect -6212 2394 -6195 2411
rect -6172 2394 -6155 2411
rect -5932 2394 -5915 2411
rect -5972 2394 -5955 2411
rect -6612 2394 -6595 2411
rect -6052 2394 -6035 2411
rect -6092 2394 -6075 2411
rect -6212 2394 -6195 2411
rect -6012 2394 -5995 2411
rect -6612 2394 -6595 2411
rect -6012 2394 -5995 2411
rect -6252 2394 -6235 2411
rect -6252 2394 -6235 2411
rect -5972 2394 -5955 2411
rect -6532 2394 -6515 2411
rect -6812 2394 -6795 2411
rect -6692 2394 -6675 2411
rect -6852 2394 -6835 2411
rect -6732 2394 -6715 2411
rect -7012 2394 -6995 2411
rect -6812 2394 -6795 2411
rect -5092 2394 -5075 2411
rect -5172 2394 -5155 2411
rect -5132 2394 -5115 2411
rect -5172 2394 -5155 2411
rect -5212 2394 -5195 2411
rect -5252 2394 -5235 2411
rect -5292 2394 -5275 2411
rect -5332 2394 -5315 2411
rect -5372 2394 -5355 2411
rect -5412 2394 -5395 2411
rect -5452 2394 -5435 2411
rect -5492 2394 -5475 2411
rect -5532 2394 -5515 2411
rect -5572 2394 -5555 2411
rect -5212 2394 -5195 2411
rect -5772 2394 -5755 2411
rect -5732 2394 -5715 2411
rect -4732 2394 -4715 2411
rect -5252 2394 -5235 2411
rect -5412 2394 -5395 2411
rect -5292 2394 -5275 2411
rect -5612 2394 -5595 2411
rect -5332 2394 -5315 2411
rect -5452 2394 -5435 2411
rect -5692 2394 -5675 2411
rect -4772 2394 -4755 2411
rect -5492 2394 -5475 2411
rect -5532 2394 -5515 2411
rect -5092 2394 -5075 2411
rect -5612 2394 -5595 2411
rect -5652 2394 -5635 2411
rect -5692 2394 -5675 2411
rect -5732 2394 -5715 2411
rect -5572 2394 -5555 2411
rect -5772 2394 -5755 2411
rect -5812 2394 -5795 2411
rect -4852 2394 -4835 2411
rect -4892 2394 -4875 2411
rect -5132 2394 -5115 2411
rect -4932 2394 -4915 2411
rect -4692 2394 -4675 2411
rect -5652 2394 -5635 2411
rect -4692 2394 -4675 2411
rect -4812 2394 -4795 2411
rect -5812 2394 -5795 2411
rect -5012 2394 -4995 2411
rect -4732 2394 -4715 2411
rect -5052 2394 -5035 2411
rect -4772 2394 -4755 2411
rect -4812 2394 -4795 2411
rect -4852 2394 -4835 2411
rect -4892 2394 -4875 2411
rect -4932 2394 -4915 2411
rect -4972 2394 -4955 2411
rect -4972 2394 -4955 2411
rect -5012 2394 -4995 2411
rect -5372 2394 -5355 2411
rect -5052 2394 -5035 2411
rect -3445 3163 -3428 3180
rect -3325 3163 -3308 3180
rect -3365 3163 -3348 3180
rect -3405 3163 -3388 3180
rect -3445 3163 -3428 3180
rect -3365 3163 -3348 3180
rect 36 3163 53 3180
rect -3365 3163 -3348 3180
rect -3765 3163 -3748 3180
rect -3685 3163 -3668 3180
rect -3685 3163 -3668 3180
rect -3405 3163 -3388 3180
rect -3605 3163 -3588 3180
rect -3445 3163 -3428 3180
rect -3445 3163 -3428 3180
rect -3725 3163 -3708 3180
rect -3325 3163 -3308 3180
rect -3405 3163 -3388 3180
rect -3325 3163 -3308 3180
rect -165 3163 -148 3180
rect -325 3163 -308 3180
rect -405 3163 -388 3180
rect -525 3163 -508 3180
rect -445 3163 -428 3180
rect -125 3163 -108 3180
rect -205 3163 -188 3180
rect -85 3163 -68 3180
rect -405 3163 -388 3180
rect -125 3163 -108 3180
rect -445 3163 -428 3180
rect -285 3163 -268 3180
rect -405 3163 -388 3180
rect -445 3163 -428 3180
rect -365 3163 -348 3180
rect -325 3163 -308 3180
rect -85 3163 -68 3180
rect -405 3163 -388 3180
rect -485 3163 -468 3180
rect -45 3163 -28 3180
rect -445 3163 -428 3180
rect -45 3163 -28 3180
rect -565 3163 -548 3180
rect -245 3163 -228 3180
rect -245 3163 -228 3180
rect -565 3163 -548 3180
rect -245 3163 -228 3180
rect -205 3163 -188 3180
rect -165 3163 -148 3180
rect -565 3163 -548 3180
rect -565 3163 -548 3180
rect -205 3163 -188 3180
rect -485 3163 -468 3180
rect -325 3163 -308 3180
rect -365 3163 -348 3180
rect -245 3163 -228 3180
rect -125 3163 -108 3180
rect -365 3163 -348 3180
rect -525 3163 -508 3180
rect -525 3163 -508 3180
rect -285 3163 -268 3180
rect -85 3163 -68 3180
rect -485 3163 -468 3180
rect -45 3163 -28 3180
rect -45 3163 -28 3180
rect -325 3163 -308 3180
rect -525 3163 -508 3180
rect -125 3163 -108 3180
rect -205 3163 -188 3180
rect -165 3163 -148 3180
rect -85 3163 -68 3180
rect -365 3163 -348 3180
rect -285 3163 -268 3180
rect -485 3163 -468 3180
rect -165 3163 -148 3180
rect -285 3163 -268 3180
rect -685 3163 -668 3180
rect -1005 3163 -988 3180
rect -685 3163 -668 3180
rect -685 3163 -668 3180
rect -1005 3163 -988 3180
rect -885 3163 -868 3180
rect -765 3163 -748 3180
rect -1045 3163 -1028 3180
rect -845 3163 -828 3180
rect -605 3163 -588 3180
rect -885 3163 -868 3180
rect -725 3163 -708 3180
rect -965 3163 -948 3180
rect -805 3163 -788 3180
rect -1045 3163 -1028 3180
rect -1085 3163 -1068 3180
rect -605 3163 -588 3180
rect -645 3163 -628 3180
rect -845 3163 -828 3180
rect -1085 3163 -1068 3180
rect -1085 3163 -1068 3180
rect -725 3163 -708 3180
rect -925 3163 -908 3180
rect -725 3163 -708 3180
rect -605 3163 -588 3180
rect -925 3163 -908 3180
rect -685 3163 -668 3180
rect -965 3163 -948 3180
rect -925 3163 -908 3180
rect -725 3163 -708 3180
rect -645 3163 -628 3180
rect -885 3163 -868 3180
rect -845 3163 -828 3180
rect -845 3163 -828 3180
rect -765 3163 -748 3180
rect -925 3163 -908 3180
rect -805 3163 -788 3180
rect -765 3163 -748 3180
rect -885 3163 -868 3180
rect -605 3163 -588 3180
rect -645 3163 -628 3180
rect -965 3163 -948 3180
rect -1045 3163 -1028 3180
rect -1005 3163 -988 3180
rect -965 3163 -948 3180
rect -645 3163 -628 3180
rect -805 3163 -788 3180
rect -1005 3163 -988 3180
rect -1045 3163 -1028 3180
rect -1085 3163 -1068 3180
rect -765 3163 -748 3180
rect -805 3163 -788 3180
rect -1645 3163 -1628 3180
rect -1325 3163 -1308 3180
rect -1485 3163 -1468 3180
rect -1205 3163 -1188 3180
rect -1245 3163 -1228 3180
rect -1565 3163 -1548 3180
rect -1405 3163 -1388 3180
rect -1525 3163 -1508 3180
rect -1485 3163 -1468 3180
rect -1485 3163 -1468 3180
rect -1325 3163 -1308 3180
rect -1125 3163 -1108 3180
rect -1445 3163 -1428 3180
rect -1645 3163 -1628 3180
rect -1325 3163 -1308 3180
rect -1605 3163 -1588 3180
rect -1365 3163 -1348 3180
rect -1565 3163 -1548 3180
rect -1405 3163 -1388 3180
rect -1245 3163 -1228 3180
rect -1205 3163 -1188 3180
rect -1285 3163 -1268 3180
rect -1525 3163 -1508 3180
rect -1645 3163 -1628 3180
rect -1605 3163 -1588 3180
rect -1525 3163 -1508 3180
rect -1205 3163 -1188 3180
rect -1525 3163 -1508 3180
rect -1325 3163 -1308 3180
rect -1285 3163 -1268 3180
rect -1165 3163 -1148 3180
rect -1565 3163 -1548 3180
rect -1565 3163 -1548 3180
rect -1245 3163 -1228 3180
rect -1285 3163 -1268 3180
rect -1445 3163 -1428 3180
rect -1285 3163 -1268 3180
rect -1205 3163 -1188 3180
rect -1605 3163 -1588 3180
rect -1405 3163 -1388 3180
rect -1365 3163 -1348 3180
rect -1125 3163 -1108 3180
rect -1365 3163 -1348 3180
rect -1165 3163 -1148 3180
rect -1245 3163 -1228 3180
rect -1605 3163 -1588 3180
rect -1125 3163 -1108 3180
rect -1485 3163 -1468 3180
rect -1405 3163 -1388 3180
rect -1365 3163 -1348 3180
rect -1125 3163 -1108 3180
rect -1445 3163 -1428 3180
rect -1445 3163 -1428 3180
rect -1165 3163 -1148 3180
rect -1645 3163 -1628 3180
rect -1165 3163 -1148 3180
rect -3645 3163 -3628 3180
rect -3325 3163 -3308 3180
rect -3365 3163 -3348 3180
rect -3525 3163 -3508 3180
rect -3405 3163 -3388 3180
rect -3805 3163 -3788 3180
rect -3485 3163 -3468 3180
rect -3565 3163 -3548 3180
rect -3485 3163 -3468 3180
rect -3485 3163 -3468 3180
rect -3525 3163 -3508 3180
rect -3525 3163 -3508 3180
rect -3565 3163 -3548 3180
rect -3605 3163 -3588 3180
rect -3645 3163 -3628 3180
rect -3605 3163 -3588 3180
rect -3685 3163 -3668 3180
rect -3725 3163 -3708 3180
rect -3765 3163 -3748 3180
rect -3805 3163 -3788 3180
rect -3725 3163 -3708 3180
rect -3565 3163 -3548 3180
rect -3645 3163 -3628 3180
rect -3605 3163 -3588 3180
rect -3685 3163 -3668 3180
rect -3565 3163 -3548 3180
rect -3645 3163 -3628 3180
rect -3765 3163 -3748 3180
rect -3725 3163 -3708 3180
rect -3805 3163 -3788 3180
rect -3525 3163 -3508 3180
rect -3765 3163 -3748 3180
rect -3485 3163 -3468 3180
rect -3805 3163 -3788 3180
rect -4365 3163 -4348 3180
rect -4365 3163 -4348 3180
rect -4365 3163 -4348 3180
rect -4365 3163 -4348 3180
rect -4325 3163 -4308 3180
rect -3885 3163 -3868 3180
rect -4205 3163 -4188 3180
rect -4125 3163 -4108 3180
rect -4245 3163 -4228 3180
rect -4085 3163 -4068 3180
rect -4125 3163 -4108 3180
rect -4165 3163 -4148 3180
rect -4205 3163 -4188 3180
rect -4245 3163 -4228 3180
rect -4285 3163 -4268 3180
rect -4325 3163 -4308 3180
rect -4085 3163 -4068 3180
rect -4325 3163 -4308 3180
rect -4205 3163 -4188 3180
rect -4125 3163 -4108 3180
rect -4285 3163 -4268 3180
rect -4285 3163 -4268 3180
rect -4085 3163 -4068 3180
rect -4165 3163 -4148 3180
rect -4165 3163 -4148 3180
rect -4245 3163 -4228 3180
rect -4245 3163 -4228 3180
rect -4165 3163 -4148 3180
rect -4325 3163 -4308 3180
rect -4085 3163 -4068 3180
rect -4205 3163 -4188 3180
rect -4125 3163 -4108 3180
rect -4285 3163 -4268 3180
rect -3885 3163 -3868 3180
rect -3925 3163 -3908 3180
rect -3925 3163 -3908 3180
rect -3925 3163 -3908 3180
rect -4045 3163 -4028 3180
rect -3845 3163 -3828 3180
rect -4045 3163 -4028 3180
rect -3965 3163 -3948 3180
rect -3885 3163 -3868 3180
rect -3885 3163 -3868 3180
rect -3965 3163 -3948 3180
rect -3925 3163 -3908 3180
rect -3845 3163 -3828 3180
rect -3965 3163 -3948 3180
rect -4005 3163 -3988 3180
rect -4005 3163 -3988 3180
rect -4045 3163 -4028 3180
rect -4005 3163 -3988 3180
rect -4045 3163 -4028 3180
rect -3965 3163 -3948 3180
rect -3845 3163 -3828 3180
rect -4005 3163 -3988 3180
rect -3845 3163 -3828 3180
rect -4405 3163 -4388 3180
rect -4565 3163 -4548 3180
rect -4565 3163 -4548 3180
rect -4445 3163 -4428 3180
rect -4565 3163 -4548 3180
rect -4405 3163 -4388 3180
rect -4445 3163 -4428 3180
rect -4445 3163 -4428 3180
rect -4605 3163 -4588 3180
rect -4525 3163 -4508 3180
rect -4525 3163 -4508 3180
rect -4485 3163 -4468 3180
rect -4485 3163 -4468 3180
rect -4485 3163 -4468 3180
rect -4405 3163 -4388 3180
rect -4485 3163 -4468 3180
rect -4605 3163 -4588 3180
rect -4645 3163 -4628 3180
rect -4525 3163 -4508 3180
rect -4605 3163 -4588 3180
rect -4605 3163 -4588 3180
rect -4645 3163 -4628 3180
rect -4525 3163 -4508 3180
rect -4645 3163 -4628 3180
rect -4645 3163 -4628 3180
rect -4445 3163 -4428 3180
rect -4565 3163 -4548 3180
rect -4405 3163 -4388 3180
rect -1965 3163 -1948 3180
rect -2005 3163 -1988 3180
rect -2045 3163 -2028 3180
rect -2085 3163 -2068 3180
rect -2125 3163 -2108 3180
rect -2165 3163 -2148 3180
rect -2205 3163 -2188 3180
rect -1685 3163 -1668 3180
rect -1725 3163 -1708 3180
rect -1765 3163 -1748 3180
rect -1805 3163 -1788 3180
rect -1845 3163 -1828 3180
rect -1885 3163 -1868 3180
rect -1925 3163 -1908 3180
rect -1965 3163 -1948 3180
rect -2005 3163 -1988 3180
rect -2045 3163 -2028 3180
rect -2085 3163 -2068 3180
rect -2125 3163 -2108 3180
rect -2165 3163 -2148 3180
rect -2205 3163 -2188 3180
rect -2205 3163 -2188 3180
rect -1765 3163 -1748 3180
rect -1805 3163 -1788 3180
rect -1845 3163 -1828 3180
rect -1885 3163 -1868 3180
rect -1925 3163 -1908 3180
rect -1965 3163 -1948 3180
rect -2005 3163 -1988 3180
rect -2045 3163 -2028 3180
rect -2085 3163 -2068 3180
rect -2125 3163 -2108 3180
rect -2205 3163 -2188 3180
rect -2165 3163 -2148 3180
rect -1685 3163 -1668 3180
rect -1725 3163 -1708 3180
rect -1685 3163 -1668 3180
rect -1725 3163 -1708 3180
rect -1765 3163 -1748 3180
rect -1805 3163 -1788 3180
rect -1845 3163 -1828 3180
rect -1885 3163 -1868 3180
rect -1925 3163 -1908 3180
rect -1685 3163 -1668 3180
rect -1725 3163 -1708 3180
rect -1765 3163 -1748 3180
rect -1805 3163 -1788 3180
rect -1845 3163 -1828 3180
rect -1885 3163 -1868 3180
rect -1925 3163 -1908 3180
rect -1965 3163 -1948 3180
rect -2005 3163 -1988 3180
rect -2045 3163 -2028 3180
rect -2085 3163 -2068 3180
rect -2125 3163 -2108 3180
rect -2165 3163 -2148 3180
rect -2565 3163 -2548 3180
rect -2285 3163 -2268 3180
rect -2485 3163 -2468 3180
rect -2285 3163 -2268 3180
rect -2605 3163 -2588 3180
rect -2325 3163 -2308 3180
rect -2405 3163 -2388 3180
rect -2285 3163 -2268 3180
rect -2725 3163 -2708 3180
rect -2365 3163 -2348 3180
rect -2365 3163 -2348 3180
rect -2325 3163 -2308 3180
rect -2365 3163 -2348 3180
rect -2405 3163 -2388 3180
rect -2405 3163 -2388 3180
rect -2685 3163 -2668 3180
rect -2445 3163 -2428 3180
rect -2445 3163 -2428 3180
rect -2445 3163 -2428 3180
rect -2725 3163 -2708 3180
rect -2245 3163 -2228 3180
rect -2485 3163 -2468 3180
rect -2485 3163 -2468 3180
rect -2365 3163 -2348 3180
rect -2525 3163 -2508 3180
rect -2525 3163 -2508 3180
rect -2525 3163 -2508 3180
rect -2645 3163 -2628 3180
rect -2245 3163 -2228 3180
rect -2565 3163 -2548 3180
rect -2565 3163 -2548 3180
rect -2405 3163 -2388 3180
rect -2245 3163 -2228 3180
rect -2605 3163 -2588 3180
rect -2605 3163 -2588 3180
rect -2245 3163 -2228 3180
rect -2645 3163 -2628 3180
rect -2325 3163 -2308 3180
rect -2445 3163 -2428 3180
rect -2685 3163 -2668 3180
rect -2725 3163 -2708 3180
rect -2605 3163 -2588 3180
rect -2485 3163 -2468 3180
rect -2565 3163 -2548 3180
rect -2645 3163 -2628 3180
rect -2685 3163 -2668 3180
rect -2725 3163 -2708 3180
rect -2645 3163 -2628 3180
rect -2285 3163 -2268 3180
rect -2325 3163 -2308 3180
rect -2525 3163 -2508 3180
rect -2685 3163 -2668 3180
rect -3005 3163 -2988 3180
rect -3045 3163 -3028 3180
rect -2845 3163 -2828 3180
rect -3085 3163 -3068 3180
rect -3125 3163 -3108 3180
rect -3165 3163 -3148 3180
rect -3205 3163 -3188 3180
rect -3245 3163 -3228 3180
rect -3285 3163 -3268 3180
rect -3045 3163 -3028 3180
rect -3085 3163 -3068 3180
rect -3125 3163 -3108 3180
rect -3165 3163 -3148 3180
rect -3205 3163 -3188 3180
rect -2885 3163 -2868 3180
rect -3245 3163 -3228 3180
rect -2925 3163 -2908 3180
rect -3285 3163 -3268 3180
rect -3005 3163 -2988 3180
rect -2885 3163 -2868 3180
rect -2925 3163 -2908 3180
rect -2885 3163 -2868 3180
rect -2965 3163 -2948 3180
rect -2925 3163 -2908 3180
rect -3005 3163 -2988 3180
rect -2965 3163 -2948 3180
rect -3045 3163 -3028 3180
rect -3005 3163 -2988 3180
rect -3085 3163 -3068 3180
rect -2885 3163 -2868 3180
rect -3125 3163 -3108 3180
rect -2925 3163 -2908 3180
rect -3165 3163 -3148 3180
rect -3205 3163 -3188 3180
rect -2805 3163 -2788 3180
rect 76 3163 93 3180
rect -2845 3163 -2828 3180
rect -3245 3163 -3228 3180
rect 76 3163 93 3180
rect -3285 3163 -3268 3180
rect -2765 3163 -2748 3180
rect -2805 3163 -2788 3180
rect -5 3163 13 3180
rect -2845 3163 -2828 3180
rect 36 3163 53 3180
rect -2965 3163 -2948 3180
rect 76 3163 93 3180
rect -3045 3163 -3028 3180
rect -5 3163 13 3180
rect -3085 3163 -3068 3180
rect -2765 3163 -2748 3180
rect 36 3163 53 3180
rect -3125 3163 -3108 3180
rect -5 3163 13 3180
rect -2805 3163 -2788 3180
rect -2765 3163 -2748 3180
rect -2805 3163 -2788 3180
rect -2845 3163 -2828 3180
rect -2765 3163 -2748 3180
rect -5 3163 13 3180
rect 36 3163 53 3180
rect -3165 3163 -3148 3180
rect -3205 3163 -3188 3180
rect -3245 3163 -3228 3180
rect -3285 3163 -3268 3180
rect 76 3163 93 3180
rect -2965 3163 -2948 3180
rect -670 3352 -653 3369
rect -4452 2394 -4435 2411
rect -4332 2394 -4315 2411
rect -4492 2394 -4475 2411
rect -4532 2394 -4515 2411
rect -4372 2394 -4355 2411
rect -4252 2394 -4235 2411
rect -4132 2394 -4115 2411
rect -4412 2394 -4395 2411
rect -4212 2394 -4195 2411
rect -4572 2394 -4555 2411
rect -3492 2394 -3475 2411
rect -3532 2394 -3515 2411
rect -4292 2394 -4275 2411
rect -3572 2394 -3555 2411
rect -4372 2394 -4355 2411
rect -3612 2394 -3595 2411
rect -4172 2394 -4155 2411
rect -4292 2394 -4275 2411
rect -3652 2394 -3635 2411
rect -4412 2394 -4395 2411
rect -3692 2394 -3675 2411
rect -4612 2394 -4595 2411
rect -3732 2394 -3715 2411
rect -4332 2394 -4315 2411
rect -3772 2394 -3755 2411
rect -3812 2394 -3795 2411
rect -3852 2394 -3835 2411
rect -3892 2394 -3875 2411
rect -3932 2394 -3915 2411
rect -3972 2394 -3955 2411
rect -4012 2394 -3995 2411
rect -4052 2394 -4035 2411
rect -4092 2394 -4075 2411
rect -4132 2394 -4115 2411
rect -4172 2394 -4155 2411
rect -3492 2394 -3475 2411
rect -3532 2394 -3515 2411
rect -3572 2394 -3555 2411
rect -3612 2394 -3595 2411
rect -3652 2394 -3635 2411
rect -3692 2394 -3675 2411
rect -3732 2394 -3715 2411
rect -4452 2394 -4435 2411
rect -3772 2394 -3755 2411
rect -3812 2394 -3795 2411
rect -4492 2394 -4475 2411
rect -4052 2394 -4035 2411
rect -4212 2394 -4195 2411
rect -3852 2394 -3835 2411
rect -4012 2394 -3995 2411
rect -3892 2394 -3875 2411
rect -4252 2394 -4235 2411
rect -3932 2394 -3915 2411
rect -4092 2394 -4075 2411
rect -3972 2394 -3955 2411
rect -4532 2394 -4515 2411
rect -4572 2394 -4555 2411
rect -4612 2394 -4595 2411
rect -3412 2394 -3395 2411
rect -2532 2394 -2515 2411
rect -2572 2394 -2555 2411
rect -2612 2394 -2595 2411
rect -2652 2394 -2635 2411
rect -2292 2394 -2275 2411
rect -2332 2394 -2315 2411
rect -2292 2394 -2275 2411
rect -2332 2394 -2315 2411
rect -2692 2394 -2675 2411
rect -2732 2394 -2715 2411
rect -2772 2394 -2755 2411
rect -2812 2394 -2795 2411
rect -2492 2394 -2475 2411
rect -2852 2394 -2835 2411
rect -2892 2394 -2875 2411
rect -2532 2394 -2515 2411
rect -2932 2394 -2915 2411
rect -2972 2394 -2955 2411
rect -3452 2394 -3435 2411
rect -3052 2394 -3035 2411
rect -3012 2394 -2995 2411
rect -3012 2394 -2995 2411
rect -2452 2394 -2435 2411
rect -2412 2394 -2395 2411
rect -2372 2394 -2355 2411
rect -2452 2394 -2435 2411
rect -2412 2394 -2395 2411
rect -2372 2394 -2355 2411
rect -3092 2394 -3075 2411
rect -2612 2394 -2595 2411
rect -3132 2394 -3115 2411
rect -3052 2394 -3035 2411
rect -3172 2394 -3155 2411
rect -2812 2394 -2795 2411
rect -3212 2394 -3195 2411
rect -3092 2394 -3075 2411
rect -3252 2394 -3235 2411
rect -3452 2394 -3435 2411
rect -2692 2394 -2675 2411
rect -3292 2394 -3275 2411
rect -3132 2394 -3115 2411
rect -3332 2394 -3315 2411
rect -2852 2394 -2835 2411
rect -3172 2394 -3155 2411
rect -2572 2394 -2555 2411
rect -3212 2394 -3195 2411
rect -2892 2394 -2875 2411
rect -3252 2394 -3235 2411
rect -2732 2394 -2715 2411
rect -3292 2394 -3275 2411
rect -2932 2394 -2915 2411
rect -3332 2394 -3315 2411
rect -2652 2394 -2635 2411
rect -3372 2394 -3355 2411
rect -2972 2394 -2955 2411
rect -3412 2394 -3395 2411
rect -2772 2394 -2755 2411
rect -3372 2394 -3355 2411
rect -2492 2394 -2475 2411
rect -1092 2394 -1075 2411
rect -1092 2394 -1075 2411
rect -1892 2394 -1875 2411
rect -2052 2394 -2035 2411
rect -1292 2394 -1275 2411
rect -2092 2394 -2075 2411
rect -1332 2394 -1315 2411
rect -2132 2394 -2115 2411
rect -1372 2394 -1355 2411
rect -2172 2394 -2155 2411
rect -1492 2394 -1475 2411
rect -1532 2394 -1515 2411
rect -1572 2394 -1555 2411
rect -1612 2394 -1595 2411
rect -1652 2394 -1635 2411
rect -1692 2394 -1675 2411
rect -1732 2394 -1715 2411
rect -1772 2394 -1755 2411
rect -1812 2394 -1795 2411
rect -1852 2394 -1835 2411
rect -1892 2394 -1875 2411
rect -1932 2394 -1915 2411
rect -1972 2394 -1955 2411
rect -2012 2394 -1995 2411
rect -2052 2394 -2035 2411
rect -2092 2394 -2075 2411
rect -2132 2394 -2115 2411
rect -2172 2394 -2155 2411
rect -2212 2394 -2195 2411
rect -2252 2394 -2235 2411
rect -1412 2394 -1395 2411
rect -2212 2394 -2195 2411
rect -1452 2394 -1435 2411
rect -2252 2394 -2235 2411
rect -1492 2394 -1475 2411
rect -1532 2394 -1515 2411
rect -1572 2394 -1555 2411
rect -1612 2394 -1595 2411
rect -1972 2394 -1955 2411
rect -1652 2394 -1635 2411
rect -1932 2394 -1915 2411
rect -1692 2394 -1675 2411
rect -2012 2394 -1995 2411
rect -1732 2394 -1715 2411
rect -1292 2394 -1275 2411
rect -1772 2394 -1755 2411
rect -1332 2394 -1315 2411
rect -1812 2394 -1795 2411
rect -1372 2394 -1355 2411
rect -1852 2394 -1835 2411
rect -1212 2394 -1195 2411
rect -1252 2394 -1235 2411
rect -1132 2394 -1115 2411
rect -1132 2394 -1115 2411
rect -1172 2394 -1155 2411
rect -1212 2394 -1195 2411
rect -1252 2394 -1235 2411
rect -1172 2394 -1155 2411
rect -1412 2394 -1395 2411
rect -1452 2394 -1435 2411
rect -572 2394 -555 2411
rect -612 2394 -595 2411
rect -652 2394 -635 2411
rect -692 2394 -675 2411
rect -732 2394 -715 2411
rect -892 2394 -875 2411
rect -932 2394 -915 2411
rect -972 2394 -955 2411
rect -1012 2394 -995 2411
rect -1052 2394 -1035 2411
rect -932 2394 -915 2411
rect -972 2394 -955 2411
rect -1012 2394 -995 2411
rect -1052 2394 -1035 2411
rect -812 2394 -795 2411
rect -252 2394 -235 2411
rect -292 2394 -275 2411
rect -332 2394 -315 2411
rect -372 2394 -355 2411
rect -412 2394 -395 2411
rect -732 2394 -715 2411
rect -852 2394 -835 2411
rect -772 2394 -755 2411
rect -212 2394 -195 2411
rect -252 2394 -235 2411
rect -292 2394 -275 2411
rect -332 2394 -315 2411
rect -372 2394 -355 2411
rect -772 2394 -755 2411
rect -412 2394 -395 2411
rect -452 2394 -435 2411
rect -212 2394 -195 2411
rect -452 2394 -435 2411
rect -492 2394 -475 2411
rect -532 2394 -515 2411
rect -572 2394 -555 2411
rect -612 2394 -595 2411
rect -652 2394 -635 2411
rect -692 2394 -675 2411
rect -812 2394 -795 2411
rect -852 2394 -835 2411
rect -892 2394 -875 2411
rect -492 2394 -475 2411
rect -532 2394 -515 2411
<< l68d20 >>
rect -701 3344 -678 3377
rect -1825 3344 -701 3377
rect 591 3959 625 3992
rect -1820 3959 591 3992
rect -971 4636 1199 4686
rect -971 4636 1199 4686
rect -971 8565 1199 8615
rect -1668 3147 516 3197
rect -1668 3147 516 3197
rect 1872 4636 4055 4686
rect 14833 4636 17016 4686
rect 12673 4636 14856 4686
rect 16993 4636 19176 4686
rect 15939 2377 18122 2427
rect 13779 2377 15962 2427
rect 11618 2377 13801 2427
rect 9458 2377 11641 2427
rect 7298 2377 9481 2427
rect 5138 2377 7321 2427
rect 2978 2377 5161 2427
rect 818 2377 3001 2427
rect 10513 4636 12696 4686
rect 10513 4636 12696 4686
rect 8353 4636 10536 4686
rect 6192 4636 8375 4686
rect 4032 4636 6215 4686
rect 1872 4636 4055 4686
rect 14833 4636 17016 4686
rect 12673 4636 14856 4686
rect 16993 4636 19176 4686
rect 8353 4636 10536 4686
rect 10513 8565 12696 8615
rect 8353 8565 10536 8615
rect 6192 8565 8375 8615
rect 4032 8565 6215 8615
rect 1872 8565 4055 8615
rect 14833 8565 17016 8615
rect 12673 8565 14856 8615
rect 16993 8565 19176 8615
rect 13454 3147 15637 3197
rect 11294 3147 13477 3197
rect 9133 3147 11316 3197
rect 6973 3147 9156 3197
rect 4813 3147 6996 3197
rect 2653 3147 4836 3197
rect 493 3147 2676 3197
rect 6192 4636 8375 4686
rect 13454 3147 15637 3197
rect 11294 3147 13477 3197
rect 9133 3147 11316 3197
rect 6973 3147 9156 3197
rect 4813 3147 6996 3197
rect 2653 3147 4836 3197
rect 493 3147 2676 3197
rect 4032 4636 6215 4686
rect 13454 3147 15637 3197
rect 11294 3147 13477 3197
rect 9133 3147 11316 3197
rect 13454 3147 15637 3197
rect 11294 3147 13477 3197
rect 9133 3147 11316 3197
rect 15614 3147 17797 3197
rect 15614 3147 17797 3197
rect 15614 3147 17797 3197
rect 15614 3147 17797 3197
rect 625 3959 658 3992
rect -16789 4636 -14606 4686
rect -2355 2377 -172 2427
rect -18949 4636 -16766 4686
rect -3828 4636 -1645 4686
rect -5988 4636 -3805 4686
rect -3828 3147 -1645 3197
rect -5988 3147 -3805 3197
rect -8148 3147 -5965 3197
rect -10308 3147 -8125 3197
rect -12468 3147 -10285 3197
rect -14629 3147 -12446 3197
rect -16789 3147 -14606 3197
rect -18949 3147 -16766 3197
rect -3828 3147 -1645 3197
rect -5988 3147 -3805 3197
rect -8148 3147 -5965 3197
rect -10308 3147 -8125 3197
rect -12468 3147 -10285 3197
rect -14629 3147 -12446 3197
rect -16789 3147 -14606 3197
rect -18949 3147 -16766 3197
rect -8149 4636 -5966 4686
rect -10309 4636 -8126 4686
rect -12469 4636 -10286 4686
rect -14629 4636 -12446 4686
rect -16789 4636 -14606 4686
rect -18949 4636 -16766 4686
rect -4515 2377 -2332 2427
rect -6675 2377 -4492 2427
rect -8835 2377 -6652 2427
rect -10995 2377 -8812 2427
rect -13156 2377 -10973 2427
rect -15316 2377 -13133 2427
rect -17476 2377 -15293 2427
rect -3828 4636 -1645 4686
rect -5988 4636 -3805 4686
rect -3828 8565 -1645 8615
rect -5988 8565 -3805 8615
rect -8149 8565 -5966 8615
rect -10309 8565 -8126 8615
rect -12469 8565 -10286 8615
rect -14629 8565 -12446 8615
rect -16789 8565 -14606 8615
rect -18949 8565 -16766 8615
rect -8149 4636 -5966 4686
rect -10309 4636 -8126 4686
rect -12469 4636 -10286 4686
rect -678 3344 -645 3377
rect -14629 4636 -12446 4686
<< l69d20 >>
rect 807 2546 847 2816
rect 801 2816 847 2946
rect -753 4355 19168 4372
rect 2051 4301 2071 4318
rect 2071 4301 19167 4318
rect 807 2350 847 2546
rect -13 2816 671 2946
<< l71d20 >>
rect -1092 4181 -992 4996
rect -10339 4996 -992 5096
rect -10339 5096 -10239 5636
rect -10339 5636 -10228 5736
rect 1697 4181 1797 5635
rect 1697 5635 9441 5735
<< l70d20 >>
rect -143 3029 -13 3247
rect -143 2946 -13 3029
rect 671 2946 801 3023
rect 671 3023 801 3247
<< l68d16 >>
rect 276 3163 333 3180
rect 236 4652 573 4669
rect -285 8581 52 8598
rect -1730 3965 -1705 3986
rect -1730 3350 -1710 3369
<< l71d44 >>
rect -119 3272 -39 3352
rect 694 3272 774 3352
rect -118 2841 -38 2921
rect 696 2841 776 2921
rect -1905 3319 -1825 3399
rect -1905 3938 -1825 4018
<< l72d20 >>
rect -174 3217 16 3407
rect 639 3217 829 3407
rect -173 2786 18 2976
rect 641 2786 831 2976
rect -1960 3264 -1770 3454
rect -1960 3883 -1770 4073
<< l76d20 >>
rect -183 2776 28 2986
rect -184 3207 26 3417
rect 629 3207 839 3417
rect 631 2776 841 2986
rect -1970 3254 -1760 3464
rect -1970 3873 -1760 4083
<< l69d16 >>
rect 2745 4357 2757 4369
rect 2745 4304 2759 4314
<< labels >>
rlabel l68d16 -1718 3974.5 -1718 3974.5 0 IN1
rlabel l68d16 -1720 3359 -1720 3359 0 IN2
rlabel l68d16 303 3170.5 303 3170.5 0 Ground
rlabel l68d16 501 4659 501 4659 0 VDD
rlabel l68d16 -133.5 8589 -133.5 8589 0 VDD
rlabel l69d16 2751.5 4361.5 2751.5 4361.5 0 OUT1
rlabel l69d16 2751 4308 2751 4308 0 OUT2
use CASCODED_nmos_1v8_lvt_4p5_10finger CASCODED_nmos_1v8_lvt_4p5_10finger_1
timestamp 1670961910
transform 1 0 243 0 1 3308
box -1795 105 -150 635
use CASCODED_nmos_1v8_lvt_4p5_10finger CASCODED_nmos_1v8_lvt_4p5_10finger_2
timestamp 1670961910
transform -1 0 412 0 1 3308
box -1795 105 -150 635
use Vdd_power_rail Vdd_power_rail_1
timestamp 1670961910
transform 1 0 -846 0 1 4056
box -815 580 -125 630
use Vdd_power_rail Vdd_power_rail_2
timestamp 1670961910
transform 1 0 2014 0 1 4056
box -815 580 -125 630
use simple_current_mirror simple_current_mirror_1
timestamp 1670961910
transform 1 0 -53 0 1 1780
box -150 -99 889 647
use Resistor_20k Resistor_20k_1
timestamp 1670961910
transform 1 0 -1206 0 1 3707
box 515 325 1119 866
use Square_Inductor_10t_2s_1w_180dout Square_Inductor_10t_2s_1w_180dout_1
timestamp 1670961910
transform 1 0 -16398 0 1 8326
box -2530 -2690 15070 14910
use Vdd_power_rail Vdd_power_rail_3
timestamp 1670961910
transform 1 0 -846 0 1 4056
box -815 580 -125 630
use Vdd_power_rail Vdd_power_rail_4
timestamp 1670961910
transform 1 0 2014 0 1 4056
box -815 580 -125 630
use Vdd_power_rail Vdd_power_rail_5
timestamp 1670961910
transform 1 0 -846 0 1 7985
box -815 580 -125 630
use Vdd_power_rail Vdd_power_rail_6
timestamp 1670961910
transform 1 0 2014 0 1 7985
box -815 580 -125 630
use M1_vias_M4 M1_vias_M4_1
timestamp 1670961910
transform 1 0 -10117 0 1 8520
box -240 -85 -110 45
use M1_vias_M4 M1_vias_M4_2
timestamp 1670961910
transform 1 0 9551 0 1 8520
box -240 -85 -110 45
use Resistor_20k Resistor_20k_2
timestamp 1670961910
transform 1 0 1567 0 1 3707
box 515 325 1119 866
use Square_Inductor_10t_2s_1w_180dout Square_Inductor_10t_2s_1w_180dout_2
timestamp 1670961910
transform 1 0 3271 0 1 8325
box -2530 -2690 15070 14910
use M1_vias_M4 M1_vias_M4_3
timestamp 1670961910
transform 1 0 1922 0 1 4136
box -240 -85 -110 45
use M1_vias_M4 M1_vias_M4_4
timestamp 1670961910
transform 1 0 -869 0 1 4136
box -240 -85 -110 45
use Via_P_Licon_Li Via_P_Licon_Li_1
timestamp 1670961910
transform 1 0 1194 0 1 3400
box 184 552 217 585
use Via_P_Licon_Li Via_P_Licon_Li_2
timestamp 1670961910
transform 1 0 -1609 0 1 3400
box 184 552 217 585
use Li_via_M2 Li_via_M2_1
timestamp 1670961910
transform 1 0 817 0 1 2320
box -10 -10 30 30
use M1_vias_M4 M1_vias_M4_5
timestamp 1670961910
transform 1 0 96 0 1 3332
box -240 -85 -110 45
use M1_vias_M4 M1_vias_M4_6
timestamp 1670961910
transform 1 0 909 0 1 3332
box -240 -85 -110 45
use M1_vias_M4 M1_vias_M4_7
timestamp 1670961910
transform 1 0 98 0 1 2901
box -240 -85 -110 45
use M1_vias_M4 M1_vias_M4_8
timestamp 1670961910
transform 1 0 911 0 1 2901
box -240 -85 -110 45
use Li_via_M2 Li_via_M2_2
timestamp 1670961910
transform 1 0 -783 0 1 4353
box -10 -10 30 30
use Li_via_M2 Li_via_M2_3
timestamp 1670961910
transform 1 0 2021 0 1 4299
box -10 -10 30 30
use Via_P_Licon_Li Via_P_Licon_Li_3
timestamp 1670961910
transform 1 0 -862 0 1 2792
box 184 552 217 585
use Via_P_Licon_Li Via_P_Licon_Li_4
timestamp 1670961910
transform 1 0 441 0 1 3407
box 184 552 217 585
use M1_vias_M4 M1_vias_M4_9
timestamp 1670961910
transform 1 0 -1690 0 1 3379
box -240 -85 -110 45
use M1_vias_M4 M1_vias_M4_10
timestamp 1670961910
transform 1 0 -1690 0 1 3998
box -240 -85 -110 45
<< end >>
