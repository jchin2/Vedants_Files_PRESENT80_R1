magic
tech sky130A
magscale 1 2
timestamp 1670553586
<< error_p >>
rect -120 0 0 1125
rect 30 0 150 1125
rect 180 0 300 1125
rect 330 0 450 1125
rect 480 0 600 1125
rect 630 0 750 1125
rect 780 0 900 1125
rect 930 0 1050 1125
rect 1080 0 1200 1125
<< nmoslvt >>
rect 0 0 30 1125
rect 150 0 180 1125
rect 300 0 330 1125
rect 450 0 480 1125
rect 600 0 630 1125
rect 750 0 780 1125
rect 900 0 930 1125
rect 1050 0 1080 1125
<< ndiff >>
rect -120 1080 0 1125
rect -120 30 -80 1080
rect -40 30 0 1080
rect -120 0 0 30
rect 30 1080 150 1125
rect 30 30 70 1080
rect 110 30 150 1080
rect 30 0 150 30
rect 180 1080 300 1125
rect 180 30 220 1080
rect 260 30 300 1080
rect 180 0 300 30
rect 330 1080 450 1125
rect 330 30 370 1080
rect 410 30 450 1080
rect 330 0 450 30
rect 480 1080 600 1125
rect 480 30 520 1080
rect 560 30 600 1080
rect 480 0 600 30
rect 630 1080 750 1125
rect 630 30 670 1080
rect 710 30 750 1080
rect 630 0 750 30
rect 780 1080 900 1125
rect 780 30 820 1080
rect 860 30 900 1080
rect 780 0 900 30
rect 930 1080 1050 1125
rect 930 30 970 1080
rect 1010 30 1050 1080
rect 930 0 1050 30
rect 1080 1080 1200 1125
rect 1080 30 1120 1080
rect 1160 30 1200 1080
rect 1080 0 1200 30
<< ndiffc >>
rect -80 30 -40 1080
rect 70 30 110 1080
rect 220 30 260 1080
rect 370 30 410 1080
rect 520 30 560 1080
rect 670 30 710 1080
rect 820 30 860 1080
rect 970 30 1010 1080
rect 1120 30 1160 1080
<< poly >>
rect 0 1125 30 1160
rect 150 1125 180 1160
rect 300 1125 330 1160
rect 450 1125 480 1160
rect 600 1125 630 1160
rect 750 1125 780 1160
rect 900 1125 930 1160
rect 1050 1125 1080 1160
rect 0 -30 30 0
rect 150 -30 180 0
rect 300 -30 330 0
rect 450 -30 480 0
rect 600 -30 630 0
rect 750 -30 780 0
rect 900 -30 930 0
rect 1050 -30 1080 0
<< locali >>
rect -100 1080 -20 1100
rect -100 30 -80 1080
rect -40 30 -20 1080
rect -100 20 -20 30
rect 50 1080 130 1100
rect 50 30 70 1080
rect 110 30 130 1080
rect 50 20 130 30
rect 200 1080 280 1100
rect 200 30 220 1080
rect 260 30 280 1080
rect 200 20 280 30
rect 350 1080 430 1100
rect 350 30 370 1080
rect 410 30 430 1080
rect 350 20 430 30
rect 500 1080 580 1100
rect 500 30 520 1080
rect 560 30 580 1080
rect 500 20 580 30
rect 650 1080 730 1100
rect 650 30 670 1080
rect 710 30 730 1080
rect 650 20 730 30
rect 800 1080 880 1100
rect 800 30 820 1080
rect 860 30 880 1080
rect 800 20 880 30
rect 950 1080 1030 1100
rect 950 30 970 1080
rect 1010 30 1030 1080
rect 950 20 1030 30
rect 1100 1080 1180 1100
rect 1100 30 1120 1080
rect 1160 30 1180 1080
rect 1100 20 1180 30
<< end >>
