* NGSPICE file created from CMOS_s3_flat.ext - technology: sky130A

.subckt CMOS_s3_flat GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar s3 VDD
X0 s3.t1 a_2442_n779# GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_2592_n1689# CMOS_AND_1/AND VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X2 VDD.t9 x3.t0 a_1735_499# VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X3 a_2592_n111# x1.t0 GND.t29 GND.t20 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_2592_499# CMOS_AND_0/A a_2592_n111# GND.t26 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 CMOS_AND_1/AND a_1380_n1689# GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_1380_n1689# x3_bar.t0 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X7 a_2742_n1689# CMOS_AND_0/AND a_2592_n1689# VDD.t34 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X8 VDD.t11 x0.t0 a_177_499# VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X9 CMOS_AND_1/A a_27_n111# VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X10 GND.t21 CMOS_AND_1/AND a_2442_n779# GND.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X11 a_2442_n779# CMOS_AND_0/AND GND.t30 GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 VDD.t36 CMOS_AND_1/A a_1380_n1689# VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X13 GND.t9 x1_bar.t0 a_177_n111# GND.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X14 a_27_n111# x0.t1 a_n123_n111# GND.t3 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X15 VDD.t13 x2_bar.t0 a_n328_n1689# VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X16 a_27_n111# x1.t1 a_n123_499# VDD.t37 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X17 CMOS_3in_OR_0/C.t1 a_n328_n1689# GND.t16 GND.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 GND.t14 CMOS_3in_OR_0/C.t2 a_2442_n779# GND.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 VDD.t1 x3.t1 a_n328_n1689# VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X20 CMOS_AND_0/AND a_2592_499# VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X21 a_1435_n111# x2.t0 GND.t2 GND.t1 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X22 a_1380_n779# x3_bar.t1 GND.t18 GND.t17 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X23 a_1380_n1689# CMOS_AND_1/A a_1380_n779# GND.t31 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X24 s3.t0 a_2442_n779# VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X25 a_1435_499# x3_bar.t2 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X26 a_n123_499# x0_bar.t0 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X27 a_n28_n779# x0.t2 a_n178_n779# GND.t5 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X28 a_n328_n1689# x2_bar.t1 a_n28_n779# GND.t4 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X29 VDD.t29 CMOS_AND_0/A a_2592_499# VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X30 a_n328_n1689# x0.t3 VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X31 CMOS_AND_1/AND a_1380_n1689# VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X32 a_1735_499# x2_bar.t2 CMOS_AND_0/A VDD.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X33 a_177_499# x1_bar.t1 a_27_n111# VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X34 CMOS_AND_0/A x3.t2 a_1435_n111# GND.t0 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X35 a_1735_n111# x3_bar.t3 CMOS_AND_0/A GND.t10 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X36 CMOS_AND_0/AND a_2592_499# GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X37 CMOS_3in_OR_0/C.t0 a_n328_n1689# VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X38 a_2442_n779# CMOS_3in_OR_0/C.t3 a_2742_n1689# VDD.t14 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X39 a_n123_n111# x1.t2 GND.t33 GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X40 a_n178_n779# x3.t3 GND.t12 GND.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X41 a_177_n111# x0_bar.t1 a_27_n111# GND.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X42 a_2592_499# x1.t3 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X43 CMOS_AND_1/A a_27_n111# GND.t25 GND.t24 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X44 GND.t7 x2_bar.t3 a_1735_n111# GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X45 CMOS_AND_0/A x2.t1 a_1435_499# VDD.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
R0 GND.n115 GND.t24 2383.33
R1 GND.n84 GND.t0 159.607
R2 GND.n116 GND.n115 150.98
R3 GND.n150 GND.t3 150.98
R4 GND.n161 GND.t32 133.725
R5 GND.n92 GND.t1 133.725
R6 GND.n142 GND.t19 125.098
R7 GND.n72 GND.t10 125.098
R8 GND.n161 GND.t11 103.529
R9 GND.n45 GND.t20 103.529
R10 GND.n92 GND.t17 103.529
R11 GND.n134 GND.t8 99.215
R12 GND.n63 GND.t6 99.215
R13 GND.n124 GND.t15 77.647
R14 GND.n169 GND.t5 77.647
R15 GND.n5 GND.t22 77.647
R16 GND.n36 GND.t26 77.647
R17 GND.n84 GND.t31 77.647
R18 GND.n146 GND.t4 51.764
R19 GND.n14 GND.t27 51.764
R20 GND.n28 GND.t13 51.764
R21 GND.n63 GND.t34 51.764
R22 GND.n154 GND 37.93
R23 GND.n160 GND.t33 30.21
R24 GND.n155 GND.t12 30.21
R25 GND.n128 GND.t16 30.21
R26 GND.n101 GND.t18 30.21
R27 GND.n67 GND.t35 30.21
R28 GND.n27 GND.t14 30.21
R29 GND.n9 GND.t23 30.21
R30 GND.n18 GND.t28 30.21
R31 GND.n53 GND.t29 30.21
R32 GND.n62 GND.t7 30.21
R33 GND.n96 GND.t2 30.21
R34 GND.n114 GND.t25 30.21
R35 GND.n133 GND.t9 30.21
R36 GND.n0 GND.t30 24
R37 GND.n0 GND.t21 24
R38 GND.n38 GND.n35 11.52
R39 GND.n86 GND.n83 11.52
R40 GND.n3 GND.n2 9.154
R41 GND.n60 GND.n59 9.154
R42 GND.n65 GND.n64 9.154
R43 GND.n64 GND.n63 9.154
R44 GND.n70 GND.n69 9.154
R45 GND.n69 GND.n68 9.154
R46 GND.n74 GND.n73 9.154
R47 GND.n73 GND.n72 9.154
R48 GND.n78 GND.n77 9.154
R49 GND.n77 GND.n76 9.154
R50 GND.n83 GND.n82 9.154
R51 GND.n82 GND.n81 9.154
R52 GND.n86 GND.n85 9.154
R53 GND.n85 GND.n84 9.154
R54 GND.n90 GND.n89 9.154
R55 GND.n89 GND.n88 9.154
R56 GND.n94 GND.n93 9.154
R57 GND.n93 GND.n92 9.154
R58 GND.n99 GND.n98 9.154
R59 GND.n7 GND.n6 9.154
R60 GND.n6 GND.n5 9.154
R61 GND.n12 GND.n11 9.154
R62 GND.n11 GND.n10 9.154
R63 GND.n16 GND.n15 9.154
R64 GND.n15 GND.n14 9.154
R65 GND.n21 GND.n20 9.154
R66 GND.n20 GND.n19 9.154
R67 GND.n25 GND.n24 9.154
R68 GND.n24 GND.n23 9.154
R69 GND.n30 GND.n29 9.154
R70 GND.n29 GND.n28 9.154
R71 GND.n35 GND.n34 9.154
R72 GND.n34 GND.n33 9.154
R73 GND.n38 GND.n37 9.154
R74 GND.n37 GND.n36 9.154
R75 GND.n42 GND.n41 9.154
R76 GND.n41 GND.n40 9.154
R77 GND.n47 GND.n46 9.154
R78 GND.n46 GND.n45 9.154
R79 GND.n51 GND.n50 9.154
R80 GND.n109 GND.n108 9.154
R81 GND.n112 GND.n111 9.154
R82 GND.n118 GND.n117 9.154
R83 GND.n117 GND.n116 9.154
R84 GND.n122 GND.n121 9.154
R85 GND.n121 GND.n120 9.154
R86 GND.n126 GND.n125 9.154
R87 GND.n125 GND.n124 9.154
R88 GND.n131 GND.n130 9.154
R89 GND.n130 GND.n129 9.154
R90 GND.n136 GND.n135 9.154
R91 GND.n135 GND.n134 9.154
R92 GND.n140 GND.n139 9.154
R93 GND.n139 GND.n138 9.154
R94 GND.n144 GND.n143 9.154
R95 GND.n143 GND.n142 9.154
R96 GND.n148 GND.n147 9.154
R97 GND.n147 GND.n146 9.154
R98 GND.n152 GND.n151 9.154
R99 GND.n151 GND.n150 9.154
R100 GND.n171 GND.n170 9.154
R101 GND.n170 GND.n169 9.154
R102 GND.n167 GND.n166 9.154
R103 GND.n166 GND.n165 9.154
R104 GND.n163 GND.n162 9.154
R105 GND.n162 GND.n161 9.154
R106 GND.n158 GND.n157 9.154
R107 GND.n2 GND.n1 8.108
R108 GND.n108 GND.n107 8.108
R109 GND.n44 GND.n0 6.21
R110 GND.n155 GND.n154 4.706
R111 GND.n103 GND.n102 4.65
R112 GND.n61 GND.n60 4.65
R113 GND.n66 GND.n65 4.65
R114 GND.n71 GND.n70 4.65
R115 GND.n75 GND.n74 4.65
R116 GND.n79 GND.n78 4.65
R117 GND.n83 GND.n80 4.65
R118 GND.n87 GND.n86 4.65
R119 GND.n91 GND.n90 4.65
R120 GND.n95 GND.n94 4.65
R121 GND.n100 GND.n99 4.65
R122 GND.n57 GND.n56 4.65
R123 GND.n55 GND.n54 4.65
R124 GND.n8 GND.n7 4.65
R125 GND.n13 GND.n12 4.65
R126 GND.n17 GND.n16 4.65
R127 GND.n22 GND.n21 4.65
R128 GND.n26 GND.n25 4.65
R129 GND.n31 GND.n30 4.65
R130 GND.n35 GND.n32 4.65
R131 GND.n39 GND.n38 4.65
R132 GND.n43 GND.n42 4.65
R133 GND.n48 GND.n47 4.65
R134 GND.n52 GND.n51 4.65
R135 GND.n110 GND.n109 4.65
R136 GND.n113 GND.n112 4.65
R137 GND.n119 GND.n118 4.65
R138 GND.n123 GND.n122 4.65
R139 GND.n127 GND.n126 4.65
R140 GND.n132 GND.n131 4.65
R141 GND.n137 GND.n136 4.65
R142 GND.n141 GND.n140 4.65
R143 GND.n145 GND.n144 4.65
R144 GND.n149 GND.n148 4.65
R145 GND.n153 GND.n152 4.65
R146 GND.n172 GND.n171 4.65
R147 GND.n168 GND.n167 4.65
R148 GND.n164 GND.n163 4.65
R149 GND.n159 GND.n158 4.65
R150 GND.n105 GND.n104 4.65
R151 GND.n50 GND.n49 2.759
R152 GND.n4 GND.n3 2.562
R153 GND.n8 GND.n4 1.145
R154 GND.n57 GND.n55 0.525
R155 GND.n107 GND.n106 0.524
R156 GND.n105 GND.n103 0.507
R157 GND.n17 GND.n13 0.09
R158 GND.n26 GND.n22 0.09
R159 GND.n32 GND.n31 0.09
R160 GND.n43 GND.n39 0.09
R161 GND.n52 GND.n48 0.09
R162 GND.n61 GND.n57 0.09
R163 GND.n75 GND.n71 0.09
R164 GND.n79 GND.n75 0.09
R165 GND.n80 GND.n79 0.09
R166 GND.n91 GND.n87 0.09
R167 GND.n95 GND.n91 0.09
R168 GND.n110 GND.n105 0.09
R169 GND.n113 GND.n110 0.09
R170 GND.n123 GND.n119 0.09
R171 GND.n127 GND.n123 0.09
R172 GND.n141 GND.n137 0.09
R173 GND.n145 GND.n141 0.09
R174 GND.n149 GND.n145 0.09
R175 GND.n153 GND.n149 0.09
R176 GND.n172 GND.n168 0.09
R177 GND.n168 GND.n164 0.09
R178 GND.n18 GND.n17 0.078
R179 GND.n31 GND.n27 0.078
R180 GND.n67 GND.n66 0.078
R181 GND.n98 GND.n97 0.074
R182 GND.n157 GND.n156 0.074
R183 GND.n9 GND.n8 0.072
R184 GND.n114 GND.n113 0.071
R185 GND.n128 GND.n127 0.071
R186 GND.n39 GND 0.065
R187 GND.n66 GND.n62 0.065
R188 GND.n87 CMOS_AND_1/GND 0.065
R189 GND.n137 GND.n133 0.065
R190 CMOS_3in_AND_0/GND GND.n172 0.065
R191 GND.n48 GND.n44 0.063
R192 GND.n55 GND.n53 0.056
R193 GND.n103 GND.n101 0.056
R194 GND.n96 GND.n95 0.055
R195 GND.n164 GND.n160 0.055
R196 GND.n59 GND.n58 0.047
R197 GND.n100 GND.n96 0.035
R198 GND.n160 GND.n159 0.035
R199 GND.n53 GND.n52 0.033
R200 GND.n101 GND.n100 0.033
R201 GND.n159 GND.n155 0.033
R202 GND.n44 GND.n43 0.026
R203 GND.n32 GND 0.025
R204 GND.n62 GND.n61 0.025
R205 GND.n80 CMOS_AND_1/GND 0.025
R206 GND.n133 GND.n132 0.025
R207 CMOS_3in_AND_0/GND GND.n153 0.025
R208 GND.n119 GND.n114 0.018
R209 GND.n132 GND.n128 0.018
R210 GND.n13 GND.n9 0.017
R211 GND.n22 GND.n18 0.011
R212 GND.n27 GND.n26 0.011
R213 GND.n71 GND.n67 0.011
R214 s3.n2 s3.t0 120.552
R215 s3.n1 s3.t1 98.438
R216 s3 s3.n2 7.84
R217 s3 s3.n1 3.68
R218 s3.n1 s3.n0 3.084
R219 s3.n0 s3 0.374
R220 VDD.n72 VDD.t7 38.206
R221 VDD.n135 VDD.t37 36.141
R222 VDD.n302 VDD.t18 32.01
R223 VDD.n80 VDD.t5 32.01
R224 VDD.n127 VDD.t4 29.945
R225 VDD.n60 VDD.t17 29.945
R226 VDD.n34 VDD.t32 24.782
R227 VDD.n181 VDD.t22 24.782
R228 VDD.n228 VDD.t2 24.782
R229 VDD.n284 VDD.t0 24.782
R230 VDD.n119 VDD.t10 23.75
R231 VDD.n52 VDD.t8 23.75
R232 VDD.n301 VDD.t19 22.029
R233 VDD.n118 VDD.t11 22.029
R234 VDD.n101 VDD.t27 22.029
R235 VDD.n84 VDD.t6 22.029
R236 VDD.n51 VDD.t9 22.029
R237 VDD.n42 VDD.t33 22.029
R238 VDD.n21 VDD.t29 22.029
R239 VDD.n8 VDD.t31 22.029
R240 VDD.n148 VDD.t25 22.029
R241 VDD.n189 VDD.t23 22.029
R242 VDD.n202 VDD.t39 22.029
R243 VDD.n215 VDD.t36 22.029
R244 VDD.n236 VDD.t3 22.029
R245 VDD.n249 VDD.t21 22.029
R246 VDD.n266 VDD.t13 22.029
R247 VDD.n139 VDD.t16 19.7
R248 VDD.n139 VDD.t1 19.7
R249 VDD.n97 VDD.t26 18.586
R250 VDD.n26 VDD.t28 18.586
R251 VDD.n144 VDD.t24 18.586
R252 VDD.n173 VDD.t34 18.586
R253 VDD.n220 VDD.t35 18.586
R254 VDD.n245 VDD.t20 18.586
R255 VDD.n275 VDD.t15 18.586
R256 VDD.n4 VDD.t30 12.391
R257 VDD.n165 VDD.t14 12.391
R258 VDD.n198 VDD.t38 12.391
R259 VDD.n267 VDD.t12 12.391
R260 VDD.n74 VDD.n71 11.52
R261 VDD.n28 VDD.n25 11.52
R262 VDD.n175 VDD.n172 11.52
R263 VDD.n222 VDD.n219 11.52
R264 VDD.n277 VDD.n274 11.52
R265 VDD.n142 VDD.n141 8.855
R266 VDD.n196 VDD.n195 8.855
R267 VDD.n243 VDD.n242 8.855
R268 VDD.n247 VDD.n246 8.855
R269 VDD.n246 VDD.n245 8.855
R270 VDD.n252 VDD.n251 8.855
R271 VDD.n251 VDD.n250 8.855
R272 VDD.n256 VDD.n255 8.855
R273 VDD.n255 VDD.n254 8.855
R274 VDD.n260 VDD.n259 8.855
R275 VDD.n259 VDD.n258 8.855
R276 VDD.n264 VDD.n263 8.855
R277 VDD.n263 VDD.n262 8.855
R278 VDD.n269 VDD.n268 8.855
R279 VDD.n268 VDD.n267 8.855
R280 VDD.n274 VDD.n273 8.855
R281 VDD.n273 VDD.n272 8.855
R282 VDD.n277 VDD.n276 8.855
R283 VDD.n276 VDD.n275 8.855
R284 VDD.n281 VDD.n280 8.855
R285 VDD.n280 VDD.n279 8.855
R286 VDD.n286 VDD.n285 8.855
R287 VDD.n285 VDD.n284 8.855
R288 VDD.n290 VDD.n289 8.855
R289 VDD.n200 VDD.n199 8.855
R290 VDD.n199 VDD.n198 8.855
R291 VDD.n205 VDD.n204 8.855
R292 VDD.n204 VDD.n203 8.855
R293 VDD.n209 VDD.n208 8.855
R294 VDD.n208 VDD.n207 8.855
R295 VDD.n213 VDD.n212 8.855
R296 VDD.n212 VDD.n211 8.855
R297 VDD.n219 VDD.n218 8.855
R298 VDD.n218 VDD.n217 8.855
R299 VDD.n222 VDD.n221 8.855
R300 VDD.n221 VDD.n220 8.855
R301 VDD.n226 VDD.n225 8.855
R302 VDD.n225 VDD.n224 8.855
R303 VDD.n230 VDD.n229 8.855
R304 VDD.n229 VDD.n228 8.855
R305 VDD.n234 VDD.n233 8.855
R306 VDD.n146 VDD.n145 8.855
R307 VDD.n145 VDD.n144 8.855
R308 VDD.n151 VDD.n150 8.855
R309 VDD.n150 VDD.n149 8.855
R310 VDD.n155 VDD.n154 8.855
R311 VDD.n154 VDD.n153 8.855
R312 VDD.n159 VDD.n158 8.855
R313 VDD.n158 VDD.n157 8.855
R314 VDD.n163 VDD.n162 8.855
R315 VDD.n162 VDD.n161 8.855
R316 VDD.n167 VDD.n166 8.855
R317 VDD.n166 VDD.n165 8.855
R318 VDD.n172 VDD.n171 8.855
R319 VDD.n171 VDD.n170 8.855
R320 VDD.n175 VDD.n174 8.855
R321 VDD.n174 VDD.n173 8.855
R322 VDD.n179 VDD.n178 8.855
R323 VDD.n178 VDD.n177 8.855
R324 VDD.n183 VDD.n182 8.855
R325 VDD.n182 VDD.n181 8.855
R326 VDD.n187 VDD.n186 8.855
R327 VDD.n2 VDD.n1 8.855
R328 VDD.n6 VDD.n5 8.855
R329 VDD.n5 VDD.n4 8.855
R330 VDD.n11 VDD.n10 8.855
R331 VDD.n10 VDD.n9 8.855
R332 VDD.n15 VDD.n14 8.855
R333 VDD.n14 VDD.n13 8.855
R334 VDD.n19 VDD.n18 8.855
R335 VDD.n18 VDD.n17 8.855
R336 VDD.n25 VDD.n24 8.855
R337 VDD.n24 VDD.n23 8.855
R338 VDD.n28 VDD.n27 8.855
R339 VDD.n27 VDD.n26 8.855
R340 VDD.n32 VDD.n31 8.855
R341 VDD.n31 VDD.n30 8.855
R342 VDD.n36 VDD.n35 8.855
R343 VDD.n35 VDD.n34 8.855
R344 VDD.n40 VDD.n39 8.855
R345 VDD.n49 VDD.n48 8.855
R346 VDD.n54 VDD.n53 8.855
R347 VDD.n53 VDD.n52 8.855
R348 VDD.n58 VDD.n57 8.855
R349 VDD.n57 VDD.n56 8.855
R350 VDD.n62 VDD.n61 8.855
R351 VDD.n61 VDD.n60 8.855
R352 VDD.n66 VDD.n65 8.855
R353 VDD.n65 VDD.n64 8.855
R354 VDD.n71 VDD.n70 8.855
R355 VDD.n70 VDD.n69 8.855
R356 VDD.n74 VDD.n73 8.855
R357 VDD.n73 VDD.n72 8.855
R358 VDD.n78 VDD.n77 8.855
R359 VDD.n77 VDD.n76 8.855
R360 VDD.n82 VDD.n81 8.855
R361 VDD.n81 VDD.n80 8.855
R362 VDD.n87 VDD.n86 8.855
R363 VDD.n95 VDD.n94 8.855
R364 VDD.n99 VDD.n98 8.855
R365 VDD.n98 VDD.n97 8.855
R366 VDD.n104 VDD.n103 8.855
R367 VDD.n103 VDD.n102 8.855
R368 VDD.n108 VDD.n107 8.855
R369 VDD.n107 VDD.n106 8.855
R370 VDD.n112 VDD.n111 8.855
R371 VDD.n111 VDD.n110 8.855
R372 VDD.n116 VDD.n115 8.855
R373 VDD.n115 VDD.n114 8.855
R374 VDD.n121 VDD.n120 8.855
R375 VDD.n120 VDD.n119 8.855
R376 VDD.n125 VDD.n124 8.855
R377 VDD.n124 VDD.n123 8.855
R378 VDD.n129 VDD.n128 8.855
R379 VDD.n128 VDD.n127 8.855
R380 VDD.n133 VDD.n132 8.855
R381 VDD.n132 VDD.n131 8.855
R382 VDD.n137 VDD.n136 8.855
R383 VDD.n136 VDD.n135 8.855
R384 VDD.n312 VDD.n311 8.855
R385 VDD.n311 VDD.n310 8.855
R386 VDD.n308 VDD.n307 8.855
R387 VDD.n307 VDD.n306 8.855
R388 VDD.n304 VDD.n303 8.855
R389 VDD.n303 VDD.n302 8.855
R390 VDD.n299 VDD.n298 8.855
R391 VDD.n294 VDD.n293 4.91
R392 VDD.n293 VDD.n292 4.65
R393 VDD.n244 VDD.n243 4.65
R394 VDD.n248 VDD.n247 4.65
R395 VDD.n253 VDD.n252 4.65
R396 VDD.n257 VDD.n256 4.65
R397 VDD.n261 VDD.n260 4.65
R398 VDD.n265 VDD.n264 4.65
R399 VDD.n270 VDD.n269 4.65
R400 VDD.n274 VDD.n271 4.65
R401 VDD.n278 VDD.n277 4.65
R402 VDD.n282 VDD.n281 4.65
R403 VDD.n287 VDD.n286 4.65
R404 VDD.n291 VDD.n290 4.65
R405 VDD.n240 VDD.n239 4.65
R406 VDD.n238 VDD.n237 4.65
R407 VDD.n197 VDD.n196 4.65
R408 VDD.n201 VDD.n200 4.65
R409 VDD.n206 VDD.n205 4.65
R410 VDD.n210 VDD.n209 4.65
R411 VDD.n214 VDD.n213 4.65
R412 VDD.n219 VDD.n216 4.65
R413 VDD.n223 VDD.n222 4.65
R414 VDD.n227 VDD.n226 4.65
R415 VDD.n231 VDD.n230 4.65
R416 VDD.n235 VDD.n234 4.65
R417 VDD.n193 VDD.n192 4.65
R418 VDD.n191 VDD.n190 4.65
R419 VDD.n147 VDD.n146 4.65
R420 VDD.n152 VDD.n151 4.65
R421 VDD.n156 VDD.n155 4.65
R422 VDD.n160 VDD.n159 4.65
R423 VDD.n164 VDD.n163 4.65
R424 VDD.n168 VDD.n167 4.65
R425 VDD.n172 VDD.n169 4.65
R426 VDD.n176 VDD.n175 4.65
R427 VDD.n180 VDD.n179 4.65
R428 VDD.n184 VDD.n183 4.65
R429 VDD.n188 VDD.n187 4.65
R430 VDD.n7 VDD.n6 4.65
R431 VDD.n12 VDD.n11 4.65
R432 VDD.n16 VDD.n15 4.65
R433 VDD.n20 VDD.n19 4.65
R434 VDD.n25 VDD.n22 4.65
R435 VDD.n29 VDD.n28 4.65
R436 VDD.n33 VDD.n32 4.65
R437 VDD.n37 VDD.n36 4.65
R438 VDD.n41 VDD.n40 4.65
R439 VDD.n44 VDD.n43 4.65
R440 VDD.n46 VDD.n45 4.65
R441 VDD.n50 VDD.n49 4.65
R442 VDD.n55 VDD.n54 4.65
R443 VDD.n59 VDD.n58 4.65
R444 VDD.n63 VDD.n62 4.65
R445 VDD.n67 VDD.n66 4.65
R446 VDD.n71 VDD.n68 4.65
R447 VDD.n75 VDD.n74 4.65
R448 VDD.n79 VDD.n78 4.65
R449 VDD.n83 VDD.n82 4.65
R450 VDD.n88 VDD.n87 4.65
R451 VDD.n90 VDD.n89 4.65
R452 VDD.n92 VDD.n91 4.65
R453 VDD.n96 VDD.n95 4.65
R454 VDD.n100 VDD.n99 4.65
R455 VDD.n105 VDD.n104 4.65
R456 VDD.n109 VDD.n108 4.65
R457 VDD.n113 VDD.n112 4.65
R458 VDD.n117 VDD.n116 4.65
R459 VDD.n122 VDD.n121 4.65
R460 VDD.n126 VDD.n125 4.65
R461 VDD.n130 VDD.n129 4.65
R462 VDD.n134 VDD.n133 4.65
R463 VDD.n138 VDD.n137 4.65
R464 VDD.n313 VDD.n312 4.65
R465 VDD.n309 VDD.n308 4.65
R466 VDD.n305 VDD.n304 4.65
R467 VDD.n300 VDD.n299 4.65
R468 VDD.n296 VDD.n295 4.65
R469 VDD.n1 VDD.n0 4.288
R470 VDD.n48 VDD.n47 4.288
R471 VDD.n94 VDD.n93 4.288
R472 VDD.n141 VDD.n140 4.288
R473 VDD.n195 VDD.n194 4.288
R474 VDD.n242 VDD.n241 4.288
R475 VDD.n289 VDD.n288 4.288
R476 VDD.n233 VDD.n232 4.288
R477 VDD.n186 VDD.n185 4.288
R478 VDD.n39 VDD.n38 4.288
R479 VDD.n86 VDD.n85 4.288
R480 VDD.n298 VDD.n297 4.288
R481 VDD.n3 VDD.n2 2.562
R482 VDD.n143 VDD.n142 2.562
R483 VDD.n283 VDD.n139 2.329
R484 VDD.n7 VDD.n3 1.145
R485 VDD.n147 VDD.n143 1.145
R486 VDD.n240 VDD.n238 0.777
R487 VDD.n193 VDD.n191 0.525
R488 VDD.n46 VDD.n44 0.525
R489 VDD.n92 VDD.n90 0.507
R490 VDD.n296 VDD.n294 0.135
R491 VDD.n156 VDD.n152 0.09
R492 VDD.n160 VDD.n156 0.09
R493 VDD.n164 VDD.n160 0.09
R494 VDD.n168 VDD.n164 0.09
R495 VDD.n169 VDD.n168 0.09
R496 VDD.n180 VDD.n176 0.09
R497 VDD.n184 VDD.n180 0.09
R498 VDD.n188 VDD.n184 0.09
R499 VDD.n197 VDD.n193 0.09
R500 VDD.n201 VDD.n197 0.09
R501 VDD.n210 VDD.n206 0.09
R502 VDD.n214 VDD.n210 0.09
R503 VDD.n216 VDD.n214 0.09
R504 VDD.n227 VDD.n223 0.09
R505 VDD.n231 VDD.n227 0.09
R506 VDD.n235 VDD.n231 0.09
R507 VDD.n244 VDD.n240 0.09
R508 VDD.n248 VDD.n244 0.09
R509 VDD.n257 VDD.n253 0.09
R510 VDD.n261 VDD.n257 0.09
R511 VDD.n265 VDD.n261 0.09
R512 VDD.n271 VDD.n270 0.09
R513 VDD.n282 VDD.n278 0.09
R514 VDD.n291 VDD.n287 0.09
R515 VDD.n293 VDD.n291 0.09
R516 VDD.n16 VDD.n12 0.09
R517 VDD.n20 VDD.n16 0.09
R518 VDD.n22 VDD.n20 0.09
R519 VDD.n33 VDD.n29 0.09
R520 VDD.n37 VDD.n33 0.09
R521 VDD.n41 VDD.n37 0.09
R522 VDD.n50 VDD.n46 0.09
R523 VDD.n59 VDD.n55 0.09
R524 VDD.n63 VDD.n59 0.09
R525 VDD.n67 VDD.n63 0.09
R526 VDD.n68 VDD.n67 0.09
R527 VDD.n79 VDD.n75 0.09
R528 VDD.n83 VDD.n79 0.09
R529 VDD.n90 VDD.n88 0.09
R530 VDD.n96 VDD.n92 0.09
R531 VDD.n100 VDD.n96 0.09
R532 VDD.n109 VDD.n105 0.09
R533 VDD.n113 VDD.n109 0.09
R534 VDD.n117 VDD.n113 0.09
R535 VDD.n126 VDD.n122 0.09
R536 VDD.n130 VDD.n126 0.09
R537 VDD.n134 VDD.n130 0.09
R538 VDD.n138 VDD.n134 0.09
R539 VDD.n313 VDD.n309 0.09
R540 VDD.n309 VDD.n305 0.09
R541 VDD.n300 VDD.n296 0.09
R542 VDD.n202 VDD.n201 0.078
R543 VDD.n270 VDD.n266 0.078
R544 VDD.n8 VDD.n7 0.078
R545 VDD.n249 VDD.n248 0.071
R546 VDD.n101 VDD.n100 0.071
R547 VDD.n148 VDD.n147 0.07
R548 VDD.n176 CMOS_3in_OR_0/VDD 0.065
R549 VDD.n223 CMOS_AND_1/VDD 0.065
R550 VDD.n278 CMOS_3in_AND_0/VDD 0.065
R551 VDD.n29 VDD 0.065
R552 VDD.n55 VDD.n51 0.065
R553 VDD.n75 CMOS_XOR_0/VDD 0.065
R554 VDD.n122 VDD.n118 0.065
R555 CMOS_XNOR_0/VDD VDD.n313 0.065
R556 VDD.n287 VDD.n283 0.063
R557 VDD.n191 VDD.n189 0.056
R558 VDD.n238 VDD.n236 0.056
R559 VDD.n44 VDD.n42 0.056
R560 VDD.n84 VDD.n83 0.055
R561 VDD.n305 VDD.n301 0.055
R562 VDD.n88 VDD.n84 0.035
R563 VDD.n301 VDD.n300 0.035
R564 VDD.n189 VDD.n188 0.033
R565 VDD.n236 VDD.n235 0.033
R566 VDD.n42 VDD.n41 0.033
R567 VDD.n294 VDD 0.027
R568 VDD.n283 VDD.n282 0.026
R569 VDD.n169 CMOS_3in_OR_0/VDD 0.025
R570 VDD.n271 CMOS_3in_AND_0/VDD 0.025
R571 VDD.n51 VDD.n50 0.025
R572 VDD.n68 CMOS_XOR_0/VDD 0.025
R573 VDD.n118 VDD.n117 0.025
R574 CMOS_XNOR_0/VDD VDD.n138 0.025
R575 VDD.n152 VDD.n148 0.02
R576 VDD.n253 VDD.n249 0.018
R577 VDD.n105 VDD.n101 0.018
R578 VDD.n216 VDD.n215 0.017
R579 VDD.n22 VDD.n21 0.017
R580 VDD.n206 VDD.n202 0.011
R581 VDD.n266 VDD.n265 0.011
R582 VDD.n12 VDD.n8 0.011
R583 VDD.n215 CMOS_AND_1/VDD 0.007
R584 VDD.n21 VDD 0.007
R585 x3.t0 x3.t2 924.95
R586 CMOS_XOR_0/B x3.t0 633.02
R587 x3.n0 x3.t3 570.366
R588 x3.n0 x3.t1 570.366
R589 x3.n1 x3 158.792
R590 x3 x3.n0 78.72
R591 CMOS_XOR_0/B x3.n1 42.894
R592 x3.n1 x3 0.157
R593 x1.n1 x1.t1 993.097
R594 x1.n0 x1.t0 579.86
R595 x1.n0 x1.t3 547.727
R596 x1.n1 x1.t2 356.59
R597 x1.n2 CMOS_XNOR_0/A 318.92
R598 CMOS_XNOR_0/A x1.n1 78.72
R599 x1.n3 x1.n2 20.984
R600 x1.n3 x1.n0 8.764
R601 x1 x1.n3 2.72
R602 x1.n2 x1 1.597
R603 x3_bar.n3 x3_bar.t2 616.084
R604 x3_bar.n0 x3_bar.t1 579.86
R605 x3_bar.n0 x3_bar.t0 547.727
R606 x3_bar.n3 x3_bar.t3 528.72
R607 x3_bar.n3 x3_bar.n2 12.411
R608 x3_bar.n2 x3_bar.n1 11.74
R609 x3_bar.n1 x3_bar.n0 8.764
R610 CMOS_XOR_0/B_bar x3_bar.n3 3.68
R611 x3_bar.n1 x3_bar 2.72
R612 x3_bar.n2 x3_bar 2.167
R613 x0.t2 x0.t3 1221.07
R614 x0.t0 x0.t1 924.95
R615 CMOS_XNOR_0/B x0.t0 633.02
R616 CMOS_XNOR_0/B x0.n0 535.88
R617 x0.n0 x0 428.025
R618 x0 x0.t2 392.02
R619 x0.n0 x0 0.152
R620 x1_bar.t0 x1_bar.t1 1345.61
R621 x1_bar x1_bar.t0 392.02
R622 x2_bar.t3 x2_bar.t2 1345.61
R623 x2_bar.t0 x2_bar.t1 1221.07
R624 x2_bar.n0 x2_bar.t0 630.3
R625 CMOS_XOR_0/A_bar x2_bar.t3 392.02
R626 CMOS_XOR_0/A_bar x2_bar.n1 44.231
R627 x2_bar.n1 x2_bar.n0 41.121
R628 x2_bar.n1 x2_bar 2.762
R629 x2_bar.n0 x2_bar 2.72
R630 CMOS_3in_OR_0/C.t3 CMOS_3in_OR_0/C.t2 1221.07
R631 CMOS_3in_OR_0/C CMOS_3in_OR_0/C.n0 787.238
R632 CMOS_3in_OR_0/C CMOS_3in_OR_0/C.t3 633.02
R633 CMOS_3in_AND_0/OUT CMOS_3in_OR_0/C.t1 117.958
R634 CMOS_3in_OR_0/C.n0 CMOS_3in_AND_0/OUT 91.717
R635 CMOS_3in_OR_0/C.n0 CMOS_3in_OR_0/C.t0 45.156
R636 x2.n0 x2.t1 993.097
R637 x2.n0 x2.t0 356.59
R638 x2.n1 x2 16.254
R639 x2.n1 x2.n0 8.764
R640 x2 x2.n1 2.72
R641 x0_bar.n0 x0_bar.t0 683.32
R642 x0_bar.n0 x0_bar.t1 528.72
R643 x0_bar x0_bar.n0 3.68
C0 CMOS_AND_0/A a_1380_n1689# 0.01fF
C1 x2 CMOS_AND_1/A 0.07fF
C2 CMOS_AND_0/AND CMOS_3in_OR_0/C 0.06fF
C3 x0 x1 0.21fF
C4 a_1380_n1689# x3 0.02fF
C5 x1 a_1735_499# 0.00fF
C6 a_n28_n779# a_27_n111# 0.00fF
C7 x2_bar x2 4.74fF
C8 x3_bar CMOS_AND_0/AND 0.00fF
C9 a_n328_n1689# a_27_n111# 0.01fF
C10 x1_bar a_n178_n779# 0.00fF
C11 x0 a_177_499# 0.02fF
C12 VDD a_27_n111# 1.04fF
C13 a_2442_n779# CMOS_AND_0/A 0.01fF
C14 CMOS_AND_0/AND s3 0.04fF
C15 x1_bar CMOS_AND_0/A 0.00fF
C16 x1 a_177_499# 0.00fF
C17 a_1380_n1689# CMOS_3in_OR_0/C 0.10fF
C18 x1_bar x3 0.04fF
C19 a_1735_n111# x1 0.01fF
C20 a_27_n111# CMOS_AND_1/A 0.08fF
C21 a_1435_n111# x1 0.01fF
C22 CMOS_AND_0/A CMOS_AND_1/AND 0.02fF
C23 a_n328_n1689# a_n178_n779# 0.01fF
C24 a_2442_n779# a_2592_499# 0.01fF
C25 x3 CMOS_AND_1/AND 0.00fF
C26 VDD a_n178_n779# 0.01fF
C27 a_1380_n1689# x3_bar 0.05fF
C28 x2_bar a_27_n111# 0.05fF
C29 a_n28_n779# x3 0.00fF
C30 a_1380_n779# x1 0.01fF
C31 VDD a_1435_499# 0.06fF
C32 x1_bar a_n123_499# 0.01fF
C33 VDD CMOS_AND_0/A 1.03fF
C34 a_2442_n779# CMOS_3in_OR_0/C 0.05fF
C35 a_n328_n1689# x3 0.09fF
C36 a_2592_n111# CMOS_AND_0/A 0.01fF
C37 a_1380_n1689# s3 0.00fF
C38 VDD x3 1.54fF
C39 x1_bar x0_bar 0.13fF
C40 x1_bar CMOS_3in_OR_0/C 0.00fF
C41 a_1735_499# CMOS_AND_0/AND 0.00fF
C42 CMOS_AND_1/A a_1435_499# 0.01fF
C43 CMOS_AND_0/A CMOS_AND_1/A 0.05fF
C44 x1 CMOS_AND_0/AND 0.06fF
C45 a_2442_n779# x3_bar 0.00fF
C46 a_2592_n1689# CMOS_AND_0/AND 0.00fF
C47 a_n123_n111# x1_bar 0.01fF
C48 CMOS_3in_OR_0/C CMOS_AND_1/AND 0.10fF
C49 x3 CMOS_AND_1/A 0.03fF
C50 x2_bar a_n178_n779# 0.01fF
C51 VDD a_2592_499# 0.78fF
C52 x1_bar x3_bar 0.09fF
C53 a_2592_n111# a_2592_499# 0.01fF
C54 a_n28_n779# x0_bar 0.00fF
C55 a_n28_n779# CMOS_3in_OR_0/C 0.00fF
C56 x2_bar a_1435_499# 0.00fF
C57 VDD a_n123_499# 0.05fF
C58 a_2442_n779# s3 0.06fF
C59 a_n328_n1689# CMOS_3in_OR_0/C 0.05fF
C60 a_n328_n1689# x0_bar 0.01fF
C61 x2_bar CMOS_AND_0/A 0.14fF
C62 x2 a_27_n111# 0.05fF
C63 VDD x0_bar 0.24fF
C64 VDD CMOS_3in_OR_0/C 2.11fF
C65 x2_bar x3 2.37fF
C66 x3_bar CMOS_AND_1/AND 0.01fF
C67 x0 a_1380_n1689# 0.00fF
C68 a_n28_n779# x3_bar 0.00fF
C69 a_1735_n111# CMOS_AND_0/AND 0.00fF
C70 a_1435_n111# CMOS_AND_0/AND 0.00fF
C71 a_n123_n111# a_n328_n1689# 0.00fF
C72 a_1380_n1689# a_1735_499# 0.00fF
C73 a_177_n111# x1_bar 0.01fF
C74 a_n123_499# CMOS_AND_1/A 0.00fF
C75 a_n123_n111# VDD 0.01fF
C76 a_n328_n1689# x3_bar 0.11fF
C77 s3 CMOS_AND_1/AND 0.01fF
C78 x0_bar CMOS_AND_1/A 0.00fF
C79 x1 a_1380_n1689# 0.03fF
C80 CMOS_3in_OR_0/C CMOS_AND_1/A 0.02fF
C81 a_1380_n1689# a_2592_n1689# 0.00fF
C82 VDD x3_bar 1.07fF
C83 x2_bar a_2592_499# 0.00fF
C84 a_2592_n111# x3_bar 0.00fF
C85 x2_bar a_n123_499# 0.00fF
C86 x2 a_n178_n779# 0.00fF
C87 a_n123_n111# CMOS_AND_1/A 0.00fF
C88 VDD s3 0.37fF
C89 x2_bar x0_bar 0.04fF
C90 x2_bar CMOS_3in_OR_0/C 0.03fF
C91 x3_bar CMOS_AND_1/A 0.12fF
C92 a_177_n111# a_n328_n1689# 0.00fF
C93 x2 CMOS_AND_0/A 0.09fF
C94 x0 x1_bar 0.20fF
C95 a_177_n111# VDD 0.01fF
C96 x2 x3 0.20fF
C97 a_1735_n111# a_1380_n1689# 0.00fF
C98 a_1435_n111# a_1380_n1689# 0.00fF
C99 a_2442_n779# x1 0.04fF
C100 x2_bar a_n123_n111# 0.00fF
C101 a_2442_n779# a_2592_n1689# 0.02fF
C102 x2_bar x3_bar 0.27fF
C103 x1_bar x1 2.81fF
C104 a_177_n111# CMOS_AND_1/A 0.00fF
C105 a_n28_n779# x0 0.00fF
C106 a_1380_n779# a_1380_n1689# 0.01fF
C107 x2 a_2592_499# 0.00fF
C108 x2_bar s3 0.00fF
C109 x1 CMOS_AND_1/AND 0.03fF
C110 a_2592_n1689# CMOS_AND_1/AND 0.01fF
C111 x0 a_n328_n1689# 0.04fF
C112 x2 a_n123_499# 0.00fF
C113 a_n28_n779# x1 0.01fF
C114 x1_bar a_177_499# 0.01fF
C115 x0 VDD 1.12fF
C116 x2_bar a_177_n111# 0.00fF
C117 a_2742_n1689# a_2592_499# 0.00fF
C118 x2 x0_bar 0.04fF
C119 x2 CMOS_3in_OR_0/C 0.03fF
C120 a_27_n111# a_1435_499# 0.00fF
C121 VDD a_1735_499# 0.06fF
C122 a_n328_n1689# x1 0.04fF
C123 CMOS_AND_0/A a_27_n111# 0.04fF
C124 x1 VDD 0.58fF
C125 a_2592_n111# x1 0.01fF
C126 VDD a_2592_n1689# 0.06fF
C127 a_1380_n1689# CMOS_AND_0/AND 0.00fF
C128 a_27_n111# x3 0.17fF
C129 a_2742_n1689# CMOS_3in_OR_0/C 0.01fF
C130 x0 CMOS_AND_1/A 0.01fF
C131 a_n123_n111# x2 0.00fF
C132 a_1380_n779# a_2442_n779# 0.00fF
C133 a_1735_499# CMOS_AND_1/A 0.00fF
C134 x2 x3_bar 0.60fF
C135 a_n328_n1689# a_177_499# 0.00fF
C136 x1 CMOS_AND_1/A 0.03fF
C137 VDD a_177_499# 0.05fF
C138 x2_bar x0 0.15fF
C139 x2_bar a_1735_499# 0.01fF
C140 a_1735_n111# VDD 0.01fF
C141 a_1380_n779# CMOS_AND_1/AND 0.00fF
C142 a_1435_n111# VDD 0.01fF
C143 a_n123_499# a_27_n111# 0.02fF
C144 a_2442_n779# CMOS_AND_0/AND 0.12fF
C145 CMOS_AND_0/A a_1435_499# 0.02fF
C146 x2_bar x1 0.86fF
C147 a_n178_n779# x3 0.00fF
C148 a_177_n111# x2 0.00fF
C149 x0_bar a_27_n111# 0.14fF
C150 a_27_n111# CMOS_3in_OR_0/C 0.01fF
C151 s3 a_2742_n1689# 0.00fF
C152 x3 a_1435_499# 0.01fF
C153 a_177_499# CMOS_AND_1/A 0.00fF
C154 a_1380_n779# a_n328_n1689# 0.00fF
C155 CMOS_AND_0/A x3 0.35fF
C156 a_1735_n111# CMOS_AND_1/A 0.00fF
C157 a_1380_n779# VDD 0.00fF
C158 a_1435_n111# CMOS_AND_1/A 0.00fF
C159 a_n123_n111# a_27_n111# 0.01fF
C160 CMOS_AND_0/AND CMOS_AND_1/AND 0.04fF
C161 x2_bar a_177_499# 0.00fF
C162 x3_bar a_27_n111# 0.25fF
C163 a_2592_499# a_1435_499# 0.00fF
C164 x2_bar a_1735_n111# 0.01fF
C165 x2_bar a_1435_n111# 0.00fF
C166 a_1380_n779# CMOS_AND_1/A 0.01fF
C167 CMOS_AND_0/A a_2592_499# 0.09fF
C168 x0_bar a_n178_n779# 0.00fF
C169 a_n178_n779# CMOS_3in_OR_0/C 0.00fF
C170 x2 x0 0.10fF
C171 x3 a_2592_499# 0.01fF
C172 a_2442_n779# a_1380_n1689# 0.01fF
C173 VDD CMOS_AND_0/AND 0.49fF
C174 a_2592_n111# CMOS_AND_0/AND 0.01fF
C175 a_n123_499# x3 0.01fF
C176 CMOS_AND_0/A x0_bar 0.00fF
C177 CMOS_AND_0/A CMOS_3in_OR_0/C 0.00fF
C178 x2 x1 0.12fF
C179 x2_bar a_1380_n779# 0.00fF
C180 a_177_n111# a_27_n111# 0.01fF
C181 x0_bar x3 0.05fF
C182 x3 CMOS_3in_OR_0/C 0.00fF
C183 x3_bar a_n178_n779# 0.00fF
C184 CMOS_AND_0/AND CMOS_AND_1/A 0.01fF
C185 a_1380_n1689# CMOS_AND_1/AND 0.07fF
C186 x3_bar a_1435_499# 0.01fF
C187 a_n28_n779# a_1380_n1689# 0.00fF
C188 CMOS_AND_0/A x3_bar 0.15fF
C189 a_n123_n111# x3 0.00fF
C190 x2 a_177_499# 0.00fF
C191 x3_bar x3 3.29fF
C192 CMOS_3in_OR_0/C a_2592_499# 0.00fF
C193 a_n328_n1689# a_1380_n1689# 0.00fF
C194 x2_bar CMOS_AND_0/AND 0.00fF
C195 x2 a_1735_n111# 0.00fF
C196 a_1435_n111# x2 0.00fF
C197 VDD a_1380_n1689# 0.75fF
C198 a_n123_499# x0_bar 0.01fF
C199 x0 a_27_n111# 0.33fF
C200 a_177_n111# CMOS_AND_0/A 0.00fF
C201 a_2442_n779# CMOS_AND_1/AND 0.10fF
C202 x3_bar a_2592_499# 0.00fF
C203 x1 a_27_n111# 0.05fF
C204 a_1380_n779# x2 0.00fF
C205 a_1380_n1689# CMOS_AND_1/A 0.05fF
C206 a_177_n111# x3 0.00fF
C207 a_n123_499# x3_bar 0.01fF
C208 a_n123_n111# x0_bar 0.00fF
C209 a_n28_n779# x1_bar 0.00fF
C210 x3_bar CMOS_3in_OR_0/C 0.05fF
C211 x3_bar x0_bar 0.06fF
C212 a_2442_n779# VDD 0.54fF
C213 a_2592_n111# a_2442_n779# 0.00fF
C214 a_n328_n1689# x1_bar 0.01fF
C215 x2_bar a_1380_n1689# 0.02fF
C216 x0 a_n178_n779# 0.01fF
C217 a_27_n111# a_177_499# 0.03fF
C218 x1_bar VDD 0.16fF
C219 x2 CMOS_AND_0/AND 0.00fF
C220 s3 CMOS_3in_OR_0/C 0.00fF
C221 a_n123_n111# x3_bar 0.01fF
C222 a_1435_n111# a_27_n111# 0.00fF
C223 x0 CMOS_AND_0/A 0.00fF
C224 x1 a_n178_n779# 0.01fF
C225 a_n328_n1689# CMOS_AND_1/AND 0.00fF
C226 a_2442_n779# CMOS_AND_1/A 0.00fF
C227 CMOS_AND_0/A a_1735_499# 0.03fF
C228 x1 a_1435_499# 0.00fF
C229 x0 x3 0.20fF
C230 a_177_n111# x0_bar 0.00fF
C231 VDD CMOS_AND_1/AND 0.52fF
C232 a_n28_n779# a_n328_n1689# 0.01fF
C233 x1_bar CMOS_AND_1/A 0.01fF
C234 CMOS_AND_0/AND a_2742_n1689# 0.00fF
C235 a_1735_499# x3 0.03fF
C236 x1 CMOS_AND_0/A 0.23fF
C237 a_n28_n779# VDD 0.01fF
C238 CMOS_AND_0/A a_2592_n1689# 0.00fF
C239 x1 x3 0.13fF
C240 a_n328_n1689# VDD 1.40fF
C241 x2_bar a_2442_n779# 0.00fF
C242 a_2592_n111# VDD 0.01fF
C243 CMOS_AND_1/AND CMOS_AND_1/A 0.00fF
C244 x2_bar x1_bar 0.05fF
C245 a_177_n111# x3_bar 0.01fF
C246 a_1735_499# a_2592_499# 0.00fF
C247 x0 a_n123_499# 0.02fF
C248 CMOS_AND_0/A a_177_499# 0.00fF
C249 x2 a_1380_n1689# 0.00fF
C250 x1 a_2592_499# 0.05fF
C251 a_n328_n1689# CMOS_AND_1/A 0.00fF
C252 x3 a_177_499# 0.01fF
C253 a_2592_n1689# a_2592_499# 0.00fF
C254 x0 CMOS_3in_OR_0/C 0.00fF
C255 x0 x0_bar 3.15fF
C256 a_1735_n111# CMOS_AND_0/A 0.01fF
C257 x2_bar CMOS_AND_1/AND 0.00fF
C258 a_1435_n111# CMOS_AND_0/A 0.01fF
C259 VDD CMOS_AND_1/A 0.51fF
C260 x1 a_n123_499# 0.00fF
C261 a_1735_n111# x3 0.01fF
C262 a_1435_n111# x3 0.01fF
C263 x2_bar a_n28_n779# 0.01fF
C264 a_1380_n1689# a_2742_n1689# 0.00fF
C265 x1 x0_bar 3.36fF
C266 x1 CMOS_3in_OR_0/C 0.03fF
C267 a_2592_n1689# CMOS_3in_OR_0/C 0.01fF
C268 x2_bar a_n328_n1689# 0.15fF
C269 a_n123_n111# x0 0.01fF
C270 x2_bar VDD 1.22fF
C271 x0 x3_bar 0.12fF
C272 x3_bar a_1735_499# 0.00fF
C273 a_1735_n111# a_2592_499# 0.00fF
C274 a_n123_n111# x1 0.01fF
C275 a_1435_n111# a_2592_499# 0.00fF
C276 x1 x3_bar 0.45fF
C277 x2 x1_bar 2.70fF
C278 x0_bar a_177_499# 0.00fF
C279 x2_bar CMOS_AND_1/A 0.04fF
C280 CMOS_AND_0/AND a_1435_499# 0.00fF
C281 a_2442_n779# a_2742_n1689# 0.02fF
C282 a_177_n111# x0 0.01fF
C283 CMOS_AND_0/A CMOS_AND_0/AND 0.04fF
C284 x1 s3 0.00fF
C285 a_2592_n1689# s3 0.00fF
C286 CMOS_AND_0/AND x3 0.00fF
C287 x3_bar a_177_499# 0.01fF
C288 a_n28_n779# x2 0.00fF
C289 a_177_n111# x1 0.00fF
C290 a_1380_n779# CMOS_3in_OR_0/C 0.01fF
C291 a_1735_n111# x3_bar 0.00fF
C292 x2 a_n328_n1689# 0.02fF
C293 a_2742_n1689# CMOS_AND_1/AND 0.00fF
C294 a_1435_n111# x3_bar 0.01fF
C295 x2 VDD 0.19fF
C296 x2 a_2592_n111# 0.00fF
C297 CMOS_AND_0/AND a_2592_499# 0.08fF
C298 a_1380_n1689# a_1435_499# 0.00fF
C299 x1_bar a_27_n111# 0.12fF
C300 VDD a_2742_n1689# 0.06fF
C301 a_1380_n779# x3_bar 0.00fF
C302 a_2742_n1689# GND 0.02fF
C303 a_2592_n1689# GND 0.02fF
C304 s3 GND 0.55fF
C305 a_1380_n779# GND 0.03fF
C306 a_n28_n779# GND 0.03fF
C307 a_n178_n779# GND 0.03fF
C308 a_2442_n779# GND 0.94fF
C309 CMOS_3in_OR_0/C GND 1.11fF $ **FLOATING
C310 CMOS_AND_1/AND GND 0.58fF
C311 a_1380_n1689# GND 0.50fF
C312 a_n328_n1689# GND 0.71fF
C313 a_2592_n111# GND 0.02fF
C314 a_1735_n111# GND 0.03fF
C315 a_1435_n111# GND 0.02fF
C316 a_177_n111# GND 0.02fF
C317 a_n123_n111# GND 0.02fF
C318 CMOS_AND_0/AND GND 1.97fF
C319 a_1735_499# GND 0.01fF
C320 a_1435_499# GND 0.01fF
C321 CMOS_AND_1/A GND 1.10fF
C322 a_177_499# GND 0.01fF
C323 a_n123_499# GND 0.01fF
C324 a_2592_499# GND 0.54fF
C325 CMOS_AND_0/A GND 1.16fF
C326 x2_bar GND 2.66fF
C327 x2 GND 6.06fF
C328 x3_bar GND 4.24fF
C329 a_27_n111# GND 0.64fF
C330 x1_bar GND 6.35fF
C331 x1 GND 2.34fF
C332 x0_bar GND 6.10fF
C333 x3 GND 1.67fF
C334 x0 GND 3.16fF
C335 VDD GND 24.56fF
C336 x0_bar.t1 GND 0.25fF
C337 x0_bar.t0 GND 0.25fF
C338 x0_bar.n0 GND 0.68fF $ **FLOATING
C339 x2.t1 GND 0.28fF
C340 x2.t0 GND 0.11fF
C341 x2.n0 GND 0.31fF $ **FLOATING
C342 x2.n1 GND 1.75fF $ **FLOATING
C343 CMOS_3in_OR_0/C.t2 GND 0.10fF
C344 CMOS_3in_OR_0/C.t3 GND 0.12fF
C345 CMOS_3in_OR_0/C.t0 GND 0.31fF
C346 CMOS_3in_OR_0/C.t1 GND 0.29fF
C347 CMOS_3in_AND_0/OUT GND 0.19fF $ **FLOATING
C348 CMOS_3in_OR_0/C.n0 GND 0.70fF $ **FLOATING
C349 x2_bar.t2 GND 0.25fF
C350 x2_bar.t3 GND 0.23fF
C351 x2_bar.t1 GND 0.18fF
C352 x2_bar.t0 GND 0.21fF
C353 x2_bar.n0 GND 0.32fF $ **FLOATING
C354 x2_bar.n1 GND 4.53fF $ **FLOATING
C355 CMOS_XOR_0/A_bar GND 0.40fF $ **FLOATING
C356 x1_bar.t1 GND 0.30fF
C357 x1_bar.t0 GND 0.27fF
C358 x0.t1 GND 0.52fF
C359 x0.t0 GND 0.35fF
C360 x0.t3 GND 0.20fF
C361 x0.t2 GND 0.16fF
C362 x0.n0 GND 3.47fF $ **FLOATING
C363 CMOS_XNOR_0/B GND 0.50fF $ **FLOATING
C364 x3_bar.t3 GND 0.17fF
C365 x3_bar.t2 GND 0.15fF
C366 x3_bar.t1 GND 0.10fF
C367 x3_bar.t0 GND 0.15fF
C368 x3_bar.n0 GND 0.20fF $ **FLOATING
C369 x3_bar.n1 GND 0.65fF $ **FLOATING
C370 x3_bar.n2 GND 3.60fF $ **FLOATING
C371 x3_bar.n3 GND 1.00fF $ **FLOATING
C372 CMOS_XOR_0/B_bar GND 0.03fF $ **FLOATING
C373 x1.t3 GND 0.13fF
C374 x1.t0 GND 0.09fF
C375 x1.n0 GND 0.18fF $ **FLOATING
C376 x1.t1 GND 0.17fF
C377 x1.t2 GND 0.07fF
C378 x1.n1 GND 0.19fF $ **FLOATING
C379 CMOS_XNOR_0/A GND 0.25fF $ **FLOATING
C380 x1.n2 GND 3.51fF $ **FLOATING
C381 x1.n3 GND 1.12fF $ **FLOATING
C382 x3.t2 GND 0.50fF
C383 x3.t0 GND 0.34fF
C384 x3.t3 GND 0.09fF
C385 x3.t1 GND 0.13fF
C386 x3.n0 GND 0.16fF $ **FLOATING
C387 x3.n1 GND 3.83fF $ **FLOATING
C388 CMOS_XOR_0/B GND 0.32fF $ **FLOATING
C389 VDD.t11 GND 0.07fF
C390 VDD.t27 GND 0.07fF
C391 VDD.t6 GND 0.07fF
C392 CMOS_XOR_0/VDD GND 0.01fF $ **FLOATING
C393 VDD.t9 GND 0.07fF
C394 VDD.t33 GND 0.07fF
C395 VDD.t31 GND 0.07fF
C396 VDD.n0 GND 0.21fF $ **FLOATING
C397 VDD.n1 GND 0.02fF $ **FLOATING
C398 VDD.n2 GND 0.02fF $ **FLOATING
C399 VDD.n3 GND 0.15fF $ **FLOATING
C400 VDD.t30 GND 0.10fF
C401 VDD.n4 GND 0.10fF $ **FLOATING
C402 VDD.n5 GND 0.02fF $ **FLOATING
C403 VDD.n6 GND 0.02fF $ **FLOATING
C404 VDD.n7 GND 0.06fF $ **FLOATING
C405 VDD.n8 GND 0.38fF $ **FLOATING
C406 VDD.n9 GND 0.17fF $ **FLOATING
C407 VDD.n10 GND 0.02fF $ **FLOATING
C408 VDD.n11 GND 0.02fF $ **FLOATING
C409 VDD.n12 GND 0.01fF $ **FLOATING
C410 VDD.n13 GND 0.17fF $ **FLOATING
C411 VDD.n14 GND 0.02fF $ **FLOATING
C412 VDD.n15 GND 0.02fF $ **FLOATING
C413 VDD.n16 GND 0.02fF $ **FLOATING
C414 VDD.n17 GND 0.17fF $ **FLOATING
C415 VDD.n18 GND 0.02fF $ **FLOATING
C416 VDD.n19 GND 0.02fF $ **FLOATING
C417 VDD.n20 GND 0.02fF $ **FLOATING
C418 VDD.t29 GND 0.07fF
C419 VDD.n21 GND 0.37fF $ **FLOATING
C420 VDD.n22 GND 0.01fF $ **FLOATING
C421 VDD.n23 GND 0.17fF $ **FLOATING
C422 VDD.n24 GND 0.02fF $ **FLOATING
C423 VDD.n25 GND 0.02fF $ **FLOATING
C424 VDD.t28 GND 0.09fF
C425 VDD.n26 GND 0.11fF $ **FLOATING
C426 VDD.n27 GND 0.02fF $ **FLOATING
C427 VDD.n28 GND 0.02fF $ **FLOATING
C428 VDD.n29 GND 0.02fF $ **FLOATING
C429 VDD.n30 GND 0.15fF $ **FLOATING
C430 VDD.n31 GND 0.02fF $ **FLOATING
C431 VDD.n32 GND 0.02fF $ **FLOATING
C432 VDD.n33 GND 0.02fF $ **FLOATING
C433 VDD.t32 GND 0.10fF
C434 VDD.n34 GND 0.12fF $ **FLOATING
C435 VDD.n35 GND 0.02fF $ **FLOATING
C436 VDD.n36 GND 0.02fF $ **FLOATING
C437 VDD.n37 GND 0.02fF $ **FLOATING
C438 VDD.n38 GND 0.19fF $ **FLOATING
C439 VDD.n39 GND 0.02fF $ **FLOATING
C440 VDD.n40 GND 0.02fF $ **FLOATING
C441 VDD.n41 GND 0.01fF $ **FLOATING
C442 VDD.n42 GND 0.38fF $ **FLOATING
C443 VDD.n43 GND 0.18fF $ **FLOATING
C444 VDD.n44 GND 0.06fF $ **FLOATING
C445 VDD.n45 GND 0.15fF $ **FLOATING
C446 VDD.n46 GND 0.06fF $ **FLOATING
C447 VDD.n47 GND 0.21fF $ **FLOATING
C448 VDD.n48 GND 0.02fF $ **FLOATING
C449 VDD.n49 GND 0.02fF $ **FLOATING
C450 VDD.n50 GND 0.01fF $ **FLOATING
C451 VDD.n51 GND 0.38fF $ **FLOATING
C452 VDD.t8 GND 0.09fF
C453 VDD.n52 GND 0.13fF $ **FLOATING
C454 VDD.n53 GND 0.02fF $ **FLOATING
C455 VDD.n54 GND 0.02fF $ **FLOATING
C456 VDD.n55 GND 0.02fF $ **FLOATING
C457 VDD.n56 GND 0.15fF $ **FLOATING
C458 VDD.n57 GND 0.02fF $ **FLOATING
C459 VDD.n58 GND 0.02fF $ **FLOATING
C460 VDD.n59 GND 0.02fF $ **FLOATING
C461 VDD.t17 GND 0.09fF
C462 VDD.n60 GND 0.12fF $ **FLOATING
C463 VDD.n61 GND 0.02fF $ **FLOATING
C464 VDD.n62 GND 0.02fF $ **FLOATING
C465 VDD.n63 GND 0.02fF $ **FLOATING
C466 VDD.n64 GND 0.14fF $ **FLOATING
C467 VDD.n65 GND 0.02fF $ **FLOATING
C468 VDD.n66 GND 0.02fF $ **FLOATING
C469 VDD.n67 GND 0.02fF $ **FLOATING
C470 VDD.n68 GND 0.01fF $ **FLOATING
C471 VDD.n69 GND 0.13fF $ **FLOATING
C472 VDD.n70 GND 0.02fF $ **FLOATING
C473 VDD.n71 GND 0.02fF $ **FLOATING
C474 VDD.t7 GND 0.09fF
C475 VDD.n72 GND 0.13fF $ **FLOATING
C476 VDD.n73 GND 0.02fF $ **FLOATING
C477 VDD.n74 GND 0.02fF $ **FLOATING
C478 VDD.n75 GND 0.02fF $ **FLOATING
C479 VDD.n76 GND 0.14fF $ **FLOATING
C480 VDD.n77 GND 0.02fF $ **FLOATING
C481 VDD.n78 GND 0.02fF $ **FLOATING
C482 VDD.n79 GND 0.02fF $ **FLOATING
C483 VDD.t5 GND 0.09fF
C484 VDD.n80 GND 0.13fF $ **FLOATING
C485 VDD.n81 GND 0.02fF $ **FLOATING
C486 VDD.n82 GND 0.02fF $ **FLOATING
C487 VDD.n83 GND 0.02fF $ **FLOATING
C488 VDD.n84 GND 0.38fF $ **FLOATING
C489 VDD.n85 GND 0.20fF $ **FLOATING
C490 VDD.n86 GND 0.02fF $ **FLOATING
C491 VDD.n87 GND 0.02fF $ **FLOATING
C492 VDD.n88 GND 0.01fF $ **FLOATING
C493 VDD.n89 GND 0.11fF $ **FLOATING
C494 VDD.n90 GND 0.06fF $ **FLOATING
C495 VDD.n91 GND 0.17fF $ **FLOATING
C496 VDD.n92 GND 0.06fF $ **FLOATING
C497 VDD.n93 GND 0.20fF $ **FLOATING
C498 VDD.n94 GND 0.02fF $ **FLOATING
C499 VDD.n95 GND 0.02fF $ **FLOATING
C500 VDD.n96 GND 0.02fF $ **FLOATING
C501 VDD.t26 GND 0.10fF
C502 VDD.n97 GND 0.11fF $ **FLOATING
C503 VDD.n98 GND 0.02fF $ **FLOATING
C504 VDD.n99 GND 0.02fF $ **FLOATING
C505 VDD.n100 GND 0.02fF $ **FLOATING
C506 VDD.n101 GND 0.38fF $ **FLOATING
C507 VDD.n102 GND 0.17fF $ **FLOATING
C508 VDD.n103 GND 0.02fF $ **FLOATING
C509 VDD.n104 GND 0.02fF $ **FLOATING
C510 VDD.n105 GND 0.01fF $ **FLOATING
C511 VDD.n106 GND 0.17fF $ **FLOATING
C512 VDD.n107 GND 0.02fF $ **FLOATING
C513 VDD.n108 GND 0.02fF $ **FLOATING
C514 VDD.n109 GND 0.02fF $ **FLOATING
C515 VDD.n110 GND 0.17fF $ **FLOATING
C516 VDD.n111 GND 0.02fF $ **FLOATING
C517 VDD.n112 GND 0.02fF $ **FLOATING
C518 VDD.n113 GND 0.02fF $ **FLOATING
C519 VDD.n114 GND 0.17fF $ **FLOATING
C520 VDD.n115 GND 0.02fF $ **FLOATING
C521 VDD.n116 GND 0.02fF $ **FLOATING
C522 VDD.n117 GND 0.01fF $ **FLOATING
C523 VDD.n118 GND 0.38fF $ **FLOATING
C524 VDD.t10 GND 0.09fF
C525 VDD.n119 GND 0.12fF $ **FLOATING
C526 VDD.n120 GND 0.02fF $ **FLOATING
C527 VDD.n121 GND 0.02fF $ **FLOATING
C528 VDD.n122 GND 0.02fF $ **FLOATING
C529 VDD.n123 GND 0.15fF $ **FLOATING
C530 VDD.n124 GND 0.02fF $ **FLOATING
C531 VDD.n125 GND 0.02fF $ **FLOATING
C532 VDD.n126 GND 0.02fF $ **FLOATING
C533 VDD.t4 GND 0.09fF
C534 VDD.n127 GND 0.12fF $ **FLOATING
C535 VDD.n128 GND 0.02fF $ **FLOATING
C536 VDD.n129 GND 0.02fF $ **FLOATING
C537 VDD.n130 GND 0.02fF $ **FLOATING
C538 VDD.n131 GND 0.14fF $ **FLOATING
C539 VDD.n132 GND 0.02fF $ **FLOATING
C540 VDD.n133 GND 0.02fF $ **FLOATING
C541 VDD.n134 GND 0.02fF $ **FLOATING
C542 VDD.t37 GND 0.09fF
C543 VDD.n135 GND 0.13fF $ **FLOATING
C544 VDD.n136 GND 0.02fF $ **FLOATING
C545 VDD.n137 GND 0.02fF $ **FLOATING
C546 VDD.n138 GND 0.01fF $ **FLOATING
C547 VDD.t19 GND 0.07fF
C548 VDD.t16 GND 0.05fF
C549 VDD.t1 GND 0.05fF
C550 VDD.n139 GND 0.19fF $ **FLOATING
C551 CMOS_3in_AND_0/VDD GND 0.01fF $ **FLOATING
C552 VDD.t13 GND 0.07fF
C553 VDD.t21 GND 0.07fF
C554 VDD.t3 GND 0.07fF
C555 CMOS_AND_1/VDD GND 0.01fF $ **FLOATING
C556 VDD.t39 GND 0.07fF
C557 VDD.t23 GND 0.07fF
C558 CMOS_3in_OR_0/VDD GND 0.01fF $ **FLOATING
C559 VDD.t25 GND 0.07fF
C560 VDD.n140 GND 0.20fF $ **FLOATING
C561 VDD.n141 GND 0.02fF $ **FLOATING
C562 VDD.n142 GND 0.02fF $ **FLOATING
C563 VDD.n143 GND 0.17fF $ **FLOATING
C564 VDD.t24 GND 0.10fF
C565 VDD.n144 GND 0.11fF $ **FLOATING
C566 VDD.n145 GND 0.02fF $ **FLOATING
C567 VDD.n146 GND 0.02fF $ **FLOATING
C568 VDD.n147 GND 0.05fF $ **FLOATING
C569 VDD.n148 GND 0.38fF $ **FLOATING
C570 VDD.n149 GND 0.17fF $ **FLOATING
C571 VDD.n150 GND 0.02fF $ **FLOATING
C572 VDD.n151 GND 0.02fF $ **FLOATING
C573 VDD.n152 GND 0.01fF $ **FLOATING
C574 VDD.n153 GND 0.17fF $ **FLOATING
C575 VDD.n154 GND 0.02fF $ **FLOATING
C576 VDD.n155 GND 0.02fF $ **FLOATING
C577 VDD.n156 GND 0.02fF $ **FLOATING
C578 VDD.n157 GND 0.17fF $ **FLOATING
C579 VDD.n158 GND 0.02fF $ **FLOATING
C580 VDD.n159 GND 0.02fF $ **FLOATING
C581 VDD.n160 GND 0.02fF $ **FLOATING
C582 VDD.n161 GND 0.17fF $ **FLOATING
C583 VDD.n162 GND 0.02fF $ **FLOATING
C584 VDD.n163 GND 0.02fF $ **FLOATING
C585 VDD.n164 GND 0.02fF $ **FLOATING
C586 VDD.t14 GND 0.09fF
C587 VDD.n165 GND 0.10fF $ **FLOATING
C588 VDD.n166 GND 0.02fF $ **FLOATING
C589 VDD.n167 GND 0.02fF $ **FLOATING
C590 VDD.n168 GND 0.02fF $ **FLOATING
C591 VDD.n169 GND 0.01fF $ **FLOATING
C592 VDD.n170 GND 0.16fF $ **FLOATING
C593 VDD.n171 GND 0.02fF $ **FLOATING
C594 VDD.n172 GND 0.02fF $ **FLOATING
C595 VDD.t34 GND 0.09fF
C596 VDD.n173 GND 0.11fF $ **FLOATING
C597 VDD.n174 GND 0.02fF $ **FLOATING
C598 VDD.n175 GND 0.02fF $ **FLOATING
C599 VDD.n176 GND 0.02fF $ **FLOATING
C600 VDD.n177 GND 0.15fF $ **FLOATING
C601 VDD.n178 GND 0.02fF $ **FLOATING
C602 VDD.n179 GND 0.02fF $ **FLOATING
C603 VDD.n180 GND 0.02fF $ **FLOATING
C604 VDD.t22 GND 0.10fF
C605 VDD.n181 GND 0.12fF $ **FLOATING
C606 VDD.n182 GND 0.02fF $ **FLOATING
C607 VDD.n183 GND 0.02fF $ **FLOATING
C608 VDD.n184 GND 0.02fF $ **FLOATING
C609 VDD.n185 GND 0.19fF $ **FLOATING
C610 VDD.n186 GND 0.02fF $ **FLOATING
C611 VDD.n187 GND 0.02fF $ **FLOATING
C612 VDD.n188 GND 0.01fF $ **FLOATING
C613 VDD.n189 GND 0.38fF $ **FLOATING
C614 VDD.n190 GND 0.18fF $ **FLOATING
C615 VDD.n191 GND 0.06fF $ **FLOATING
C616 VDD.n192 GND 0.16fF $ **FLOATING
C617 VDD.n193 GND 0.06fF $ **FLOATING
C618 VDD.n194 GND 0.20fF $ **FLOATING
C619 VDD.n195 GND 0.02fF $ **FLOATING
C620 VDD.n196 GND 0.02fF $ **FLOATING
C621 VDD.n197 GND 0.02fF $ **FLOATING
C622 VDD.t38 GND 0.10fF
C623 VDD.n198 GND 0.10fF $ **FLOATING
C624 VDD.n199 GND 0.02fF $ **FLOATING
C625 VDD.n200 GND 0.02fF $ **FLOATING
C626 VDD.n201 GND 0.02fF $ **FLOATING
C627 VDD.n202 GND 0.38fF $ **FLOATING
C628 VDD.n203 GND 0.17fF $ **FLOATING
C629 VDD.n204 GND 0.02fF $ **FLOATING
C630 VDD.n205 GND 0.02fF $ **FLOATING
C631 VDD.n206 GND 0.01fF $ **FLOATING
C632 VDD.n207 GND 0.17fF $ **FLOATING
C633 VDD.n208 GND 0.02fF $ **FLOATING
C634 VDD.n209 GND 0.02fF $ **FLOATING
C635 VDD.n210 GND 0.02fF $ **FLOATING
C636 VDD.n211 GND 0.17fF $ **FLOATING
C637 VDD.n212 GND 0.02fF $ **FLOATING
C638 VDD.n213 GND 0.02fF $ **FLOATING
C639 VDD.n214 GND 0.02fF $ **FLOATING
C640 VDD.t36 GND 0.07fF
C641 VDD.n215 GND 0.37fF $ **FLOATING
C642 VDD.n216 GND 0.01fF $ **FLOATING
C643 VDD.n217 GND 0.17fF $ **FLOATING
C644 VDD.n218 GND 0.02fF $ **FLOATING
C645 VDD.n219 GND 0.02fF $ **FLOATING
C646 VDD.t35 GND 0.09fF
C647 VDD.n220 GND 0.11fF $ **FLOATING
C648 VDD.n221 GND 0.02fF $ **FLOATING
C649 VDD.n222 GND 0.02fF $ **FLOATING
C650 VDD.n223 GND 0.02fF $ **FLOATING
C651 VDD.n224 GND 0.15fF $ **FLOATING
C652 VDD.n225 GND 0.02fF $ **FLOATING
C653 VDD.n226 GND 0.02fF $ **FLOATING
C654 VDD.n227 GND 0.02fF $ **FLOATING
C655 VDD.t2 GND 0.10fF
C656 VDD.n228 GND 0.12fF $ **FLOATING
C657 VDD.n229 GND 0.02fF $ **FLOATING
C658 VDD.n230 GND 0.02fF $ **FLOATING
C659 VDD.n231 GND 0.02fF $ **FLOATING
C660 VDD.n232 GND 0.19fF $ **FLOATING
C661 VDD.n233 GND 0.02fF $ **FLOATING
C662 VDD.n234 GND 0.02fF $ **FLOATING
C663 VDD.n235 GND 0.01fF $ **FLOATING
C664 VDD.n236 GND 0.38fF $ **FLOATING
C665 VDD.n237 GND 0.18fF $ **FLOATING
C666 VDD.n238 GND 0.09fF $ **FLOATING
C667 VDD.n239 GND 0.17fF $ **FLOATING
C668 VDD.n240 GND 0.09fF $ **FLOATING
C669 VDD.n241 GND 0.20fF $ **FLOATING
C670 VDD.n242 GND 0.02fF $ **FLOATING
C671 VDD.n243 GND 0.02fF $ **FLOATING
C672 VDD.n244 GND 0.02fF $ **FLOATING
C673 VDD.t20 GND 0.10fF
C674 VDD.n245 GND 0.11fF $ **FLOATING
C675 VDD.n246 GND 0.02fF $ **FLOATING
C676 VDD.n247 GND 0.02fF $ **FLOATING
C677 VDD.n248 GND 0.02fF $ **FLOATING
C678 VDD.n249 GND 0.38fF $ **FLOATING
C679 VDD.n250 GND 0.17fF $ **FLOATING
C680 VDD.n251 GND 0.02fF $ **FLOATING
C681 VDD.n252 GND 0.02fF $ **FLOATING
C682 VDD.n253 GND 0.01fF $ **FLOATING
C683 VDD.n254 GND 0.17fF $ **FLOATING
C684 VDD.n255 GND 0.02fF $ **FLOATING
C685 VDD.n256 GND 0.02fF $ **FLOATING
C686 VDD.n257 GND 0.02fF $ **FLOATING
C687 VDD.n258 GND 0.17fF $ **FLOATING
C688 VDD.n259 GND 0.02fF $ **FLOATING
C689 VDD.n260 GND 0.02fF $ **FLOATING
C690 VDD.n261 GND 0.02fF $ **FLOATING
C691 VDD.n262 GND 0.17fF $ **FLOATING
C692 VDD.n263 GND 0.02fF $ **FLOATING
C693 VDD.n264 GND 0.02fF $ **FLOATING
C694 VDD.n265 GND 0.01fF $ **FLOATING
C695 VDD.n266 GND 0.38fF $ **FLOATING
C696 VDD.t12 GND 0.09fF
C697 VDD.n267 GND 0.10fF $ **FLOATING
C698 VDD.n268 GND 0.02fF $ **FLOATING
C699 VDD.n269 GND 0.02fF $ **FLOATING
C700 VDD.n270 GND 0.02fF $ **FLOATING
C701 VDD.n271 GND 0.01fF $ **FLOATING
C702 VDD.n272 GND 0.16fF $ **FLOATING
C703 VDD.n273 GND 0.02fF $ **FLOATING
C704 VDD.n274 GND 0.02fF $ **FLOATING
C705 VDD.t15 GND 0.09fF
C706 VDD.n275 GND 0.11fF $ **FLOATING
C707 VDD.n276 GND 0.02fF $ **FLOATING
C708 VDD.n277 GND 0.02fF $ **FLOATING
C709 VDD.n278 GND 0.02fF $ **FLOATING
C710 VDD.n279 GND 0.15fF $ **FLOATING
C711 VDD.n280 GND 0.02fF $ **FLOATING
C712 VDD.n281 GND 0.02fF $ **FLOATING
C713 VDD.n282 GND 0.01fF $ **FLOATING
C714 VDD.n283 GND 0.16fF $ **FLOATING
C715 VDD.t0 GND 0.10fF
C716 VDD.n284 GND 0.12fF $ **FLOATING
C717 VDD.n285 GND 0.02fF $ **FLOATING
C718 VDD.n286 GND 0.02fF $ **FLOATING
C719 VDD.n287 GND 0.02fF $ **FLOATING
C720 VDD.n288 GND 0.19fF $ **FLOATING
C721 VDD.n289 GND 0.02fF $ **FLOATING
C722 VDD.n290 GND 0.02fF $ **FLOATING
C723 VDD.n291 GND 0.02fF $ **FLOATING
C724 VDD.n292 GND 0.18fF $ **FLOATING
C725 VDD.n293 GND 0.36fF $ **FLOATING
C726 VDD.n294 GND 0.35fF $ **FLOATING
C727 VDD.n295 GND 0.11fF $ **FLOATING
C728 VDD.n296 GND 0.02fF $ **FLOATING
C729 VDD.n297 GND 0.20fF $ **FLOATING
C730 VDD.n298 GND 0.02fF $ **FLOATING
C731 VDD.n299 GND 0.02fF $ **FLOATING
C732 VDD.n300 GND 0.01fF $ **FLOATING
C733 VDD.n301 GND 0.38fF $ **FLOATING
C734 VDD.t18 GND 0.09fF
C735 VDD.n302 GND 0.13fF $ **FLOATING
C736 VDD.n303 GND 0.02fF $ **FLOATING
C737 VDD.n304 GND 0.02fF $ **FLOATING
C738 VDD.n305 GND 0.02fF $ **FLOATING
C739 VDD.n306 GND 0.14fF $ **FLOATING
C740 VDD.n307 GND 0.02fF $ **FLOATING
C741 VDD.n308 GND 0.02fF $ **FLOATING
C742 VDD.n309 GND 0.02fF $ **FLOATING
C743 VDD.n310 GND 0.13fF $ **FLOATING
C744 VDD.n311 GND 0.02fF $ **FLOATING
C745 VDD.n312 GND 0.02fF $ **FLOATING
C746 VDD.n313 GND 0.02fF $ **FLOATING
C747 CMOS_XNOR_0/VDD GND 0.01fF $ **FLOATING
.ends

