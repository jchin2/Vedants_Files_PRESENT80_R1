magic
tech sky130A
magscale 1 2
timestamp 1671058898
<< xpolycontact >>
rect -512 69 -442 501
rect -512 -501 -442 -69
rect -194 69 -124 501
rect -194 -501 -124 -69
rect 124 69 194 501
rect 124 -501 194 -69
rect 442 69 512 501
rect 442 -501 512 -69
<< xpolyres >>
rect -512 -69 -442 69
rect -194 -69 -124 69
rect 124 -69 194 69
rect 442 -69 512 69
<< viali >>
rect -494 447 -460 481
rect -494 375 -460 409
rect -494 303 -460 337
rect -494 231 -460 265
rect -494 159 -460 193
rect -494 87 -460 121
rect -176 447 -142 481
rect -176 375 -142 409
rect -176 303 -142 337
rect -176 231 -142 265
rect -176 159 -142 193
rect -176 87 -142 121
rect 142 447 176 481
rect 142 375 176 409
rect 142 303 176 337
rect 142 231 176 265
rect 142 159 176 193
rect 142 87 176 121
rect 460 447 494 481
rect 460 375 494 409
rect 460 303 494 337
rect 460 231 494 265
rect 460 159 494 193
rect 460 87 494 121
rect -494 -122 -460 -88
rect -494 -194 -460 -160
rect -494 -266 -460 -232
rect -494 -338 -460 -304
rect -494 -410 -460 -376
rect -494 -482 -460 -448
rect -176 -122 -142 -88
rect -176 -194 -142 -160
rect -176 -266 -142 -232
rect -176 -338 -142 -304
rect -176 -410 -142 -376
rect -176 -482 -142 -448
rect 142 -122 176 -88
rect 142 -194 176 -160
rect 142 -266 176 -232
rect 142 -338 176 -304
rect 142 -410 176 -376
rect 142 -482 176 -448
rect 460 -122 494 -88
rect 460 -194 494 -160
rect 460 -266 494 -232
rect 460 -338 494 -304
rect 460 -410 494 -376
rect 460 -482 494 -448
<< metal1 >>
rect -502 481 -452 495
rect -502 447 -494 481
rect -460 447 -452 481
rect -502 409 -452 447
rect -502 375 -494 409
rect -460 375 -452 409
rect -502 337 -452 375
rect -502 303 -494 337
rect -460 303 -452 337
rect -502 265 -452 303
rect -502 231 -494 265
rect -460 231 -452 265
rect -502 193 -452 231
rect -502 159 -494 193
rect -460 159 -452 193
rect -502 121 -452 159
rect -502 87 -494 121
rect -460 87 -452 121
rect -502 74 -452 87
rect -184 481 -134 495
rect -184 447 -176 481
rect -142 447 -134 481
rect -184 409 -134 447
rect -184 375 -176 409
rect -142 375 -134 409
rect -184 337 -134 375
rect -184 303 -176 337
rect -142 303 -134 337
rect -184 265 -134 303
rect -184 231 -176 265
rect -142 231 -134 265
rect -184 193 -134 231
rect -184 159 -176 193
rect -142 159 -134 193
rect -184 121 -134 159
rect -184 87 -176 121
rect -142 87 -134 121
rect -184 74 -134 87
rect 134 481 184 495
rect 134 447 142 481
rect 176 447 184 481
rect 134 409 184 447
rect 134 375 142 409
rect 176 375 184 409
rect 134 337 184 375
rect 134 303 142 337
rect 176 303 184 337
rect 134 265 184 303
rect 134 231 142 265
rect 176 231 184 265
rect 134 193 184 231
rect 134 159 142 193
rect 176 159 184 193
rect 134 121 184 159
rect 134 87 142 121
rect 176 87 184 121
rect 134 74 184 87
rect 452 481 502 495
rect 452 447 460 481
rect 494 447 502 481
rect 452 409 502 447
rect 452 375 460 409
rect 494 375 502 409
rect 452 337 502 375
rect 452 303 460 337
rect 494 303 502 337
rect 452 265 502 303
rect 452 231 460 265
rect 494 231 502 265
rect 452 193 502 231
rect 452 159 460 193
rect 494 159 502 193
rect 452 121 502 159
rect 452 87 460 121
rect 494 87 502 121
rect 452 74 502 87
rect -502 -88 -452 -74
rect -502 -122 -494 -88
rect -460 -122 -452 -88
rect -502 -160 -452 -122
rect -502 -194 -494 -160
rect -460 -194 -452 -160
rect -502 -232 -452 -194
rect -502 -266 -494 -232
rect -460 -266 -452 -232
rect -502 -304 -452 -266
rect -502 -338 -494 -304
rect -460 -338 -452 -304
rect -502 -376 -452 -338
rect -502 -410 -494 -376
rect -460 -410 -452 -376
rect -502 -448 -452 -410
rect -502 -482 -494 -448
rect -460 -482 -452 -448
rect -502 -495 -452 -482
rect -184 -88 -134 -74
rect -184 -122 -176 -88
rect -142 -122 -134 -88
rect -184 -160 -134 -122
rect -184 -194 -176 -160
rect -142 -194 -134 -160
rect -184 -232 -134 -194
rect -184 -266 -176 -232
rect -142 -266 -134 -232
rect -184 -304 -134 -266
rect -184 -338 -176 -304
rect -142 -338 -134 -304
rect -184 -376 -134 -338
rect -184 -410 -176 -376
rect -142 -410 -134 -376
rect -184 -448 -134 -410
rect -184 -482 -176 -448
rect -142 -482 -134 -448
rect -184 -495 -134 -482
rect 134 -88 184 -74
rect 134 -122 142 -88
rect 176 -122 184 -88
rect 134 -160 184 -122
rect 134 -194 142 -160
rect 176 -194 184 -160
rect 134 -232 184 -194
rect 134 -266 142 -232
rect 176 -266 184 -232
rect 134 -304 184 -266
rect 134 -338 142 -304
rect 176 -338 184 -304
rect 134 -376 184 -338
rect 134 -410 142 -376
rect 176 -410 184 -376
rect 134 -448 184 -410
rect 134 -482 142 -448
rect 176 -482 184 -448
rect 134 -495 184 -482
rect 452 -88 502 -74
rect 452 -122 460 -88
rect 494 -122 502 -88
rect 452 -160 502 -122
rect 452 -194 460 -160
rect 494 -194 502 -160
rect 452 -232 502 -194
rect 452 -266 460 -232
rect 494 -266 502 -232
rect 452 -304 502 -266
rect 452 -338 460 -304
rect 494 -338 502 -304
rect 452 -376 502 -338
rect 452 -410 460 -376
rect 494 -410 502 -376
rect 452 -448 502 -410
rect 452 -482 460 -448
rect 494 -482 502 -448
rect 452 -495 502 -482
<< end >>
