magic
tech sky130A
timestamp 1666994426
<< nwell >>
rect -170 760 710 855
rect 65 565 475 760
<< nmos >>
rect -90 205 -75 355
rect -15 205 0 355
rect 150 205 165 355
rect 225 205 240 355
rect 300 205 315 355
rect 375 205 390 355
rect 540 205 555 355
rect 615 205 630 355
<< pmos >>
rect 150 590 165 740
rect 225 590 240 740
rect 300 590 315 740
rect 375 590 390 740
<< ndiff >>
rect -150 320 -90 355
rect -150 300 -130 320
rect -110 300 -90 320
rect -150 280 -90 300
rect -150 260 -130 280
rect -110 260 -90 280
rect -150 240 -90 260
rect -150 220 -130 240
rect -110 220 -90 240
rect -150 205 -90 220
rect -75 320 -15 355
rect -75 300 -55 320
rect -35 300 -15 320
rect -75 280 -15 300
rect -75 260 -55 280
rect -35 260 -15 280
rect -75 240 -15 260
rect -75 220 -55 240
rect -35 220 -15 240
rect -75 205 -15 220
rect 0 320 60 355
rect 0 300 20 320
rect 40 300 60 320
rect 0 280 60 300
rect 0 260 20 280
rect 40 260 60 280
rect 0 240 60 260
rect 0 220 20 240
rect 40 220 60 240
rect 0 205 60 220
rect 90 320 150 355
rect 90 300 110 320
rect 130 300 150 320
rect 90 280 150 300
rect 90 260 110 280
rect 130 260 150 280
rect 90 240 150 260
rect 90 220 110 240
rect 130 220 150 240
rect 90 205 150 220
rect 165 320 225 355
rect 165 300 185 320
rect 205 300 225 320
rect 165 280 225 300
rect 165 260 185 280
rect 205 260 225 280
rect 165 240 225 260
rect 165 220 185 240
rect 205 220 225 240
rect 165 205 225 220
rect 240 320 300 355
rect 240 300 260 320
rect 280 300 300 320
rect 240 280 300 300
rect 240 260 260 280
rect 280 260 300 280
rect 240 240 300 260
rect 240 220 260 240
rect 280 220 300 240
rect 240 205 300 220
rect 315 320 375 355
rect 315 300 335 320
rect 355 300 375 320
rect 315 280 375 300
rect 315 260 335 280
rect 355 260 375 280
rect 315 240 375 260
rect 315 220 335 240
rect 355 220 375 240
rect 315 205 375 220
rect 390 320 450 355
rect 390 300 410 320
rect 430 300 450 320
rect 390 280 450 300
rect 390 260 410 280
rect 430 260 450 280
rect 390 240 450 260
rect 390 220 410 240
rect 430 220 450 240
rect 390 205 450 220
rect 480 320 540 355
rect 480 300 500 320
rect 520 300 540 320
rect 480 280 540 300
rect 480 260 500 280
rect 520 260 540 280
rect 480 240 540 260
rect 480 220 500 240
rect 520 220 540 240
rect 480 205 540 220
rect 555 205 615 355
rect 630 320 690 355
rect 630 300 650 320
rect 670 300 690 320
rect 630 280 690 300
rect 630 260 650 280
rect 670 260 690 280
rect 630 240 690 260
rect 630 220 650 240
rect 670 220 690 240
rect 630 205 690 220
<< pdiff >>
rect 90 705 150 740
rect 90 685 110 705
rect 130 685 150 705
rect 90 665 150 685
rect 90 645 110 665
rect 130 645 150 665
rect 90 625 150 645
rect 90 605 110 625
rect 130 605 150 625
rect 90 590 150 605
rect 165 705 225 740
rect 165 685 185 705
rect 205 685 225 705
rect 165 665 225 685
rect 165 645 185 665
rect 205 645 225 665
rect 165 625 225 645
rect 165 605 185 625
rect 205 605 225 625
rect 165 590 225 605
rect 240 705 300 740
rect 240 685 260 705
rect 280 685 300 705
rect 240 665 300 685
rect 240 645 260 665
rect 280 645 300 665
rect 240 625 300 645
rect 240 605 260 625
rect 280 605 300 625
rect 240 590 300 605
rect 315 705 375 740
rect 315 685 335 705
rect 355 685 375 705
rect 315 665 375 685
rect 315 645 335 665
rect 355 645 375 665
rect 315 625 375 645
rect 315 605 335 625
rect 355 605 375 625
rect 315 590 375 605
rect 390 705 450 740
rect 390 685 410 705
rect 430 685 450 705
rect 390 665 450 685
rect 390 645 410 665
rect 430 645 450 665
rect 390 625 450 645
rect 390 605 410 625
rect 430 605 450 625
rect 390 590 450 605
<< ndiffc >>
rect -130 300 -110 320
rect -130 260 -110 280
rect -130 220 -110 240
rect -55 300 -35 320
rect -55 260 -35 280
rect -55 220 -35 240
rect 20 300 40 320
rect 20 260 40 280
rect 20 220 40 240
rect 110 300 130 320
rect 110 260 130 280
rect 110 220 130 240
rect 185 300 205 320
rect 185 260 205 280
rect 185 220 205 240
rect 260 300 280 320
rect 260 260 280 280
rect 260 220 280 240
rect 335 300 355 320
rect 335 260 355 280
rect 335 220 355 240
rect 410 300 430 320
rect 410 260 430 280
rect 410 220 430 240
rect 500 300 520 320
rect 500 260 520 280
rect 500 220 520 240
rect 650 300 670 320
rect 650 260 670 280
rect 650 220 670 240
<< pdiffc >>
rect 110 685 130 705
rect 110 645 130 665
rect 110 605 130 625
rect 185 685 205 705
rect 185 645 205 665
rect 185 605 205 625
rect 260 685 280 705
rect 260 645 280 665
rect 260 605 280 625
rect 335 685 355 705
rect 335 645 355 665
rect 335 605 355 625
rect 410 685 430 705
rect 410 645 430 665
rect 410 605 430 625
<< psubdiff >>
rect -150 120 690 135
rect -150 100 -140 120
rect -120 100 -100 120
rect -80 100 -60 120
rect -40 100 -20 120
rect 0 100 20 120
rect 40 100 60 120
rect 80 100 100 120
rect 120 100 140 120
rect 160 100 180 120
rect 200 100 220 120
rect 240 100 260 120
rect 280 100 300 120
rect 320 100 340 120
rect 360 100 380 120
rect 400 100 420 120
rect 440 100 460 120
rect 480 100 500 120
rect 520 100 540 120
rect 560 100 580 120
rect 600 100 620 120
rect 640 100 660 120
rect 680 100 690 120
rect -150 85 690 100
<< nsubdiff >>
rect -150 815 690 830
rect -150 795 -140 815
rect -120 795 -100 815
rect -80 795 -60 815
rect -40 795 -20 815
rect 0 795 20 815
rect 40 795 60 815
rect 80 795 100 815
rect 120 795 140 815
rect 160 795 180 815
rect 200 795 220 815
rect 240 795 260 815
rect 280 795 300 815
rect 320 795 340 815
rect 360 795 380 815
rect 400 795 420 815
rect 440 795 460 815
rect 480 795 500 815
rect 520 795 540 815
rect 560 795 580 815
rect 600 795 620 815
rect 640 795 660 815
rect 680 795 690 815
rect -150 780 690 795
<< psubdiffcont >>
rect -140 100 -120 120
rect -100 100 -80 120
rect -60 100 -40 120
rect -20 100 0 120
rect 20 100 40 120
rect 60 100 80 120
rect 100 100 120 120
rect 140 100 160 120
rect 180 100 200 120
rect 220 100 240 120
rect 260 100 280 120
rect 300 100 320 120
rect 340 100 360 120
rect 380 100 400 120
rect 420 100 440 120
rect 460 100 480 120
rect 500 100 520 120
rect 540 100 560 120
rect 580 100 600 120
rect 620 100 640 120
rect 660 100 680 120
<< nsubdiffcont >>
rect -140 795 -120 815
rect -100 795 -80 815
rect -60 795 -40 815
rect -20 795 0 815
rect 20 795 40 815
rect 60 795 80 815
rect 100 795 120 815
rect 140 795 160 815
rect 180 795 200 815
rect 220 795 240 815
rect 260 795 280 815
rect 300 795 320 815
rect 340 795 360 815
rect 380 795 400 815
rect 420 795 440 815
rect 460 795 480 815
rect 500 795 520 815
rect 540 795 560 815
rect 580 795 600 815
rect 620 795 640 815
rect 660 795 680 815
<< poly >>
rect 150 755 240 770
rect 150 740 165 755
rect 225 740 240 755
rect 300 755 390 770
rect 300 740 315 755
rect 375 740 390 755
rect 150 575 165 590
rect 225 515 240 590
rect 300 575 315 590
rect 375 575 390 590
rect 275 565 315 575
rect 275 545 285 565
rect 305 545 315 565
rect 275 535 315 545
rect 225 505 265 515
rect 225 485 235 505
rect 255 485 265 505
rect 225 475 265 485
rect -115 425 -75 435
rect -115 405 -105 425
rect -85 405 -75 425
rect -115 395 -75 405
rect -40 425 0 435
rect -40 405 -30 425
rect -10 405 0 425
rect -40 395 0 405
rect -90 355 -75 395
rect -15 355 0 395
rect 150 355 165 370
rect 225 355 240 475
rect 300 355 315 535
rect 590 455 630 465
rect 590 435 600 455
rect 620 435 630 455
rect 590 425 630 435
rect 530 405 570 415
rect 530 385 540 405
rect 560 385 570 405
rect 530 375 570 385
rect 375 355 390 370
rect 540 355 555 375
rect 615 355 630 425
rect -90 190 -75 205
rect -15 190 0 205
rect 150 190 165 205
rect 225 190 240 205
rect 300 190 315 205
rect 375 190 390 205
rect 540 190 555 205
rect 615 190 630 205
rect 150 180 190 190
rect 150 160 160 180
rect 180 160 190 180
rect 150 150 190 160
rect 350 180 390 190
rect 350 160 360 180
rect 380 160 390 180
rect 350 150 390 160
<< polycont >>
rect 285 545 305 565
rect 235 485 255 505
rect -105 405 -85 425
rect -30 405 -10 425
rect 600 435 620 455
rect 540 385 560 405
rect 160 160 180 180
rect 360 160 380 180
<< locali >>
rect -150 815 690 825
rect -150 795 -140 815
rect -120 795 -100 815
rect -80 795 -60 815
rect -40 795 -20 815
rect 0 795 20 815
rect 40 795 60 815
rect 80 795 100 815
rect 120 795 140 815
rect 160 795 180 815
rect 200 795 220 815
rect 240 795 260 815
rect 280 795 300 815
rect 320 795 340 815
rect 360 795 380 815
rect 400 795 420 815
rect 440 795 460 815
rect 480 795 500 815
rect 520 795 540 815
rect 560 795 580 815
rect 600 795 620 815
rect 640 795 660 815
rect 680 795 690 815
rect -150 785 690 795
rect 100 705 140 720
rect 100 685 110 705
rect 130 685 140 705
rect 100 665 140 685
rect 100 645 110 665
rect 130 645 140 665
rect 100 625 140 645
rect 100 605 110 625
rect 130 605 140 625
rect 100 595 140 605
rect 175 705 215 720
rect 175 685 185 705
rect 205 685 215 705
rect 175 665 215 685
rect 175 645 185 665
rect 205 645 215 665
rect 175 625 215 645
rect 175 605 185 625
rect 205 605 215 625
rect 175 590 215 605
rect 250 705 290 720
rect 250 685 260 705
rect 280 685 290 705
rect 250 665 290 685
rect 250 645 260 665
rect 280 645 290 665
rect 250 625 290 645
rect 250 605 260 625
rect 280 605 290 625
rect 250 595 290 605
rect 325 705 365 720
rect 325 685 335 705
rect 355 685 365 705
rect 325 665 365 685
rect 325 645 335 665
rect 355 645 365 665
rect 325 625 365 645
rect 325 605 335 625
rect 355 605 365 625
rect 325 590 365 605
rect 400 705 440 720
rect 400 685 410 705
rect 430 685 440 705
rect 400 665 440 685
rect 400 645 410 665
rect 430 645 440 665
rect 400 625 440 645
rect 400 605 410 625
rect 430 605 440 625
rect 400 595 440 605
rect 185 565 205 590
rect 275 565 315 575
rect -150 545 110 565
rect 70 535 110 545
rect 10 515 50 525
rect -150 495 20 515
rect 40 495 50 515
rect 70 515 80 535
rect 100 515 110 535
rect 70 505 110 515
rect 185 545 285 565
rect 305 545 315 565
rect 10 485 50 495
rect -150 455 -10 475
rect -30 435 -10 455
rect -115 425 -75 435
rect -150 405 -105 425
rect -85 405 -75 425
rect -115 395 -75 405
rect -40 425 0 435
rect -40 405 -30 425
rect -10 405 0 425
rect -40 395 0 405
rect 185 375 205 545
rect 275 535 315 545
rect 225 505 265 515
rect 335 505 355 590
rect 475 565 515 575
rect 475 545 485 565
rect 505 545 690 565
rect 475 535 515 545
rect 225 485 235 505
rect 255 485 690 505
rect 225 475 265 485
rect 335 375 355 485
rect 590 455 630 465
rect 590 435 600 455
rect 620 435 630 455
rect 590 425 630 435
rect 530 405 570 415
rect 530 385 540 405
rect 560 385 570 405
rect 530 375 570 385
rect -130 355 215 375
rect -130 335 -110 355
rect 20 335 40 355
rect -140 320 -100 335
rect -140 300 -130 320
rect -110 300 -100 320
rect -140 280 -100 300
rect -140 260 -130 280
rect -110 260 -100 280
rect -140 240 -100 260
rect -140 220 -130 240
rect -110 220 -100 240
rect -140 210 -100 220
rect -65 320 -25 335
rect -65 300 -55 320
rect -35 300 -25 320
rect -65 280 -25 300
rect -65 260 -55 280
rect -35 260 -25 280
rect -65 240 -25 260
rect -65 220 -55 240
rect -35 220 -25 240
rect -65 210 -25 220
rect 10 320 50 335
rect 10 300 20 320
rect 40 300 50 320
rect 10 280 50 300
rect 10 260 20 280
rect 40 260 50 280
rect 10 240 50 260
rect 10 220 20 240
rect 40 220 50 240
rect 10 210 50 220
rect 100 320 140 335
rect 100 300 110 320
rect 130 300 140 320
rect 100 280 140 300
rect 100 260 110 280
rect 130 260 140 280
rect 100 240 140 260
rect 100 220 110 240
rect 130 220 140 240
rect 100 210 140 220
rect 175 320 215 355
rect 325 355 510 375
rect 175 300 185 320
rect 205 300 215 320
rect 175 280 215 300
rect 175 260 185 280
rect 205 260 215 280
rect 175 240 215 260
rect 175 220 185 240
rect 205 220 215 240
rect 175 210 215 220
rect 250 320 290 335
rect 250 300 260 320
rect 280 300 290 320
rect 250 280 290 300
rect 250 260 260 280
rect 280 260 290 280
rect 250 240 290 260
rect 250 220 260 240
rect 280 220 290 240
rect 250 210 290 220
rect 325 320 365 355
rect 490 335 510 355
rect 325 300 335 320
rect 355 300 365 320
rect 325 280 365 300
rect 325 260 335 280
rect 355 260 365 280
rect 325 240 365 260
rect 325 220 335 240
rect 355 220 365 240
rect 325 210 365 220
rect 400 320 440 335
rect 400 300 410 320
rect 430 300 440 320
rect 400 280 440 300
rect 400 260 410 280
rect 430 260 440 280
rect 400 240 440 260
rect 400 220 410 240
rect 430 220 440 240
rect 400 210 440 220
rect 490 320 530 335
rect 490 300 500 320
rect 520 300 530 320
rect 490 280 530 300
rect 490 260 500 280
rect 520 260 530 280
rect 490 240 530 260
rect 490 220 500 240
rect 520 220 530 240
rect 490 210 530 220
rect 640 320 680 335
rect 640 300 650 320
rect 670 300 680 320
rect 640 280 680 300
rect 640 260 650 280
rect 670 260 680 280
rect 640 240 680 260
rect 640 220 650 240
rect 670 220 680 240
rect 640 210 680 220
rect 150 180 190 190
rect 350 180 390 190
rect -150 160 160 180
rect 180 160 360 180
rect 380 160 390 180
rect 150 150 190 160
rect 350 150 390 160
rect -150 120 690 130
rect -150 100 -140 120
rect -120 100 -100 120
rect -80 100 -60 120
rect -40 100 -20 120
rect 0 100 20 120
rect 40 100 60 120
rect 80 100 100 120
rect 120 100 140 120
rect 160 100 180 120
rect 200 100 220 120
rect 240 100 260 120
rect 280 100 300 120
rect 320 100 340 120
rect 360 100 380 120
rect 400 100 420 120
rect 440 100 460 120
rect 480 100 500 120
rect 520 100 540 120
rect 560 100 580 120
rect 600 100 620 120
rect 640 100 660 120
rect 680 100 690 120
rect -150 90 690 100
<< viali >>
rect -140 795 -120 815
rect -100 795 -80 815
rect -60 795 -40 815
rect -20 795 0 815
rect 20 795 40 815
rect 60 795 80 815
rect 100 795 120 815
rect 140 795 160 815
rect 180 795 200 815
rect 220 795 240 815
rect 260 795 280 815
rect 300 795 320 815
rect 340 795 360 815
rect 380 795 400 815
rect 420 795 440 815
rect 460 795 480 815
rect 500 795 520 815
rect 540 795 560 815
rect 580 795 600 815
rect 620 795 640 815
rect 660 795 680 815
rect 110 685 130 705
rect 110 645 130 665
rect 110 605 130 625
rect 260 685 280 705
rect 260 645 280 665
rect 260 605 280 625
rect 410 685 430 705
rect 410 645 430 665
rect 410 605 430 625
rect 20 495 40 515
rect 80 515 100 535
rect 285 545 305 565
rect 485 545 505 565
rect 600 435 620 455
rect 540 385 560 405
rect -55 300 -35 320
rect -55 260 -35 280
rect -55 220 -35 240
rect 110 300 130 320
rect 110 260 130 280
rect 110 220 130 240
rect 260 300 280 320
rect 260 260 280 280
rect 260 220 280 240
rect 410 300 430 320
rect 410 260 430 280
rect 410 220 430 240
rect 650 300 670 320
rect 650 260 670 280
rect 650 220 670 240
rect -140 100 -120 120
rect -100 100 -80 120
rect -60 100 -40 120
rect -20 100 0 120
rect 20 100 40 120
rect 60 100 80 120
rect 100 100 120 120
rect 140 100 160 120
rect 180 100 200 120
rect 220 100 240 120
rect 260 100 280 120
rect 300 100 320 120
rect 340 100 360 120
rect 380 100 400 120
rect 420 100 440 120
rect 460 100 480 120
rect 500 100 520 120
rect 540 100 560 120
rect 580 100 600 120
rect 620 100 640 120
rect 660 100 680 120
<< metal1 >>
rect -150 815 690 830
rect -150 795 -140 815
rect -120 795 -100 815
rect -80 795 -60 815
rect -40 795 -20 815
rect 0 795 20 815
rect 40 795 60 815
rect 80 795 100 815
rect 120 795 140 815
rect 160 795 180 815
rect 200 795 220 815
rect 240 795 260 815
rect 280 795 300 815
rect 320 795 340 815
rect 360 795 380 815
rect 400 795 420 815
rect 440 795 460 815
rect 480 795 500 815
rect 520 795 540 815
rect 560 795 580 815
rect 600 795 620 815
rect 640 795 660 815
rect 680 795 690 815
rect -150 780 690 795
rect -55 335 -35 780
rect 100 705 140 780
rect 100 685 110 705
rect 130 685 140 705
rect 100 665 140 685
rect 100 645 110 665
rect 130 645 140 665
rect 100 625 140 645
rect 100 605 110 625
rect 130 605 140 625
rect 100 595 140 605
rect 250 705 290 780
rect 250 685 260 705
rect 280 685 290 705
rect 250 665 290 685
rect 250 645 260 665
rect 280 645 290 665
rect 250 625 290 645
rect 250 605 260 625
rect 280 605 290 625
rect 250 595 290 605
rect 400 705 440 780
rect 400 685 410 705
rect 430 685 440 705
rect 400 665 440 685
rect 400 645 410 665
rect 430 645 440 665
rect 400 625 440 645
rect 400 605 410 625
rect 430 605 440 625
rect 400 595 440 605
rect 275 565 315 575
rect 475 565 515 575
rect 275 545 285 565
rect 305 545 485 565
rect 505 545 515 565
rect 70 535 110 545
rect 275 535 315 545
rect 475 535 515 545
rect 10 515 50 525
rect 10 495 20 515
rect 40 495 50 515
rect 70 515 80 535
rect 100 515 110 535
rect 70 505 110 515
rect 10 485 50 495
rect 20 405 40 485
rect 80 455 100 505
rect 590 455 630 465
rect 80 435 600 455
rect 620 435 630 455
rect 590 425 630 435
rect 530 405 570 415
rect 20 385 540 405
rect 560 385 570 405
rect 530 375 570 385
rect 650 335 670 780
rect -65 320 -25 335
rect -65 300 -55 320
rect -35 300 -25 320
rect -65 280 -25 300
rect -65 260 -55 280
rect -35 260 -25 280
rect -65 240 -25 260
rect -65 220 -55 240
rect -35 220 -25 240
rect -65 210 -25 220
rect 100 320 140 335
rect 100 300 110 320
rect 130 300 140 320
rect 100 280 140 300
rect 100 260 110 280
rect 130 260 140 280
rect 100 240 140 260
rect 100 220 110 240
rect 130 220 140 240
rect 100 210 140 220
rect 250 320 290 335
rect 250 300 260 320
rect 280 300 290 320
rect 250 280 290 300
rect 250 260 260 280
rect 280 260 290 280
rect 250 240 290 260
rect 250 220 260 240
rect 280 220 290 240
rect 250 210 290 220
rect 400 320 440 335
rect 400 300 410 320
rect 430 300 440 320
rect 400 280 440 300
rect 400 260 410 280
rect 430 260 440 280
rect 400 240 440 260
rect 400 220 410 240
rect 430 220 440 240
rect 400 210 440 220
rect 640 320 680 335
rect 640 300 650 320
rect 670 300 680 320
rect 640 280 680 300
rect 640 260 650 280
rect 670 260 680 280
rect 640 240 680 260
rect 640 220 650 240
rect 670 220 680 240
rect 640 210 680 220
rect 110 135 130 210
rect 260 135 280 210
rect 410 135 430 210
rect -150 120 690 135
rect -150 100 -140 120
rect -120 100 -100 120
rect -80 100 -60 120
rect -40 100 -20 120
rect 0 100 20 120
rect 40 100 60 120
rect 80 100 100 120
rect 120 100 140 120
rect 160 100 180 120
rect 200 100 220 120
rect 240 100 260 120
rect 280 100 300 120
rect 320 100 340 120
rect 360 100 380 120
rect 400 100 420 120
rect 440 100 460 120
rect 480 100 500 120
rect 520 100 540 120
rect 560 100 580 120
rect 600 100 620 120
rect 640 100 660 120
rect 680 100 690 120
rect -150 85 690 100
<< labels >>
rlabel locali -145 550 -135 560 7 A
port 1 w
rlabel locali -145 500 -135 510 7 B
port 3 w
rlabel locali -145 410 -135 420 7 B_bar
port 4 w
rlabel locali -145 460 -135 470 7 A_bar
port 2 w
rlabel viali 285 545 305 565 7 OUT_bar
port 6 w
rlabel locali 235 485 255 505 7 OUT
port 5 w
rlabel locali 160 160 180 180 7 Dis
port 7 w
rlabel metal1 260 795 280 815 7 CLK
port 9 w
rlabel metal1 260 100 280 120 7 GND!
port 8 w
<< end >>
