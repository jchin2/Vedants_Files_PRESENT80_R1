magic
tech sky130A
timestamp 1676417541
<< nwell >>
rect -695 250 -175 595
<< nmos >>
rect -615 45 -600 195
rect -540 45 -525 195
rect -465 45 -450 195
rect -270 45 -255 195
<< pmos >>
rect -615 275 -600 575
rect -540 275 -525 575
rect -465 275 -450 575
rect -270 275 -255 575
<< ndiff >>
rect -675 180 -615 195
rect -675 60 -655 180
rect -635 60 -615 180
rect -675 45 -615 60
rect -600 45 -540 195
rect -525 45 -465 195
rect -450 180 -390 195
rect -450 60 -430 180
rect -410 60 -390 180
rect -450 45 -390 60
rect -330 180 -270 195
rect -330 60 -310 180
rect -290 60 -270 180
rect -330 45 -270 60
rect -255 180 -195 195
rect -255 60 -235 180
rect -215 60 -195 180
rect -255 45 -195 60
<< pdiff >>
rect -675 560 -615 575
rect -675 290 -655 560
rect -635 290 -615 560
rect -675 275 -615 290
rect -600 560 -540 575
rect -600 290 -580 560
rect -560 290 -540 560
rect -600 275 -540 290
rect -525 560 -465 575
rect -525 290 -505 560
rect -485 290 -465 560
rect -525 275 -465 290
rect -450 560 -390 575
rect -450 290 -430 560
rect -410 290 -390 560
rect -450 275 -390 290
rect -330 560 -270 575
rect -330 290 -310 560
rect -290 290 -270 560
rect -330 275 -270 290
rect -255 555 -195 575
rect -255 295 -235 555
rect -215 295 -195 555
rect -255 275 -195 295
<< ndiffc >>
rect -655 60 -635 180
rect -430 60 -410 180
rect -310 60 -290 180
rect -235 60 -215 180
<< pdiffc >>
rect -655 290 -635 560
rect -580 290 -560 560
rect -505 290 -485 560
rect -430 290 -410 560
rect -310 290 -290 560
rect -235 295 -215 555
<< poly >>
rect -615 575 -600 590
rect -540 575 -525 590
rect -465 575 -450 590
rect -270 575 -255 590
rect -615 255 -600 275
rect -640 245 -600 255
rect -640 225 -630 245
rect -610 225 -600 245
rect -640 215 -600 225
rect -615 195 -600 215
rect -540 195 -525 275
rect -465 195 -450 275
rect -270 260 -255 275
rect -310 250 -255 260
rect -310 230 -300 250
rect -280 230 -255 250
rect -310 220 -255 230
rect -270 195 -255 220
rect -615 30 -600 45
rect -540 30 -525 45
rect -565 20 -525 30
rect -565 0 -555 20
rect -535 0 -525 20
rect -565 -10 -525 0
rect -465 -20 -450 45
rect -270 30 -255 45
rect -480 -30 -440 -20
rect -480 -50 -470 -30
rect -450 -50 -440 -30
rect -480 -60 -440 -50
<< polycont >>
rect -630 225 -610 245
rect -300 230 -280 250
rect -555 0 -535 20
rect -470 -50 -450 -30
<< locali >>
rect -655 585 -485 605
rect -655 565 -635 585
rect -505 565 -485 585
rect -665 560 -625 565
rect -665 290 -655 560
rect -635 290 -625 560
rect -665 285 -625 290
rect -590 560 -550 565
rect -590 290 -580 560
rect -560 290 -550 560
rect -590 285 -550 290
rect -515 560 -475 565
rect -515 290 -505 560
rect -485 290 -475 560
rect -515 285 -475 290
rect -440 560 -400 565
rect -440 290 -430 560
rect -410 290 -400 560
rect -440 285 -400 290
rect -320 560 -280 565
rect -320 290 -310 560
rect -290 290 -280 560
rect -320 285 -280 290
rect -245 555 -205 565
rect -245 295 -235 555
rect -215 295 -205 555
rect -245 285 -205 295
rect -640 245 -600 255
rect -640 225 -630 245
rect -610 225 -600 245
rect -505 250 -485 285
rect -310 250 -270 260
rect -505 230 -300 250
rect -280 230 -270 250
rect -640 215 -600 225
rect -430 185 -410 230
rect -310 220 -270 230
rect -235 185 -215 285
rect -665 180 -625 185
rect -665 60 -655 180
rect -635 60 -625 180
rect -665 55 -625 60
rect -440 180 -400 185
rect -440 60 -430 180
rect -410 60 -400 180
rect -440 55 -400 60
rect -320 180 -280 185
rect -320 60 -310 180
rect -290 60 -280 180
rect -320 55 -280 60
rect -245 180 -205 185
rect -245 60 -235 180
rect -215 60 -205 180
rect -245 55 -205 60
rect -565 20 -525 30
rect -565 0 -555 20
rect -535 0 -525 20
rect -565 -10 -525 0
rect -480 -30 -440 -20
rect -480 -50 -470 -30
rect -450 -50 -440 -30
rect -480 -60 -440 -50
<< viali >>
rect -580 290 -560 560
rect -430 290 -410 560
rect -310 290 -290 560
rect -655 60 -635 180
rect -310 60 -290 180
<< metal1 >>
rect -590 560 -550 565
rect -590 290 -580 560
rect -560 290 -550 560
rect -590 285 -550 290
rect -440 560 -400 565
rect -440 290 -430 560
rect -410 290 -400 560
rect -440 285 -400 290
rect -320 560 -280 565
rect -320 290 -310 560
rect -290 290 -280 560
rect -320 285 -280 290
rect -665 180 -625 185
rect -665 60 -655 180
rect -635 60 -625 180
rect -665 55 -625 60
rect -320 180 -280 185
rect -320 60 -310 180
rect -290 60 -280 180
rect -320 55 -280 60
<< end >>
