magic
tech sky130A
timestamp 1670967604
<< error_p >>
rect 192 582 200 585
rect 201 582 209 585
rect 184 569 187 577
rect 214 569 217 577
rect 184 560 187 568
rect 214 560 217 568
rect 192 552 200 555
rect 201 552 209 555
<< poly >>
rect 187 577 214 582
rect 187 560 192 577
rect 209 560 214 577
rect 187 555 214 560
<< polycont >>
rect 192 560 209 577
<< locali >>
rect 184 577 217 585
rect 184 560 192 577
rect 209 560 217 577
rect 184 552 217 560
<< end >>
