* NGSPICE file created from EESPFAL_XOR_v3_flat.ext - technology: sky130A

.subckt EESPFAL_XOR_v3_flat OUT A A_bar B B_bar Dis OUT_bar GND CLK
X0 CLK.t7 OUT.t6 OUT_bar.t1 CLK.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 OUT_bar.t5 Dis.t0 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n840_410# A.t0 CLK.t9 GND.t13 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n1140_410# B_bar.t0 OUT_bar.t3 GND.t9 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_420_410# B_bar.t1 OUT.t3 GND.t8 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 GND.t1 Dis.t1 OUT.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 OUT.t5 OUT_bar.t6 CLK.t3 CLK.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_720_410# A_bar.t0 CLK.t11 GND.t15 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar.t2 OUT.t7 CLK.t5 CLK.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 CLK.t1 OUT_bar.t7 OUT.t0 CLK.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 OUT_bar.t4 B.t0 a_n840_410# GND.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 GND.t7 OUT.t8 OUT_bar.t0 GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK.t10 A_bar.t1 a_n1140_410# GND.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 OUT.t2 OUT_bar.t8 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 CLK.t8 A.t1 a_420_410# GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 OUT.t4 B.t1 a_720_410# GND.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
R0 OUT.t6 OUT.t7 819.4
R1 OUT.n4 OUT.t6 514.133
R2 OUT.n4 OUT.t8 305.266
R3 OUT.n2 OUT.t4 289.936
R4 OUT.n3 OUT.n0 166.734
R5 OUT.n3 OUT.n2 105.6
R6 OUT.n2 OUT.t3 97.937
R7 OUT.n5 OUT.n4 76
R8 OUT.n3 OUT.n1 73.937
R9 OUT.n5 OUT.n3 57.6
R10 OUT.n0 OUT.t0 39.4
R11 OUT.n0 OUT.t5 39.4
R12 OUT.n1 OUT.t1 24
R13 OUT.n1 OUT.t2 24
R14 OUT OUT.n5 3.2
R15 OUT_bar.t6 OUT_bar.t7 819.4
R16 OUT_bar.n0 OUT_bar.t8 506.1
R17 OUT_bar.n0 OUT_bar.t6 313.3
R18 OUT_bar.n3 OUT_bar.t3 273.936
R19 OUT_bar.n5 OUT_bar.n1 128.334
R20 OUT_bar.n4 OUT_bar.n3 105.6
R21 OUT_bar.n3 OUT_bar.t4 81.937
R22 OUT_bar.n4 OUT_bar.n2 57.937
R23 OUT_bar.n6 OUT_bar.n5 57.6
R24 OUT_bar.n5 OUT_bar.n4 41.6
R25 OUT_bar.n1 OUT_bar.t1 39.4
R26 OUT_bar.n1 OUT_bar.t2 39.4
R27 OUT_bar.n2 OUT_bar.t0 24
R28 OUT_bar.n2 OUT_bar.t5 24
R29 OUT_bar.n6 OUT_bar.n0 8.764
R30 OUT_bar OUT_bar.n6 4.681
R31 CLK.n94 CLK.t5 44.337
R32 CLK.n39 CLK.t1 44.337
R33 CLK.n0 CLK.t3 39.4
R34 CLK.n0 CLK.t7 39.4
R35 CLK.n40 CLK.t0 24.568
R36 CLK.n95 CLK.t4 24.568
R37 CLK.n56 CLK.t9 24
R38 CLK.n56 CLK.t10 24
R39 CLK.n1 CLK.t11 24
R40 CLK.n1 CLK.t8 24
R41 CLK.n4 CLK.n3 8.855
R42 CLK.n8 CLK.n7 8.855
R43 CLK.n7 CLK.n6 8.855
R44 CLK.n12 CLK.n11 8.855
R45 CLK.n11 CLK.n10 8.855
R46 CLK.n17 CLK.n16 8.855
R47 CLK.n16 CLK.n15 8.855
R48 CLK.n21 CLK.n20 8.855
R49 CLK.n20 CLK.n19 8.855
R50 CLK.n25 CLK.n24 8.855
R51 CLK.n24 CLK.n23 8.855
R52 CLK.n29 CLK.n28 8.855
R53 CLK.n28 CLK.n27 8.855
R54 CLK.n33 CLK.n32 8.855
R55 CLK.n32 CLK.n31 8.855
R56 CLK.n37 CLK.n36 8.855
R57 CLK.n36 CLK.n35 8.855
R58 CLK.n42 CLK.n41 8.855
R59 CLK.n41 CLK.n40 8.855
R60 CLK.n46 CLK.n45 8.855
R61 CLK.n45 CLK.n44 8.855
R62 CLK.n50 CLK.n49 8.855
R63 CLK.n49 CLK.n48 8.855
R64 CLK.n54 CLK.n53 8.855
R65 CLK.n53 CLK.n52 8.855
R66 CLK.n105 CLK.n104 8.855
R67 CLK.n104 CLK.n103 8.855
R68 CLK.n101 CLK.n100 8.855
R69 CLK.n100 CLK.n99 8.855
R70 CLK.n97 CLK.n96 8.855
R71 CLK.n96 CLK.n95 8.855
R72 CLK.n92 CLK.n91 8.855
R73 CLK.n91 CLK.n90 8.855
R74 CLK.n88 CLK.n87 8.855
R75 CLK.n87 CLK.n86 8.855
R76 CLK.n84 CLK.n83 8.855
R77 CLK.n83 CLK.n82 8.855
R78 CLK.n80 CLK.n79 8.855
R79 CLK.n79 CLK.n78 8.855
R80 CLK.n76 CLK.n75 8.855
R81 CLK.n75 CLK.n74 8.855
R82 CLK.n72 CLK.n71 8.855
R83 CLK.n71 CLK.n70 8.855
R84 CLK.n67 CLK.n66 8.855
R85 CLK.n66 CLK.n65 8.855
R86 CLK.n63 CLK.n62 8.855
R87 CLK.n62 CLK.n61 8.855
R88 CLK.n59 CLK.n58 8.855
R89 CLK.n48 CLK.t2 8.189
R90 CLK.n103 CLK.t6 8.189
R91 CLK.n69 CLK.n56 6.776
R92 CLK.n14 CLK.n1 6.776
R93 CLK.n55 CLK.n0 4.938
R94 CLK.n9 CLK.n8 4.65
R95 CLK.n13 CLK.n12 4.65
R96 CLK.n18 CLK.n17 4.65
R97 CLK.n22 CLK.n21 4.65
R98 CLK.n26 CLK.n25 4.65
R99 CLK.n30 CLK.n29 4.65
R100 CLK.n34 CLK.n33 4.65
R101 CLK.n38 CLK.n37 4.65
R102 CLK.n43 CLK.n42 4.65
R103 CLK.n47 CLK.n46 4.65
R104 CLK.n51 CLK.n50 4.65
R105 CLK.n55 CLK.n54 4.65
R106 CLK.n106 CLK.n105 4.65
R107 CLK.n102 CLK.n101 4.65
R108 CLK.n98 CLK.n97 4.65
R109 CLK.n93 CLK.n92 4.65
R110 CLK.n89 CLK.n88 4.65
R111 CLK.n85 CLK.n84 4.65
R112 CLK.n81 CLK.n80 4.65
R113 CLK.n77 CLK.n76 4.65
R114 CLK.n73 CLK.n72 4.65
R115 CLK.n68 CLK.n67 4.65
R116 CLK.n64 CLK.n63 4.65
R117 CLK.n5 CLK.n4 2.682
R118 CLK.n60 CLK.n59 2.682
R119 CLK.n3 CLK.n2 1.655
R120 CLK.n58 CLK.n57 1.655
R121 CLK.n9 CLK.n5 1.096
R122 CLK.n64 CLK.n60 1.095
R123 CLK.n13 CLK.n9 0.1
R124 CLK.n22 CLK.n18 0.1
R125 CLK.n26 CLK.n22 0.1
R126 CLK.n30 CLK.n26 0.1
R127 CLK.n34 CLK.n30 0.1
R128 CLK.n38 CLK.n34 0.1
R129 CLK.n47 CLK.n43 0.1
R130 CLK.n51 CLK.n47 0.1
R131 CLK.n55 CLK.n51 0.1
R132 CLK.n106 CLK.n102 0.1
R133 CLK.n102 CLK.n98 0.1
R134 CLK.n93 CLK.n89 0.1
R135 CLK.n89 CLK.n85 0.1
R136 CLK.n85 CLK.n81 0.1
R137 CLK.n81 CLK.n77 0.1
R138 CLK.n77 CLK.n73 0.1
R139 CLK.n68 CLK.n64 0.1
R140 CLK.n18 CLK.n14 0.075
R141 CLK.n43 CLK.n39 0.075
R142 CLK CLK.n106 0.075
R143 CLK.n98 CLK.n94 0.075
R144 CLK.n73 CLK.n69 0.075
R145 CLK.n14 CLK.n13 0.025
R146 CLK.n39 CLK.n38 0.025
R147 CLK CLK.n55 0.025
R148 CLK.n94 CLK.n93 0.025
R149 CLK.n69 CLK.n68 0.025
R150 Dis.n0 Dis.t1 504.5
R151 Dis.n0 Dis.t0 389.3
R152 Dis Dis.n0 3.2
R153 GND.n1 GND.t10 269.289
R154 GND.n55 GND.t9 269.289
R155 GND.n6 GND.t15 185.81
R156 GND.n60 GND.t14 185.81
R157 GND.n14 GND.t12 111.486
R158 GND.n39 GND.t0 111.486
R159 GND.n93 GND.t2 111.486
R160 GND.n68 GND.t13 111.486
R161 GND.n22 GND.t8 37.162
R162 GND.n47 GND.t4 37.162
R163 GND.n101 GND.t6 37.162
R164 GND.n76 GND.t11 37.162
R165 GND.n38 GND.t1 29.103
R166 GND.n92 GND.t3 29.103
R167 GND.n0 GND.t5 24
R168 GND.n0 GND.t7 24
R169 GND.n59 GND.n55 11.894
R170 GND.n5 GND.n1 11.894
R171 GND.n4 GND.n3 9.154
R172 GND.n3 GND.n2 9.154
R173 GND.n8 GND.n7 9.154
R174 GND.n7 GND.n6 9.154
R175 GND.n12 GND.n11 9.154
R176 GND.n11 GND.n10 9.154
R177 GND.n16 GND.n15 9.154
R178 GND.n15 GND.n14 9.154
R179 GND.n20 GND.n19 9.154
R180 GND.n19 GND.n18 9.154
R181 GND.n24 GND.n23 9.154
R182 GND.n23 GND.n22 9.154
R183 GND.n28 GND.n27 9.154
R184 GND.n27 GND.n26 9.154
R185 GND.n32 GND.n31 9.154
R186 GND.n31 GND.n30 9.154
R187 GND.n36 GND.n35 9.154
R188 GND.n35 GND.n34 9.154
R189 GND.n41 GND.n40 9.154
R190 GND.n40 GND.n39 9.154
R191 GND.n45 GND.n44 9.154
R192 GND.n44 GND.n43 9.154
R193 GND.n49 GND.n48 9.154
R194 GND.n48 GND.n47 9.154
R195 GND.n53 GND.n52 9.154
R196 GND.n52 GND.n51 9.154
R197 GND.n103 GND.n102 9.154
R198 GND.n102 GND.n101 9.154
R199 GND.n99 GND.n98 9.154
R200 GND.n98 GND.n97 9.154
R201 GND.n95 GND.n94 9.154
R202 GND.n94 GND.n93 9.154
R203 GND.n90 GND.n89 9.154
R204 GND.n89 GND.n88 9.154
R205 GND.n86 GND.n85 9.154
R206 GND.n85 GND.n84 9.154
R207 GND.n82 GND.n81 9.154
R208 GND.n81 GND.n80 9.154
R209 GND.n78 GND.n77 9.154
R210 GND.n77 GND.n76 9.154
R211 GND.n74 GND.n73 9.154
R212 GND.n73 GND.n72 9.154
R213 GND.n70 GND.n69 9.154
R214 GND.n69 GND.n68 9.154
R215 GND.n66 GND.n65 9.154
R216 GND.n65 GND.n64 9.154
R217 GND.n62 GND.n61 9.154
R218 GND.n61 GND.n60 9.154
R219 GND.n58 GND.n57 9.154
R220 GND.n57 GND.n56 9.154
R221 GND.n54 GND.n0 5.103
R222 GND.n9 GND.n8 4.65
R223 GND.n13 GND.n12 4.65
R224 GND.n17 GND.n16 4.65
R225 GND.n21 GND.n20 4.65
R226 GND.n25 GND.n24 4.65
R227 GND.n29 GND.n28 4.65
R228 GND.n33 GND.n32 4.65
R229 GND.n37 GND.n36 4.65
R230 GND.n42 GND.n41 4.65
R231 GND.n46 GND.n45 4.65
R232 GND.n50 GND.n49 4.65
R233 GND.n54 GND.n53 4.65
R234 GND.n104 GND.n103 4.65
R235 GND.n100 GND.n99 4.65
R236 GND.n96 GND.n95 4.65
R237 GND.n91 GND.n90 4.65
R238 GND.n87 GND.n86 4.65
R239 GND.n83 GND.n82 4.65
R240 GND.n79 GND.n78 4.65
R241 GND.n75 GND.n74 4.65
R242 GND.n71 GND.n70 4.65
R243 GND.n67 GND.n66 4.65
R244 GND.n63 GND.n62 4.65
R245 GND.n5 GND.n4 2.682
R246 GND.n59 GND.n58 2.682
R247 GND.n9 GND.n5 1.095
R248 GND.n63 GND.n59 1.095
R249 GND.n13 GND.n9 0.1
R250 GND.n17 GND.n13 0.1
R251 GND.n21 GND.n17 0.1
R252 GND.n25 GND.n21 0.1
R253 GND.n29 GND.n25 0.1
R254 GND.n33 GND.n29 0.1
R255 GND.n37 GND.n33 0.1
R256 GND.n46 GND.n42 0.1
R257 GND.n50 GND.n46 0.1
R258 GND.n54 GND.n50 0.1
R259 GND.n104 GND.n100 0.1
R260 GND.n100 GND.n96 0.1
R261 GND.n91 GND.n87 0.1
R262 GND.n87 GND.n83 0.1
R263 GND.n83 GND.n79 0.1
R264 GND.n79 GND.n75 0.1
R265 GND.n75 GND.n71 0.1
R266 GND.n71 GND.n67 0.1
R267 GND.n67 GND.n63 0.1
R268 GND.n42 GND.n38 0.075
R269 GND GND.n104 0.075
R270 GND.n96 GND.n92 0.075
R271 GND.n38 GND.n37 0.025
R272 GND GND.n54 0.025
R273 GND.n92 GND.n91 0.025
R274 A.n0 A.t0 1176.57
R275 A.n0 A.t1 1149.49
R276 A A.n0 128
R277 B_bar.n0 B_bar.t1 810.772
R278 B_bar.n0 B_bar.t0 694.566
R279 B_bar B_bar.n0 25.6
R280 A_bar.n0 A_bar.t0 1069.04
R281 A_bar.n0 A_bar.t1 1015.9
R282 A_bar A_bar.n0 89.6
R283 B.n0 B.t1 800.452
R284 B.n0 B.t0 787.997
R285 B B.n0 169.6
C0 CLK OUT_bar 0.98fF
C1 B A 0.15fF
C2 OUT_bar A_bar 0.05fF
C3 a_n1140_410# B_bar 0.00fF
C4 a_n1140_410# OUT_bar 0.01fF
C5 CLK OUT 0.65fF
C6 OUT_bar B_bar 0.30fF
C7 OUT A_bar 0.03fF
C8 a_n840_410# A 0.00fF
C9 a_420_410# A 0.00fF
C10 a_n1140_410# OUT 0.00fF
C11 CLK Dis 0.14fF
C12 Dis A_bar 0.00fF
C13 OUT B_bar 0.07fF
C14 CLK B 0.32fF
C15 B A_bar 1.50fF
C16 OUT_bar OUT 0.78fF
C17 a_n1140_410# Dis 0.00fF
C18 B a_n1140_410# 0.00fF
C19 CLK a_720_410# 0.02fF
C20 Dis B_bar 0.02fF
C21 a_720_410# A_bar 0.00fF
C22 B B_bar 1.24fF
C23 CLK a_n840_410# 0.01fF
C24 OUT_bar Dis 0.25fF
C25 CLK a_420_410# 0.01fF
C26 A_bar a_n840_410# 0.00fF
C27 a_420_410# A_bar 0.00fF
C28 CLK A 1.11fF
C29 B OUT_bar 0.07fF
C30 A_bar A 1.51fF
C31 a_n1140_410# A 0.00fF
C32 Dis OUT 0.08fF
C33 a_720_410# OUT_bar 0.00fF
C34 a_n840_410# B_bar 0.00fF
C35 a_420_410# B_bar 0.00fF
C36 B OUT 0.05fF
C37 A B_bar 0.06fF
C38 OUT_bar a_n840_410# 0.01fF
C39 OUT_bar a_420_410# 0.00fF
C40 OUT_bar A 0.05fF
C41 a_720_410# OUT 0.01fF
C42 B Dis 0.01fF
C43 OUT a_n840_410# 0.00fF
C44 CLK A_bar 0.48fF
C45 OUT a_420_410# 0.01fF
C46 OUT A 0.03fF
C47 CLK a_n1140_410# 0.02fF
C48 a_n1140_410# A_bar 0.00fF
C49 a_720_410# B 0.00fF
C50 Dis a_n840_410# 0.00fF
C51 CLK B_bar 0.24fF
C52 B a_n840_410# 0.00fF
C53 Dis A 0.01fF
C54 A_bar B_bar 0.10fF
C55 B a_420_410# 0.00fF
.ends

