* NGSPICE file created from INV_sanity_check.ext - technology: sky130A

.subckt INV_sanity_check B C D A
X0 C B D D sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X1 C B A A sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
.ends

