* NGSPICE file created from EESPFAL_4in_Buffer.ext - technology: sky130A

.subckt EESPFAL_INV4 A A_bar OUT OUT_bar Dis GND CLK
X0 OUT A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=5.25e+12p ps=2.32e+07u w=1.5e+06u l=150000u
X1 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X2 GND Dis OUT_bar GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X3 GND OUT_bar OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X5 OUT_bar OUT GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 CLK A OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT Dis GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_4in_Buffer A A_bar B B_bar C C_bar D D_bar OUT0 OUT0_bar OUT1 OUT1_bar
+ OUT2 OUT2_bar OUT3 OUT3_bar Dis GND CLK
XEESPFAL_INV4_0 A A_bar OUT0 OUT0_bar Dis GND CLK EESPFAL_INV4
XEESPFAL_INV4_1 B B_bar OUT1 OUT1_bar Dis GND CLK EESPFAL_INV4
XEESPFAL_INV4_2 C C_bar OUT2 OUT2_bar Dis GND CLK EESPFAL_INV4
XEESPFAL_INV4_3 D D_bar OUT3 OUT3_bar Dis GND CLK EESPFAL_INV4
.ends

