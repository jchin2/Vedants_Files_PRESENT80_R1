magic
tech sky130A
magscale 1 2
timestamp 1671306811
<< metal3 >>
rect -1355 1272 1354 1305
rect -1355 1208 1270 1272
rect 1334 1208 1354 1272
rect -1355 1192 1354 1208
rect -1355 1128 1270 1192
rect 1334 1128 1354 1192
rect -1355 1112 1354 1128
rect -1355 1048 1270 1112
rect 1334 1048 1354 1112
rect -1355 1032 1354 1048
rect -1355 968 1270 1032
rect 1334 968 1354 1032
rect -1355 952 1354 968
rect -1355 888 1270 952
rect 1334 888 1354 952
rect -1355 872 1354 888
rect -1355 808 1270 872
rect 1334 808 1354 872
rect -1355 792 1354 808
rect -1355 728 1270 792
rect 1334 728 1354 792
rect -1355 712 1354 728
rect -1355 648 1270 712
rect 1334 648 1354 712
rect -1355 632 1354 648
rect -1355 568 1270 632
rect 1334 568 1354 632
rect -1355 552 1354 568
rect -1355 488 1270 552
rect 1334 488 1354 552
rect -1355 472 1354 488
rect -1355 408 1270 472
rect 1334 408 1354 472
rect -1355 392 1354 408
rect -1355 328 1270 392
rect 1334 328 1354 392
rect -1355 312 1354 328
rect -1355 248 1270 312
rect 1334 248 1354 312
rect -1355 232 1354 248
rect -1355 168 1270 232
rect 1334 168 1354 232
rect -1355 152 1354 168
rect -1355 88 1270 152
rect 1334 88 1354 152
rect -1355 72 1354 88
rect -1355 8 1270 72
rect 1334 8 1354 72
rect -1355 -8 1354 8
rect -1355 -72 1270 -8
rect 1334 -72 1354 -8
rect -1355 -88 1354 -72
rect -1355 -152 1270 -88
rect 1334 -152 1354 -88
rect -1355 -168 1354 -152
rect -1355 -232 1270 -168
rect 1334 -232 1354 -168
rect -1355 -248 1354 -232
rect -1355 -312 1270 -248
rect 1334 -312 1354 -248
rect -1355 -328 1354 -312
rect -1355 -392 1270 -328
rect 1334 -392 1354 -328
rect -1355 -408 1354 -392
rect -1355 -472 1270 -408
rect 1334 -472 1354 -408
rect -1355 -488 1354 -472
rect -1355 -552 1270 -488
rect 1334 -552 1354 -488
rect -1355 -568 1354 -552
rect -1355 -632 1270 -568
rect 1334 -632 1354 -568
rect -1355 -648 1354 -632
rect -1355 -712 1270 -648
rect 1334 -712 1354 -648
rect -1355 -728 1354 -712
rect -1355 -792 1270 -728
rect 1334 -792 1354 -728
rect -1355 -808 1354 -792
rect -1355 -872 1270 -808
rect 1334 -872 1354 -808
rect -1355 -888 1354 -872
rect -1355 -952 1270 -888
rect 1334 -952 1354 -888
rect -1355 -968 1354 -952
rect -1355 -1032 1270 -968
rect 1334 -1032 1354 -968
rect -1355 -1048 1354 -1032
rect -1355 -1112 1270 -1048
rect 1334 -1112 1354 -1048
rect -1355 -1128 1354 -1112
rect -1355 -1192 1270 -1128
rect 1334 -1192 1354 -1128
rect -1355 -1208 1354 -1192
rect -1355 -1272 1270 -1208
rect 1334 -1272 1354 -1208
rect -1355 -1305 1354 -1272
<< via3 >>
rect 1270 1208 1334 1272
rect 1270 1128 1334 1192
rect 1270 1048 1334 1112
rect 1270 968 1334 1032
rect 1270 888 1334 952
rect 1270 808 1334 872
rect 1270 728 1334 792
rect 1270 648 1334 712
rect 1270 568 1334 632
rect 1270 488 1334 552
rect 1270 408 1334 472
rect 1270 328 1334 392
rect 1270 248 1334 312
rect 1270 168 1334 232
rect 1270 88 1334 152
rect 1270 8 1334 72
rect 1270 -72 1334 -8
rect 1270 -152 1334 -88
rect 1270 -232 1334 -168
rect 1270 -312 1334 -248
rect 1270 -392 1334 -328
rect 1270 -472 1334 -408
rect 1270 -552 1334 -488
rect 1270 -632 1334 -568
rect 1270 -712 1334 -648
rect 1270 -792 1334 -728
rect 1270 -872 1334 -808
rect 1270 -952 1334 -888
rect 1270 -1032 1334 -968
rect 1270 -1112 1334 -1048
rect 1270 -1192 1334 -1128
rect 1270 -1272 1334 -1208
<< mimcap >>
rect -1255 1152 1155 1205
rect -1255 -1152 -1202 1152
rect 1102 -1152 1155 1152
rect -1255 -1205 1155 -1152
<< mimcapcontact >>
rect -1202 -1152 1102 1152
<< metal4 >>
rect 1254 1272 1350 1293
rect 1254 1208 1270 1272
rect 1334 1208 1350 1272
rect 1254 1192 1350 1208
rect -1216 1152 1116 1166
rect -1216 -1152 -1202 1152
rect 1102 -1152 1116 1152
rect -1216 -1166 1116 -1152
rect 1254 1128 1270 1192
rect 1334 1128 1350 1192
rect 1254 1112 1350 1128
rect 1254 1048 1270 1112
rect 1334 1048 1350 1112
rect 1254 1032 1350 1048
rect 1254 968 1270 1032
rect 1334 968 1350 1032
rect 1254 952 1350 968
rect 1254 888 1270 952
rect 1334 888 1350 952
rect 1254 872 1350 888
rect 1254 808 1270 872
rect 1334 808 1350 872
rect 1254 792 1350 808
rect 1254 728 1270 792
rect 1334 728 1350 792
rect 1254 712 1350 728
rect 1254 648 1270 712
rect 1334 648 1350 712
rect 1254 632 1350 648
rect 1254 568 1270 632
rect 1334 568 1350 632
rect 1254 552 1350 568
rect 1254 488 1270 552
rect 1334 488 1350 552
rect 1254 472 1350 488
rect 1254 408 1270 472
rect 1334 408 1350 472
rect 1254 392 1350 408
rect 1254 328 1270 392
rect 1334 328 1350 392
rect 1254 312 1350 328
rect 1254 248 1270 312
rect 1334 248 1350 312
rect 1254 232 1350 248
rect 1254 168 1270 232
rect 1334 168 1350 232
rect 1254 152 1350 168
rect 1254 88 1270 152
rect 1334 88 1350 152
rect 1254 72 1350 88
rect 1254 8 1270 72
rect 1334 8 1350 72
rect 1254 -8 1350 8
rect 1254 -72 1270 -8
rect 1334 -72 1350 -8
rect 1254 -88 1350 -72
rect 1254 -152 1270 -88
rect 1334 -152 1350 -88
rect 1254 -168 1350 -152
rect 1254 -232 1270 -168
rect 1334 -232 1350 -168
rect 1254 -248 1350 -232
rect 1254 -312 1270 -248
rect 1334 -312 1350 -248
rect 1254 -328 1350 -312
rect 1254 -392 1270 -328
rect 1334 -392 1350 -328
rect 1254 -408 1350 -392
rect 1254 -472 1270 -408
rect 1334 -472 1350 -408
rect 1254 -488 1350 -472
rect 1254 -552 1270 -488
rect 1334 -552 1350 -488
rect 1254 -568 1350 -552
rect 1254 -632 1270 -568
rect 1334 -632 1350 -568
rect 1254 -648 1350 -632
rect 1254 -712 1270 -648
rect 1334 -712 1350 -648
rect 1254 -728 1350 -712
rect 1254 -792 1270 -728
rect 1334 -792 1350 -728
rect 1254 -808 1350 -792
rect 1254 -872 1270 -808
rect 1334 -872 1350 -808
rect 1254 -888 1350 -872
rect 1254 -952 1270 -888
rect 1334 -952 1350 -888
rect 1254 -968 1350 -952
rect 1254 -1032 1270 -968
rect 1334 -1032 1350 -968
rect 1254 -1048 1350 -1032
rect 1254 -1112 1270 -1048
rect 1334 -1112 1350 -1048
rect 1254 -1128 1350 -1112
rect 1254 -1192 1270 -1128
rect 1334 -1192 1350 -1128
rect 1254 -1208 1350 -1192
rect 1254 -1272 1270 -1208
rect 1334 -1272 1350 -1208
rect 1254 -1293 1350 -1272
<< properties >>
string FIXED_BBOX -1355 -1305 1255 1305
<< end >>
