magic
tech sky130A
timestamp 1670531611
<< error_p >>
rect 120 525 180 1650
rect 195 525 255 1650
rect 270 525 330 1650
rect 345 525 405 1650
rect 420 525 480 1650
<< nmoslvt >>
rect 180 525 195 1650
rect 255 525 270 1650
rect 330 525 345 1650
rect 405 525 420 1650
<< ndiff >>
rect 120 1630 180 1650
rect 120 545 140 1630
rect 160 545 180 1630
rect 120 525 180 545
rect 195 1630 255 1650
rect 195 545 215 1630
rect 235 545 255 1630
rect 195 525 255 545
rect 270 1630 330 1650
rect 270 545 290 1630
rect 310 545 330 1630
rect 270 525 330 545
rect 345 1630 405 1650
rect 345 545 365 1630
rect 385 545 405 1630
rect 345 525 405 545
rect 420 1630 480 1650
rect 420 545 440 1630
rect 460 545 480 1630
rect 420 525 480 545
<< ndiffc >>
rect 140 545 160 1630
rect 215 545 235 1630
rect 290 545 310 1630
rect 365 545 385 1630
rect 440 545 460 1630
<< poly >>
rect 180 1650 195 1665
rect 255 1650 270 1665
rect 330 1650 345 1665
rect 405 1650 420 1665
rect 180 510 195 525
rect 255 510 270 525
rect 330 510 345 525
rect 405 510 420 525
<< locali >>
rect 130 1630 170 1640
rect 130 545 140 1630
rect 160 545 170 1630
rect 130 535 170 545
rect 205 1630 245 1640
rect 205 545 215 1630
rect 235 545 245 1630
rect 205 535 245 545
rect 280 1630 320 1640
rect 280 545 290 1630
rect 310 545 320 1630
rect 280 535 320 545
rect 355 1630 395 1640
rect 355 545 365 1630
rect 385 545 395 1630
rect 355 535 395 545
rect 430 1630 470 1640
rect 430 545 440 1630
rect 460 545 470 1630
rect 430 535 470 545
<< end >>
