magic
tech sky130A
magscale 1 2
timestamp 1675786016
<< nwell >>
rect -1330 1310 1030 1500
rect -560 920 260 1310
<< pwell >>
rect -1316 144 1016 736
<< nmos >>
rect -1170 410 -1140 710
rect -1020 410 -990 710
rect -870 410 -840 710
rect -720 410 -690 710
rect -390 410 -360 710
rect -240 410 -210 710
rect -90 410 -60 710
rect 60 410 90 710
rect 390 410 420 710
rect 540 410 570 710
rect 690 410 720 710
rect 840 410 870 710
<< pmos >>
rect -390 970 -360 1270
rect -240 970 -210 1270
rect -90 970 -60 1270
rect 60 970 90 1270
<< ndiff >>
rect -1290 637 -1170 710
rect -1290 603 -1247 637
rect -1213 603 -1170 637
rect -1290 557 -1170 603
rect -1290 523 -1247 557
rect -1213 523 -1170 557
rect -1290 477 -1170 523
rect -1290 443 -1247 477
rect -1213 443 -1170 477
rect -1290 410 -1170 443
rect -1140 410 -1020 710
rect -990 637 -870 710
rect -990 603 -947 637
rect -913 603 -870 637
rect -990 557 -870 603
rect -990 523 -947 557
rect -913 523 -870 557
rect -990 477 -870 523
rect -990 443 -947 477
rect -913 443 -870 477
rect -990 410 -870 443
rect -840 410 -720 710
rect -690 637 -570 710
rect -690 603 -647 637
rect -613 603 -570 637
rect -690 557 -570 603
rect -690 523 -647 557
rect -613 523 -570 557
rect -690 477 -570 523
rect -690 443 -647 477
rect -613 443 -570 477
rect -690 410 -570 443
rect -510 637 -390 710
rect -510 603 -467 637
rect -433 603 -390 637
rect -510 557 -390 603
rect -510 523 -467 557
rect -433 523 -390 557
rect -510 477 -390 523
rect -510 443 -467 477
rect -433 443 -390 477
rect -510 410 -390 443
rect -360 637 -240 710
rect -360 603 -317 637
rect -283 603 -240 637
rect -360 557 -240 603
rect -360 523 -317 557
rect -283 523 -240 557
rect -360 477 -240 523
rect -360 443 -317 477
rect -283 443 -240 477
rect -360 410 -240 443
rect -210 637 -90 710
rect -210 603 -167 637
rect -133 603 -90 637
rect -210 557 -90 603
rect -210 523 -167 557
rect -133 523 -90 557
rect -210 477 -90 523
rect -210 443 -167 477
rect -133 443 -90 477
rect -210 410 -90 443
rect -60 637 60 710
rect -60 603 -17 637
rect 17 603 60 637
rect -60 557 60 603
rect -60 523 -17 557
rect 17 523 60 557
rect -60 477 60 523
rect -60 443 -17 477
rect 17 443 60 477
rect -60 410 60 443
rect 90 637 210 710
rect 90 603 133 637
rect 167 603 210 637
rect 90 557 210 603
rect 90 523 133 557
rect 167 523 210 557
rect 90 477 210 523
rect 90 443 133 477
rect 167 443 210 477
rect 90 410 210 443
rect 270 637 390 710
rect 270 603 313 637
rect 347 603 390 637
rect 270 557 390 603
rect 270 523 313 557
rect 347 523 390 557
rect 270 477 390 523
rect 270 443 313 477
rect 347 443 390 477
rect 270 410 390 443
rect 420 410 540 710
rect 570 637 690 710
rect 570 603 613 637
rect 647 603 690 637
rect 570 557 690 603
rect 570 523 613 557
rect 647 523 690 557
rect 570 477 690 523
rect 570 443 613 477
rect 647 443 690 477
rect 570 410 690 443
rect 720 410 840 710
rect 870 637 990 710
rect 870 603 913 637
rect 947 603 990 637
rect 870 557 990 603
rect 870 523 913 557
rect 947 523 990 557
rect 870 477 990 523
rect 870 443 913 477
rect 947 443 990 477
rect 870 410 990 443
<< pdiff >>
rect -510 1197 -390 1270
rect -510 1163 -467 1197
rect -433 1163 -390 1197
rect -510 1117 -390 1163
rect -510 1083 -467 1117
rect -433 1083 -390 1117
rect -510 1037 -390 1083
rect -510 1003 -467 1037
rect -433 1003 -390 1037
rect -510 970 -390 1003
rect -360 1197 -240 1270
rect -360 1163 -317 1197
rect -283 1163 -240 1197
rect -360 1117 -240 1163
rect -360 1083 -317 1117
rect -283 1083 -240 1117
rect -360 1037 -240 1083
rect -360 1003 -317 1037
rect -283 1003 -240 1037
rect -360 970 -240 1003
rect -210 1197 -90 1270
rect -210 1163 -167 1197
rect -133 1163 -90 1197
rect -210 1117 -90 1163
rect -210 1083 -167 1117
rect -133 1083 -90 1117
rect -210 1037 -90 1083
rect -210 1003 -167 1037
rect -133 1003 -90 1037
rect -210 970 -90 1003
rect -60 1197 60 1270
rect -60 1163 -17 1197
rect 17 1163 60 1197
rect -60 1117 60 1163
rect -60 1083 -17 1117
rect 17 1083 60 1117
rect -60 1037 60 1083
rect -60 1003 -17 1037
rect 17 1003 60 1037
rect -60 970 60 1003
rect 90 1197 210 1270
rect 90 1163 133 1197
rect 167 1163 210 1197
rect 90 1117 210 1163
rect 90 1083 133 1117
rect 167 1083 210 1117
rect 90 1037 210 1083
rect 90 1003 133 1037
rect 167 1003 210 1037
rect 90 970 210 1003
<< ndiffc >>
rect -1247 603 -1213 637
rect -1247 523 -1213 557
rect -1247 443 -1213 477
rect -947 603 -913 637
rect -947 523 -913 557
rect -947 443 -913 477
rect -647 603 -613 637
rect -647 523 -613 557
rect -647 443 -613 477
rect -467 603 -433 637
rect -467 523 -433 557
rect -467 443 -433 477
rect -317 603 -283 637
rect -317 523 -283 557
rect -317 443 -283 477
rect -167 603 -133 637
rect -167 523 -133 557
rect -167 443 -133 477
rect -17 603 17 637
rect -17 523 17 557
rect -17 443 17 477
rect 133 603 167 637
rect 133 523 167 557
rect 133 443 167 477
rect 313 603 347 637
rect 313 523 347 557
rect 313 443 347 477
rect 613 603 647 637
rect 613 523 647 557
rect 613 443 647 477
rect 913 603 947 637
rect 913 523 947 557
rect 913 443 947 477
<< pdiffc >>
rect -467 1163 -433 1197
rect -467 1083 -433 1117
rect -467 1003 -433 1037
rect -317 1163 -283 1197
rect -317 1083 -283 1117
rect -317 1003 -283 1037
rect -167 1163 -133 1197
rect -167 1083 -133 1117
rect -167 1003 -133 1037
rect -17 1163 17 1197
rect -17 1083 17 1117
rect -17 1003 17 1037
rect 133 1163 167 1197
rect 133 1083 167 1117
rect 133 1003 167 1037
<< psubdiff >>
rect -1290 237 990 270
rect -1290 203 -1207 237
rect -1173 203 -1127 237
rect -1093 203 -1047 237
rect -1013 203 -967 237
rect -933 203 -887 237
rect -853 203 -807 237
rect -773 203 -727 237
rect -693 203 -647 237
rect -613 203 -567 237
rect -533 203 -487 237
rect -453 203 -407 237
rect -373 203 -327 237
rect -293 203 -247 237
rect -213 203 -167 237
rect -133 203 -87 237
rect -53 203 -7 237
rect 27 203 73 237
rect 107 203 153 237
rect 187 203 233 237
rect 267 203 313 237
rect 347 203 393 237
rect 427 203 473 237
rect 507 203 553 237
rect 587 203 633 237
rect 667 203 713 237
rect 747 203 793 237
rect 827 203 873 237
rect 907 203 990 237
rect -1290 170 990 203
<< nsubdiff >>
rect -1290 1417 990 1450
rect -1290 1383 -1207 1417
rect -1173 1383 -1127 1417
rect -1093 1383 -1047 1417
rect -1013 1383 -967 1417
rect -933 1383 -887 1417
rect -853 1383 -807 1417
rect -773 1383 -727 1417
rect -693 1383 -647 1417
rect -613 1383 -567 1417
rect -533 1383 -487 1417
rect -453 1383 -407 1417
rect -373 1383 -327 1417
rect -293 1383 -247 1417
rect -213 1383 -167 1417
rect -133 1383 -87 1417
rect -53 1383 -7 1417
rect 27 1383 73 1417
rect 107 1383 153 1417
rect 187 1383 233 1417
rect 267 1383 313 1417
rect 347 1383 393 1417
rect 427 1383 473 1417
rect 507 1383 553 1417
rect 587 1383 633 1417
rect 667 1383 713 1417
rect 747 1383 793 1417
rect 827 1383 873 1417
rect 907 1383 990 1417
rect -1290 1350 990 1383
<< psubdiffcont >>
rect -1207 203 -1173 237
rect -1127 203 -1093 237
rect -1047 203 -1013 237
rect -967 203 -933 237
rect -887 203 -853 237
rect -807 203 -773 237
rect -727 203 -693 237
rect -647 203 -613 237
rect -567 203 -533 237
rect -487 203 -453 237
rect -407 203 -373 237
rect -327 203 -293 237
rect -247 203 -213 237
rect -167 203 -133 237
rect -87 203 -53 237
rect -7 203 27 237
rect 73 203 107 237
rect 153 203 187 237
rect 233 203 267 237
rect 313 203 347 237
rect 393 203 427 237
rect 473 203 507 237
rect 553 203 587 237
rect 633 203 667 237
rect 713 203 747 237
rect 793 203 827 237
rect 873 203 907 237
<< nsubdiffcont >>
rect -1207 1383 -1173 1417
rect -1127 1383 -1093 1417
rect -1047 1383 -1013 1417
rect -967 1383 -933 1417
rect -887 1383 -853 1417
rect -807 1383 -773 1417
rect -727 1383 -693 1417
rect -647 1383 -613 1417
rect -567 1383 -533 1417
rect -487 1383 -453 1417
rect -407 1383 -373 1417
rect -327 1383 -293 1417
rect -247 1383 -213 1417
rect -167 1383 -133 1417
rect -87 1383 -53 1417
rect -7 1383 27 1417
rect 73 1383 107 1417
rect 153 1383 187 1417
rect 233 1383 267 1417
rect 313 1383 347 1417
rect 393 1383 427 1417
rect 473 1383 507 1417
rect 553 1383 587 1417
rect 633 1383 667 1417
rect 713 1383 747 1417
rect 793 1383 827 1417
rect 873 1383 907 1417
<< poly >>
rect -900 1287 -820 1310
rect -900 1253 -877 1287
rect -843 1253 -820 1287
rect -390 1300 -210 1330
rect -390 1270 -360 1300
rect -240 1270 -210 1300
rect -90 1300 90 1330
rect -90 1270 -60 1300
rect 60 1270 90 1300
rect 490 1287 570 1310
rect -900 1230 -820 1253
rect -1045 1187 -965 1210
rect -1045 1153 -1022 1187
rect -988 1153 -965 1187
rect -1045 1130 -965 1153
rect -1220 987 -1140 1010
rect -1220 953 -1197 987
rect -1163 953 -1140 987
rect -1220 930 -1140 953
rect -1170 710 -1140 930
rect -1020 710 -990 1130
rect -870 710 -840 1230
rect -770 1087 -690 1110
rect -770 1053 -747 1087
rect -713 1053 -690 1087
rect -770 1030 -690 1053
rect -720 710 -690 1030
rect 490 1253 513 1287
rect 547 1253 570 1287
rect 490 1230 570 1253
rect 390 987 470 1010
rect -390 940 -360 970
rect -240 815 -210 970
rect -90 940 -60 970
rect 60 940 90 970
rect 390 953 413 987
rect 447 953 470 987
rect -140 917 -60 940
rect -140 883 -117 917
rect -83 883 -60 917
rect -140 860 -60 883
rect -240 792 -160 815
rect -240 758 -217 792
rect -183 758 -160 792
rect -390 710 -360 740
rect -240 735 -160 758
rect -240 710 -210 735
rect -90 710 -60 860
rect 390 930 470 953
rect 60 710 90 740
rect 390 710 420 930
rect 540 710 570 1230
rect 690 1187 770 1210
rect 690 1153 713 1187
rect 747 1153 770 1187
rect 690 1130 770 1153
rect 690 710 720 1130
rect 840 1087 920 1110
rect 840 1053 863 1087
rect 897 1053 920 1087
rect 840 1030 920 1053
rect 840 710 870 1030
rect -1170 380 -1140 410
rect -1020 380 -990 410
rect -870 380 -840 410
rect -720 380 -690 410
rect -390 380 -360 410
rect -240 380 -210 410
rect -90 380 -60 410
rect 60 380 90 410
rect 390 380 420 410
rect -390 357 -310 380
rect -390 323 -367 357
rect -333 323 -310 357
rect -390 300 -310 323
rect 10 357 90 380
rect 540 370 570 410
rect 690 370 720 410
rect 840 370 870 410
rect 10 323 33 357
rect 67 323 90 357
rect 10 300 90 323
<< polycont >>
rect -877 1253 -843 1287
rect -1022 1153 -988 1187
rect -1197 953 -1163 987
rect -747 1053 -713 1087
rect 513 1253 547 1287
rect 413 953 447 987
rect -117 883 -83 917
rect -217 758 -183 792
rect 713 1153 747 1187
rect 863 1053 897 1087
rect -367 323 -333 357
rect 33 323 67 357
<< locali >>
rect -1290 1417 990 1440
rect -1290 1383 -1207 1417
rect -1173 1383 -1127 1417
rect -1093 1383 -1047 1417
rect -1013 1383 -967 1417
rect -933 1383 -887 1417
rect -853 1383 -807 1417
rect -773 1383 -727 1417
rect -693 1383 -647 1417
rect -613 1383 -567 1417
rect -533 1383 -487 1417
rect -453 1383 -407 1417
rect -373 1383 -327 1417
rect -293 1383 -247 1417
rect -213 1383 -167 1417
rect -133 1383 -87 1417
rect -53 1383 -7 1417
rect 27 1383 73 1417
rect 107 1383 153 1417
rect 187 1383 233 1417
rect 267 1383 313 1417
rect 347 1383 393 1417
rect 427 1383 473 1417
rect 507 1383 553 1417
rect 587 1383 633 1417
rect 667 1383 713 1417
rect 747 1383 793 1417
rect 827 1383 873 1417
rect 907 1383 990 1417
rect -1290 1360 990 1383
rect -900 1290 -820 1310
rect -770 1290 -690 1310
rect -1290 1287 -690 1290
rect -1290 1253 -877 1287
rect -843 1253 -747 1287
rect -713 1253 -690 1287
rect -1290 1250 -690 1253
rect -900 1230 -820 1250
rect -770 1230 -690 1250
rect 490 1287 570 1310
rect 490 1253 513 1287
rect 547 1253 570 1287
rect 490 1230 570 1253
rect -1045 1190 -965 1210
rect -640 1190 -560 1210
rect -1290 1187 -560 1190
rect -1290 1153 -1022 1187
rect -988 1153 -617 1187
rect -583 1153 -560 1187
rect -1290 1150 -560 1153
rect -1045 1130 -965 1150
rect -640 1130 -560 1150
rect -490 1197 -410 1230
rect -490 1163 -467 1197
rect -433 1163 -410 1197
rect -490 1117 -410 1163
rect -770 1090 -690 1110
rect -1290 1087 -690 1090
rect -1290 1053 -747 1087
rect -713 1053 -690 1087
rect -1290 1050 -690 1053
rect -770 1030 -690 1050
rect -490 1083 -467 1117
rect -433 1083 -410 1117
rect -490 1037 -410 1083
rect -1220 990 -1140 1010
rect -640 990 -560 1010
rect -1290 987 -560 990
rect -1290 953 -1197 987
rect -1163 953 -617 987
rect -583 953 -560 987
rect -490 1003 -467 1037
rect -433 1003 -410 1037
rect -490 980 -410 1003
rect -340 1197 -260 1230
rect -340 1163 -317 1197
rect -283 1163 -260 1197
rect -340 1117 -260 1163
rect -340 1083 -317 1117
rect -283 1083 -260 1117
rect -340 1037 -260 1083
rect -340 1003 -317 1037
rect -283 1003 -260 1037
rect -340 970 -260 1003
rect -190 1197 -110 1230
rect -190 1163 -167 1197
rect -133 1163 -110 1197
rect -190 1117 -110 1163
rect -190 1083 -167 1117
rect -133 1083 -110 1117
rect -190 1037 -110 1083
rect -190 1003 -167 1037
rect -133 1003 -110 1037
rect -190 980 -110 1003
rect -40 1197 40 1230
rect -40 1163 -17 1197
rect 17 1163 40 1197
rect -40 1117 40 1163
rect -40 1083 -17 1117
rect 17 1083 40 1117
rect -40 1037 40 1083
rect -40 1003 -17 1037
rect 17 1003 40 1037
rect -40 970 40 1003
rect 110 1197 190 1230
rect 110 1163 133 1197
rect 167 1163 190 1197
rect 110 1117 190 1163
rect 690 1187 770 1210
rect 690 1153 713 1187
rect 747 1153 770 1187
rect 690 1130 770 1153
rect 110 1083 133 1117
rect 167 1083 190 1117
rect 110 1037 190 1083
rect 110 1003 133 1037
rect 167 1003 190 1037
rect 840 1087 920 1110
rect 840 1053 863 1087
rect 897 1053 920 1087
rect 840 1030 920 1053
rect 110 980 190 1003
rect 390 987 470 1010
rect -1290 950 -560 953
rect -1220 930 -1140 950
rect -640 930 -560 950
rect -320 920 -280 970
rect -140 920 -60 940
rect -320 917 -60 920
rect -320 883 -117 917
rect -83 883 -60 917
rect -320 880 -60 883
rect -320 750 -280 880
rect -140 860 -60 880
rect -1250 710 -280 750
rect -240 800 -160 815
rect -20 800 20 970
rect 390 953 413 987
rect 447 953 470 987
rect 390 930 470 953
rect 230 907 310 930
rect 230 873 253 907
rect 287 890 310 907
rect 287 873 990 890
rect 230 850 990 873
rect -240 792 990 800
rect -240 758 -217 792
rect -183 760 990 792
rect -183 758 -160 760
rect -240 735 -160 758
rect -1250 670 -1210 710
rect -650 670 -610 710
rect -320 670 -280 710
rect -20 670 20 760
rect 310 670 350 760
rect 910 670 950 760
rect -1270 637 -1190 670
rect -1270 603 -1247 637
rect -1213 603 -1190 637
rect -1270 557 -1190 603
rect -1270 523 -1247 557
rect -1213 523 -1190 557
rect -1270 477 -1190 523
rect -1270 443 -1247 477
rect -1213 443 -1190 477
rect -1270 420 -1190 443
rect -970 637 -890 670
rect -970 603 -947 637
rect -913 603 -890 637
rect -970 557 -890 603
rect -970 523 -947 557
rect -913 523 -890 557
rect -970 477 -890 523
rect -970 443 -947 477
rect -913 443 -890 477
rect -970 420 -890 443
rect -670 637 -590 670
rect -670 603 -647 637
rect -613 603 -590 637
rect -670 557 -590 603
rect -670 523 -647 557
rect -613 523 -590 557
rect -670 477 -590 523
rect -670 443 -647 477
rect -613 443 -590 477
rect -670 420 -590 443
rect -490 637 -410 670
rect -490 603 -467 637
rect -433 603 -410 637
rect -490 557 -410 603
rect -490 523 -467 557
rect -433 523 -410 557
rect -490 477 -410 523
rect -490 443 -467 477
rect -433 443 -410 477
rect -490 420 -410 443
rect -340 637 -260 670
rect -340 603 -317 637
rect -283 603 -260 637
rect -340 557 -260 603
rect -340 523 -317 557
rect -283 523 -260 557
rect -340 477 -260 523
rect -340 443 -317 477
rect -283 443 -260 477
rect -340 420 -260 443
rect -190 637 -110 670
rect -190 603 -167 637
rect -133 603 -110 637
rect -190 557 -110 603
rect -190 523 -167 557
rect -133 523 -110 557
rect -190 477 -110 523
rect -190 443 -167 477
rect -133 443 -110 477
rect -190 420 -110 443
rect -40 637 40 670
rect -40 603 -17 637
rect 17 603 40 637
rect -40 557 40 603
rect -40 523 -17 557
rect 17 523 40 557
rect -40 477 40 523
rect -40 443 -17 477
rect 17 443 40 477
rect -40 420 40 443
rect 110 637 190 670
rect 110 603 133 637
rect 167 603 190 637
rect 110 557 190 603
rect 110 523 133 557
rect 167 523 190 557
rect 110 477 190 523
rect 110 443 133 477
rect 167 443 190 477
rect 110 420 190 443
rect 290 637 370 670
rect 290 603 313 637
rect 347 603 370 637
rect 290 557 370 603
rect 290 523 313 557
rect 347 523 370 557
rect 290 477 370 523
rect 290 443 313 477
rect 347 443 370 477
rect 290 420 370 443
rect 590 637 670 670
rect 590 603 613 637
rect 647 603 670 637
rect 590 557 670 603
rect 590 523 613 557
rect 647 523 670 557
rect 590 477 670 523
rect 590 443 613 477
rect 647 443 670 477
rect 590 420 670 443
rect 890 637 970 670
rect 890 603 913 637
rect 947 603 970 637
rect 890 557 970 603
rect 890 523 913 557
rect 947 523 970 557
rect 890 477 970 523
rect 890 443 913 477
rect 947 443 970 477
rect 890 420 970 443
rect -390 360 -310 380
rect 10 360 90 380
rect -1290 357 90 360
rect -1290 323 -367 357
rect -333 323 33 357
rect 67 323 90 357
rect -1290 320 90 323
rect -390 300 -310 320
rect 10 300 90 320
rect -1290 237 990 260
rect -1290 203 -1207 237
rect -1173 203 -1127 237
rect -1093 203 -1047 237
rect -1013 203 -967 237
rect -933 203 -887 237
rect -853 203 -807 237
rect -773 203 -727 237
rect -693 203 -647 237
rect -613 203 -567 237
rect -533 203 -487 237
rect -453 203 -407 237
rect -373 203 -327 237
rect -293 203 -247 237
rect -213 203 -167 237
rect -133 203 -87 237
rect -53 203 -7 237
rect 27 203 73 237
rect 107 203 153 237
rect 187 203 233 237
rect 267 203 313 237
rect 347 203 393 237
rect 427 203 473 237
rect 507 203 553 237
rect 587 203 633 237
rect 667 203 713 237
rect 747 203 793 237
rect 827 203 873 237
rect 907 203 990 237
rect -1290 180 990 203
<< viali >>
rect -1207 1383 -1173 1417
rect -1127 1383 -1093 1417
rect -1047 1383 -1013 1417
rect -967 1383 -933 1417
rect -887 1383 -853 1417
rect -807 1383 -773 1417
rect -727 1383 -693 1417
rect -647 1383 -613 1417
rect -567 1383 -533 1417
rect -487 1383 -453 1417
rect -407 1383 -373 1417
rect -327 1383 -293 1417
rect -247 1383 -213 1417
rect -167 1383 -133 1417
rect -87 1383 -53 1417
rect -7 1383 27 1417
rect 73 1383 107 1417
rect 153 1383 187 1417
rect 233 1383 267 1417
rect 313 1383 347 1417
rect 393 1383 427 1417
rect 473 1383 507 1417
rect 553 1383 587 1417
rect 633 1383 667 1417
rect 713 1383 747 1417
rect 793 1383 827 1417
rect 873 1383 907 1417
rect -747 1253 -713 1287
rect 513 1253 547 1287
rect -617 1153 -583 1187
rect -467 1163 -433 1197
rect -747 1053 -713 1087
rect -467 1083 -433 1117
rect -617 953 -583 987
rect -467 1003 -433 1037
rect -167 1163 -133 1197
rect -167 1083 -133 1117
rect -167 1003 -133 1037
rect 133 1163 167 1197
rect 713 1153 747 1187
rect 133 1083 167 1117
rect 133 1003 167 1037
rect 863 1053 897 1087
rect -117 883 -83 917
rect 413 953 447 987
rect 253 873 287 907
rect -947 603 -913 637
rect -947 523 -913 557
rect -947 443 -913 477
rect -467 603 -433 637
rect -467 523 -433 557
rect -467 443 -433 477
rect -167 603 -133 637
rect -167 523 -133 557
rect -167 443 -133 477
rect 133 603 167 637
rect 133 523 167 557
rect 133 443 167 477
rect 613 603 647 637
rect 613 523 647 557
rect 613 443 647 477
rect -1207 203 -1173 237
rect -1127 203 -1093 237
rect -1047 203 -1013 237
rect -967 203 -933 237
rect -887 203 -853 237
rect -807 203 -773 237
rect -727 203 -693 237
rect -647 203 -613 237
rect -567 203 -533 237
rect -487 203 -453 237
rect -407 203 -373 237
rect -327 203 -293 237
rect -247 203 -213 237
rect -167 203 -133 237
rect -87 203 -53 237
rect -7 203 27 237
rect 73 203 107 237
rect 153 203 187 237
rect 233 203 267 237
rect 313 203 347 237
rect 393 203 427 237
rect 473 203 507 237
rect 553 203 587 237
rect 633 203 667 237
rect 713 203 747 237
rect 793 203 827 237
rect 873 203 907 237
<< metal1 >>
rect -1290 1417 990 1450
rect -1290 1383 -1207 1417
rect -1173 1383 -1127 1417
rect -1093 1383 -1047 1417
rect -1013 1383 -967 1417
rect -933 1383 -887 1417
rect -853 1383 -807 1417
rect -773 1383 -727 1417
rect -693 1383 -647 1417
rect -613 1383 -567 1417
rect -533 1383 -487 1417
rect -453 1383 -407 1417
rect -373 1383 -327 1417
rect -293 1383 -247 1417
rect -213 1383 -167 1417
rect -133 1383 -87 1417
rect -53 1383 -7 1417
rect 27 1383 73 1417
rect 107 1383 153 1417
rect 187 1383 233 1417
rect 267 1383 313 1417
rect 347 1383 393 1417
rect 427 1383 473 1417
rect 507 1383 553 1417
rect 587 1383 633 1417
rect 667 1383 713 1417
rect 747 1383 793 1417
rect 827 1383 873 1417
rect 907 1383 990 1417
rect -1290 1350 990 1383
rect -950 670 -910 1350
rect -770 1296 -690 1310
rect -770 1244 -756 1296
rect -704 1244 -690 1296
rect -770 1230 -690 1244
rect -640 1196 -560 1210
rect -640 1144 -626 1196
rect -574 1144 -560 1196
rect -640 1130 -560 1144
rect -490 1197 -410 1350
rect -490 1163 -467 1197
rect -433 1163 -410 1197
rect -490 1117 -410 1163
rect -770 1096 -690 1110
rect -770 1044 -756 1096
rect -704 1044 -690 1096
rect -770 1030 -690 1044
rect -490 1083 -467 1117
rect -433 1083 -410 1117
rect -490 1037 -410 1083
rect -640 996 -560 1010
rect -640 944 -626 996
rect -574 944 -560 996
rect -490 1003 -467 1037
rect -433 1003 -410 1037
rect -490 980 -410 1003
rect -190 1197 -110 1350
rect -190 1163 -167 1197
rect -133 1163 -110 1197
rect -190 1117 -110 1163
rect -190 1083 -167 1117
rect -133 1083 -110 1117
rect -190 1037 -110 1083
rect -190 1003 -167 1037
rect -133 1003 -110 1037
rect -190 980 -110 1003
rect 110 1197 190 1350
rect 490 1296 570 1310
rect 490 1244 504 1296
rect 556 1244 570 1296
rect 490 1230 570 1244
rect 110 1163 133 1197
rect 167 1163 190 1197
rect 110 1117 190 1163
rect 110 1083 133 1117
rect 167 1083 190 1117
rect 110 1037 190 1083
rect 110 1003 133 1037
rect 167 1003 190 1037
rect 110 980 190 1003
rect 390 996 470 1010
rect -640 930 -560 944
rect 390 944 404 996
rect 456 944 470 996
rect -140 917 -60 940
rect 390 930 470 944
rect -140 883 -117 917
rect -83 900 -60 917
rect 230 907 310 930
rect 230 900 253 907
rect -83 883 253 900
rect -140 873 253 883
rect 287 873 310 907
rect -140 860 310 873
rect 230 850 310 860
rect 610 670 650 1350
rect 690 1196 770 1210
rect 690 1144 704 1196
rect 756 1144 770 1196
rect 690 1130 770 1144
rect 840 1096 920 1110
rect 840 1044 854 1096
rect 906 1044 920 1096
rect 840 1030 920 1044
rect -970 637 -890 670
rect -970 603 -947 637
rect -913 603 -890 637
rect -970 557 -890 603
rect -970 523 -947 557
rect -913 523 -890 557
rect -970 477 -890 523
rect -970 443 -947 477
rect -913 443 -890 477
rect -970 420 -890 443
rect -490 637 -410 670
rect -490 603 -467 637
rect -433 603 -410 637
rect -490 557 -410 603
rect -490 523 -467 557
rect -433 523 -410 557
rect -490 477 -410 523
rect -490 443 -467 477
rect -433 443 -410 477
rect -490 420 -410 443
rect -190 637 -110 670
rect -190 603 -167 637
rect -133 603 -110 637
rect -190 557 -110 603
rect -190 523 -167 557
rect -133 523 -110 557
rect -190 477 -110 523
rect -190 443 -167 477
rect -133 443 -110 477
rect -190 420 -110 443
rect 110 637 190 670
rect 110 603 133 637
rect 167 603 190 637
rect 110 557 190 603
rect 110 523 133 557
rect 167 523 190 557
rect 110 477 190 523
rect 110 443 133 477
rect 167 443 190 477
rect 110 420 190 443
rect 590 637 670 670
rect 590 603 613 637
rect 647 603 670 637
rect 590 557 670 603
rect 590 523 613 557
rect 647 523 670 557
rect 590 477 670 523
rect 590 443 613 477
rect 647 443 670 477
rect 590 420 670 443
rect -470 270 -430 420
rect -170 270 -130 420
rect 130 270 170 420
rect -1290 237 990 270
rect -1290 203 -1207 237
rect -1173 203 -1127 237
rect -1093 203 -1047 237
rect -1013 203 -967 237
rect -933 203 -887 237
rect -853 203 -807 237
rect -773 203 -727 237
rect -693 203 -647 237
rect -613 203 -567 237
rect -533 203 -487 237
rect -453 203 -407 237
rect -373 203 -327 237
rect -293 203 -247 237
rect -213 203 -167 237
rect -133 203 -87 237
rect -53 203 -7 237
rect 27 203 73 237
rect 107 203 153 237
rect 187 203 233 237
rect 267 203 313 237
rect 347 203 393 237
rect 427 203 473 237
rect 507 203 553 237
rect 587 203 633 237
rect 667 203 713 237
rect 747 203 793 237
rect 827 203 873 237
rect 907 203 990 237
rect -1290 170 990 203
<< via1 >>
rect -756 1287 -704 1296
rect -756 1253 -747 1287
rect -747 1253 -713 1287
rect -713 1253 -704 1287
rect -756 1244 -704 1253
rect -626 1187 -574 1196
rect -626 1153 -617 1187
rect -617 1153 -583 1187
rect -583 1153 -574 1187
rect -626 1144 -574 1153
rect -756 1087 -704 1096
rect -756 1053 -747 1087
rect -747 1053 -713 1087
rect -713 1053 -704 1087
rect -756 1044 -704 1053
rect -626 987 -574 996
rect -626 953 -617 987
rect -617 953 -583 987
rect -583 953 -574 987
rect -626 944 -574 953
rect 504 1287 556 1296
rect 504 1253 513 1287
rect 513 1253 547 1287
rect 547 1253 556 1287
rect 504 1244 556 1253
rect 404 987 456 996
rect 404 953 413 987
rect 413 953 447 987
rect 447 953 456 987
rect 404 944 456 953
rect 704 1187 756 1196
rect 704 1153 713 1187
rect 713 1153 747 1187
rect 747 1153 756 1187
rect 704 1144 756 1153
rect 854 1087 906 1096
rect 854 1053 863 1087
rect 863 1053 897 1087
rect 897 1053 906 1087
rect 854 1044 906 1053
<< metal2 >>
rect -770 1296 -690 1310
rect -770 1244 -756 1296
rect -704 1290 -690 1296
rect 490 1296 570 1310
rect 490 1290 504 1296
rect -704 1250 504 1290
rect -704 1244 -690 1250
rect -770 1230 -690 1244
rect 490 1244 504 1250
rect 556 1244 570 1296
rect 490 1230 570 1244
rect -640 1196 -560 1210
rect -640 1144 -626 1196
rect -574 1190 -560 1196
rect 690 1196 770 1210
rect 690 1190 704 1196
rect -574 1150 704 1190
rect -574 1144 -560 1150
rect -640 1130 -560 1144
rect 690 1144 704 1150
rect 756 1144 770 1196
rect 690 1130 770 1144
rect -770 1096 -690 1110
rect -770 1044 -756 1096
rect -704 1090 -690 1096
rect 840 1096 920 1110
rect 840 1090 854 1096
rect -704 1050 854 1090
rect -704 1044 -690 1050
rect -770 1030 -690 1044
rect 840 1044 854 1050
rect 906 1044 920 1096
rect 840 1030 920 1044
rect -640 996 -560 1010
rect -640 944 -626 996
rect -574 990 -560 996
rect 390 996 470 1010
rect 390 990 404 996
rect -574 950 404 990
rect -574 944 -560 950
rect -640 930 -560 944
rect 390 944 404 950
rect 456 944 470 996
rect 390 930 470 944
<< labels >>
rlabel metal1 s -120 880 -80 920 4 OUT_bar
port 1 nsew
rlabel metal1 s -170 200 -130 240 4 GND!
port 2 nsew
rlabel metal1 s -170 1380 -130 1420 4 CLK
port 3 nsew
rlabel locali s -220 755 -180 795 4 OUT
port 4 nsew
rlabel locali s -1280 1260 -1260 1280 4 A
port 5 nsew
rlabel locali s -1280 1160 -1260 1180 4 A_bar
port 6 nsew
rlabel locali s -1280 1060 -1260 1080 4 B
port 7 nsew
rlabel locali s -1280 960 -1260 980 4 B_bar
port 8 nsew
rlabel locali s -370 320 -330 360 4 Dis
port 9 nsew
<< end >>
