* NGSPICE file created from EESPFAL_4in_XOR.ext - technology: sky130A

.subckt EESPFAL_XOR_v3 OUT A A_bar B B_bar Dis OUT_bar GND CLK
X0 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 OUT_bar B a_n690_n412# GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X2 a_570_n412# B_bar OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X3 a_n690_n412# A CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.5e+12p ps=3.22e+07u w=1.5e+06u l=150000u
X4 OUT_bar OUT CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X5 CLK A a_570_n412# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 CLK A_bar a_n990_n412# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X7 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X8 a_870_n412# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n990_n412# B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 OUT B a_870_n412# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_4in_XOR x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar x2 x2_bar k2 k2_bar
+ x3 x3_bar k3 k3_bar XOR0_bar XOR0 XOR1_bar XOR1 XOR2_bar XOR2 XOR3_bar XOR3 GND
+ CLK Dis
XEESPFAL_XOR_v3_0 XOR3 x3 x3_bar k3 k3_bar Dis XOR3_bar GND CLK EESPFAL_XOR_v3
XEESPFAL_XOR_v3_1 XOR2 x2 x2_bar k2 k2_bar Dis XOR2_bar GND CLK EESPFAL_XOR_v3
XEESPFAL_XOR_v3_2 XOR1 x1 x1_bar k1 k1_bar Dis XOR1_bar GND CLK EESPFAL_XOR_v3
XEESPFAL_XOR_v3_3 XOR0 x0 x0_bar k0 k0_bar Dis XOR0_bar GND CLK EESPFAL_XOR_v3
.ends

