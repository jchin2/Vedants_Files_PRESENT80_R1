magic
tech sky130A
magscale 1 2
timestamp 1671306811
<< metal3 >>
rect -1030 952 1029 1000
rect -1030 888 945 952
rect 1009 888 1029 952
rect -1030 872 1029 888
rect -1030 808 945 872
rect 1009 808 1029 872
rect -1030 792 1029 808
rect -1030 728 945 792
rect 1009 728 1029 792
rect -1030 712 1029 728
rect -1030 648 945 712
rect 1009 648 1029 712
rect -1030 632 1029 648
rect -1030 568 945 632
rect 1009 568 1029 632
rect -1030 552 1029 568
rect -1030 488 945 552
rect 1009 488 1029 552
rect -1030 472 1029 488
rect -1030 408 945 472
rect 1009 408 1029 472
rect -1030 392 1029 408
rect -1030 328 945 392
rect 1009 328 1029 392
rect -1030 312 1029 328
rect -1030 248 945 312
rect 1009 248 1029 312
rect -1030 232 1029 248
rect -1030 168 945 232
rect 1009 168 1029 232
rect -1030 152 1029 168
rect -1030 88 945 152
rect 1009 88 1029 152
rect -1030 72 1029 88
rect -1030 8 945 72
rect 1009 8 1029 72
rect -1030 -8 1029 8
rect -1030 -72 945 -8
rect 1009 -72 1029 -8
rect -1030 -88 1029 -72
rect -1030 -152 945 -88
rect 1009 -152 1029 -88
rect -1030 -168 1029 -152
rect -1030 -232 945 -168
rect 1009 -232 1029 -168
rect -1030 -248 1029 -232
rect -1030 -312 945 -248
rect 1009 -312 1029 -248
rect -1030 -328 1029 -312
rect -1030 -392 945 -328
rect 1009 -392 1029 -328
rect -1030 -408 1029 -392
rect -1030 -472 945 -408
rect 1009 -472 1029 -408
rect -1030 -488 1029 -472
rect -1030 -552 945 -488
rect 1009 -552 1029 -488
rect -1030 -568 1029 -552
rect -1030 -632 945 -568
rect 1009 -632 1029 -568
rect -1030 -648 1029 -632
rect -1030 -712 945 -648
rect 1009 -712 1029 -648
rect -1030 -728 1029 -712
rect -1030 -792 945 -728
rect 1009 -792 1029 -728
rect -1030 -808 1029 -792
rect -1030 -872 945 -808
rect 1009 -872 1029 -808
rect -1030 -888 1029 -872
rect -1030 -952 945 -888
rect 1009 -952 1029 -888
rect -1030 -1000 1029 -952
<< via3 >>
rect 945 888 1009 952
rect 945 808 1009 872
rect 945 728 1009 792
rect 945 648 1009 712
rect 945 568 1009 632
rect 945 488 1009 552
rect 945 408 1009 472
rect 945 328 1009 392
rect 945 248 1009 312
rect 945 168 1009 232
rect 945 88 1009 152
rect 945 8 1009 72
rect 945 -72 1009 -8
rect 945 -152 1009 -88
rect 945 -232 1009 -168
rect 945 -312 1009 -248
rect 945 -392 1009 -328
rect 945 -472 1009 -408
rect 945 -552 1009 -488
rect 945 -632 1009 -568
rect 945 -712 1009 -648
rect 945 -792 1009 -728
rect 945 -872 1009 -808
rect 945 -952 1009 -888
<< mimcap >>
rect -930 832 830 900
rect -930 -832 -882 832
rect 782 -832 830 832
rect -930 -900 830 -832
<< mimcapcontact >>
rect -882 -832 782 832
<< metal4 >>
rect 929 952 1025 988
rect 929 888 945 952
rect 1009 888 1025 952
rect 929 872 1025 888
rect -891 832 791 861
rect -891 -832 -882 832
rect 782 -832 791 832
rect -891 -861 791 -832
rect 929 808 945 872
rect 1009 808 1025 872
rect 929 792 1025 808
rect 929 728 945 792
rect 1009 728 1025 792
rect 929 712 1025 728
rect 929 648 945 712
rect 1009 648 1025 712
rect 929 632 1025 648
rect 929 568 945 632
rect 1009 568 1025 632
rect 929 552 1025 568
rect 929 488 945 552
rect 1009 488 1025 552
rect 929 472 1025 488
rect 929 408 945 472
rect 1009 408 1025 472
rect 929 392 1025 408
rect 929 328 945 392
rect 1009 328 1025 392
rect 929 312 1025 328
rect 929 248 945 312
rect 1009 248 1025 312
rect 929 232 1025 248
rect 929 168 945 232
rect 1009 168 1025 232
rect 929 152 1025 168
rect 929 88 945 152
rect 1009 88 1025 152
rect 929 72 1025 88
rect 929 8 945 72
rect 1009 8 1025 72
rect 929 -8 1025 8
rect 929 -72 945 -8
rect 1009 -72 1025 -8
rect 929 -88 1025 -72
rect 929 -152 945 -88
rect 1009 -152 1025 -88
rect 929 -168 1025 -152
rect 929 -232 945 -168
rect 1009 -232 1025 -168
rect 929 -248 1025 -232
rect 929 -312 945 -248
rect 1009 -312 1025 -248
rect 929 -328 1025 -312
rect 929 -392 945 -328
rect 1009 -392 1025 -328
rect 929 -408 1025 -392
rect 929 -472 945 -408
rect 1009 -472 1025 -408
rect 929 -488 1025 -472
rect 929 -552 945 -488
rect 1009 -552 1025 -488
rect 929 -568 1025 -552
rect 929 -632 945 -568
rect 1009 -632 1025 -568
rect 929 -648 1025 -632
rect 929 -712 945 -648
rect 1009 -712 1025 -648
rect 929 -728 1025 -712
rect 929 -792 945 -728
rect 1009 -792 1025 -728
rect 929 -808 1025 -792
rect 929 -872 945 -808
rect 1009 -872 1025 -808
rect 929 -888 1025 -872
rect 929 -952 945 -888
rect 1009 -952 1025 -888
rect 929 -988 1025 -952
<< properties >>
string FIXED_BBOX -1030 -1000 930 1000
<< end >>
