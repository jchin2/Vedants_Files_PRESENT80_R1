magic
tech sky130A
magscale 1 2
timestamp 1671058898
<< error_p >>
rect -1110 20 -990 1020
rect -960 20 -840 1020
rect -810 20 -690 1020
rect -660 20 -540 1020
rect -510 20 -390 1020
<< pwell >>
rect -1136 -6 -364 1046
<< nmoslvt >>
rect -990 20 -960 1020
rect -840 20 -810 1020
rect -690 20 -660 1020
rect -540 20 -510 1020
<< ndiff >>
rect -1110 962 -990 1020
rect -1110 928 -1067 962
rect -1033 928 -990 962
rect -1110 861 -990 928
rect -1110 827 -1067 861
rect -1033 827 -990 861
rect -1110 793 -990 827
rect -1110 759 -1067 793
rect -1033 759 -990 793
rect -1110 725 -990 759
rect -1110 691 -1067 725
rect -1033 691 -990 725
rect -1110 657 -990 691
rect -1110 623 -1067 657
rect -1033 623 -990 657
rect -1110 589 -990 623
rect -1110 555 -1067 589
rect -1033 555 -990 589
rect -1110 521 -990 555
rect -1110 487 -1067 521
rect -1033 487 -990 521
rect -1110 453 -990 487
rect -1110 419 -1067 453
rect -1033 419 -990 453
rect -1110 385 -990 419
rect -1110 351 -1067 385
rect -1033 351 -990 385
rect -1110 317 -990 351
rect -1110 283 -1067 317
rect -1033 283 -990 317
rect -1110 249 -990 283
rect -1110 215 -1067 249
rect -1033 215 -990 249
rect -1110 181 -990 215
rect -1110 147 -1067 181
rect -1033 147 -990 181
rect -1110 113 -990 147
rect -1110 79 -1067 113
rect -1033 79 -990 113
rect -1110 20 -990 79
rect -960 962 -840 1020
rect -960 928 -917 962
rect -883 928 -840 962
rect -960 851 -840 928
rect -960 817 -917 851
rect -883 817 -840 851
rect -960 783 -840 817
rect -960 749 -917 783
rect -883 749 -840 783
rect -960 715 -840 749
rect -960 681 -917 715
rect -883 681 -840 715
rect -960 647 -840 681
rect -960 613 -917 647
rect -883 613 -840 647
rect -960 579 -840 613
rect -960 545 -917 579
rect -883 545 -840 579
rect -960 511 -840 545
rect -960 477 -917 511
rect -883 477 -840 511
rect -960 443 -840 477
rect -960 409 -917 443
rect -883 409 -840 443
rect -960 375 -840 409
rect -960 341 -917 375
rect -883 341 -840 375
rect -960 307 -840 341
rect -960 273 -917 307
rect -883 273 -840 307
rect -960 239 -840 273
rect -960 205 -917 239
rect -883 205 -840 239
rect -960 171 -840 205
rect -960 137 -917 171
rect -883 137 -840 171
rect -960 103 -840 137
rect -960 69 -917 103
rect -883 69 -840 103
rect -960 20 -840 69
rect -810 962 -690 1020
rect -810 928 -767 962
rect -733 928 -690 962
rect -810 861 -690 928
rect -810 827 -767 861
rect -733 827 -690 861
rect -810 793 -690 827
rect -810 759 -767 793
rect -733 759 -690 793
rect -810 725 -690 759
rect -810 691 -767 725
rect -733 691 -690 725
rect -810 657 -690 691
rect -810 623 -767 657
rect -733 623 -690 657
rect -810 589 -690 623
rect -810 555 -767 589
rect -733 555 -690 589
rect -810 521 -690 555
rect -810 487 -767 521
rect -733 487 -690 521
rect -810 453 -690 487
rect -810 419 -767 453
rect -733 419 -690 453
rect -810 385 -690 419
rect -810 351 -767 385
rect -733 351 -690 385
rect -810 317 -690 351
rect -810 283 -767 317
rect -733 283 -690 317
rect -810 249 -690 283
rect -810 215 -767 249
rect -733 215 -690 249
rect -810 181 -690 215
rect -810 147 -767 181
rect -733 147 -690 181
rect -810 113 -690 147
rect -810 79 -767 113
rect -733 79 -690 113
rect -810 20 -690 79
rect -660 962 -540 1020
rect -660 928 -617 962
rect -583 928 -540 962
rect -660 861 -540 928
rect -660 827 -617 861
rect -583 827 -540 861
rect -660 793 -540 827
rect -660 759 -617 793
rect -583 759 -540 793
rect -660 725 -540 759
rect -660 691 -617 725
rect -583 691 -540 725
rect -660 657 -540 691
rect -660 623 -617 657
rect -583 623 -540 657
rect -660 589 -540 623
rect -660 555 -617 589
rect -583 555 -540 589
rect -660 521 -540 555
rect -660 487 -617 521
rect -583 487 -540 521
rect -660 453 -540 487
rect -660 419 -617 453
rect -583 419 -540 453
rect -660 385 -540 419
rect -660 351 -617 385
rect -583 351 -540 385
rect -660 317 -540 351
rect -660 283 -617 317
rect -583 283 -540 317
rect -660 249 -540 283
rect -660 215 -617 249
rect -583 215 -540 249
rect -660 181 -540 215
rect -660 147 -617 181
rect -583 147 -540 181
rect -660 113 -540 147
rect -660 79 -617 113
rect -583 79 -540 113
rect -660 20 -540 79
rect -510 962 -390 1020
rect -510 928 -467 962
rect -433 928 -390 962
rect -510 861 -390 928
rect -510 827 -467 861
rect -433 827 -390 861
rect -510 793 -390 827
rect -510 759 -467 793
rect -433 759 -390 793
rect -510 725 -390 759
rect -510 691 -467 725
rect -433 691 -390 725
rect -510 657 -390 691
rect -510 623 -467 657
rect -433 623 -390 657
rect -510 589 -390 623
rect -510 555 -467 589
rect -433 555 -390 589
rect -510 521 -390 555
rect -510 487 -467 521
rect -433 487 -390 521
rect -510 453 -390 487
rect -510 419 -467 453
rect -433 419 -390 453
rect -510 385 -390 419
rect -510 351 -467 385
rect -433 351 -390 385
rect -510 317 -390 351
rect -510 283 -467 317
rect -433 283 -390 317
rect -510 249 -390 283
rect -510 215 -467 249
rect -433 215 -390 249
rect -510 181 -390 215
rect -510 147 -467 181
rect -433 147 -390 181
rect -510 113 -390 147
rect -510 79 -467 113
rect -433 79 -390 113
rect -510 20 -390 79
<< ndiffc >>
rect -1067 928 -1033 962
rect -1067 827 -1033 861
rect -1067 759 -1033 793
rect -1067 691 -1033 725
rect -1067 623 -1033 657
rect -1067 555 -1033 589
rect -1067 487 -1033 521
rect -1067 419 -1033 453
rect -1067 351 -1033 385
rect -1067 283 -1033 317
rect -1067 215 -1033 249
rect -1067 147 -1033 181
rect -1067 79 -1033 113
rect -917 928 -883 962
rect -917 817 -883 851
rect -917 749 -883 783
rect -917 681 -883 715
rect -917 613 -883 647
rect -917 545 -883 579
rect -917 477 -883 511
rect -917 409 -883 443
rect -917 341 -883 375
rect -917 273 -883 307
rect -917 205 -883 239
rect -917 137 -883 171
rect -917 69 -883 103
rect -767 928 -733 962
rect -767 827 -733 861
rect -767 759 -733 793
rect -767 691 -733 725
rect -767 623 -733 657
rect -767 555 -733 589
rect -767 487 -733 521
rect -767 419 -733 453
rect -767 351 -733 385
rect -767 283 -733 317
rect -767 215 -733 249
rect -767 147 -733 181
rect -767 79 -733 113
rect -617 928 -583 962
rect -617 827 -583 861
rect -617 759 -583 793
rect -617 691 -583 725
rect -617 623 -583 657
rect -617 555 -583 589
rect -617 487 -583 521
rect -617 419 -583 453
rect -617 351 -583 385
rect -617 283 -583 317
rect -617 215 -583 249
rect -617 147 -583 181
rect -617 79 -583 113
rect -467 928 -433 962
rect -467 827 -433 861
rect -467 759 -433 793
rect -467 691 -433 725
rect -467 623 -433 657
rect -467 555 -433 589
rect -467 487 -433 521
rect -467 419 -433 453
rect -467 351 -433 385
rect -467 283 -433 317
rect -467 215 -433 249
rect -467 147 -433 181
rect -467 79 -433 113
<< poly >>
rect -990 1070 -510 1100
rect -990 1020 -960 1070
rect -840 1020 -810 1070
rect -690 1020 -660 1070
rect -540 1020 -510 1070
rect -990 -10 -960 20
rect -840 -10 -810 20
rect -690 -10 -660 20
rect -540 -10 -510 20
<< locali >>
rect -920 1040 -580 1080
rect -920 1000 -880 1040
rect -620 1000 -580 1040
rect -1090 962 -1010 1000
rect -1090 928 -1067 962
rect -1033 928 -1010 962
rect -1090 861 -1010 928
rect -1090 827 -1067 861
rect -1033 827 -1010 861
rect -1090 793 -1010 827
rect -1090 759 -1067 793
rect -1033 759 -1010 793
rect -1090 725 -1010 759
rect -1090 691 -1067 725
rect -1033 691 -1010 725
rect -1090 657 -1010 691
rect -1090 623 -1067 657
rect -1033 623 -1010 657
rect -1090 589 -1010 623
rect -1090 555 -1067 589
rect -1033 555 -1010 589
rect -1090 521 -1010 555
rect -1090 487 -1067 521
rect -1033 487 -1010 521
rect -1090 453 -1010 487
rect -1090 419 -1067 453
rect -1033 419 -1010 453
rect -1090 385 -1010 419
rect -1090 351 -1067 385
rect -1033 351 -1010 385
rect -1090 317 -1010 351
rect -1090 283 -1067 317
rect -1033 283 -1010 317
rect -1090 249 -1010 283
rect -1090 215 -1067 249
rect -1033 215 -1010 249
rect -1090 181 -1010 215
rect -1090 147 -1067 181
rect -1033 147 -1010 181
rect -1090 113 -1010 147
rect -1090 79 -1067 113
rect -1033 79 -1010 113
rect -1090 40 -1010 79
rect -940 962 -860 1000
rect -940 928 -917 962
rect -883 928 -860 962
rect -940 851 -860 928
rect -940 817 -917 851
rect -883 817 -860 851
rect -940 783 -860 817
rect -940 749 -917 783
rect -883 749 -860 783
rect -940 715 -860 749
rect -940 681 -917 715
rect -883 681 -860 715
rect -940 647 -860 681
rect -940 613 -917 647
rect -883 613 -860 647
rect -940 579 -860 613
rect -940 545 -917 579
rect -883 545 -860 579
rect -940 511 -860 545
rect -940 477 -917 511
rect -883 477 -860 511
rect -940 443 -860 477
rect -940 409 -917 443
rect -883 409 -860 443
rect -940 375 -860 409
rect -940 341 -917 375
rect -883 341 -860 375
rect -940 307 -860 341
rect -940 273 -917 307
rect -883 273 -860 307
rect -940 239 -860 273
rect -940 205 -917 239
rect -883 205 -860 239
rect -940 171 -860 205
rect -940 137 -917 171
rect -883 137 -860 171
rect -940 103 -860 137
rect -940 69 -917 103
rect -883 69 -860 103
rect -940 40 -860 69
rect -790 962 -710 1000
rect -790 928 -767 962
rect -733 928 -710 962
rect -790 861 -710 928
rect -790 827 -767 861
rect -733 827 -710 861
rect -790 793 -710 827
rect -790 759 -767 793
rect -733 759 -710 793
rect -790 725 -710 759
rect -790 691 -767 725
rect -733 691 -710 725
rect -790 657 -710 691
rect -790 623 -767 657
rect -733 623 -710 657
rect -790 589 -710 623
rect -790 555 -767 589
rect -733 555 -710 589
rect -790 521 -710 555
rect -790 487 -767 521
rect -733 487 -710 521
rect -790 453 -710 487
rect -790 419 -767 453
rect -733 419 -710 453
rect -790 385 -710 419
rect -790 351 -767 385
rect -733 351 -710 385
rect -790 317 -710 351
rect -790 283 -767 317
rect -733 283 -710 317
rect -790 249 -710 283
rect -790 215 -767 249
rect -733 215 -710 249
rect -790 181 -710 215
rect -790 147 -767 181
rect -733 147 -710 181
rect -790 113 -710 147
rect -790 79 -767 113
rect -733 79 -710 113
rect -790 40 -710 79
rect -640 962 -560 1000
rect -640 928 -617 962
rect -583 928 -560 962
rect -640 861 -560 928
rect -640 827 -617 861
rect -583 827 -560 861
rect -640 793 -560 827
rect -640 759 -617 793
rect -583 759 -560 793
rect -640 725 -560 759
rect -640 691 -617 725
rect -583 691 -560 725
rect -640 657 -560 691
rect -640 623 -617 657
rect -583 623 -560 657
rect -640 589 -560 623
rect -640 555 -617 589
rect -583 555 -560 589
rect -640 521 -560 555
rect -640 487 -617 521
rect -583 487 -560 521
rect -640 453 -560 487
rect -640 419 -617 453
rect -583 419 -560 453
rect -640 385 -560 419
rect -640 351 -617 385
rect -583 351 -560 385
rect -640 317 -560 351
rect -640 283 -617 317
rect -583 283 -560 317
rect -640 249 -560 283
rect -640 215 -617 249
rect -583 215 -560 249
rect -640 181 -560 215
rect -640 147 -617 181
rect -583 147 -560 181
rect -640 113 -560 147
rect -640 79 -617 113
rect -583 79 -560 113
rect -640 40 -560 79
rect -490 962 -410 1000
rect -490 928 -467 962
rect -433 928 -410 962
rect -490 861 -410 928
rect -490 827 -467 861
rect -433 827 -410 861
rect -490 793 -410 827
rect -490 759 -467 793
rect -433 759 -410 793
rect -490 725 -410 759
rect -490 691 -467 725
rect -433 691 -410 725
rect -490 657 -410 691
rect -490 623 -467 657
rect -433 623 -410 657
rect -490 589 -410 623
rect -490 555 -467 589
rect -433 555 -410 589
rect -490 521 -410 555
rect -490 487 -467 521
rect -433 487 -410 521
rect -490 453 -410 487
rect -490 419 -467 453
rect -433 419 -410 453
rect -490 385 -410 419
rect -490 351 -467 385
rect -433 351 -410 385
rect -490 317 -410 351
rect -490 283 -467 317
rect -433 283 -410 317
rect -490 249 -410 283
rect -490 215 -467 249
rect -433 215 -410 249
rect -490 181 -410 215
rect -490 147 -467 181
rect -433 147 -410 181
rect -490 113 -410 147
rect -490 79 -467 113
rect -433 79 -410 113
rect -490 40 -410 79
rect -1070 0 -1030 40
rect -770 0 -730 40
rect -470 0 -430 40
rect -1070 -40 -430 0
<< end >>
