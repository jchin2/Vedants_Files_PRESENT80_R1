magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -150 -99 889 647
<< l67d20 >>
rect -130 -94 876 -54
rect -119 585 -102 602
rect 109 -54 126 0
rect 654 540 888 560
rect -150 602 889 642
<< l66d20 >>
rect 389 555 449 570
<< l66d44 >>
rect -100 -82 -83 -65
rect -66 -82 -49 -65
rect -32 -82 -15 -65
rect 3 -82 20 -65
rect 37 -82 54 -65
rect 71 -82 88 -65
rect 105 -82 122 -65
rect 139 -82 156 -65
rect 173 -82 190 -65
rect 207 -82 224 -65
rect 241 -82 258 -65
rect 275 -82 292 -65
rect 309 -82 326 -65
rect 343 -82 360 -65
rect 377 -82 394 -65
rect 411 -82 428 -65
rect 445 -82 462 -65
rect 479 -82 496 -65
rect 513 -82 530 -65
rect 549 -83 566 -66
rect 583 -83 600 -66
rect 617 -83 634 -66
rect 651 -83 668 -66
rect 685 -83 702 -66
rect 719 -83 736 -66
rect 753 -83 770 -66
rect 787 -83 804 -66
rect 821 -83 838 -66
<< l125d44 >>
rect 407 12 431 548
<< l67d44 >>
rect -119 614 -102 631
rect -83 614 -66 631
rect -47 614 -30 631
rect -11 614 6 631
rect 25 614 42 631
rect 61 614 78 631
rect 97 614 114 631
rect 133 614 150 631
rect 169 614 186 631
rect 205 614 222 631
rect 241 614 258 631
rect 277 614 294 631
rect 313 614 330 631
rect 349 614 366 631
rect 385 614 402 631
rect 421 614 438 631
rect 457 614 474 631
rect 493 614 510 631
rect 313 614 330 631
rect 349 614 366 631
rect 385 614 402 631
rect 421 614 438 631
rect 457 614 474 631
rect 493 614 510 631
rect 529 614 546 631
rect 565 614 582 631
rect 601 614 618 631
rect 637 614 654 631
rect 673 614 690 631
rect 709 614 726 631
rect 745 614 762 631
rect 781 614 798 631
rect 817 614 834 631
rect 853 614 870 631
rect 673 614 690 631
rect 709 614 726 631
rect 745 614 762 631
rect 781 614 798 631
rect 817 614 834 631
rect 853 614 870 631
rect -100 -82 -83 -65
rect -64 -82 -47 -65
rect -28 -82 -11 -65
rect 9 -82 26 -65
rect 45 -82 62 -65
rect 81 -82 98 -65
rect 117 -82 134 -65
rect 153 -82 170 -65
rect 189 -82 206 -65
rect 225 -82 242 -65
rect 261 -82 278 -65
rect 297 -82 314 -65
rect 333 -82 350 -65
rect 369 -82 386 -65
rect 405 -82 422 -65
rect 441 -82 458 -65
rect 477 -82 494 -65
rect 513 -82 530 -65
rect 549 -83 566 -66
rect 585 -83 602 -66
rect 621 -83 638 -66
rect 657 -83 674 -66
rect 693 -83 710 -66
rect 729 -83 746 -66
rect 765 -83 782 -66
rect 801 -83 818 -66
rect 837 -83 854 -66
<< l68d20 >>
rect -150 597 889 647
rect -130 -99 876 -49
<< l68d16 >>
rect 332 -82 350 -65
rect 313 614 330 631
<< l67d16 >>
rect 875 545 886 555
<< labels >>
rlabel l67d20 373 -74 373 -74 0 Ground
rlabel l68d16 341 -73.5 341 -73.5 0 Ground
rlabel l68d16 321.5 622 321.5 622 0 VDD
rlabel l67d16 880 550 880 550 0 Mirror_out
use nmos_1v8_lvt_5p0_body_4finger nmos_1v8_lvt_5p0_body_4finger_1
timestamp 1670961910
transform 1 0 644 0 1 20
box -628 -20 -183 550
use nmos_1v8_lvt_5p0_4finger nmos_1v8_lvt_5p0_4finger_1
timestamp 1670961910
transform 1 0 944 0 1 20
box -568 -20 -183 550
use Via_P_Licon_Li Via_P_Licon_Li_1
timestamp 1670961910
transform 1 0 0 0 1 0
box 184 552 217 585
use Li_res_185p223ohm Li_res_185p223ohm_1
timestamp 1670961910
transform 0 1 -239 -1 0 455
box -130 120 -113 423
<< end >>
