magic
tech sky130A
magscale 1 2
timestamp 1670967604
<< locali >>
rect -1630 1227 -250 1250
rect -1630 1193 -1597 1227
rect -1563 1193 -1517 1227
rect -1483 1193 -1437 1227
rect -1403 1193 -1357 1227
rect -1323 1193 -1277 1227
rect -1243 1193 -1197 1227
rect -1163 1193 -1117 1227
rect -1083 1193 -1037 1227
rect -1003 1193 -957 1227
rect -923 1193 -877 1227
rect -843 1193 -797 1227
rect -763 1193 -717 1227
rect -683 1193 -637 1227
rect -603 1193 -557 1227
rect -523 1193 -477 1227
rect -443 1193 -397 1227
rect -363 1193 -317 1227
rect -283 1193 -250 1227
rect -1630 1170 -250 1193
<< viali >>
rect -1597 1193 -1563 1227
rect -1517 1193 -1483 1227
rect -1437 1193 -1403 1227
rect -1357 1193 -1323 1227
rect -1277 1193 -1243 1227
rect -1197 1193 -1163 1227
rect -1117 1193 -1083 1227
rect -1037 1193 -1003 1227
rect -957 1193 -923 1227
rect -877 1193 -843 1227
rect -797 1193 -763 1227
rect -717 1193 -683 1227
rect -637 1193 -603 1227
rect -557 1193 -523 1227
rect -477 1193 -443 1227
rect -397 1193 -363 1227
rect -317 1193 -283 1227
<< metal1 >>
rect -1630 1227 -250 1260
rect -1630 1193 -1597 1227
rect -1563 1193 -1517 1227
rect -1483 1193 -1437 1227
rect -1403 1193 -1357 1227
rect -1323 1193 -1277 1227
rect -1243 1193 -1197 1227
rect -1163 1193 -1117 1227
rect -1083 1193 -1037 1227
rect -1003 1193 -957 1227
rect -923 1193 -877 1227
rect -843 1193 -797 1227
rect -763 1193 -717 1227
rect -683 1193 -637 1227
rect -603 1193 -557 1227
rect -523 1193 -477 1227
rect -443 1193 -397 1227
rect -363 1193 -317 1227
rect -283 1193 -250 1227
rect -1630 1160 -250 1193
<< end >>
