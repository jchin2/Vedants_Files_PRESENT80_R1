magic
tech sky130A
magscale 1 2
timestamp 1671080489
<< poly >>
rect -151 712 -3 714
rect -2606 -2003 -2506 -1939
rect -1726 -2099 -1626 -1939
rect -152 -2249 -52 -1971
rect 1388 -2171 1488 -1971
rect 2302 -2085 2402 -1939
rect 3182 -2003 3282 -1939
<< locali >>
rect -4865 1059 5702 1082
rect -4865 1025 -4804 1059
rect -4770 1025 -4732 1059
rect -4698 1025 -4660 1059
rect -4626 1025 -4588 1059
rect -4554 1025 -4516 1059
rect -4482 1025 -4444 1059
rect -4410 1025 -4372 1059
rect -4338 1025 -4300 1059
rect -4266 1025 -4228 1059
rect -4194 1025 -4156 1059
rect -4122 1025 -4084 1059
rect -4050 1025 -4012 1059
rect -3978 1025 -3940 1059
rect -3906 1025 -3868 1059
rect -3834 1025 -3796 1059
rect -3762 1025 -3724 1059
rect -3690 1025 -3652 1059
rect -3618 1025 -3580 1059
rect -3546 1025 -3485 1059
rect -3451 1025 -3413 1059
rect -3379 1025 -3341 1059
rect -3307 1025 -3269 1059
rect -3235 1025 -3197 1059
rect -3163 1025 -3125 1059
rect -3091 1025 -3053 1059
rect -3019 1025 -2981 1059
rect -2947 1025 -2909 1059
rect -2875 1025 -2837 1059
rect -2803 1025 -2765 1059
rect -2731 1025 -2693 1059
rect -2659 1025 -2621 1059
rect -2587 1025 -2549 1059
rect -2515 1025 -2477 1059
rect -2443 1025 -2405 1059
rect -2371 1025 -2333 1059
rect -2299 1025 -2261 1059
rect -2227 1025 -2189 1059
rect -2155 1025 -2117 1059
rect -2083 1025 -2045 1059
rect -2011 1025 -1973 1059
rect -1939 1025 -1901 1059
rect -1867 1025 -1829 1059
rect -1795 1025 -1757 1059
rect -1723 1025 -1685 1059
rect -1651 1025 -1613 1059
rect -1579 1025 -1541 1059
rect -1507 1025 -1469 1059
rect -1435 1025 -1397 1059
rect -1363 1025 -1325 1059
rect -1291 1025 -1253 1059
rect -1219 1025 -1181 1059
rect -1147 1025 -1109 1059
rect -1075 1025 -1037 1059
rect -1003 1025 -965 1059
rect -931 1025 -870 1059
rect -836 1025 -798 1059
rect -764 1025 -726 1059
rect -692 1025 -654 1059
rect -620 1025 -582 1059
rect -548 1025 -510 1059
rect -476 1025 -438 1059
rect -404 1025 -366 1059
rect -332 1025 -294 1059
rect -260 1025 -222 1059
rect -188 1025 -150 1059
rect -116 1025 -78 1059
rect -44 1025 -6 1059
rect 28 1025 66 1059
rect 100 1025 138 1059
rect 172 1025 210 1059
rect 244 1025 282 1059
rect 316 1025 354 1059
rect 388 1025 426 1059
rect 460 1025 498 1059
rect 532 1025 570 1059
rect 604 1025 642 1059
rect 676 1025 714 1059
rect 748 1025 786 1059
rect 820 1025 858 1059
rect 892 1025 930 1059
rect 964 1025 1002 1059
rect 1036 1025 1074 1059
rect 1108 1025 1146 1059
rect 1180 1025 1218 1059
rect 1252 1025 1290 1059
rect 1324 1025 1362 1059
rect 1396 1025 1434 1059
rect 1468 1025 1506 1059
rect 1540 1025 1578 1059
rect 1612 1025 1650 1059
rect 1684 1025 1745 1059
rect 1779 1025 1817 1059
rect 1851 1025 1889 1059
rect 1923 1025 1961 1059
rect 1995 1025 2033 1059
rect 2067 1025 2105 1059
rect 2139 1025 2177 1059
rect 2211 1025 2249 1059
rect 2283 1025 2321 1059
rect 2355 1025 2393 1059
rect 2427 1025 2465 1059
rect 2499 1025 2537 1059
rect 2571 1025 2609 1059
rect 2643 1025 2681 1059
rect 2715 1025 2753 1059
rect 2787 1025 2825 1059
rect 2859 1025 2897 1059
rect 2931 1025 2969 1059
rect 3003 1025 3041 1059
rect 3075 1025 3113 1059
rect 3147 1025 3185 1059
rect 3219 1025 3257 1059
rect 3291 1025 3329 1059
rect 3363 1025 3401 1059
rect 3435 1025 3473 1059
rect 3507 1025 3545 1059
rect 3579 1025 3617 1059
rect 3651 1025 3689 1059
rect 3723 1025 3761 1059
rect 3795 1025 3833 1059
rect 3867 1025 3905 1059
rect 3939 1025 3977 1059
rect 4011 1025 4049 1059
rect 4083 1025 4121 1059
rect 4155 1025 4193 1059
rect 4227 1025 4265 1059
rect 4299 1025 4360 1059
rect 4394 1025 4432 1059
rect 4466 1025 4504 1059
rect 4538 1025 4576 1059
rect 4610 1025 4648 1059
rect 4682 1025 4720 1059
rect 4754 1025 4792 1059
rect 4826 1025 4864 1059
rect 4898 1025 4936 1059
rect 4970 1025 5008 1059
rect 5042 1025 5080 1059
rect 5114 1025 5152 1059
rect 5186 1025 5224 1059
rect 5258 1025 5296 1059
rect 5330 1025 5368 1059
rect 5402 1025 5440 1059
rect 5474 1025 5512 1059
rect 5546 1025 5584 1059
rect 5618 1025 5702 1059
rect -4865 1002 5702 1025
rect -2500 714 -151 794
rect 596 564 744 1002
rect -2259 -1009 -2189 -511
rect -1186 -1009 -1106 -798
rect 196 -931 264 -396
rect 1075 -931 1143 -396
rect -923 -965 -12 -931
rect 1348 -965 2259 -931
rect -923 -1089 -889 -965
rect -2826 -2454 -2746 -1889
rect -826 -2454 -746 -1889
rect -292 -1921 -252 -1011
rect 1588 -1921 1628 -1011
rect 2225 -1093 2259 -965
rect 2442 -1009 2522 -907
rect 3527 -1009 3597 -511
rect 270 -2454 1070 -2001
rect 2082 -2454 2162 -1889
rect 4082 -2454 4162 -1889
rect -4866 -2477 5701 -2454
rect -4866 -2511 -4805 -2477
rect -4771 -2511 -4733 -2477
rect -4699 -2511 -4661 -2477
rect -4627 -2511 -4589 -2477
rect -4555 -2511 -4517 -2477
rect -4483 -2511 -4445 -2477
rect -4411 -2511 -4373 -2477
rect -4339 -2511 -4301 -2477
rect -4267 -2511 -4229 -2477
rect -4195 -2511 -4157 -2477
rect -4123 -2511 -4085 -2477
rect -4051 -2511 -4013 -2477
rect -3979 -2511 -3941 -2477
rect -3907 -2511 -3869 -2477
rect -3835 -2511 -3797 -2477
rect -3763 -2511 -3725 -2477
rect -3691 -2511 -3653 -2477
rect -3619 -2511 -3581 -2477
rect -3547 -2511 -3486 -2477
rect -3452 -2511 -3414 -2477
rect -3380 -2511 -3342 -2477
rect -3308 -2511 -3270 -2477
rect -3236 -2511 -3198 -2477
rect -3164 -2511 -3126 -2477
rect -3092 -2511 -3054 -2477
rect -3020 -2511 -2982 -2477
rect -2948 -2511 -2910 -2477
rect -2876 -2511 -2838 -2477
rect -2804 -2511 -2766 -2477
rect -2732 -2511 -2694 -2477
rect -2660 -2511 -2622 -2477
rect -2588 -2511 -2550 -2477
rect -2516 -2511 -2478 -2477
rect -2444 -2511 -2406 -2477
rect -2372 -2511 -2334 -2477
rect -2300 -2511 -2262 -2477
rect -2228 -2511 -2190 -2477
rect -2156 -2511 -2118 -2477
rect -2084 -2511 -2046 -2477
rect -2012 -2511 -1974 -2477
rect -1940 -2511 -1902 -2477
rect -1868 -2511 -1830 -2477
rect -1796 -2511 -1758 -2477
rect -1724 -2511 -1686 -2477
rect -1652 -2511 -1614 -2477
rect -1580 -2511 -1542 -2477
rect -1508 -2511 -1470 -2477
rect -1436 -2511 -1398 -2477
rect -1364 -2511 -1326 -2477
rect -1292 -2511 -1254 -2477
rect -1220 -2511 -1182 -2477
rect -1148 -2511 -1110 -2477
rect -1076 -2511 -1038 -2477
rect -1004 -2511 -966 -2477
rect -932 -2511 -871 -2477
rect -837 -2511 -799 -2477
rect -765 -2511 -727 -2477
rect -693 -2511 -655 -2477
rect -621 -2511 -583 -2477
rect -549 -2511 -511 -2477
rect -477 -2511 -439 -2477
rect -405 -2511 -367 -2477
rect -333 -2511 -295 -2477
rect -261 -2511 -223 -2477
rect -189 -2511 -151 -2477
rect -117 -2511 -79 -2477
rect -45 -2511 -7 -2477
rect 27 -2511 65 -2477
rect 99 -2511 137 -2477
rect 171 -2511 209 -2477
rect 243 -2511 281 -2477
rect 315 -2511 353 -2477
rect 387 -2511 425 -2477
rect 459 -2511 497 -2477
rect 531 -2511 569 -2477
rect 603 -2511 641 -2477
rect 675 -2511 713 -2477
rect 747 -2511 785 -2477
rect 819 -2511 857 -2477
rect 891 -2511 929 -2477
rect 963 -2511 1001 -2477
rect 1035 -2511 1073 -2477
rect 1107 -2511 1145 -2477
rect 1179 -2511 1217 -2477
rect 1251 -2511 1289 -2477
rect 1323 -2511 1361 -2477
rect 1395 -2511 1433 -2477
rect 1467 -2511 1505 -2477
rect 1539 -2511 1577 -2477
rect 1611 -2511 1649 -2477
rect 1683 -2511 1744 -2477
rect 1778 -2511 1816 -2477
rect 1850 -2511 1888 -2477
rect 1922 -2511 1960 -2477
rect 1994 -2511 2032 -2477
rect 2066 -2511 2104 -2477
rect 2138 -2511 2176 -2477
rect 2210 -2511 2248 -2477
rect 2282 -2511 2320 -2477
rect 2354 -2511 2392 -2477
rect 2426 -2511 2464 -2477
rect 2498 -2511 2536 -2477
rect 2570 -2511 2608 -2477
rect 2642 -2511 2680 -2477
rect 2714 -2511 2752 -2477
rect 2786 -2511 2824 -2477
rect 2858 -2511 2896 -2477
rect 2930 -2511 2968 -2477
rect 3002 -2511 3040 -2477
rect 3074 -2511 3112 -2477
rect 3146 -2511 3184 -2477
rect 3218 -2511 3256 -2477
rect 3290 -2511 3328 -2477
rect 3362 -2511 3400 -2477
rect 3434 -2511 3472 -2477
rect 3506 -2511 3544 -2477
rect 3578 -2511 3616 -2477
rect 3650 -2511 3688 -2477
rect 3722 -2511 3760 -2477
rect 3794 -2511 3832 -2477
rect 3866 -2511 3904 -2477
rect 3938 -2511 3976 -2477
rect 4010 -2511 4048 -2477
rect 4082 -2511 4120 -2477
rect 4154 -2511 4192 -2477
rect 4226 -2511 4264 -2477
rect 4298 -2511 4359 -2477
rect 4393 -2511 4431 -2477
rect 4465 -2511 4503 -2477
rect 4537 -2511 4575 -2477
rect 4609 -2511 4647 -2477
rect 4681 -2511 4719 -2477
rect 4753 -2511 4791 -2477
rect 4825 -2511 4863 -2477
rect 4897 -2511 4935 -2477
rect 4969 -2511 5007 -2477
rect 5041 -2511 5079 -2477
rect 5113 -2511 5151 -2477
rect 5185 -2511 5223 -2477
rect 5257 -2511 5295 -2477
rect 5329 -2511 5367 -2477
rect 5401 -2511 5439 -2477
rect 5473 -2511 5511 -2477
rect 5545 -2511 5583 -2477
rect 5617 -2511 5701 -2477
rect -4866 -2534 5701 -2511
<< viali >>
rect -4804 1025 -4770 1059
rect -4732 1025 -4698 1059
rect -4660 1025 -4626 1059
rect -4588 1025 -4554 1059
rect -4516 1025 -4482 1059
rect -4444 1025 -4410 1059
rect -4372 1025 -4338 1059
rect -4300 1025 -4266 1059
rect -4228 1025 -4194 1059
rect -4156 1025 -4122 1059
rect -4084 1025 -4050 1059
rect -4012 1025 -3978 1059
rect -3940 1025 -3906 1059
rect -3868 1025 -3834 1059
rect -3796 1025 -3762 1059
rect -3724 1025 -3690 1059
rect -3652 1025 -3618 1059
rect -3580 1025 -3546 1059
rect -3485 1025 -3451 1059
rect -3413 1025 -3379 1059
rect -3341 1025 -3307 1059
rect -3269 1025 -3235 1059
rect -3197 1025 -3163 1059
rect -3125 1025 -3091 1059
rect -3053 1025 -3019 1059
rect -2981 1025 -2947 1059
rect -2909 1025 -2875 1059
rect -2837 1025 -2803 1059
rect -2765 1025 -2731 1059
rect -2693 1025 -2659 1059
rect -2621 1025 -2587 1059
rect -2549 1025 -2515 1059
rect -2477 1025 -2443 1059
rect -2405 1025 -2371 1059
rect -2333 1025 -2299 1059
rect -2261 1025 -2227 1059
rect -2189 1025 -2155 1059
rect -2117 1025 -2083 1059
rect -2045 1025 -2011 1059
rect -1973 1025 -1939 1059
rect -1901 1025 -1867 1059
rect -1829 1025 -1795 1059
rect -1757 1025 -1723 1059
rect -1685 1025 -1651 1059
rect -1613 1025 -1579 1059
rect -1541 1025 -1507 1059
rect -1469 1025 -1435 1059
rect -1397 1025 -1363 1059
rect -1325 1025 -1291 1059
rect -1253 1025 -1219 1059
rect -1181 1025 -1147 1059
rect -1109 1025 -1075 1059
rect -1037 1025 -1003 1059
rect -965 1025 -931 1059
rect -870 1025 -836 1059
rect -798 1025 -764 1059
rect -726 1025 -692 1059
rect -654 1025 -620 1059
rect -582 1025 -548 1059
rect -510 1025 -476 1059
rect -438 1025 -404 1059
rect -366 1025 -332 1059
rect -294 1025 -260 1059
rect -222 1025 -188 1059
rect -150 1025 -116 1059
rect -78 1025 -44 1059
rect -6 1025 28 1059
rect 66 1025 100 1059
rect 138 1025 172 1059
rect 210 1025 244 1059
rect 282 1025 316 1059
rect 354 1025 388 1059
rect 426 1025 460 1059
rect 498 1025 532 1059
rect 570 1025 604 1059
rect 642 1025 676 1059
rect 714 1025 748 1059
rect 786 1025 820 1059
rect 858 1025 892 1059
rect 930 1025 964 1059
rect 1002 1025 1036 1059
rect 1074 1025 1108 1059
rect 1146 1025 1180 1059
rect 1218 1025 1252 1059
rect 1290 1025 1324 1059
rect 1362 1025 1396 1059
rect 1434 1025 1468 1059
rect 1506 1025 1540 1059
rect 1578 1025 1612 1059
rect 1650 1025 1684 1059
rect 1745 1025 1779 1059
rect 1817 1025 1851 1059
rect 1889 1025 1923 1059
rect 1961 1025 1995 1059
rect 2033 1025 2067 1059
rect 2105 1025 2139 1059
rect 2177 1025 2211 1059
rect 2249 1025 2283 1059
rect 2321 1025 2355 1059
rect 2393 1025 2427 1059
rect 2465 1025 2499 1059
rect 2537 1025 2571 1059
rect 2609 1025 2643 1059
rect 2681 1025 2715 1059
rect 2753 1025 2787 1059
rect 2825 1025 2859 1059
rect 2897 1025 2931 1059
rect 2969 1025 3003 1059
rect 3041 1025 3075 1059
rect 3113 1025 3147 1059
rect 3185 1025 3219 1059
rect 3257 1025 3291 1059
rect 3329 1025 3363 1059
rect 3401 1025 3435 1059
rect 3473 1025 3507 1059
rect 3545 1025 3579 1059
rect 3617 1025 3651 1059
rect 3689 1025 3723 1059
rect 3761 1025 3795 1059
rect 3833 1025 3867 1059
rect 3905 1025 3939 1059
rect 3977 1025 4011 1059
rect 4049 1025 4083 1059
rect 4121 1025 4155 1059
rect 4193 1025 4227 1059
rect 4265 1025 4299 1059
rect 4360 1025 4394 1059
rect 4432 1025 4466 1059
rect 4504 1025 4538 1059
rect 4576 1025 4610 1059
rect 4648 1025 4682 1059
rect 4720 1025 4754 1059
rect 4792 1025 4826 1059
rect 4864 1025 4898 1059
rect 4936 1025 4970 1059
rect 5008 1025 5042 1059
rect 5080 1025 5114 1059
rect 5152 1025 5186 1059
rect 5224 1025 5258 1059
rect 5296 1025 5330 1059
rect 5368 1025 5402 1059
rect 5440 1025 5474 1059
rect 5512 1025 5546 1059
rect 5584 1025 5618 1059
rect -2583 -966 -2549 -932
rect -1703 -966 -1669 -932
rect -2573 -2060 -2539 -2026
rect -1693 -2142 -1659 -2108
rect -119 -2306 -85 -2272
rect 1420 -2224 1454 -2190
rect 3212 -2060 3246 -2026
rect 2335 -2142 2369 -2108
rect -4805 -2511 -4771 -2477
rect -4733 -2511 -4699 -2477
rect -4661 -2511 -4627 -2477
rect -4589 -2511 -4555 -2477
rect -4517 -2511 -4483 -2477
rect -4445 -2511 -4411 -2477
rect -4373 -2511 -4339 -2477
rect -4301 -2511 -4267 -2477
rect -4229 -2511 -4195 -2477
rect -4157 -2511 -4123 -2477
rect -4085 -2511 -4051 -2477
rect -4013 -2511 -3979 -2477
rect -3941 -2511 -3907 -2477
rect -3869 -2511 -3835 -2477
rect -3797 -2511 -3763 -2477
rect -3725 -2511 -3691 -2477
rect -3653 -2511 -3619 -2477
rect -3581 -2511 -3547 -2477
rect -3486 -2511 -3452 -2477
rect -3414 -2511 -3380 -2477
rect -3342 -2511 -3308 -2477
rect -3270 -2511 -3236 -2477
rect -3198 -2511 -3164 -2477
rect -3126 -2511 -3092 -2477
rect -3054 -2511 -3020 -2477
rect -2982 -2511 -2948 -2477
rect -2910 -2511 -2876 -2477
rect -2838 -2511 -2804 -2477
rect -2766 -2511 -2732 -2477
rect -2694 -2511 -2660 -2477
rect -2622 -2511 -2588 -2477
rect -2550 -2511 -2516 -2477
rect -2478 -2511 -2444 -2477
rect -2406 -2511 -2372 -2477
rect -2334 -2511 -2300 -2477
rect -2262 -2511 -2228 -2477
rect -2190 -2511 -2156 -2477
rect -2118 -2511 -2084 -2477
rect -2046 -2511 -2012 -2477
rect -1974 -2511 -1940 -2477
rect -1902 -2511 -1868 -2477
rect -1830 -2511 -1796 -2477
rect -1758 -2511 -1724 -2477
rect -1686 -2511 -1652 -2477
rect -1614 -2511 -1580 -2477
rect -1542 -2511 -1508 -2477
rect -1470 -2511 -1436 -2477
rect -1398 -2511 -1364 -2477
rect -1326 -2511 -1292 -2477
rect -1254 -2511 -1220 -2477
rect -1182 -2511 -1148 -2477
rect -1110 -2511 -1076 -2477
rect -1038 -2511 -1004 -2477
rect -966 -2511 -932 -2477
rect -871 -2511 -837 -2477
rect -799 -2511 -765 -2477
rect -727 -2511 -693 -2477
rect -655 -2511 -621 -2477
rect -583 -2511 -549 -2477
rect -511 -2511 -477 -2477
rect -439 -2511 -405 -2477
rect -367 -2511 -333 -2477
rect -295 -2511 -261 -2477
rect -223 -2511 -189 -2477
rect -151 -2511 -117 -2477
rect -79 -2511 -45 -2477
rect -7 -2511 27 -2477
rect 65 -2511 99 -2477
rect 137 -2511 171 -2477
rect 209 -2511 243 -2477
rect 281 -2511 315 -2477
rect 353 -2511 387 -2477
rect 425 -2511 459 -2477
rect 497 -2511 531 -2477
rect 569 -2511 603 -2477
rect 641 -2511 675 -2477
rect 713 -2511 747 -2477
rect 785 -2511 819 -2477
rect 857 -2511 891 -2477
rect 929 -2511 963 -2477
rect 1001 -2511 1035 -2477
rect 1073 -2511 1107 -2477
rect 1145 -2511 1179 -2477
rect 1217 -2511 1251 -2477
rect 1289 -2511 1323 -2477
rect 1361 -2511 1395 -2477
rect 1433 -2511 1467 -2477
rect 1505 -2511 1539 -2477
rect 1577 -2511 1611 -2477
rect 1649 -2511 1683 -2477
rect 1744 -2511 1778 -2477
rect 1816 -2511 1850 -2477
rect 1888 -2511 1922 -2477
rect 1960 -2511 1994 -2477
rect 2032 -2511 2066 -2477
rect 2104 -2511 2138 -2477
rect 2176 -2511 2210 -2477
rect 2248 -2511 2282 -2477
rect 2320 -2511 2354 -2477
rect 2392 -2511 2426 -2477
rect 2464 -2511 2498 -2477
rect 2536 -2511 2570 -2477
rect 2608 -2511 2642 -2477
rect 2680 -2511 2714 -2477
rect 2752 -2511 2786 -2477
rect 2824 -2511 2858 -2477
rect 2896 -2511 2930 -2477
rect 2968 -2511 3002 -2477
rect 3040 -2511 3074 -2477
rect 3112 -2511 3146 -2477
rect 3184 -2511 3218 -2477
rect 3256 -2511 3290 -2477
rect 3328 -2511 3362 -2477
rect 3400 -2511 3434 -2477
rect 3472 -2511 3506 -2477
rect 3544 -2511 3578 -2477
rect 3616 -2511 3650 -2477
rect 3688 -2511 3722 -2477
rect 3760 -2511 3794 -2477
rect 3832 -2511 3866 -2477
rect 3904 -2511 3938 -2477
rect 3976 -2511 4010 -2477
rect 4048 -2511 4082 -2477
rect 4120 -2511 4154 -2477
rect 4192 -2511 4226 -2477
rect 4264 -2511 4298 -2477
rect 4359 -2511 4393 -2477
rect 4431 -2511 4465 -2477
rect 4503 -2511 4537 -2477
rect 4575 -2511 4609 -2477
rect 4647 -2511 4681 -2477
rect 4719 -2511 4753 -2477
rect 4791 -2511 4825 -2477
rect 4863 -2511 4897 -2477
rect 4935 -2511 4969 -2477
rect 5007 -2511 5041 -2477
rect 5079 -2511 5113 -2477
rect 5151 -2511 5185 -2477
rect 5223 -2511 5257 -2477
rect 5295 -2511 5329 -2477
rect 5367 -2511 5401 -2477
rect 5439 -2511 5473 -2477
rect 5511 -2511 5545 -2477
rect 5583 -2511 5617 -2477
<< metal1 >>
rect -4865 1059 5702 1092
rect -4865 1025 -4804 1059
rect -4770 1025 -4732 1059
rect -4698 1025 -4660 1059
rect -4626 1025 -4588 1059
rect -4554 1025 -4516 1059
rect -4482 1025 -4444 1059
rect -4410 1025 -4372 1059
rect -4338 1025 -4300 1059
rect -4266 1025 -4228 1059
rect -4194 1025 -4156 1059
rect -4122 1025 -4084 1059
rect -4050 1025 -4012 1059
rect -3978 1025 -3940 1059
rect -3906 1025 -3868 1059
rect -3834 1025 -3796 1059
rect -3762 1025 -3724 1059
rect -3690 1025 -3652 1059
rect -3618 1025 -3580 1059
rect -3546 1025 -3485 1059
rect -3451 1025 -3413 1059
rect -3379 1025 -3341 1059
rect -3307 1025 -3269 1059
rect -3235 1025 -3197 1059
rect -3163 1025 -3125 1059
rect -3091 1025 -3053 1059
rect -3019 1025 -2981 1059
rect -2947 1025 -2909 1059
rect -2875 1025 -2837 1059
rect -2803 1025 -2765 1059
rect -2731 1025 -2693 1059
rect -2659 1025 -2621 1059
rect -2587 1025 -2549 1059
rect -2515 1025 -2477 1059
rect -2443 1025 -2405 1059
rect -2371 1025 -2333 1059
rect -2299 1025 -2261 1059
rect -2227 1025 -2189 1059
rect -2155 1025 -2117 1059
rect -2083 1025 -2045 1059
rect -2011 1025 -1973 1059
rect -1939 1025 -1901 1059
rect -1867 1025 -1829 1059
rect -1795 1025 -1757 1059
rect -1723 1025 -1685 1059
rect -1651 1025 -1613 1059
rect -1579 1025 -1541 1059
rect -1507 1025 -1469 1059
rect -1435 1025 -1397 1059
rect -1363 1025 -1325 1059
rect -1291 1025 -1253 1059
rect -1219 1025 -1181 1059
rect -1147 1025 -1109 1059
rect -1075 1025 -1037 1059
rect -1003 1025 -965 1059
rect -931 1025 -870 1059
rect -836 1025 -798 1059
rect -764 1025 -726 1059
rect -692 1025 -654 1059
rect -620 1025 -582 1059
rect -548 1025 -510 1059
rect -476 1025 -438 1059
rect -404 1025 -366 1059
rect -332 1025 -294 1059
rect -260 1025 -222 1059
rect -188 1025 -150 1059
rect -116 1025 -78 1059
rect -44 1025 -6 1059
rect 28 1025 66 1059
rect 100 1025 138 1059
rect 172 1025 210 1059
rect 244 1025 282 1059
rect 316 1025 354 1059
rect 388 1025 426 1059
rect 460 1025 498 1059
rect 532 1025 570 1059
rect 604 1025 642 1059
rect 676 1025 714 1059
rect 748 1025 786 1059
rect 820 1025 858 1059
rect 892 1025 930 1059
rect 964 1025 1002 1059
rect 1036 1025 1074 1059
rect 1108 1025 1146 1059
rect 1180 1025 1218 1059
rect 1252 1025 1290 1059
rect 1324 1025 1362 1059
rect 1396 1025 1434 1059
rect 1468 1025 1506 1059
rect 1540 1025 1578 1059
rect 1612 1025 1650 1059
rect 1684 1025 1745 1059
rect 1779 1025 1817 1059
rect 1851 1025 1889 1059
rect 1923 1025 1961 1059
rect 1995 1025 2033 1059
rect 2067 1025 2105 1059
rect 2139 1025 2177 1059
rect 2211 1025 2249 1059
rect 2283 1025 2321 1059
rect 2355 1025 2393 1059
rect 2427 1025 2465 1059
rect 2499 1025 2537 1059
rect 2571 1025 2609 1059
rect 2643 1025 2681 1059
rect 2715 1025 2753 1059
rect 2787 1025 2825 1059
rect 2859 1025 2897 1059
rect 2931 1025 2969 1059
rect 3003 1025 3041 1059
rect 3075 1025 3113 1059
rect 3147 1025 3185 1059
rect 3219 1025 3257 1059
rect 3291 1025 3329 1059
rect 3363 1025 3401 1059
rect 3435 1025 3473 1059
rect 3507 1025 3545 1059
rect 3579 1025 3617 1059
rect 3651 1025 3689 1059
rect 3723 1025 3761 1059
rect 3795 1025 3833 1059
rect 3867 1025 3905 1059
rect 3939 1025 3977 1059
rect 4011 1025 4049 1059
rect 4083 1025 4121 1059
rect 4155 1025 4193 1059
rect 4227 1025 4265 1059
rect 4299 1025 4360 1059
rect 4394 1025 4432 1059
rect 4466 1025 4504 1059
rect 4538 1025 4576 1059
rect 4610 1025 4648 1059
rect 4682 1025 4720 1059
rect 4754 1025 4792 1059
rect 4826 1025 4864 1059
rect 4898 1025 4936 1059
rect 4970 1025 5008 1059
rect 5042 1025 5080 1059
rect 5114 1025 5152 1059
rect 5186 1025 5224 1059
rect 5258 1025 5296 1059
rect 5330 1025 5368 1059
rect 5402 1025 5440 1059
rect 5474 1025 5512 1059
rect 5546 1025 5584 1059
rect 5618 1025 5702 1059
rect -4865 992 5702 1025
rect -2962 740 -2580 768
rect -2249 485 -2199 992
rect 3537 485 3587 992
rect -1106 -774 3522 -746
rect -2962 -881 -2470 -853
rect -2184 -881 2442 -853
rect -2606 -932 -2526 -909
rect -2606 -936 -2583 -932
rect -2962 -964 -2583 -936
rect -2606 -966 -2583 -964
rect -2549 -966 -2526 -932
rect -2498 -937 -2470 -881
rect -1726 -932 -1646 -909
rect -1726 -937 -1703 -932
rect -2498 -965 -1703 -937
rect -2606 -989 -2526 -966
rect -1726 -966 -1703 -965
rect -1669 -966 -1646 -932
rect -1726 -989 -1646 -966
rect -2596 -2026 -2516 -2003
rect -2596 -2060 -2573 -2026
rect -2539 -2029 -2516 -2026
rect 3189 -2026 3269 -2003
rect 3189 -2029 3212 -2026
rect -2539 -2057 3212 -2029
rect -2539 -2060 -2516 -2057
rect -2596 -2083 -2516 -2060
rect 3189 -2060 3212 -2057
rect 3246 -2060 3269 -2026
rect 3189 -2083 3269 -2060
rect -1716 -2108 -1636 -2085
rect -1716 -2142 -1693 -2108
rect -1659 -2111 -1636 -2108
rect 2312 -2108 2392 -2085
rect 2312 -2111 2335 -2108
rect -1659 -2139 2335 -2111
rect -1659 -2142 -1636 -2139
rect -1716 -2165 -1636 -2142
rect 2312 -2142 2335 -2139
rect 2369 -2142 2392 -2108
rect 2312 -2165 2392 -2142
rect 1397 -2190 1477 -2167
rect 1397 -2193 1420 -2190
rect -2962 -2221 1420 -2193
rect 1397 -2224 1420 -2221
rect 1454 -2224 1477 -2190
rect 1397 -2247 1477 -2224
rect -142 -2272 -62 -2249
rect -142 -2276 -119 -2272
rect -2962 -2304 -119 -2276
rect -142 -2306 -119 -2304
rect -85 -2306 -62 -2272
rect -142 -2329 -62 -2306
rect -4866 -2477 5701 -2444
rect -4866 -2511 -4805 -2477
rect -4771 -2511 -4733 -2477
rect -4699 -2511 -4661 -2477
rect -4627 -2511 -4589 -2477
rect -4555 -2511 -4517 -2477
rect -4483 -2511 -4445 -2477
rect -4411 -2511 -4373 -2477
rect -4339 -2511 -4301 -2477
rect -4267 -2511 -4229 -2477
rect -4195 -2511 -4157 -2477
rect -4123 -2511 -4085 -2477
rect -4051 -2511 -4013 -2477
rect -3979 -2511 -3941 -2477
rect -3907 -2511 -3869 -2477
rect -3835 -2511 -3797 -2477
rect -3763 -2511 -3725 -2477
rect -3691 -2511 -3653 -2477
rect -3619 -2511 -3581 -2477
rect -3547 -2511 -3486 -2477
rect -3452 -2511 -3414 -2477
rect -3380 -2511 -3342 -2477
rect -3308 -2511 -3270 -2477
rect -3236 -2511 -3198 -2477
rect -3164 -2511 -3126 -2477
rect -3092 -2511 -3054 -2477
rect -3020 -2511 -2982 -2477
rect -2948 -2511 -2910 -2477
rect -2876 -2511 -2838 -2477
rect -2804 -2511 -2766 -2477
rect -2732 -2511 -2694 -2477
rect -2660 -2511 -2622 -2477
rect -2588 -2511 -2550 -2477
rect -2516 -2511 -2478 -2477
rect -2444 -2511 -2406 -2477
rect -2372 -2511 -2334 -2477
rect -2300 -2511 -2262 -2477
rect -2228 -2511 -2190 -2477
rect -2156 -2511 -2118 -2477
rect -2084 -2511 -2046 -2477
rect -2012 -2511 -1974 -2477
rect -1940 -2511 -1902 -2477
rect -1868 -2511 -1830 -2477
rect -1796 -2511 -1758 -2477
rect -1724 -2511 -1686 -2477
rect -1652 -2511 -1614 -2477
rect -1580 -2511 -1542 -2477
rect -1508 -2511 -1470 -2477
rect -1436 -2511 -1398 -2477
rect -1364 -2511 -1326 -2477
rect -1292 -2511 -1254 -2477
rect -1220 -2511 -1182 -2477
rect -1148 -2511 -1110 -2477
rect -1076 -2511 -1038 -2477
rect -1004 -2511 -966 -2477
rect -932 -2511 -871 -2477
rect -837 -2511 -799 -2477
rect -765 -2511 -727 -2477
rect -693 -2511 -655 -2477
rect -621 -2511 -583 -2477
rect -549 -2511 -511 -2477
rect -477 -2511 -439 -2477
rect -405 -2511 -367 -2477
rect -333 -2511 -295 -2477
rect -261 -2511 -223 -2477
rect -189 -2511 -151 -2477
rect -117 -2511 -79 -2477
rect -45 -2511 -7 -2477
rect 27 -2511 65 -2477
rect 99 -2511 137 -2477
rect 171 -2511 209 -2477
rect 243 -2511 281 -2477
rect 315 -2511 353 -2477
rect 387 -2511 425 -2477
rect 459 -2511 497 -2477
rect 531 -2511 569 -2477
rect 603 -2511 641 -2477
rect 675 -2511 713 -2477
rect 747 -2511 785 -2477
rect 819 -2511 857 -2477
rect 891 -2511 929 -2477
rect 963 -2511 1001 -2477
rect 1035 -2511 1073 -2477
rect 1107 -2511 1145 -2477
rect 1179 -2511 1217 -2477
rect 1251 -2511 1289 -2477
rect 1323 -2511 1361 -2477
rect 1395 -2511 1433 -2477
rect 1467 -2511 1505 -2477
rect 1539 -2511 1577 -2477
rect 1611 -2511 1649 -2477
rect 1683 -2511 1744 -2477
rect 1778 -2511 1816 -2477
rect 1850 -2511 1888 -2477
rect 1922 -2511 1960 -2477
rect 1994 -2511 2032 -2477
rect 2066 -2511 2104 -2477
rect 2138 -2511 2176 -2477
rect 2210 -2511 2248 -2477
rect 2282 -2511 2320 -2477
rect 2354 -2511 2392 -2477
rect 2426 -2511 2464 -2477
rect 2498 -2511 2536 -2477
rect 2570 -2511 2608 -2477
rect 2642 -2511 2680 -2477
rect 2714 -2511 2752 -2477
rect 2786 -2511 2824 -2477
rect 2858 -2511 2896 -2477
rect 2930 -2511 2968 -2477
rect 3002 -2511 3040 -2477
rect 3074 -2511 3112 -2477
rect 3146 -2511 3184 -2477
rect 3218 -2511 3256 -2477
rect 3290 -2511 3328 -2477
rect 3362 -2511 3400 -2477
rect 3434 -2511 3472 -2477
rect 3506 -2511 3544 -2477
rect 3578 -2511 3616 -2477
rect 3650 -2511 3688 -2477
rect 3722 -2511 3760 -2477
rect 3794 -2511 3832 -2477
rect 3866 -2511 3904 -2477
rect 3938 -2511 3976 -2477
rect 4010 -2511 4048 -2477
rect 4082 -2511 4120 -2477
rect 4154 -2511 4192 -2477
rect 4226 -2511 4264 -2477
rect 4298 -2511 4359 -2477
rect 4393 -2511 4431 -2477
rect 4465 -2511 4503 -2477
rect 4537 -2511 4575 -2477
rect 4609 -2511 4647 -2477
rect 4681 -2511 4719 -2477
rect 4753 -2511 4791 -2477
rect 4825 -2511 4863 -2477
rect 4897 -2511 4935 -2477
rect 4969 -2511 5007 -2477
rect 5041 -2511 5079 -2477
rect 5113 -2511 5151 -2477
rect 5185 -2511 5223 -2477
rect 5257 -2511 5295 -2477
rect 5329 -2511 5367 -2477
rect 5401 -2511 5439 -2477
rect 5473 -2511 5511 -2477
rect 5545 -2511 5583 -2477
rect 5617 -2511 5701 -2477
rect -4866 -2544 5701 -2511
<< via1 >>
rect -2250 -675 -2198 -623
rect 3536 -785 3588 -733
<< metal2 >>
rect -2432 -635 -2404 1150
rect -2432 -663 -2264 -635
rect 3522 -733 3602 -719
rect 3522 -785 3536 -733
rect 3588 -745 3602 -733
rect 3742 -745 3770 1150
rect 3588 -773 3770 -745
rect 3588 -785 3602 -773
rect 3522 -799 3602 -785
use CASCODE_pmos_1v8_lvt_4p75_4finger  CASCODE_pmos_1v8_lvt_4p75_4finger_0
timestamp 1671080489
transform 1 0 270 0 1 -443
box -753 -28 1549 1232
use Li_via_M1  Li_via_M1_0
timestamp 1671080489
transform 1 0 -2560 0 1 734
box -20 -20 60 60
use Li_via_M1  Li_via_M1_1
timestamp 1671080489
transform 1 0 3542 0 1 -779
box -20 -20 60 60
use Li_via_M1  Li_via_M1_2
timestamp 1671080489
transform 1 0 -1166 0 1 -779
box -20 -20 60 60
use Li_via_M1  Li_via_M1_3
timestamp 1671080489
transform 1 0 2462 0 1 -887
box -20 -20 60 60
use Li_via_M1  Li_via_M1_4
timestamp 1671080489
transform 1 0 -2244 0 1 -887
box -20 -20 60 60
use Li_via_M2  Li_via_M2_0
timestamp 1671080489
transform 1 0 -2244 0 1 -669
box -20 -20 60 60
use P_pcon_li_single  P_pcon_li_single_0
timestamp 1671080489
transform 1 0 -122 0 1 -2309
box -20 -20 60 60
use P_pcon_li_single  P_pcon_li_single_1
timestamp 1671080489
transform 1 0 1417 0 1 -2227
box -20 -20 60 60
use P_pcon_li_single  P_pcon_li_single_2
timestamp 1671080489
transform 1 0 -1706 0 1 -969
box -20 -20 60 60
use P_pcon_li_single  P_pcon_li_single_3
timestamp 1671080489
transform 1 0 2332 0 1 -2145
box -20 -20 60 60
use P_pcon_li_single  P_pcon_li_single_4
timestamp 1671080489
transform 1 0 -1696 0 1 -2145
box -20 -20 60 60
use P_pcon_li_single  P_pcon_li_single_5
timestamp 1671080489
transform 1 0 3209 0 1 -2063
box -20 -20 60 60
use P_pcon_li_single  P_pcon_li_single_6
timestamp 1671080489
transform 1 0 -2576 0 1 -2063
box -20 -20 60 60
use P_pcon_li_single  P_pcon_li_single_7
timestamp 1671080489
transform 1 0 -2586 0 1 -969
box -20 -20 60 60
use Poly_pcon_Li_double  Poly_pcon_Li_double_0
timestamp 1671080489
transform 1 0 -131 0 1 734
box -20 -20 128 60
use fuckthisresistor3  fuckthisresistor3_0
timestamp 1671080489
transform 1 0 4039 0 1 -10
box -512 -501 -442 501
use fuckthisresistor3  fuckthisresistor3_1
timestamp 1671080489
transform 1 0 -1747 0 1 -10
box -512 -501 -442 501
use nmos_1v8_lvt_4p2_body_4finger  nmos_1v8_lvt_4p2_body_4finger_0
timestamp 1671080489
transform -1 0 2412 0 1 -1969
box -1796 0 -624 980
use nmos_1v8_lvt_4p2_body_4finger  nmos_1v8_lvt_4p2_body_4finger_1
timestamp 1671080489
transform 1 0 3832 0 1 -1969
box -1796 0 -624 980
use nmos_1v8_lvt_4p2_body_4finger  nmos_1v8_lvt_4p2_body_4finger_2
timestamp 1671080489
transform -1 0 -2496 0 1 -1969
box -1796 0 -624 980
use nmos_1v8_lvt_4p2_body_4finger  nmos_1v8_lvt_4p2_body_4finger_3
timestamp 1671080489
transform 1 0 -1076 0 1 -1969
box -1796 0 -624 980
use nmos_1v8_lvt_4p75_body_4finger  nmos_1v8_lvt_4p75_body_4finger_0
timestamp 1671080489
transform -1 0 -382 0 1 -1961
box -2136 -40 -964 1050
use nmos_1v8_lvt_4p75_body_4finger  nmos_1v8_lvt_4p75_body_4finger_1
timestamp 1671080489
transform 1 0 1718 0 1 -1961
box -2136 -40 -964 1050
<< labels >>
flabel metal1 s -2949 746 -2934 759 2 FreeSans 100000 0 0 0 v_bias_p
port 1 nsew
flabel metal1 s 569 -2511 748 -2477 2 FreeSans 100000 0 0 0 Ground
port 2 nsew
flabel metal1 s 604 1025 642 1059 2 FreeSans 100000 0 0 0 VDD
port 3 nsew
flabel metal1 s -2953 -2298 -2938 -2282 2 FreeSans 100000 0 0 0 RFP
port 4 nsew
flabel metal1 s -2953 -2215 -2938 -2199 2 FreeSans 100000 0 0 0 RFN
port 5 nsew
flabel metal1 s -2949 -959 -2931 -942 2 FreeSans 100000 0 0 0 LOP
port 6 nsew
flabel metal1 s -2948 -876 -2930 -859 2 FreeSans 100000 0 0 0 LON
port 7 nsew
flabel metal2 s -2383 -655 -2367 -642 2 FreeSans 100000 0 0 0 VoutP
port 8 nsew
flabel metal2 s 3684 -767 3703 -750 2 FreeSans 100000 0 0 0 VoutN
port 9 nsew
<< properties >>
string path 18.780 -3.635 18.780 5.750 
<< end >>
