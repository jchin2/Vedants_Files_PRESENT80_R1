magic
tech sky130A
timestamp 1670863536
<< error_p >>
rect -680 225 -620 675
rect -605 225 -545 675
rect -530 225 -470 675
rect -455 225 -395 675
rect -380 225 -320 675
rect -305 225 -245 675
rect -230 225 -170 675
rect -155 225 -95 675
rect -80 225 -20 675
rect -5 225 55 675
rect 70 225 130 675
rect 145 225 205 675
rect 220 225 280 675
rect 295 225 355 675
rect 370 225 430 675
rect 445 225 505 675
rect 520 225 580 675
rect 595 225 655 675
rect 670 225 730 675
rect 745 225 805 675
rect 820 225 880 675
<< nmoslvt >>
rect -620 225 -605 675
rect -545 225 -530 675
rect -470 225 -455 675
rect -395 225 -380 675
rect -320 225 -305 675
rect -245 225 -230 675
rect -170 225 -155 675
rect -95 225 -80 675
rect -20 225 -5 675
rect 55 225 70 675
rect 130 225 145 675
rect 205 225 220 675
rect 280 225 295 675
rect 355 225 370 675
rect 430 225 445 675
rect 505 225 520 675
rect 580 225 595 675
rect 655 225 670 675
rect 730 225 745 675
rect 805 225 820 675
<< ndiff >>
rect -680 660 -620 675
rect -680 240 -660 660
rect -640 240 -620 660
rect -680 225 -620 240
rect -605 650 -545 675
rect -605 240 -585 650
rect -565 240 -545 650
rect -605 225 -545 240
rect -530 660 -470 675
rect -530 240 -510 660
rect -490 240 -470 660
rect -530 225 -470 240
rect -455 660 -395 675
rect -455 240 -435 660
rect -415 240 -395 660
rect -455 225 -395 240
rect -380 660 -320 675
rect -380 240 -360 660
rect -340 240 -320 660
rect -380 225 -320 240
rect -305 660 -245 675
rect -305 240 -285 660
rect -265 240 -245 660
rect -305 225 -245 240
rect -230 660 -170 675
rect -230 240 -210 660
rect -190 240 -170 660
rect -230 225 -170 240
rect -155 660 -95 675
rect -155 240 -135 660
rect -115 240 -95 660
rect -155 225 -95 240
rect -80 660 -20 675
rect -80 240 -60 660
rect -40 240 -20 660
rect -80 225 -20 240
rect -5 660 55 675
rect -5 240 15 660
rect 35 240 55 660
rect -5 225 55 240
rect 70 660 130 675
rect 70 240 90 660
rect 110 240 130 660
rect 70 225 130 240
rect 145 660 205 675
rect 145 250 165 660
rect 185 250 205 660
rect 145 225 205 250
rect 220 660 280 675
rect 220 240 240 660
rect 260 240 280 660
rect 220 225 280 240
rect 295 660 355 675
rect 295 240 315 660
rect 335 240 355 660
rect 295 225 355 240
rect 370 660 430 675
rect 370 240 390 660
rect 410 240 430 660
rect 370 225 430 240
rect 445 660 505 675
rect 445 240 465 660
rect 485 240 505 660
rect 445 225 505 240
rect 520 660 580 675
rect 520 240 540 660
rect 560 240 580 660
rect 520 225 580 240
rect 595 660 655 675
rect 595 240 615 660
rect 635 240 655 660
rect 595 225 655 240
rect 670 660 730 675
rect 670 240 690 660
rect 710 240 730 660
rect 670 225 730 240
rect 745 660 805 675
rect 745 240 765 660
rect 785 240 805 660
rect 745 225 805 240
rect 820 660 880 675
rect 820 240 840 660
rect 860 240 880 660
rect 820 225 880 240
<< ndiffc >>
rect -660 240 -640 660
rect -585 240 -565 650
rect -510 240 -490 660
rect -435 240 -415 660
rect -360 240 -340 660
rect -285 240 -265 660
rect -210 240 -190 660
rect -135 240 -115 660
rect -60 240 -40 660
rect 15 240 35 660
rect 90 240 110 660
rect 165 250 185 660
rect 240 240 260 660
rect 315 240 335 660
rect 390 240 410 660
rect 465 240 485 660
rect 540 240 560 660
rect 615 240 635 660
rect 690 240 710 660
rect 765 240 785 660
rect 840 240 860 660
<< poly >>
rect -620 700 70 715
rect -620 675 -605 700
rect -545 675 -530 700
rect -470 675 -455 700
rect -395 675 -380 700
rect -320 675 -305 700
rect -245 675 -230 700
rect -170 675 -155 700
rect -95 675 -80 700
rect -20 675 -5 700
rect 55 675 70 700
rect 130 675 145 690
rect 205 675 220 690
rect 280 675 295 690
rect 355 675 370 690
rect 430 675 445 690
rect 505 675 520 690
rect 580 675 595 690
rect 655 675 670 690
rect 730 675 745 690
rect 805 675 820 690
rect -620 210 -605 225
rect -545 210 -530 225
rect -470 210 -455 225
rect -395 210 -380 225
rect -320 210 -305 225
rect -245 210 -230 225
rect -170 210 -155 225
rect -95 210 -80 225
rect -20 210 -5 225
rect 55 210 70 225
rect 130 200 145 225
rect 205 200 220 225
rect 280 200 295 225
rect 355 200 370 225
rect 430 200 445 225
rect 505 200 520 225
rect 580 200 595 225
rect 655 200 670 225
rect 730 200 745 225
rect 805 200 820 225
rect 130 185 820 200
<< locali >>
rect -585 685 35 705
rect -585 665 -565 685
rect -435 665 -415 685
rect -285 665 -265 685
rect -135 665 -115 685
rect 15 665 35 685
rect 90 685 860 705
rect 90 665 110 685
rect 240 665 260 685
rect 390 665 410 685
rect 540 665 560 685
rect 690 665 710 685
rect 840 665 860 685
rect -670 660 -630 665
rect -670 240 -660 660
rect -640 240 -630 660
rect -670 235 -630 240
rect -595 650 -555 665
rect -595 240 -585 650
rect -565 240 -555 650
rect -595 235 -555 240
rect -520 660 -480 665
rect -520 240 -510 660
rect -490 240 -480 660
rect -520 235 -480 240
rect -445 660 -405 665
rect -445 240 -435 660
rect -415 240 -405 660
rect -445 235 -405 240
rect -370 660 -330 665
rect -370 240 -360 660
rect -340 240 -330 660
rect -370 235 -330 240
rect -295 660 -255 665
rect -295 240 -285 660
rect -265 240 -255 660
rect -295 235 -255 240
rect -220 660 -180 665
rect -220 240 -210 660
rect -190 240 -180 660
rect -220 235 -180 240
rect -145 660 -105 665
rect -145 240 -135 660
rect -115 240 -105 660
rect -145 235 -105 240
rect -70 660 -30 665
rect -70 240 -60 660
rect -40 240 -30 660
rect -70 235 -30 240
rect 5 660 45 665
rect 5 240 15 660
rect 35 240 45 660
rect 5 235 45 240
rect 80 660 120 665
rect 80 240 90 660
rect 110 240 120 660
rect 80 235 120 240
rect 155 660 195 665
rect 155 250 165 660
rect 185 250 195 660
rect 155 235 195 250
rect 230 660 270 665
rect 230 240 240 660
rect 260 240 270 660
rect 230 235 270 240
rect 305 660 345 665
rect 305 240 315 660
rect 335 240 345 660
rect 305 235 345 240
rect 380 660 420 665
rect 380 240 390 660
rect 410 240 420 660
rect 380 235 420 240
rect 455 660 495 665
rect 455 240 465 660
rect 485 240 495 660
rect 455 235 495 240
rect 530 660 570 665
rect 530 240 540 660
rect 560 240 570 660
rect 530 235 570 240
rect 605 660 645 665
rect 605 240 615 660
rect 635 240 645 660
rect 605 235 645 240
rect 680 660 720 665
rect 680 240 690 660
rect 710 240 720 660
rect 680 235 720 240
rect 755 660 795 665
rect 755 240 765 660
rect 785 240 795 660
rect 755 235 795 240
rect 830 660 870 665
rect 830 240 840 660
rect 860 240 870 660
rect 830 235 870 240
rect -660 215 -640 235
rect -510 215 -490 235
rect -360 215 -340 235
rect -210 215 -190 235
rect -60 215 -40 235
rect 90 215 110 235
rect -660 195 110 215
rect 165 215 185 235
rect 315 215 335 235
rect 465 215 485 235
rect 615 215 635 235
rect 765 215 785 235
rect 165 195 785 215
<< end >>
