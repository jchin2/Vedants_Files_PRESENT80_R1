magic
tech sky130A
magscale 1 2
timestamp 1672696580
<< nwell >>
rect -3110 1400 -710 1590
rect -2320 1010 -1500 1400
<< pwell >>
rect -3076 66 -744 506
rect -3096 -86 -724 66
<< nmos >>
rect -2930 180 -2900 480
rect -2780 180 -2750 480
rect -2630 180 -2600 480
rect -2480 180 -2450 480
rect -2150 180 -2120 480
rect -2000 180 -1970 480
rect -1850 180 -1820 480
rect -1700 180 -1670 480
rect -1370 180 -1340 480
rect -1220 180 -1190 480
rect -1070 180 -1040 480
rect -920 180 -890 480
<< pmos >>
rect -2150 1060 -2120 1360
rect -2000 1060 -1970 1360
rect -1850 1060 -1820 1360
rect -1700 1060 -1670 1360
<< ndiff >>
rect -3050 407 -2930 480
rect -3050 373 -3007 407
rect -2973 373 -2930 407
rect -3050 327 -2930 373
rect -3050 293 -3007 327
rect -2973 293 -2930 327
rect -3050 247 -2930 293
rect -3050 213 -3007 247
rect -2973 213 -2930 247
rect -3050 180 -2930 213
rect -2900 407 -2780 480
rect -2900 373 -2857 407
rect -2823 373 -2780 407
rect -2900 327 -2780 373
rect -2900 293 -2857 327
rect -2823 293 -2780 327
rect -2900 247 -2780 293
rect -2900 213 -2857 247
rect -2823 213 -2780 247
rect -2900 180 -2780 213
rect -2750 407 -2630 480
rect -2750 373 -2707 407
rect -2673 373 -2630 407
rect -2750 327 -2630 373
rect -2750 293 -2707 327
rect -2673 293 -2630 327
rect -2750 247 -2630 293
rect -2750 213 -2707 247
rect -2673 213 -2630 247
rect -2750 180 -2630 213
rect -2600 407 -2480 480
rect -2600 373 -2557 407
rect -2523 373 -2480 407
rect -2600 327 -2480 373
rect -2600 293 -2557 327
rect -2523 293 -2480 327
rect -2600 247 -2480 293
rect -2600 213 -2557 247
rect -2523 213 -2480 247
rect -2600 180 -2480 213
rect -2450 407 -2330 480
rect -2450 373 -2407 407
rect -2373 373 -2330 407
rect -2450 327 -2330 373
rect -2450 293 -2407 327
rect -2373 293 -2330 327
rect -2450 247 -2330 293
rect -2450 213 -2407 247
rect -2373 213 -2330 247
rect -2450 180 -2330 213
rect -2270 407 -2150 480
rect -2270 373 -2227 407
rect -2193 373 -2150 407
rect -2270 327 -2150 373
rect -2270 293 -2227 327
rect -2193 293 -2150 327
rect -2270 247 -2150 293
rect -2270 213 -2227 247
rect -2193 213 -2150 247
rect -2270 180 -2150 213
rect -2120 407 -2000 480
rect -2120 373 -2077 407
rect -2043 373 -2000 407
rect -2120 327 -2000 373
rect -2120 293 -2077 327
rect -2043 293 -2000 327
rect -2120 247 -2000 293
rect -2120 213 -2077 247
rect -2043 213 -2000 247
rect -2120 180 -2000 213
rect -1970 407 -1850 480
rect -1970 373 -1927 407
rect -1893 373 -1850 407
rect -1970 327 -1850 373
rect -1970 293 -1927 327
rect -1893 293 -1850 327
rect -1970 247 -1850 293
rect -1970 213 -1927 247
rect -1893 213 -1850 247
rect -1970 180 -1850 213
rect -1820 407 -1700 480
rect -1820 373 -1777 407
rect -1743 373 -1700 407
rect -1820 327 -1700 373
rect -1820 293 -1777 327
rect -1743 293 -1700 327
rect -1820 247 -1700 293
rect -1820 213 -1777 247
rect -1743 213 -1700 247
rect -1820 180 -1700 213
rect -1670 407 -1550 480
rect -1670 373 -1627 407
rect -1593 373 -1550 407
rect -1670 327 -1550 373
rect -1670 293 -1627 327
rect -1593 293 -1550 327
rect -1670 247 -1550 293
rect -1670 213 -1627 247
rect -1593 213 -1550 247
rect -1670 180 -1550 213
rect -1490 407 -1370 480
rect -1490 373 -1447 407
rect -1413 373 -1370 407
rect -1490 327 -1370 373
rect -1490 293 -1447 327
rect -1413 293 -1370 327
rect -1490 247 -1370 293
rect -1490 213 -1447 247
rect -1413 213 -1370 247
rect -1490 180 -1370 213
rect -1340 180 -1220 480
rect -1190 180 -1070 480
rect -1040 180 -920 480
rect -890 407 -770 480
rect -890 373 -847 407
rect -813 373 -770 407
rect -890 327 -770 373
rect -890 293 -847 327
rect -813 293 -770 327
rect -890 247 -770 293
rect -890 213 -847 247
rect -813 213 -770 247
rect -890 180 -770 213
<< pdiff >>
rect -2270 1287 -2150 1360
rect -2270 1253 -2227 1287
rect -2193 1253 -2150 1287
rect -2270 1207 -2150 1253
rect -2270 1173 -2227 1207
rect -2193 1173 -2150 1207
rect -2270 1127 -2150 1173
rect -2270 1093 -2227 1127
rect -2193 1093 -2150 1127
rect -2270 1060 -2150 1093
rect -2120 1287 -2000 1360
rect -2120 1253 -2077 1287
rect -2043 1253 -2000 1287
rect -2120 1207 -2000 1253
rect -2120 1173 -2077 1207
rect -2043 1173 -2000 1207
rect -2120 1127 -2000 1173
rect -2120 1093 -2077 1127
rect -2043 1093 -2000 1127
rect -2120 1060 -2000 1093
rect -1970 1287 -1850 1360
rect -1970 1253 -1927 1287
rect -1893 1253 -1850 1287
rect -1970 1207 -1850 1253
rect -1970 1173 -1927 1207
rect -1893 1173 -1850 1207
rect -1970 1127 -1850 1173
rect -1970 1093 -1927 1127
rect -1893 1093 -1850 1127
rect -1970 1060 -1850 1093
rect -1820 1287 -1700 1360
rect -1820 1253 -1777 1287
rect -1743 1253 -1700 1287
rect -1820 1207 -1700 1253
rect -1820 1173 -1777 1207
rect -1743 1173 -1700 1207
rect -1820 1127 -1700 1173
rect -1820 1093 -1777 1127
rect -1743 1093 -1700 1127
rect -1820 1060 -1700 1093
rect -1670 1287 -1550 1360
rect -1670 1253 -1627 1287
rect -1593 1253 -1550 1287
rect -1670 1207 -1550 1253
rect -1670 1173 -1627 1207
rect -1593 1173 -1550 1207
rect -1670 1127 -1550 1173
rect -1670 1093 -1627 1127
rect -1593 1093 -1550 1127
rect -1670 1060 -1550 1093
<< ndiffc >>
rect -3007 373 -2973 407
rect -3007 293 -2973 327
rect -3007 213 -2973 247
rect -2857 373 -2823 407
rect -2857 293 -2823 327
rect -2857 213 -2823 247
rect -2707 373 -2673 407
rect -2707 293 -2673 327
rect -2707 213 -2673 247
rect -2557 373 -2523 407
rect -2557 293 -2523 327
rect -2557 213 -2523 247
rect -2407 373 -2373 407
rect -2407 293 -2373 327
rect -2407 213 -2373 247
rect -2227 373 -2193 407
rect -2227 293 -2193 327
rect -2227 213 -2193 247
rect -2077 373 -2043 407
rect -2077 293 -2043 327
rect -2077 213 -2043 247
rect -1927 373 -1893 407
rect -1927 293 -1893 327
rect -1927 213 -1893 247
rect -1777 373 -1743 407
rect -1777 293 -1743 327
rect -1777 213 -1743 247
rect -1627 373 -1593 407
rect -1627 293 -1593 327
rect -1627 213 -1593 247
rect -1447 373 -1413 407
rect -1447 293 -1413 327
rect -1447 213 -1413 247
rect -847 373 -813 407
rect -847 293 -813 327
rect -847 213 -813 247
<< pdiffc >>
rect -2227 1253 -2193 1287
rect -2227 1173 -2193 1207
rect -2227 1093 -2193 1127
rect -2077 1253 -2043 1287
rect -2077 1173 -2043 1207
rect -2077 1093 -2043 1127
rect -1927 1253 -1893 1287
rect -1927 1173 -1893 1207
rect -1927 1093 -1893 1127
rect -1777 1253 -1743 1287
rect -1777 1173 -1743 1207
rect -1777 1093 -1743 1127
rect -1627 1253 -1593 1287
rect -1627 1173 -1593 1207
rect -1627 1093 -1593 1127
<< psubdiff >>
rect -3070 7 -750 40
rect -3070 -27 -3047 7
rect -3013 -27 -2967 7
rect -2933 -27 -2887 7
rect -2853 -27 -2807 7
rect -2773 -27 -2727 7
rect -2693 -27 -2647 7
rect -2613 -27 -2567 7
rect -2533 -27 -2487 7
rect -2453 -27 -2407 7
rect -2373 -27 -2327 7
rect -2293 -27 -2247 7
rect -2213 -27 -2167 7
rect -2133 -27 -2087 7
rect -2053 -27 -2007 7
rect -1973 -27 -1927 7
rect -1893 -27 -1847 7
rect -1813 -27 -1767 7
rect -1733 -27 -1687 7
rect -1653 -27 -1607 7
rect -1573 -27 -1527 7
rect -1493 -27 -1447 7
rect -1413 -27 -1367 7
rect -1333 -27 -1287 7
rect -1253 -27 -1207 7
rect -1173 -27 -1127 7
rect -1093 -27 -1047 7
rect -1013 -27 -967 7
rect -933 -27 -887 7
rect -853 -27 -807 7
rect -773 -27 -750 7
rect -3070 -60 -750 -27
<< nsubdiff >>
rect -3070 1507 -750 1540
rect -3070 1473 -3047 1507
rect -3013 1473 -2967 1507
rect -2933 1473 -2887 1507
rect -2853 1473 -2807 1507
rect -2773 1473 -2727 1507
rect -2693 1473 -2647 1507
rect -2613 1473 -2567 1507
rect -2533 1473 -2487 1507
rect -2453 1473 -2407 1507
rect -2373 1473 -2327 1507
rect -2293 1473 -2247 1507
rect -2213 1473 -2167 1507
rect -2133 1473 -2087 1507
rect -2053 1473 -2007 1507
rect -1973 1473 -1927 1507
rect -1893 1473 -1847 1507
rect -1813 1473 -1767 1507
rect -1733 1473 -1687 1507
rect -1653 1473 -1607 1507
rect -1573 1473 -1527 1507
rect -1493 1473 -1447 1507
rect -1413 1473 -1367 1507
rect -1333 1473 -1287 1507
rect -1253 1473 -1207 1507
rect -1173 1473 -1127 1507
rect -1093 1473 -1047 1507
rect -1013 1473 -967 1507
rect -933 1473 -887 1507
rect -853 1473 -807 1507
rect -773 1473 -750 1507
rect -3070 1440 -750 1473
<< psubdiffcont >>
rect -3047 -27 -3013 7
rect -2967 -27 -2933 7
rect -2887 -27 -2853 7
rect -2807 -27 -2773 7
rect -2727 -27 -2693 7
rect -2647 -27 -2613 7
rect -2567 -27 -2533 7
rect -2487 -27 -2453 7
rect -2407 -27 -2373 7
rect -2327 -27 -2293 7
rect -2247 -27 -2213 7
rect -2167 -27 -2133 7
rect -2087 -27 -2053 7
rect -2007 -27 -1973 7
rect -1927 -27 -1893 7
rect -1847 -27 -1813 7
rect -1767 -27 -1733 7
rect -1687 -27 -1653 7
rect -1607 -27 -1573 7
rect -1527 -27 -1493 7
rect -1447 -27 -1413 7
rect -1367 -27 -1333 7
rect -1287 -27 -1253 7
rect -1207 -27 -1173 7
rect -1127 -27 -1093 7
rect -1047 -27 -1013 7
rect -967 -27 -933 7
rect -887 -27 -853 7
rect -807 -27 -773 7
<< nsubdiffcont >>
rect -3047 1473 -3013 1507
rect -2967 1473 -2933 1507
rect -2887 1473 -2853 1507
rect -2807 1473 -2773 1507
rect -2727 1473 -2693 1507
rect -2647 1473 -2613 1507
rect -2567 1473 -2533 1507
rect -2487 1473 -2453 1507
rect -2407 1473 -2373 1507
rect -2327 1473 -2293 1507
rect -2247 1473 -2213 1507
rect -2167 1473 -2133 1507
rect -2087 1473 -2053 1507
rect -2007 1473 -1973 1507
rect -1927 1473 -1893 1507
rect -1847 1473 -1813 1507
rect -1767 1473 -1733 1507
rect -1687 1473 -1653 1507
rect -1607 1473 -1573 1507
rect -1527 1473 -1493 1507
rect -1447 1473 -1413 1507
rect -1367 1473 -1333 1507
rect -1287 1473 -1253 1507
rect -1207 1473 -1173 1507
rect -1127 1473 -1093 1507
rect -1047 1473 -1013 1507
rect -967 1473 -933 1507
rect -887 1473 -853 1507
rect -807 1473 -773 1507
<< poly >>
rect -2150 1390 -1970 1420
rect -2150 1360 -2120 1390
rect -2000 1360 -1970 1390
rect -1850 1390 -1670 1420
rect -1850 1360 -1820 1390
rect -1700 1360 -1670 1390
rect -2150 1030 -2120 1060
rect -2530 917 -2450 940
rect -2530 883 -2507 917
rect -2473 883 -2450 917
rect -2530 860 -2450 883
rect -2680 817 -2600 840
rect -2680 783 -2657 817
rect -2623 783 -2600 817
rect -2680 760 -2600 783
rect -2830 717 -2750 740
rect -2830 683 -2807 717
rect -2773 683 -2750 717
rect -2830 660 -2750 683
rect -2980 617 -2900 640
rect -2980 583 -2957 617
rect -2923 583 -2900 617
rect -2980 560 -2900 583
rect -2930 480 -2900 560
rect -2780 480 -2750 660
rect -2630 480 -2600 760
rect -2480 480 -2450 860
rect -2000 810 -1970 1060
rect -1850 940 -1820 1060
rect -1700 1030 -1670 1060
rect -1900 917 -1820 940
rect -1900 883 -1877 917
rect -1843 883 -1820 917
rect -1900 860 -1820 883
rect -2000 787 -1920 810
rect -2000 753 -1977 787
rect -1943 753 -1920 787
rect -2000 730 -1920 753
rect -2150 480 -2120 510
rect -2000 480 -1970 730
rect -1850 480 -1820 860
rect -1420 617 -1340 640
rect -1420 583 -1397 617
rect -1363 583 -1340 617
rect -1420 560 -1340 583
rect -1270 617 -1190 640
rect -1270 583 -1247 617
rect -1213 583 -1190 617
rect -1270 560 -1190 583
rect -1120 617 -1040 640
rect -1120 583 -1097 617
rect -1063 583 -1040 617
rect -1120 560 -1040 583
rect -970 617 -890 640
rect -970 583 -947 617
rect -913 583 -890 617
rect -970 560 -890 583
rect -1700 480 -1670 510
rect -1370 480 -1340 560
rect -1220 480 -1190 560
rect -1070 480 -1040 560
rect -920 480 -890 560
rect -2930 150 -2900 180
rect -2780 150 -2750 180
rect -2630 150 -2600 180
rect -2480 150 -2450 180
rect -2150 150 -2120 180
rect -2000 150 -1970 180
rect -1850 150 -1820 180
rect -1700 150 -1670 180
rect -1370 150 -1340 180
rect -1220 150 -1190 180
rect -1070 150 -1040 180
rect -920 150 -890 180
rect -2150 127 -2070 150
rect -2150 93 -2127 127
rect -2093 93 -2070 127
rect -2150 70 -2070 93
rect -1750 127 -1670 150
rect -1750 93 -1727 127
rect -1693 93 -1670 127
rect -1750 70 -1670 93
<< polycont >>
rect -2507 883 -2473 917
rect -2657 783 -2623 817
rect -2807 683 -2773 717
rect -2957 583 -2923 617
rect -1877 883 -1843 917
rect -1977 753 -1943 787
rect -1397 583 -1363 617
rect -1247 583 -1213 617
rect -1097 583 -1063 617
rect -947 583 -913 617
rect -2127 93 -2093 127
rect -1727 93 -1693 127
<< locali >>
rect -3070 1507 -750 1530
rect -3070 1473 -3047 1507
rect -3013 1473 -2967 1507
rect -2933 1473 -2887 1507
rect -2853 1473 -2807 1507
rect -2773 1473 -2727 1507
rect -2693 1473 -2647 1507
rect -2613 1473 -2567 1507
rect -2533 1473 -2487 1507
rect -2453 1473 -2407 1507
rect -2373 1473 -2327 1507
rect -2293 1473 -2247 1507
rect -2213 1473 -2167 1507
rect -2133 1473 -2087 1507
rect -2053 1473 -2007 1507
rect -1973 1473 -1927 1507
rect -1893 1473 -1847 1507
rect -1813 1473 -1767 1507
rect -1733 1473 -1687 1507
rect -1653 1473 -1607 1507
rect -1573 1473 -1527 1507
rect -1493 1473 -1447 1507
rect -1413 1473 -1367 1507
rect -1333 1473 -1287 1507
rect -1253 1473 -1207 1507
rect -1173 1473 -1127 1507
rect -1093 1473 -1047 1507
rect -1013 1473 -967 1507
rect -933 1473 -887 1507
rect -853 1473 -807 1507
rect -773 1473 -750 1507
rect -3070 1450 -750 1473
rect -2980 1380 -2900 1400
rect -3050 1377 -2900 1380
rect -3050 1343 -2957 1377
rect -2923 1343 -2900 1377
rect -3050 1340 -2900 1343
rect -2980 1320 -2900 1340
rect -2250 1287 -2170 1320
rect -2980 1260 -2900 1280
rect -3050 1257 -2900 1260
rect -3050 1223 -2957 1257
rect -2923 1223 -2900 1257
rect -3050 1220 -2900 1223
rect -2980 1200 -2900 1220
rect -2250 1253 -2227 1287
rect -2193 1253 -2170 1287
rect -2250 1207 -2170 1253
rect -2250 1173 -2227 1207
rect -2193 1173 -2170 1207
rect -2980 1140 -2900 1160
rect -3050 1137 -2900 1140
rect -3050 1103 -2957 1137
rect -2923 1103 -2900 1137
rect -3050 1100 -2900 1103
rect -2980 1080 -2900 1100
rect -2250 1127 -2170 1173
rect -2250 1093 -2227 1127
rect -2193 1093 -2170 1127
rect -2250 1070 -2170 1093
rect -2100 1287 -2020 1320
rect -2100 1253 -2077 1287
rect -2043 1253 -2020 1287
rect -2100 1207 -2020 1253
rect -2100 1173 -2077 1207
rect -2043 1173 -2020 1207
rect -2100 1127 -2020 1173
rect -2100 1093 -2077 1127
rect -2043 1093 -2020 1127
rect -2100 1060 -2020 1093
rect -1950 1287 -1870 1320
rect -1950 1253 -1927 1287
rect -1893 1253 -1870 1287
rect -1950 1207 -1870 1253
rect -1950 1173 -1927 1207
rect -1893 1173 -1870 1207
rect -1950 1127 -1870 1173
rect -1950 1093 -1927 1127
rect -1893 1093 -1870 1127
rect -1950 1070 -1870 1093
rect -1800 1287 -1720 1320
rect -1800 1253 -1777 1287
rect -1743 1253 -1720 1287
rect -1800 1207 -1720 1253
rect -1800 1173 -1777 1207
rect -1743 1173 -1720 1207
rect -1800 1127 -1720 1173
rect -1800 1093 -1777 1127
rect -1743 1093 -1720 1127
rect -1800 1060 -1720 1093
rect -1650 1287 -1570 1320
rect -1650 1253 -1627 1287
rect -1593 1253 -1570 1287
rect -1650 1207 -1570 1253
rect -1650 1173 -1627 1207
rect -1593 1173 -1570 1207
rect -1650 1127 -1570 1173
rect -1650 1093 -1627 1127
rect -1593 1093 -1570 1127
rect -1650 1070 -1570 1093
rect -2980 1020 -2900 1040
rect -3050 1017 -2900 1020
rect -3050 983 -2957 1017
rect -2923 983 -2900 1017
rect -3050 980 -2900 983
rect -2980 960 -2900 980
rect -2530 920 -2450 940
rect -3050 917 -2450 920
rect -3050 883 -2507 917
rect -2473 883 -2450 917
rect -3050 880 -2450 883
rect -2530 860 -2450 880
rect -2080 920 -2040 1060
rect -1900 920 -1820 940
rect -2080 917 -1820 920
rect -2080 883 -1877 917
rect -1843 883 -1820 917
rect -2080 880 -1820 883
rect -2680 820 -2600 840
rect -3050 817 -2600 820
rect -3050 783 -2657 817
rect -2623 783 -2600 817
rect -3050 780 -2600 783
rect -2680 760 -2600 780
rect -2830 720 -2750 740
rect -3050 717 -2750 720
rect -3050 683 -2807 717
rect -2773 683 -2750 717
rect -3050 680 -2750 683
rect -2830 660 -2750 680
rect -2980 620 -2900 640
rect -3050 617 -2900 620
rect -3050 583 -2957 617
rect -2923 583 -2900 617
rect -3050 580 -2900 583
rect -2980 560 -2900 580
rect -2080 520 -2040 880
rect -1900 860 -1820 880
rect -2000 800 -1920 810
rect -1780 800 -1740 1060
rect -1700 920 -1620 940
rect -1700 917 -770 920
rect -1700 883 -1677 917
rect -1643 883 -770 917
rect -1700 880 -770 883
rect -1700 860 -1620 880
rect -2000 787 -770 800
rect -2000 753 -1977 787
rect -1943 760 -770 787
rect -1943 753 -1920 760
rect -2000 730 -1920 753
rect -3010 480 -2040 520
rect -3010 440 -2970 480
rect -2710 440 -2670 480
rect -2410 440 -2370 480
rect -2080 440 -2040 480
rect -1780 520 -1740 760
rect -1420 617 -1340 640
rect -1420 583 -1397 617
rect -1363 583 -1340 617
rect -1420 560 -1340 583
rect -1270 617 -1190 640
rect -1270 583 -1247 617
rect -1213 583 -1190 617
rect -1270 560 -1190 583
rect -1120 617 -1040 640
rect -1120 583 -1097 617
rect -1063 583 -1040 617
rect -1120 560 -1040 583
rect -970 617 -890 640
rect -970 583 -947 617
rect -913 583 -890 617
rect -970 560 -890 583
rect -1780 480 -1430 520
rect -1780 440 -1740 480
rect -1470 440 -1430 480
rect -3030 407 -2950 440
rect -3030 373 -3007 407
rect -2973 373 -2950 407
rect -3030 327 -2950 373
rect -3030 293 -3007 327
rect -2973 293 -2950 327
rect -3030 247 -2950 293
rect -3030 213 -3007 247
rect -2973 213 -2950 247
rect -3030 190 -2950 213
rect -2880 407 -2800 440
rect -2880 373 -2857 407
rect -2823 373 -2800 407
rect -2880 327 -2800 373
rect -2880 293 -2857 327
rect -2823 293 -2800 327
rect -2880 247 -2800 293
rect -2880 213 -2857 247
rect -2823 213 -2800 247
rect -2880 190 -2800 213
rect -2730 407 -2650 440
rect -2730 373 -2707 407
rect -2673 373 -2650 407
rect -2730 327 -2650 373
rect -2730 293 -2707 327
rect -2673 293 -2650 327
rect -2730 247 -2650 293
rect -2730 213 -2707 247
rect -2673 213 -2650 247
rect -2730 190 -2650 213
rect -2580 407 -2500 440
rect -2580 373 -2557 407
rect -2523 373 -2500 407
rect -2580 327 -2500 373
rect -2580 293 -2557 327
rect -2523 293 -2500 327
rect -2580 247 -2500 293
rect -2580 213 -2557 247
rect -2523 213 -2500 247
rect -2580 190 -2500 213
rect -2430 407 -2350 440
rect -2430 373 -2407 407
rect -2373 373 -2350 407
rect -2430 327 -2350 373
rect -2430 293 -2407 327
rect -2373 293 -2350 327
rect -2430 247 -2350 293
rect -2430 213 -2407 247
rect -2373 213 -2350 247
rect -2430 190 -2350 213
rect -2250 407 -2170 440
rect -2250 373 -2227 407
rect -2193 373 -2170 407
rect -2250 327 -2170 373
rect -2250 293 -2227 327
rect -2193 293 -2170 327
rect -2250 247 -2170 293
rect -2250 213 -2227 247
rect -2193 213 -2170 247
rect -2250 190 -2170 213
rect -2100 407 -2020 440
rect -2100 373 -2077 407
rect -2043 373 -2020 407
rect -2100 327 -2020 373
rect -2100 293 -2077 327
rect -2043 293 -2020 327
rect -2100 247 -2020 293
rect -2100 213 -2077 247
rect -2043 213 -2020 247
rect -2100 190 -2020 213
rect -1950 407 -1870 440
rect -1950 373 -1927 407
rect -1893 373 -1870 407
rect -1950 327 -1870 373
rect -1950 293 -1927 327
rect -1893 293 -1870 327
rect -1950 247 -1870 293
rect -1950 213 -1927 247
rect -1893 213 -1870 247
rect -1950 190 -1870 213
rect -1800 407 -1720 440
rect -1800 373 -1777 407
rect -1743 373 -1720 407
rect -1800 327 -1720 373
rect -1800 293 -1777 327
rect -1743 293 -1720 327
rect -1800 247 -1720 293
rect -1800 213 -1777 247
rect -1743 213 -1720 247
rect -1800 190 -1720 213
rect -1650 407 -1570 440
rect -1650 373 -1627 407
rect -1593 373 -1570 407
rect -1650 327 -1570 373
rect -1650 293 -1627 327
rect -1593 293 -1570 327
rect -1650 247 -1570 293
rect -1650 213 -1627 247
rect -1593 213 -1570 247
rect -1650 190 -1570 213
rect -1470 407 -1390 440
rect -1470 373 -1447 407
rect -1413 373 -1390 407
rect -1470 327 -1390 373
rect -1470 293 -1447 327
rect -1413 293 -1390 327
rect -1470 247 -1390 293
rect -1470 213 -1447 247
rect -1413 213 -1390 247
rect -1470 190 -1390 213
rect -870 407 -790 440
rect -870 373 -847 407
rect -813 373 -790 407
rect -870 327 -790 373
rect -870 293 -847 327
rect -813 293 -790 327
rect -870 247 -790 293
rect -870 213 -847 247
rect -813 213 -790 247
rect -870 190 -790 213
rect -2150 130 -2070 150
rect -1750 130 -1670 150
rect -3050 127 -1670 130
rect -3050 93 -2127 127
rect -2093 93 -1727 127
rect -1693 93 -1670 127
rect -3050 90 -1670 93
rect -2150 70 -2070 90
rect -1750 70 -1670 90
rect -3070 7 -750 30
rect -3070 -27 -3047 7
rect -3013 -27 -2967 7
rect -2933 -27 -2887 7
rect -2853 -27 -2807 7
rect -2773 -27 -2727 7
rect -2693 -27 -2647 7
rect -2613 -27 -2567 7
rect -2533 -27 -2487 7
rect -2453 -27 -2407 7
rect -2373 -27 -2327 7
rect -2293 -27 -2247 7
rect -2213 -27 -2167 7
rect -2133 -27 -2087 7
rect -2053 -27 -2007 7
rect -1973 -27 -1927 7
rect -1893 -27 -1847 7
rect -1813 -27 -1767 7
rect -1733 -27 -1687 7
rect -1653 -27 -1607 7
rect -1573 -27 -1527 7
rect -1493 -27 -1447 7
rect -1413 -27 -1367 7
rect -1333 -27 -1287 7
rect -1253 -27 -1207 7
rect -1173 -27 -1127 7
rect -1093 -27 -1047 7
rect -1013 -27 -967 7
rect -933 -27 -887 7
rect -853 -27 -807 7
rect -773 -27 -750 7
rect -3070 -50 -750 -27
<< viali >>
rect -3047 1473 -3013 1507
rect -2967 1473 -2933 1507
rect -2887 1473 -2853 1507
rect -2807 1473 -2773 1507
rect -2727 1473 -2693 1507
rect -2647 1473 -2613 1507
rect -2567 1473 -2533 1507
rect -2487 1473 -2453 1507
rect -2407 1473 -2373 1507
rect -2327 1473 -2293 1507
rect -2247 1473 -2213 1507
rect -2167 1473 -2133 1507
rect -2087 1473 -2053 1507
rect -2007 1473 -1973 1507
rect -1927 1473 -1893 1507
rect -1847 1473 -1813 1507
rect -1767 1473 -1733 1507
rect -1687 1473 -1653 1507
rect -1607 1473 -1573 1507
rect -1527 1473 -1493 1507
rect -1447 1473 -1413 1507
rect -1367 1473 -1333 1507
rect -1287 1473 -1253 1507
rect -1207 1473 -1173 1507
rect -1127 1473 -1093 1507
rect -1047 1473 -1013 1507
rect -967 1473 -933 1507
rect -887 1473 -853 1507
rect -807 1473 -773 1507
rect -2957 1343 -2923 1377
rect -2957 1223 -2923 1257
rect -2227 1253 -2193 1287
rect -2227 1173 -2193 1207
rect -2957 1103 -2923 1137
rect -2227 1093 -2193 1127
rect -1927 1253 -1893 1287
rect -1927 1173 -1893 1207
rect -1927 1093 -1893 1127
rect -1627 1253 -1593 1287
rect -1627 1173 -1593 1207
rect -1627 1093 -1593 1127
rect -2957 983 -2923 1017
rect -1877 883 -1843 917
rect -1677 883 -1643 917
rect -1397 583 -1363 617
rect -1247 583 -1213 617
rect -1097 583 -1063 617
rect -947 583 -913 617
rect -2857 373 -2823 407
rect -2857 293 -2823 327
rect -2857 213 -2823 247
rect -2557 373 -2523 407
rect -2557 293 -2523 327
rect -2557 213 -2523 247
rect -2227 373 -2193 407
rect -2227 293 -2193 327
rect -2227 213 -2193 247
rect -1927 373 -1893 407
rect -1927 293 -1893 327
rect -1927 213 -1893 247
rect -1627 373 -1593 407
rect -1627 293 -1593 327
rect -1627 213 -1593 247
rect -847 373 -813 407
rect -847 293 -813 327
rect -847 213 -813 247
rect -3047 -27 -3013 7
rect -2967 -27 -2933 7
rect -2887 -27 -2853 7
rect -2807 -27 -2773 7
rect -2727 -27 -2693 7
rect -2647 -27 -2613 7
rect -2567 -27 -2533 7
rect -2487 -27 -2453 7
rect -2407 -27 -2373 7
rect -2327 -27 -2293 7
rect -2247 -27 -2213 7
rect -2167 -27 -2133 7
rect -2087 -27 -2053 7
rect -2007 -27 -1973 7
rect -1927 -27 -1893 7
rect -1847 -27 -1813 7
rect -1767 -27 -1733 7
rect -1687 -27 -1653 7
rect -1607 -27 -1573 7
rect -1527 -27 -1493 7
rect -1447 -27 -1413 7
rect -1367 -27 -1333 7
rect -1287 -27 -1253 7
rect -1207 -27 -1173 7
rect -1127 -27 -1093 7
rect -1047 -27 -1013 7
rect -967 -27 -933 7
rect -887 -27 -853 7
rect -807 -27 -773 7
<< metal1 >>
rect -3070 1507 -750 1540
rect -3070 1473 -3047 1507
rect -3013 1473 -2967 1507
rect -2933 1473 -2887 1507
rect -2853 1473 -2807 1507
rect -2773 1473 -2727 1507
rect -2693 1473 -2647 1507
rect -2613 1473 -2567 1507
rect -2533 1473 -2487 1507
rect -2453 1473 -2407 1507
rect -2373 1473 -2327 1507
rect -2293 1473 -2247 1507
rect -2213 1473 -2167 1507
rect -2133 1473 -2087 1507
rect -2053 1473 -2007 1507
rect -1973 1473 -1927 1507
rect -1893 1473 -1847 1507
rect -1813 1473 -1767 1507
rect -1733 1473 -1687 1507
rect -1653 1473 -1607 1507
rect -1573 1473 -1527 1507
rect -1493 1473 -1447 1507
rect -1413 1473 -1367 1507
rect -1333 1473 -1287 1507
rect -1253 1473 -1207 1507
rect -1173 1473 -1127 1507
rect -1093 1473 -1047 1507
rect -1013 1473 -967 1507
rect -933 1473 -887 1507
rect -853 1473 -807 1507
rect -773 1473 -750 1507
rect -3070 1440 -750 1473
rect -2980 1386 -2900 1400
rect -2980 1334 -2966 1386
rect -2914 1334 -2900 1386
rect -2980 1320 -2900 1334
rect -2980 1266 -2900 1280
rect -2980 1214 -2966 1266
rect -2914 1214 -2900 1266
rect -2980 1200 -2900 1214
rect -2980 1146 -2900 1160
rect -2980 1094 -2966 1146
rect -2914 1094 -2900 1146
rect -2980 1080 -2900 1094
rect -2980 1026 -2900 1040
rect -2980 974 -2966 1026
rect -2914 974 -2900 1026
rect -2980 960 -2900 974
rect -2860 440 -2820 1440
rect -2560 440 -2520 1440
rect -2250 1287 -2170 1440
rect -2250 1253 -2227 1287
rect -2193 1253 -2170 1287
rect -2250 1207 -2170 1253
rect -2250 1173 -2227 1207
rect -2193 1173 -2170 1207
rect -2250 1127 -2170 1173
rect -2250 1093 -2227 1127
rect -2193 1093 -2170 1127
rect -2250 1070 -2170 1093
rect -1950 1287 -1870 1440
rect -1950 1253 -1927 1287
rect -1893 1253 -1870 1287
rect -1950 1207 -1870 1253
rect -1950 1173 -1927 1207
rect -1893 1173 -1870 1207
rect -1950 1127 -1870 1173
rect -1950 1093 -1927 1127
rect -1893 1093 -1870 1127
rect -1950 1070 -1870 1093
rect -1650 1287 -1570 1440
rect -970 1386 -890 1400
rect -970 1334 -956 1386
rect -904 1334 -890 1386
rect -970 1320 -890 1334
rect -1650 1253 -1627 1287
rect -1593 1253 -1570 1287
rect -1650 1207 -1570 1253
rect -1650 1173 -1627 1207
rect -1593 1173 -1570 1207
rect -1120 1266 -1040 1280
rect -1120 1214 -1106 1266
rect -1054 1214 -1040 1266
rect -1120 1200 -1040 1214
rect -1650 1127 -1570 1173
rect -1650 1093 -1627 1127
rect -1593 1093 -1570 1127
rect -1650 1070 -1570 1093
rect -1270 1146 -1190 1160
rect -1270 1094 -1256 1146
rect -1204 1094 -1190 1146
rect -1270 1080 -1190 1094
rect -1420 1026 -1340 1040
rect -1420 974 -1406 1026
rect -1354 974 -1340 1026
rect -1420 960 -1340 974
rect -1900 920 -1820 940
rect -1700 920 -1620 940
rect -1900 917 -1620 920
rect -1900 883 -1877 917
rect -1843 883 -1677 917
rect -1643 883 -1620 917
rect -1900 880 -1620 883
rect -1900 860 -1820 880
rect -1700 860 -1620 880
rect -1400 640 -1360 960
rect -1250 640 -1210 1080
rect -1100 640 -1060 1200
rect -950 640 -910 1320
rect -1420 617 -1340 640
rect -1420 583 -1397 617
rect -1363 583 -1340 617
rect -1420 560 -1340 583
rect -1270 617 -1190 640
rect -1270 583 -1247 617
rect -1213 583 -1190 617
rect -1270 560 -1190 583
rect -1120 617 -1040 640
rect -1120 583 -1097 617
rect -1063 583 -1040 617
rect -1120 560 -1040 583
rect -970 617 -890 640
rect -970 583 -947 617
rect -913 583 -890 617
rect -970 560 -890 583
rect -850 440 -810 1440
rect -2880 407 -2800 440
rect -2880 373 -2857 407
rect -2823 373 -2800 407
rect -2880 327 -2800 373
rect -2880 293 -2857 327
rect -2823 293 -2800 327
rect -2880 247 -2800 293
rect -2880 213 -2857 247
rect -2823 213 -2800 247
rect -2880 190 -2800 213
rect -2580 407 -2500 440
rect -2580 373 -2557 407
rect -2523 373 -2500 407
rect -2580 327 -2500 373
rect -2580 293 -2557 327
rect -2523 293 -2500 327
rect -2580 247 -2500 293
rect -2580 213 -2557 247
rect -2523 213 -2500 247
rect -2580 190 -2500 213
rect -2250 407 -2170 440
rect -2250 373 -2227 407
rect -2193 373 -2170 407
rect -2250 327 -2170 373
rect -2250 293 -2227 327
rect -2193 293 -2170 327
rect -2250 247 -2170 293
rect -2250 213 -2227 247
rect -2193 213 -2170 247
rect -2250 190 -2170 213
rect -1950 407 -1870 440
rect -1950 373 -1927 407
rect -1893 373 -1870 407
rect -1950 327 -1870 373
rect -1950 293 -1927 327
rect -1893 293 -1870 327
rect -1950 247 -1870 293
rect -1950 213 -1927 247
rect -1893 213 -1870 247
rect -1950 190 -1870 213
rect -1650 407 -1570 440
rect -1650 373 -1627 407
rect -1593 373 -1570 407
rect -1650 327 -1570 373
rect -1650 293 -1627 327
rect -1593 293 -1570 327
rect -1650 247 -1570 293
rect -1650 213 -1627 247
rect -1593 213 -1570 247
rect -1650 190 -1570 213
rect -870 407 -790 440
rect -870 373 -847 407
rect -813 373 -790 407
rect -870 327 -790 373
rect -870 293 -847 327
rect -813 293 -790 327
rect -870 247 -790 293
rect -870 213 -847 247
rect -813 213 -790 247
rect -870 190 -790 213
rect -2230 40 -2190 190
rect -1930 40 -1890 190
rect -1630 40 -1590 190
rect -3070 7 -750 40
rect -3070 -27 -3047 7
rect -3013 -27 -2967 7
rect -2933 -27 -2887 7
rect -2853 -27 -2807 7
rect -2773 -27 -2727 7
rect -2693 -27 -2647 7
rect -2613 -27 -2567 7
rect -2533 -27 -2487 7
rect -2453 -27 -2407 7
rect -2373 -27 -2327 7
rect -2293 -27 -2247 7
rect -2213 -27 -2167 7
rect -2133 -27 -2087 7
rect -2053 -27 -2007 7
rect -1973 -27 -1927 7
rect -1893 -27 -1847 7
rect -1813 -27 -1767 7
rect -1733 -27 -1687 7
rect -1653 -27 -1607 7
rect -1573 -27 -1527 7
rect -1493 -27 -1447 7
rect -1413 -27 -1367 7
rect -1333 -27 -1287 7
rect -1253 -27 -1207 7
rect -1173 -27 -1127 7
rect -1093 -27 -1047 7
rect -1013 -27 -967 7
rect -933 -27 -887 7
rect -853 -27 -807 7
rect -773 -27 -750 7
rect -3070 -60 -750 -27
<< via1 >>
rect -2966 1377 -2914 1386
rect -2966 1343 -2957 1377
rect -2957 1343 -2923 1377
rect -2923 1343 -2914 1377
rect -2966 1334 -2914 1343
rect -2966 1257 -2914 1266
rect -2966 1223 -2957 1257
rect -2957 1223 -2923 1257
rect -2923 1223 -2914 1257
rect -2966 1214 -2914 1223
rect -2966 1137 -2914 1146
rect -2966 1103 -2957 1137
rect -2957 1103 -2923 1137
rect -2923 1103 -2914 1137
rect -2966 1094 -2914 1103
rect -2966 1017 -2914 1026
rect -2966 983 -2957 1017
rect -2957 983 -2923 1017
rect -2923 983 -2914 1017
rect -2966 974 -2914 983
rect -956 1334 -904 1386
rect -1106 1214 -1054 1266
rect -1256 1094 -1204 1146
rect -1406 974 -1354 1026
<< metal2 >>
rect -2980 1386 -2900 1400
rect -2980 1334 -2966 1386
rect -2914 1380 -2900 1386
rect -970 1386 -890 1400
rect -970 1380 -956 1386
rect -2914 1340 -956 1380
rect -2914 1334 -2900 1340
rect -2980 1320 -2900 1334
rect -970 1334 -956 1340
rect -904 1334 -890 1386
rect -970 1320 -890 1334
rect -2980 1266 -2900 1280
rect -2980 1214 -2966 1266
rect -2914 1260 -2900 1266
rect -1120 1266 -1040 1280
rect -1120 1260 -1106 1266
rect -2914 1220 -1106 1260
rect -2914 1214 -2900 1220
rect -2980 1200 -2900 1214
rect -1120 1214 -1106 1220
rect -1054 1214 -1040 1266
rect -1120 1200 -1040 1214
rect -2980 1146 -2900 1160
rect -2980 1094 -2966 1146
rect -2914 1140 -2900 1146
rect -1270 1146 -1190 1160
rect -1270 1140 -1256 1146
rect -2914 1100 -1256 1140
rect -2914 1094 -2900 1100
rect -2980 1080 -2900 1094
rect -1270 1094 -1256 1100
rect -1204 1094 -1190 1146
rect -1270 1080 -1190 1094
rect -2980 1026 -2900 1040
rect -2980 974 -2966 1026
rect -2914 1020 -2900 1026
rect -1420 1026 -1340 1040
rect -1420 1020 -1406 1026
rect -2914 980 -1406 1020
rect -2914 974 -2900 980
rect -2980 960 -2900 974
rect -1420 974 -1406 980
rect -1354 974 -1340 1026
rect -1420 960 -1340 974
<< labels >>
rlabel locali s -1980 750 -1940 790 4 OUT
port 1 nsew
rlabel locali s -3040 1350 -3020 1370 4 A
port 2 nsew
rlabel locali s -3040 890 -3020 910 4 A_bar
port 3 nsew
rlabel locali s -3040 1230 -3020 1250 4 B
port 4 nsew
rlabel locali s -3040 790 -3020 810 4 B_bar
port 5 nsew
rlabel locali s -3040 1110 -3020 1130 4 C
port 6 nsew
rlabel locali s -3040 690 -3020 710 4 C_bar
port 7 nsew
rlabel locali s -3040 990 -3020 1010 4 D
port 8 nsew
rlabel locali s -3040 590 -3020 610 4 D_bar
port 9 nsew
rlabel locali s -2130 90 -2090 130 4 Dis
port 10 nsew
rlabel metal1 s -1880 880 -1840 920 4 OUT_bar
port 11 nsew
rlabel metal1 s -1930 -30 -1890 10 4 GND!
port 12 nsew
rlabel metal1 s -1930 1470 -1890 1510 4 CLK
port 13 nsew
<< properties >>
string path -8.800 2.200 -8.800 2.400 
<< end >>
