magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect 0 0 38125 45587
use CASCODED_nmos_1v8_lvt_4p5_10finger CASCODED_nmos_1v8_lvt_4p5_10finger_1
timestamp 1670961910
transform 1 0 1795 0 1 -105
box -1795 105 -150 635
use Ground_rail Ground_rail_1
timestamp 1670961910
transform 1 0 805 0 1 531
box -805 0 -115 50
use Li_res_185p223ohm Li_res_185p223ohm_1
timestamp 1670961910
transform 1 0 130 0 1 461
box -130 120 -113 423
use Li_via_M2 Li_via_M2_1
timestamp 1670961910
transform 1 0 10 0 1 894
box -10 -10 30 30
use M1_vias_M4 M1_vias_M4_1
timestamp 1670961910
transform 1 0 240 0 1 1009
box -240 -85 -110 45
use Resistor_20k Resistor_20k_1
timestamp 1670961910
transform 1 0 -515 0 1 729
box 515 325 1119 866
use Square_Inductor_10t_2s_1w_180dout Square_Inductor_10t_2s_1w_180dout_1
timestamp 1670961910
transform 1 0 2530 0 1 4285
box -2530 -2690 15070 14910
use TOP TOP_1
timestamp 1670961910
transform 1 0 18949 0 1 17513
box -18949 1682 19176 23236
use Vdd_power_rail Vdd_power_rail_1
timestamp 1670961910
transform 1 0 815 0 1 40169
box -815 580 -125 630
use Via_P_Licon_Li Via_P_Licon_Li_1
timestamp 1670961910
transform 1 0 -184 0 1 40247
box 184 552 217 585
use nmos_1v8_lvt_4p5_10finger nmos_1v8_lvt_4p5_10finger_1
timestamp 1670961910
transform 1 0 -28 0 1 40847
box 28 -15 863 505
use nmos_1v8_lvt_4p5_10fingerx241 nmos_1v8_lvt_4p5_10fingerx241_1
timestamp 1670961910
transform 1 0 -28 0 1 41355
box 28 -3 863 490
use nmos_1v8_lvt_4p5_10fingerx241x241 nmos_1v8_lvt_4p5_10fingerx241x241_1
timestamp 1670961910
transform 1 0 -28 0 1 41848
box 28 -3 863 490
use nmos_1v8_lvt_4p5_body_10fingerx242 nmos_1v8_lvt_4p5_body_10fingerx242_1
timestamp 1670961910
transform 1 0 33 0 1 42353
box -33 -15 863 505
use nmos_1v8_lvt_5p0_4finger nmos_1v8_lvt_5p0_4finger_1
timestamp 1670961910
transform 1 0 568 0 1 42878
box -568 -20 -183 550
use nmos_1v8_lvt_5p0_body_4finger nmos_1v8_lvt_5p0_body_4finger_1
timestamp 1670961910
transform 1 0 628 0 1 43448
box -628 -20 -183 550
use simple_current_mirror simple_current_mirror_1
timestamp 1670961910
transform 1 0 150 0 1 44096
box -150 -99 889 647
use sky130_fd_pr__res_generic_l1_PK88MT sky130_fd_pr__res_generic_l1_PK88MT_1
timestamp 1670961910
transform 1 0 9 0 1 44895
box -9 -152 9 152
use sky130_fd_pr__res_xhigh_po_0p35_2RLX6B sky130_fd_pr__res_xhigh_po_0p35_2RLX6B_1
timestamp 1670961910
transform 1 0 302 0 1 45317
box -302 -271 302 271
<< end >>
