magic
tech sky130A
magscale 1 2
timestamp 1675457615
<< nwell >>
rect 980 2371 3340 2561
rect 3600 2371 5360 2561
rect 5620 2371 7380 2561
rect 1750 1981 2570 2371
rect 4070 1981 4890 2371
rect 6090 1981 6910 2371
rect 1750 191 2570 581
rect 4070 191 4890 581
rect 6090 191 6910 581
rect 1280 1 3040 191
rect 3600 1 5360 191
rect 5620 1 7380 191
rect 980 -449 3340 -259
rect 3600 -449 5090 -259
rect 5350 -449 7110 -259
rect 1750 -839 2570 -449
rect 3940 -839 4760 -449
rect 5820 -839 6640 -449
rect 1750 -2629 2570 -2239
rect 3940 -2629 4760 -2239
rect 5820 -2629 6640 -2239
rect 980 -2819 3340 -2629
rect 3600 -2819 5090 -2629
rect 5350 -2819 7110 -2629
rect 1121 -3269 3201 -3079
rect 3461 -3269 4951 -3079
rect 1751 -3659 2571 -3269
rect 3801 -3659 4621 -3269
rect 5211 -3270 7291 -3080
rect 5841 -3660 6661 -3270
rect 1790 -5849 2610 -5459
rect 4001 -5530 4821 -5140
rect 6060 -5530 6880 -5140
rect 3661 -5720 5151 -5530
rect 5430 -5720 7510 -5530
rect 980 -6170 3400 -5849
rect 3660 -6170 5150 -5980
rect 5409 -6170 7169 -5980
rect 1790 -6560 2610 -6170
rect 4000 -6560 4820 -6170
rect 5879 -6560 6699 -6170
rect 1790 -8350 2610 -7960
rect 4000 -8350 4820 -7960
rect 5879 -8350 6699 -7960
rect 1020 -8540 3380 -8350
rect 3660 -8540 5150 -8350
rect 5409 -8540 7169 -8350
rect 980 -8990 3340 -8800
rect 3600 -8990 5090 -8800
rect 5350 -8990 7110 -8800
rect 1750 -9380 2570 -8990
rect 3940 -9380 4760 -8990
rect 5820 -9380 6640 -8990
rect 1750 -11170 2570 -10780
rect 3940 -11170 4760 -10780
rect 5820 -11170 6640 -10780
rect 980 -11360 3340 -11170
rect 3600 -11360 5090 -11170
rect 5350 -11360 7110 -11170
rect 1121 -11810 3201 -11620
rect 3461 -11810 4951 -11620
rect 1751 -12200 2571 -11810
rect 3801 -12200 4621 -11810
rect 5211 -11811 7291 -11621
rect 5841 -12201 6661 -11811
<< pwell >>
rect 994 1205 3326 1797
rect 1294 765 3026 1205
rect 3614 765 5346 1797
rect 5634 765 7366 1797
rect 994 -2055 3326 -1023
rect 3634 -2055 5066 -1023
rect 5364 -2055 7096 -1023
rect 1145 -4283 3177 -3843
rect 3495 -4283 4927 -3843
rect 5235 -4283 7267 -3844
rect 1014 -4383 3386 -4283
rect 3495 -4383 5127 -4283
rect 5235 -4284 7496 -4283
rect 5225 -4383 7496 -4284
rect 1014 -4415 7496 -4383
rect 1014 -4515 3386 -4415
rect 3495 -4416 7496 -4415
rect 1034 -4955 3366 -4515
rect 3495 -4516 5127 -4416
rect 5225 -4516 7496 -4416
rect 3695 -4956 5127 -4516
rect 5454 -4956 7486 -4516
rect 1034 -7776 3366 -6744
rect 3694 -7776 5126 -6744
rect 5423 -7776 7155 -6744
rect 994 -10596 3326 -9564
rect 3634 -10596 5066 -9564
rect 5364 -10596 7096 -9564
rect 1145 -12824 3177 -12384
rect 1135 -12976 3187 -12824
rect 3495 -12976 4927 -12384
rect 5235 -12825 7267 -12385
rect 5225 -12977 7277 -12825
<< nmos >>
rect 1140 1471 1170 1771
rect 1290 1471 1320 1771
rect 1440 1471 1470 1771
rect 1590 1471 1620 1771
rect 1920 1471 1950 1771
rect 2070 1471 2100 1771
rect 2220 1471 2250 1771
rect 2370 1471 2400 1771
rect 2700 1471 2730 1771
rect 2850 1471 2880 1771
rect 3000 1471 3030 1771
rect 3150 1471 3180 1771
rect 3760 1471 3790 1771
rect 3910 1471 3940 1771
rect 4240 1471 4270 1771
rect 4390 1471 4420 1771
rect 4540 1471 4570 1771
rect 4690 1471 4720 1771
rect 5020 1471 5050 1771
rect 5170 1471 5200 1771
rect 5780 1471 5810 1771
rect 5930 1471 5960 1771
rect 6260 1471 6290 1771
rect 6410 1471 6440 1771
rect 6560 1471 6590 1771
rect 6710 1471 6740 1771
rect 7040 1471 7070 1771
rect 7190 1471 7220 1771
rect 1440 791 1470 1091
rect 1590 791 1620 1091
rect 1920 791 1950 1091
rect 2070 791 2100 1091
rect 2220 791 2250 1091
rect 2370 791 2400 1091
rect 2700 791 2730 1091
rect 2850 791 2880 1091
rect 3760 791 3790 1091
rect 3910 791 3940 1091
rect 4240 791 4270 1091
rect 4390 791 4420 1091
rect 4540 791 4570 1091
rect 4690 791 4720 1091
rect 5020 791 5050 1091
rect 5170 791 5200 1091
rect 5780 791 5810 1091
rect 5930 791 5960 1091
rect 6260 791 6290 1091
rect 6410 791 6440 1091
rect 6560 791 6590 1091
rect 6710 791 6740 1091
rect 7040 791 7070 1091
rect 7190 791 7220 1091
rect 1140 -1349 1170 -1049
rect 1290 -1349 1320 -1049
rect 1440 -1349 1470 -1049
rect 1590 -1349 1620 -1049
rect 1920 -1349 1950 -1049
rect 2070 -1349 2100 -1049
rect 2220 -1349 2250 -1049
rect 2370 -1349 2400 -1049
rect 2700 -1349 2730 -1049
rect 2850 -1349 2880 -1049
rect 3000 -1349 3030 -1049
rect 3150 -1349 3180 -1049
rect 3780 -1349 3810 -1049
rect 4110 -1349 4140 -1049
rect 4260 -1349 4290 -1049
rect 4410 -1349 4440 -1049
rect 4560 -1349 4590 -1049
rect 4890 -1349 4920 -1049
rect 5510 -1349 5540 -1049
rect 5660 -1349 5690 -1049
rect 5990 -1349 6020 -1049
rect 6140 -1349 6170 -1049
rect 6290 -1349 6320 -1049
rect 6440 -1349 6470 -1049
rect 6770 -1349 6800 -1049
rect 6920 -1349 6950 -1049
rect 1140 -2029 1170 -1729
rect 1290 -2029 1320 -1729
rect 1440 -2029 1470 -1729
rect 1590 -2029 1620 -1729
rect 1920 -2029 1950 -1729
rect 2070 -2029 2100 -1729
rect 2220 -2029 2250 -1729
rect 2370 -2029 2400 -1729
rect 2700 -2029 2730 -1729
rect 2850 -2029 2880 -1729
rect 3000 -2029 3030 -1729
rect 3150 -2029 3180 -1729
rect 3780 -2029 3810 -1729
rect 4110 -2029 4140 -1729
rect 4260 -2029 4290 -1729
rect 4410 -2029 4440 -1729
rect 4560 -2029 4590 -1729
rect 4890 -2029 4920 -1729
rect 5510 -2029 5540 -1729
rect 5660 -2029 5690 -1729
rect 5990 -2029 6020 -1729
rect 6140 -2029 6170 -1729
rect 6290 -2029 6320 -1729
rect 6440 -2029 6470 -1729
rect 6770 -2029 6800 -1729
rect 6920 -2029 6950 -1729
rect 1291 -4169 1321 -3869
rect 1441 -4169 1471 -3869
rect 1591 -4169 1621 -3869
rect 1921 -4169 1951 -3869
rect 2071 -4169 2101 -3869
rect 2221 -4169 2251 -3869
rect 2371 -4169 2401 -3869
rect 2701 -4169 2731 -3869
rect 2851 -4169 2881 -3869
rect 3001 -4169 3031 -3869
rect 3641 -4169 3671 -3869
rect 3971 -4169 4001 -3869
rect 4121 -4169 4151 -3869
rect 4271 -4169 4301 -3869
rect 4421 -4169 4451 -3869
rect 4751 -4169 4781 -3869
rect 5381 -4170 5411 -3870
rect 5531 -4170 5561 -3870
rect 5681 -4170 5711 -3870
rect 6011 -4170 6041 -3870
rect 6161 -4170 6191 -3870
rect 6311 -4170 6341 -3870
rect 6461 -4170 6491 -3870
rect 6791 -4170 6821 -3870
rect 6941 -4170 6971 -3870
rect 7091 -4170 7121 -3870
rect 1180 -4929 1210 -4629
rect 1330 -4929 1360 -4629
rect 1480 -4929 1510 -4629
rect 1630 -4929 1660 -4629
rect 1960 -4929 1990 -4629
rect 2110 -4929 2140 -4629
rect 2260 -4929 2290 -4629
rect 2410 -4929 2440 -4629
rect 2740 -4929 2770 -4629
rect 2890 -4929 2920 -4629
rect 3040 -4929 3070 -4629
rect 3190 -4929 3220 -4629
rect 3841 -4930 3871 -4630
rect 4171 -4930 4201 -4630
rect 4321 -4930 4351 -4630
rect 4471 -4930 4501 -4630
rect 4621 -4930 4651 -4630
rect 4951 -4930 4981 -4630
rect 5600 -4930 5630 -4630
rect 5750 -4930 5780 -4630
rect 5900 -4930 5930 -4630
rect 6230 -4930 6260 -4630
rect 6380 -4930 6410 -4630
rect 6530 -4930 6560 -4630
rect 6680 -4930 6710 -4630
rect 7010 -4930 7040 -4630
rect 7160 -4930 7190 -4630
rect 7310 -4930 7340 -4630
rect 1180 -7070 1210 -6770
rect 1330 -7070 1360 -6770
rect 1480 -7070 1510 -6770
rect 1630 -7070 1660 -6770
rect 1960 -7070 1990 -6770
rect 2110 -7070 2140 -6770
rect 2260 -7070 2290 -6770
rect 2410 -7070 2440 -6770
rect 2740 -7070 2770 -6770
rect 2890 -7070 2920 -6770
rect 3040 -7070 3070 -6770
rect 3190 -7070 3220 -6770
rect 3840 -7070 3870 -6770
rect 4170 -7070 4200 -6770
rect 4320 -7070 4350 -6770
rect 4470 -7070 4500 -6770
rect 4620 -7070 4650 -6770
rect 4950 -7070 4980 -6770
rect 5569 -7070 5599 -6770
rect 5719 -7070 5749 -6770
rect 6049 -7070 6079 -6770
rect 6199 -7070 6229 -6770
rect 6349 -7070 6379 -6770
rect 6499 -7070 6529 -6770
rect 6829 -7070 6859 -6770
rect 6979 -7070 7009 -6770
rect 1180 -7750 1210 -7450
rect 1330 -7750 1360 -7450
rect 1480 -7750 1510 -7450
rect 1630 -7750 1660 -7450
rect 1960 -7750 1990 -7450
rect 2110 -7750 2140 -7450
rect 2260 -7750 2290 -7450
rect 2410 -7750 2440 -7450
rect 2740 -7750 2770 -7450
rect 2890 -7750 2920 -7450
rect 3040 -7750 3070 -7450
rect 3190 -7750 3220 -7450
rect 3840 -7750 3870 -7450
rect 4170 -7750 4200 -7450
rect 4320 -7750 4350 -7450
rect 4470 -7750 4500 -7450
rect 4620 -7750 4650 -7450
rect 4950 -7750 4980 -7450
rect 5569 -7750 5599 -7450
rect 5719 -7750 5749 -7450
rect 6049 -7750 6079 -7450
rect 6199 -7750 6229 -7450
rect 6349 -7750 6379 -7450
rect 6499 -7750 6529 -7450
rect 6829 -7750 6859 -7450
rect 6979 -7750 7009 -7450
rect 1140 -9890 1170 -9590
rect 1290 -9890 1320 -9590
rect 1440 -9890 1470 -9590
rect 1590 -9890 1620 -9590
rect 1920 -9890 1950 -9590
rect 2070 -9890 2100 -9590
rect 2220 -9890 2250 -9590
rect 2370 -9890 2400 -9590
rect 2700 -9890 2730 -9590
rect 2850 -9890 2880 -9590
rect 3000 -9890 3030 -9590
rect 3150 -9890 3180 -9590
rect 3780 -9890 3810 -9590
rect 4110 -9890 4140 -9590
rect 4260 -9890 4290 -9590
rect 4410 -9890 4440 -9590
rect 4560 -9890 4590 -9590
rect 4890 -9890 4920 -9590
rect 5510 -9890 5540 -9590
rect 5660 -9890 5690 -9590
rect 5990 -9890 6020 -9590
rect 6140 -9890 6170 -9590
rect 6290 -9890 6320 -9590
rect 6440 -9890 6470 -9590
rect 6770 -9890 6800 -9590
rect 6920 -9890 6950 -9590
rect 1140 -10570 1170 -10270
rect 1290 -10570 1320 -10270
rect 1440 -10570 1470 -10270
rect 1590 -10570 1620 -10270
rect 1920 -10570 1950 -10270
rect 2070 -10570 2100 -10270
rect 2220 -10570 2250 -10270
rect 2370 -10570 2400 -10270
rect 2700 -10570 2730 -10270
rect 2850 -10570 2880 -10270
rect 3000 -10570 3030 -10270
rect 3150 -10570 3180 -10270
rect 3780 -10570 3810 -10270
rect 4110 -10570 4140 -10270
rect 4260 -10570 4290 -10270
rect 4410 -10570 4440 -10270
rect 4560 -10570 4590 -10270
rect 4890 -10570 4920 -10270
rect 5510 -10570 5540 -10270
rect 5660 -10570 5690 -10270
rect 5990 -10570 6020 -10270
rect 6140 -10570 6170 -10270
rect 6290 -10570 6320 -10270
rect 6440 -10570 6470 -10270
rect 6770 -10570 6800 -10270
rect 6920 -10570 6950 -10270
rect 1291 -12710 1321 -12410
rect 1441 -12710 1471 -12410
rect 1591 -12710 1621 -12410
rect 1921 -12710 1951 -12410
rect 2071 -12710 2101 -12410
rect 2221 -12710 2251 -12410
rect 2371 -12710 2401 -12410
rect 2701 -12710 2731 -12410
rect 2851 -12710 2881 -12410
rect 3001 -12710 3031 -12410
rect 3641 -12710 3671 -12410
rect 3971 -12710 4001 -12410
rect 4121 -12710 4151 -12410
rect 4271 -12710 4301 -12410
rect 4421 -12710 4451 -12410
rect 4751 -12710 4781 -12410
rect 5381 -12711 5411 -12411
rect 5531 -12711 5561 -12411
rect 5681 -12711 5711 -12411
rect 6011 -12711 6041 -12411
rect 6161 -12711 6191 -12411
rect 6311 -12711 6341 -12411
rect 6461 -12711 6491 -12411
rect 6791 -12711 6821 -12411
rect 6941 -12711 6971 -12411
rect 7091 -12711 7121 -12411
<< pmos >>
rect 1920 2031 1950 2331
rect 2070 2031 2100 2331
rect 2220 2031 2250 2331
rect 2370 2031 2400 2331
rect 4240 2031 4270 2331
rect 4390 2031 4420 2331
rect 4540 2031 4570 2331
rect 4690 2031 4720 2331
rect 6260 2031 6290 2331
rect 6410 2031 6440 2331
rect 6560 2031 6590 2331
rect 6710 2031 6740 2331
rect 1920 231 1950 531
rect 2070 231 2100 531
rect 2220 231 2250 531
rect 2370 231 2400 531
rect 4240 231 4270 531
rect 4390 231 4420 531
rect 4540 231 4570 531
rect 4690 231 4720 531
rect 6260 231 6290 531
rect 6410 231 6440 531
rect 6560 231 6590 531
rect 6710 231 6740 531
rect 1920 -789 1950 -489
rect 2070 -789 2100 -489
rect 2220 -789 2250 -489
rect 2370 -789 2400 -489
rect 4110 -789 4140 -489
rect 4260 -789 4290 -489
rect 4410 -789 4440 -489
rect 4560 -789 4590 -489
rect 5990 -789 6020 -489
rect 6140 -789 6170 -489
rect 6290 -789 6320 -489
rect 6440 -789 6470 -489
rect 1920 -2589 1950 -2289
rect 2070 -2589 2100 -2289
rect 2220 -2589 2250 -2289
rect 2370 -2589 2400 -2289
rect 4110 -2589 4140 -2289
rect 4260 -2589 4290 -2289
rect 4410 -2589 4440 -2289
rect 4560 -2589 4590 -2289
rect 5990 -2589 6020 -2289
rect 6140 -2589 6170 -2289
rect 6290 -2589 6320 -2289
rect 6440 -2589 6470 -2289
rect 1921 -3609 1951 -3309
rect 2071 -3609 2101 -3309
rect 2221 -3609 2251 -3309
rect 2371 -3609 2401 -3309
rect 3971 -3609 4001 -3309
rect 4121 -3609 4151 -3309
rect 4271 -3609 4301 -3309
rect 4421 -3609 4451 -3309
rect 6011 -3610 6041 -3310
rect 6161 -3610 6191 -3310
rect 6311 -3610 6341 -3310
rect 6461 -3610 6491 -3310
rect 4171 -5490 4201 -5190
rect 4321 -5490 4351 -5190
rect 4471 -5490 4501 -5190
rect 4621 -5490 4651 -5190
rect 1960 -5809 1990 -5509
rect 2110 -5809 2140 -5509
rect 2260 -5809 2290 -5509
rect 2410 -5809 2440 -5509
rect 6230 -5490 6260 -5190
rect 6380 -5490 6410 -5190
rect 6530 -5490 6560 -5190
rect 6680 -5490 6710 -5190
rect 1960 -6510 1990 -6210
rect 2110 -6510 2140 -6210
rect 2260 -6510 2290 -6210
rect 2410 -6510 2440 -6210
rect 4170 -6510 4200 -6210
rect 4320 -6510 4350 -6210
rect 4470 -6510 4500 -6210
rect 4620 -6510 4650 -6210
rect 6049 -6510 6079 -6210
rect 6199 -6510 6229 -6210
rect 6349 -6510 6379 -6210
rect 6499 -6510 6529 -6210
rect 1960 -8310 1990 -8010
rect 2110 -8310 2140 -8010
rect 2260 -8310 2290 -8010
rect 2410 -8310 2440 -8010
rect 4170 -8310 4200 -8010
rect 4320 -8310 4350 -8010
rect 4470 -8310 4500 -8010
rect 4620 -8310 4650 -8010
rect 6049 -8310 6079 -8010
rect 6199 -8310 6229 -8010
rect 6349 -8310 6379 -8010
rect 6499 -8310 6529 -8010
rect 1920 -9330 1950 -9030
rect 2070 -9330 2100 -9030
rect 2220 -9330 2250 -9030
rect 2370 -9330 2400 -9030
rect 4110 -9330 4140 -9030
rect 4260 -9330 4290 -9030
rect 4410 -9330 4440 -9030
rect 4560 -9330 4590 -9030
rect 5990 -9330 6020 -9030
rect 6140 -9330 6170 -9030
rect 6290 -9330 6320 -9030
rect 6440 -9330 6470 -9030
rect 1920 -11130 1950 -10830
rect 2070 -11130 2100 -10830
rect 2220 -11130 2250 -10830
rect 2370 -11130 2400 -10830
rect 4110 -11130 4140 -10830
rect 4260 -11130 4290 -10830
rect 4410 -11130 4440 -10830
rect 4560 -11130 4590 -10830
rect 5990 -11130 6020 -10830
rect 6140 -11130 6170 -10830
rect 6290 -11130 6320 -10830
rect 6440 -11130 6470 -10830
rect 1921 -12150 1951 -11850
rect 2071 -12150 2101 -11850
rect 2221 -12150 2251 -11850
rect 2371 -12150 2401 -11850
rect 3971 -12150 4001 -11850
rect 4121 -12150 4151 -11850
rect 4271 -12150 4301 -11850
rect 4421 -12150 4451 -11850
rect 6011 -12151 6041 -11851
rect 6161 -12151 6191 -11851
rect 6311 -12151 6341 -11851
rect 6461 -12151 6491 -11851
<< ndiff >>
rect 1020 1698 1140 1771
rect 1020 1664 1063 1698
rect 1097 1664 1140 1698
rect 1020 1618 1140 1664
rect 1020 1584 1063 1618
rect 1097 1584 1140 1618
rect 1020 1538 1140 1584
rect 1020 1504 1063 1538
rect 1097 1504 1140 1538
rect 1020 1471 1140 1504
rect 1170 1471 1290 1771
rect 1320 1698 1440 1771
rect 1320 1664 1363 1698
rect 1397 1664 1440 1698
rect 1320 1618 1440 1664
rect 1320 1584 1363 1618
rect 1397 1584 1440 1618
rect 1320 1538 1440 1584
rect 1320 1504 1363 1538
rect 1397 1504 1440 1538
rect 1320 1471 1440 1504
rect 1470 1471 1590 1771
rect 1620 1698 1740 1771
rect 1620 1664 1663 1698
rect 1697 1664 1740 1698
rect 1620 1618 1740 1664
rect 1620 1584 1663 1618
rect 1697 1584 1740 1618
rect 1620 1538 1740 1584
rect 1620 1504 1663 1538
rect 1697 1504 1740 1538
rect 1620 1471 1740 1504
rect 1800 1698 1920 1771
rect 1800 1664 1843 1698
rect 1877 1664 1920 1698
rect 1800 1618 1920 1664
rect 1800 1584 1843 1618
rect 1877 1584 1920 1618
rect 1800 1538 1920 1584
rect 1800 1504 1843 1538
rect 1877 1504 1920 1538
rect 1800 1471 1920 1504
rect 1950 1698 2070 1771
rect 1950 1664 1993 1698
rect 2027 1664 2070 1698
rect 1950 1618 2070 1664
rect 1950 1584 1993 1618
rect 2027 1584 2070 1618
rect 1950 1538 2070 1584
rect 1950 1504 1993 1538
rect 2027 1504 2070 1538
rect 1950 1471 2070 1504
rect 2100 1698 2220 1771
rect 2100 1664 2143 1698
rect 2177 1664 2220 1698
rect 2100 1618 2220 1664
rect 2100 1584 2143 1618
rect 2177 1584 2220 1618
rect 2100 1538 2220 1584
rect 2100 1504 2143 1538
rect 2177 1504 2220 1538
rect 2100 1471 2220 1504
rect 2250 1698 2370 1771
rect 2250 1664 2293 1698
rect 2327 1664 2370 1698
rect 2250 1618 2370 1664
rect 2250 1584 2293 1618
rect 2327 1584 2370 1618
rect 2250 1538 2370 1584
rect 2250 1504 2293 1538
rect 2327 1504 2370 1538
rect 2250 1471 2370 1504
rect 2400 1698 2520 1771
rect 2400 1664 2443 1698
rect 2477 1664 2520 1698
rect 2400 1618 2520 1664
rect 2400 1584 2443 1618
rect 2477 1584 2520 1618
rect 2400 1538 2520 1584
rect 2400 1504 2443 1538
rect 2477 1504 2520 1538
rect 2400 1471 2520 1504
rect 2580 1698 2700 1771
rect 2580 1664 2623 1698
rect 2657 1664 2700 1698
rect 2580 1618 2700 1664
rect 2580 1584 2623 1618
rect 2657 1584 2700 1618
rect 2580 1538 2700 1584
rect 2580 1504 2623 1538
rect 2657 1504 2700 1538
rect 2580 1471 2700 1504
rect 2730 1471 2850 1771
rect 2880 1698 3000 1771
rect 2880 1664 2923 1698
rect 2957 1664 3000 1698
rect 2880 1618 3000 1664
rect 2880 1584 2923 1618
rect 2957 1584 3000 1618
rect 2880 1538 3000 1584
rect 2880 1504 2923 1538
rect 2957 1504 3000 1538
rect 2880 1471 3000 1504
rect 3030 1471 3150 1771
rect 3180 1698 3300 1771
rect 3180 1664 3223 1698
rect 3257 1664 3300 1698
rect 3180 1618 3300 1664
rect 3180 1584 3223 1618
rect 3257 1584 3300 1618
rect 3180 1538 3300 1584
rect 3180 1504 3223 1538
rect 3257 1504 3300 1538
rect 3180 1471 3300 1504
rect 3640 1698 3760 1771
rect 3640 1664 3683 1698
rect 3717 1664 3760 1698
rect 3640 1618 3760 1664
rect 3640 1584 3683 1618
rect 3717 1584 3760 1618
rect 3640 1538 3760 1584
rect 3640 1504 3683 1538
rect 3717 1504 3760 1538
rect 3640 1471 3760 1504
rect 3790 1471 3910 1771
rect 3940 1698 4060 1771
rect 3940 1664 3983 1698
rect 4017 1664 4060 1698
rect 3940 1618 4060 1664
rect 3940 1584 3983 1618
rect 4017 1584 4060 1618
rect 3940 1538 4060 1584
rect 3940 1504 3983 1538
rect 4017 1504 4060 1538
rect 3940 1471 4060 1504
rect 4120 1698 4240 1771
rect 4120 1664 4163 1698
rect 4197 1664 4240 1698
rect 4120 1618 4240 1664
rect 4120 1584 4163 1618
rect 4197 1584 4240 1618
rect 4120 1538 4240 1584
rect 4120 1504 4163 1538
rect 4197 1504 4240 1538
rect 4120 1471 4240 1504
rect 4270 1698 4390 1771
rect 4270 1664 4313 1698
rect 4347 1664 4390 1698
rect 4270 1618 4390 1664
rect 4270 1584 4313 1618
rect 4347 1584 4390 1618
rect 4270 1538 4390 1584
rect 4270 1504 4313 1538
rect 4347 1504 4390 1538
rect 4270 1471 4390 1504
rect 4420 1698 4540 1771
rect 4420 1664 4463 1698
rect 4497 1664 4540 1698
rect 4420 1618 4540 1664
rect 4420 1584 4463 1618
rect 4497 1584 4540 1618
rect 4420 1538 4540 1584
rect 4420 1504 4463 1538
rect 4497 1504 4540 1538
rect 4420 1471 4540 1504
rect 4570 1698 4690 1771
rect 4570 1664 4613 1698
rect 4647 1664 4690 1698
rect 4570 1618 4690 1664
rect 4570 1584 4613 1618
rect 4647 1584 4690 1618
rect 4570 1538 4690 1584
rect 4570 1504 4613 1538
rect 4647 1504 4690 1538
rect 4570 1471 4690 1504
rect 4720 1698 4840 1771
rect 4720 1664 4763 1698
rect 4797 1664 4840 1698
rect 4720 1618 4840 1664
rect 4720 1584 4763 1618
rect 4797 1584 4840 1618
rect 4720 1538 4840 1584
rect 4720 1504 4763 1538
rect 4797 1504 4840 1538
rect 4720 1471 4840 1504
rect 4900 1698 5020 1771
rect 4900 1664 4943 1698
rect 4977 1664 5020 1698
rect 4900 1618 5020 1664
rect 4900 1584 4943 1618
rect 4977 1584 5020 1618
rect 4900 1538 5020 1584
rect 4900 1504 4943 1538
rect 4977 1504 5020 1538
rect 4900 1471 5020 1504
rect 5050 1698 5170 1771
rect 5050 1664 5093 1698
rect 5127 1664 5170 1698
rect 5050 1618 5170 1664
rect 5050 1584 5093 1618
rect 5127 1584 5170 1618
rect 5050 1538 5170 1584
rect 5050 1504 5093 1538
rect 5127 1504 5170 1538
rect 5050 1471 5170 1504
rect 5200 1698 5320 1771
rect 5200 1664 5243 1698
rect 5277 1664 5320 1698
rect 5200 1618 5320 1664
rect 5200 1584 5243 1618
rect 5277 1584 5320 1618
rect 5200 1538 5320 1584
rect 5200 1504 5243 1538
rect 5277 1504 5320 1538
rect 5200 1471 5320 1504
rect 5660 1698 5780 1771
rect 5660 1664 5703 1698
rect 5737 1664 5780 1698
rect 5660 1618 5780 1664
rect 5660 1584 5703 1618
rect 5737 1584 5780 1618
rect 5660 1538 5780 1584
rect 5660 1504 5703 1538
rect 5737 1504 5780 1538
rect 5660 1471 5780 1504
rect 5810 1698 5930 1771
rect 5810 1664 5853 1698
rect 5887 1664 5930 1698
rect 5810 1618 5930 1664
rect 5810 1584 5853 1618
rect 5887 1584 5930 1618
rect 5810 1538 5930 1584
rect 5810 1504 5853 1538
rect 5887 1504 5930 1538
rect 5810 1471 5930 1504
rect 5960 1698 6080 1771
rect 5960 1664 6003 1698
rect 6037 1664 6080 1698
rect 5960 1618 6080 1664
rect 5960 1584 6003 1618
rect 6037 1584 6080 1618
rect 5960 1538 6080 1584
rect 5960 1504 6003 1538
rect 6037 1504 6080 1538
rect 5960 1471 6080 1504
rect 6140 1698 6260 1771
rect 6140 1664 6183 1698
rect 6217 1664 6260 1698
rect 6140 1618 6260 1664
rect 6140 1584 6183 1618
rect 6217 1584 6260 1618
rect 6140 1538 6260 1584
rect 6140 1504 6183 1538
rect 6217 1504 6260 1538
rect 6140 1471 6260 1504
rect 6290 1698 6410 1771
rect 6290 1664 6333 1698
rect 6367 1664 6410 1698
rect 6290 1618 6410 1664
rect 6290 1584 6333 1618
rect 6367 1584 6410 1618
rect 6290 1538 6410 1584
rect 6290 1504 6333 1538
rect 6367 1504 6410 1538
rect 6290 1471 6410 1504
rect 6440 1698 6560 1771
rect 6440 1664 6483 1698
rect 6517 1664 6560 1698
rect 6440 1618 6560 1664
rect 6440 1584 6483 1618
rect 6517 1584 6560 1618
rect 6440 1538 6560 1584
rect 6440 1504 6483 1538
rect 6517 1504 6560 1538
rect 6440 1471 6560 1504
rect 6590 1698 6710 1771
rect 6590 1664 6633 1698
rect 6667 1664 6710 1698
rect 6590 1618 6710 1664
rect 6590 1584 6633 1618
rect 6667 1584 6710 1618
rect 6590 1538 6710 1584
rect 6590 1504 6633 1538
rect 6667 1504 6710 1538
rect 6590 1471 6710 1504
rect 6740 1698 6860 1771
rect 6740 1664 6783 1698
rect 6817 1664 6860 1698
rect 6740 1618 6860 1664
rect 6740 1584 6783 1618
rect 6817 1584 6860 1618
rect 6740 1538 6860 1584
rect 6740 1504 6783 1538
rect 6817 1504 6860 1538
rect 6740 1471 6860 1504
rect 6920 1698 7040 1771
rect 6920 1664 6963 1698
rect 6997 1664 7040 1698
rect 6920 1618 7040 1664
rect 6920 1584 6963 1618
rect 6997 1584 7040 1618
rect 6920 1538 7040 1584
rect 6920 1504 6963 1538
rect 6997 1504 7040 1538
rect 6920 1471 7040 1504
rect 7070 1471 7190 1771
rect 7220 1698 7340 1771
rect 7220 1664 7263 1698
rect 7297 1664 7340 1698
rect 7220 1618 7340 1664
rect 7220 1584 7263 1618
rect 7297 1584 7340 1618
rect 7220 1538 7340 1584
rect 7220 1504 7263 1538
rect 7297 1504 7340 1538
rect 7220 1471 7340 1504
rect 1320 1058 1440 1091
rect 1320 1024 1363 1058
rect 1397 1024 1440 1058
rect 1320 978 1440 1024
rect 1320 944 1363 978
rect 1397 944 1440 978
rect 1320 898 1440 944
rect 1320 864 1363 898
rect 1397 864 1440 898
rect 1320 791 1440 864
rect 1470 1058 1590 1091
rect 1470 1024 1513 1058
rect 1547 1024 1590 1058
rect 1470 978 1590 1024
rect 1470 944 1513 978
rect 1547 944 1590 978
rect 1470 898 1590 944
rect 1470 864 1513 898
rect 1547 864 1590 898
rect 1470 791 1590 864
rect 1620 1058 1740 1091
rect 1620 1024 1663 1058
rect 1697 1024 1740 1058
rect 1620 978 1740 1024
rect 1620 944 1663 978
rect 1697 944 1740 978
rect 1620 898 1740 944
rect 1620 864 1663 898
rect 1697 864 1740 898
rect 1620 791 1740 864
rect 1800 1058 1920 1091
rect 1800 1024 1843 1058
rect 1877 1024 1920 1058
rect 1800 978 1920 1024
rect 1800 944 1843 978
rect 1877 944 1920 978
rect 1800 898 1920 944
rect 1800 864 1843 898
rect 1877 864 1920 898
rect 1800 791 1920 864
rect 1950 1058 2070 1091
rect 1950 1024 1993 1058
rect 2027 1024 2070 1058
rect 1950 978 2070 1024
rect 1950 944 1993 978
rect 2027 944 2070 978
rect 1950 898 2070 944
rect 1950 864 1993 898
rect 2027 864 2070 898
rect 1950 791 2070 864
rect 2100 1058 2220 1091
rect 2100 1024 2143 1058
rect 2177 1024 2220 1058
rect 2100 978 2220 1024
rect 2100 944 2143 978
rect 2177 944 2220 978
rect 2100 898 2220 944
rect 2100 864 2143 898
rect 2177 864 2220 898
rect 2100 791 2220 864
rect 2250 1058 2370 1091
rect 2250 1024 2293 1058
rect 2327 1024 2370 1058
rect 2250 978 2370 1024
rect 2250 944 2293 978
rect 2327 944 2370 978
rect 2250 898 2370 944
rect 2250 864 2293 898
rect 2327 864 2370 898
rect 2250 791 2370 864
rect 2400 1058 2520 1091
rect 2400 1024 2443 1058
rect 2477 1024 2520 1058
rect 2400 978 2520 1024
rect 2400 944 2443 978
rect 2477 944 2520 978
rect 2400 898 2520 944
rect 2400 864 2443 898
rect 2477 864 2520 898
rect 2400 791 2520 864
rect 2580 1058 2700 1091
rect 2580 1024 2623 1058
rect 2657 1024 2700 1058
rect 2580 978 2700 1024
rect 2580 944 2623 978
rect 2657 944 2700 978
rect 2580 898 2700 944
rect 2580 864 2623 898
rect 2657 864 2700 898
rect 2580 791 2700 864
rect 2730 791 2850 1091
rect 2880 1058 3000 1091
rect 2880 1024 2923 1058
rect 2957 1024 3000 1058
rect 2880 978 3000 1024
rect 2880 944 2923 978
rect 2957 944 3000 978
rect 2880 898 3000 944
rect 2880 864 2923 898
rect 2957 864 3000 898
rect 2880 791 3000 864
rect 3640 1058 3760 1091
rect 3640 1024 3683 1058
rect 3717 1024 3760 1058
rect 3640 978 3760 1024
rect 3640 944 3683 978
rect 3717 944 3760 978
rect 3640 898 3760 944
rect 3640 864 3683 898
rect 3717 864 3760 898
rect 3640 791 3760 864
rect 3790 1058 3910 1091
rect 3790 1024 3833 1058
rect 3867 1024 3910 1058
rect 3790 978 3910 1024
rect 3790 944 3833 978
rect 3867 944 3910 978
rect 3790 898 3910 944
rect 3790 864 3833 898
rect 3867 864 3910 898
rect 3790 791 3910 864
rect 3940 1058 4060 1091
rect 3940 1024 3983 1058
rect 4017 1024 4060 1058
rect 3940 978 4060 1024
rect 3940 944 3983 978
rect 4017 944 4060 978
rect 3940 898 4060 944
rect 3940 864 3983 898
rect 4017 864 4060 898
rect 3940 791 4060 864
rect 4120 1058 4240 1091
rect 4120 1024 4163 1058
rect 4197 1024 4240 1058
rect 4120 978 4240 1024
rect 4120 944 4163 978
rect 4197 944 4240 978
rect 4120 898 4240 944
rect 4120 864 4163 898
rect 4197 864 4240 898
rect 4120 791 4240 864
rect 4270 1058 4390 1091
rect 4270 1024 4313 1058
rect 4347 1024 4390 1058
rect 4270 978 4390 1024
rect 4270 944 4313 978
rect 4347 944 4390 978
rect 4270 898 4390 944
rect 4270 864 4313 898
rect 4347 864 4390 898
rect 4270 791 4390 864
rect 4420 1058 4540 1091
rect 4420 1024 4463 1058
rect 4497 1024 4540 1058
rect 4420 978 4540 1024
rect 4420 944 4463 978
rect 4497 944 4540 978
rect 4420 898 4540 944
rect 4420 864 4463 898
rect 4497 864 4540 898
rect 4420 791 4540 864
rect 4570 1058 4690 1091
rect 4570 1024 4613 1058
rect 4647 1024 4690 1058
rect 4570 978 4690 1024
rect 4570 944 4613 978
rect 4647 944 4690 978
rect 4570 898 4690 944
rect 4570 864 4613 898
rect 4647 864 4690 898
rect 4570 791 4690 864
rect 4720 1058 4840 1091
rect 4720 1024 4763 1058
rect 4797 1024 4840 1058
rect 4720 978 4840 1024
rect 4720 944 4763 978
rect 4797 944 4840 978
rect 4720 898 4840 944
rect 4720 864 4763 898
rect 4797 864 4840 898
rect 4720 791 4840 864
rect 4900 1058 5020 1091
rect 4900 1024 4943 1058
rect 4977 1024 5020 1058
rect 4900 978 5020 1024
rect 4900 944 4943 978
rect 4977 944 5020 978
rect 4900 898 5020 944
rect 4900 864 4943 898
rect 4977 864 5020 898
rect 4900 791 5020 864
rect 5050 791 5170 1091
rect 5200 1058 5320 1091
rect 5200 1024 5243 1058
rect 5277 1024 5320 1058
rect 5200 978 5320 1024
rect 5200 944 5243 978
rect 5277 944 5320 978
rect 5200 898 5320 944
rect 5200 864 5243 898
rect 5277 864 5320 898
rect 5200 791 5320 864
rect 5660 1058 5780 1091
rect 5660 1024 5703 1058
rect 5737 1024 5780 1058
rect 5660 978 5780 1024
rect 5660 944 5703 978
rect 5737 944 5780 978
rect 5660 898 5780 944
rect 5660 864 5703 898
rect 5737 864 5780 898
rect 5660 791 5780 864
rect 5810 1058 5930 1091
rect 5810 1024 5853 1058
rect 5887 1024 5930 1058
rect 5810 978 5930 1024
rect 5810 944 5853 978
rect 5887 944 5930 978
rect 5810 898 5930 944
rect 5810 864 5853 898
rect 5887 864 5930 898
rect 5810 791 5930 864
rect 5960 1058 6080 1091
rect 5960 1024 6003 1058
rect 6037 1024 6080 1058
rect 5960 978 6080 1024
rect 5960 944 6003 978
rect 6037 944 6080 978
rect 5960 898 6080 944
rect 5960 864 6003 898
rect 6037 864 6080 898
rect 5960 791 6080 864
rect 6140 1058 6260 1091
rect 6140 1024 6183 1058
rect 6217 1024 6260 1058
rect 6140 978 6260 1024
rect 6140 944 6183 978
rect 6217 944 6260 978
rect 6140 898 6260 944
rect 6140 864 6183 898
rect 6217 864 6260 898
rect 6140 791 6260 864
rect 6290 1058 6410 1091
rect 6290 1024 6333 1058
rect 6367 1024 6410 1058
rect 6290 978 6410 1024
rect 6290 944 6333 978
rect 6367 944 6410 978
rect 6290 898 6410 944
rect 6290 864 6333 898
rect 6367 864 6410 898
rect 6290 791 6410 864
rect 6440 1058 6560 1091
rect 6440 1024 6483 1058
rect 6517 1024 6560 1058
rect 6440 978 6560 1024
rect 6440 944 6483 978
rect 6517 944 6560 978
rect 6440 898 6560 944
rect 6440 864 6483 898
rect 6517 864 6560 898
rect 6440 791 6560 864
rect 6590 1058 6710 1091
rect 6590 1024 6633 1058
rect 6667 1024 6710 1058
rect 6590 978 6710 1024
rect 6590 944 6633 978
rect 6667 944 6710 978
rect 6590 898 6710 944
rect 6590 864 6633 898
rect 6667 864 6710 898
rect 6590 791 6710 864
rect 6740 1058 6860 1091
rect 6740 1024 6783 1058
rect 6817 1024 6860 1058
rect 6740 978 6860 1024
rect 6740 944 6783 978
rect 6817 944 6860 978
rect 6740 898 6860 944
rect 6740 864 6783 898
rect 6817 864 6860 898
rect 6740 791 6860 864
rect 6920 1058 7040 1091
rect 6920 1024 6963 1058
rect 6997 1024 7040 1058
rect 6920 978 7040 1024
rect 6920 944 6963 978
rect 6997 944 7040 978
rect 6920 898 7040 944
rect 6920 864 6963 898
rect 6997 864 7040 898
rect 6920 791 7040 864
rect 7070 791 7190 1091
rect 7220 1058 7340 1091
rect 7220 1024 7263 1058
rect 7297 1024 7340 1058
rect 7220 978 7340 1024
rect 7220 944 7263 978
rect 7297 944 7340 978
rect 7220 898 7340 944
rect 7220 864 7263 898
rect 7297 864 7340 898
rect 7220 791 7340 864
rect 1020 -1122 1140 -1049
rect 1020 -1156 1063 -1122
rect 1097 -1156 1140 -1122
rect 1020 -1202 1140 -1156
rect 1020 -1236 1063 -1202
rect 1097 -1236 1140 -1202
rect 1020 -1282 1140 -1236
rect 1020 -1316 1063 -1282
rect 1097 -1316 1140 -1282
rect 1020 -1349 1140 -1316
rect 1170 -1349 1290 -1049
rect 1320 -1122 1440 -1049
rect 1320 -1156 1363 -1122
rect 1397 -1156 1440 -1122
rect 1320 -1202 1440 -1156
rect 1320 -1236 1363 -1202
rect 1397 -1236 1440 -1202
rect 1320 -1282 1440 -1236
rect 1320 -1316 1363 -1282
rect 1397 -1316 1440 -1282
rect 1320 -1349 1440 -1316
rect 1470 -1349 1590 -1049
rect 1620 -1122 1740 -1049
rect 1620 -1156 1663 -1122
rect 1697 -1156 1740 -1122
rect 1620 -1202 1740 -1156
rect 1620 -1236 1663 -1202
rect 1697 -1236 1740 -1202
rect 1620 -1282 1740 -1236
rect 1620 -1316 1663 -1282
rect 1697 -1316 1740 -1282
rect 1620 -1349 1740 -1316
rect 1800 -1122 1920 -1049
rect 1800 -1156 1843 -1122
rect 1877 -1156 1920 -1122
rect 1800 -1202 1920 -1156
rect 1800 -1236 1843 -1202
rect 1877 -1236 1920 -1202
rect 1800 -1282 1920 -1236
rect 1800 -1316 1843 -1282
rect 1877 -1316 1920 -1282
rect 1800 -1349 1920 -1316
rect 1950 -1122 2070 -1049
rect 1950 -1156 1993 -1122
rect 2027 -1156 2070 -1122
rect 1950 -1202 2070 -1156
rect 1950 -1236 1993 -1202
rect 2027 -1236 2070 -1202
rect 1950 -1282 2070 -1236
rect 1950 -1316 1993 -1282
rect 2027 -1316 2070 -1282
rect 1950 -1349 2070 -1316
rect 2100 -1122 2220 -1049
rect 2100 -1156 2143 -1122
rect 2177 -1156 2220 -1122
rect 2100 -1202 2220 -1156
rect 2100 -1236 2143 -1202
rect 2177 -1236 2220 -1202
rect 2100 -1282 2220 -1236
rect 2100 -1316 2143 -1282
rect 2177 -1316 2220 -1282
rect 2100 -1349 2220 -1316
rect 2250 -1122 2370 -1049
rect 2250 -1156 2293 -1122
rect 2327 -1156 2370 -1122
rect 2250 -1202 2370 -1156
rect 2250 -1236 2293 -1202
rect 2327 -1236 2370 -1202
rect 2250 -1282 2370 -1236
rect 2250 -1316 2293 -1282
rect 2327 -1316 2370 -1282
rect 2250 -1349 2370 -1316
rect 2400 -1122 2520 -1049
rect 2400 -1156 2443 -1122
rect 2477 -1156 2520 -1122
rect 2400 -1202 2520 -1156
rect 2400 -1236 2443 -1202
rect 2477 -1236 2520 -1202
rect 2400 -1282 2520 -1236
rect 2400 -1316 2443 -1282
rect 2477 -1316 2520 -1282
rect 2400 -1349 2520 -1316
rect 2580 -1122 2700 -1049
rect 2580 -1156 2623 -1122
rect 2657 -1156 2700 -1122
rect 2580 -1202 2700 -1156
rect 2580 -1236 2623 -1202
rect 2657 -1236 2700 -1202
rect 2580 -1282 2700 -1236
rect 2580 -1316 2623 -1282
rect 2657 -1316 2700 -1282
rect 2580 -1349 2700 -1316
rect 2730 -1349 2850 -1049
rect 2880 -1122 3000 -1049
rect 2880 -1156 2923 -1122
rect 2957 -1156 3000 -1122
rect 2880 -1202 3000 -1156
rect 2880 -1236 2923 -1202
rect 2957 -1236 3000 -1202
rect 2880 -1282 3000 -1236
rect 2880 -1316 2923 -1282
rect 2957 -1316 3000 -1282
rect 2880 -1349 3000 -1316
rect 3030 -1349 3150 -1049
rect 3180 -1122 3300 -1049
rect 3180 -1156 3223 -1122
rect 3257 -1156 3300 -1122
rect 3180 -1202 3300 -1156
rect 3180 -1236 3223 -1202
rect 3257 -1236 3300 -1202
rect 3180 -1282 3300 -1236
rect 3180 -1316 3223 -1282
rect 3257 -1316 3300 -1282
rect 3180 -1349 3300 -1316
rect 3660 -1122 3780 -1049
rect 3660 -1156 3703 -1122
rect 3737 -1156 3780 -1122
rect 3660 -1202 3780 -1156
rect 3660 -1236 3703 -1202
rect 3737 -1236 3780 -1202
rect 3660 -1282 3780 -1236
rect 3660 -1316 3703 -1282
rect 3737 -1316 3780 -1282
rect 3660 -1349 3780 -1316
rect 3810 -1122 3930 -1049
rect 3810 -1156 3853 -1122
rect 3887 -1156 3930 -1122
rect 3810 -1202 3930 -1156
rect 3810 -1236 3853 -1202
rect 3887 -1236 3930 -1202
rect 3810 -1282 3930 -1236
rect 3810 -1316 3853 -1282
rect 3887 -1316 3930 -1282
rect 3810 -1349 3930 -1316
rect 3990 -1122 4110 -1049
rect 3990 -1156 4033 -1122
rect 4067 -1156 4110 -1122
rect 3990 -1202 4110 -1156
rect 3990 -1236 4033 -1202
rect 4067 -1236 4110 -1202
rect 3990 -1282 4110 -1236
rect 3990 -1316 4033 -1282
rect 4067 -1316 4110 -1282
rect 3990 -1349 4110 -1316
rect 4140 -1122 4260 -1049
rect 4140 -1156 4183 -1122
rect 4217 -1156 4260 -1122
rect 4140 -1202 4260 -1156
rect 4140 -1236 4183 -1202
rect 4217 -1236 4260 -1202
rect 4140 -1282 4260 -1236
rect 4140 -1316 4183 -1282
rect 4217 -1316 4260 -1282
rect 4140 -1349 4260 -1316
rect 4290 -1122 4410 -1049
rect 4290 -1156 4333 -1122
rect 4367 -1156 4410 -1122
rect 4290 -1202 4410 -1156
rect 4290 -1236 4333 -1202
rect 4367 -1236 4410 -1202
rect 4290 -1282 4410 -1236
rect 4290 -1316 4333 -1282
rect 4367 -1316 4410 -1282
rect 4290 -1349 4410 -1316
rect 4440 -1122 4560 -1049
rect 4440 -1156 4483 -1122
rect 4517 -1156 4560 -1122
rect 4440 -1202 4560 -1156
rect 4440 -1236 4483 -1202
rect 4517 -1236 4560 -1202
rect 4440 -1282 4560 -1236
rect 4440 -1316 4483 -1282
rect 4517 -1316 4560 -1282
rect 4440 -1349 4560 -1316
rect 4590 -1122 4710 -1049
rect 4590 -1156 4633 -1122
rect 4667 -1156 4710 -1122
rect 4590 -1202 4710 -1156
rect 4590 -1236 4633 -1202
rect 4667 -1236 4710 -1202
rect 4590 -1282 4710 -1236
rect 4590 -1316 4633 -1282
rect 4667 -1316 4710 -1282
rect 4590 -1349 4710 -1316
rect 4770 -1122 4890 -1049
rect 4770 -1156 4813 -1122
rect 4847 -1156 4890 -1122
rect 4770 -1202 4890 -1156
rect 4770 -1236 4813 -1202
rect 4847 -1236 4890 -1202
rect 4770 -1282 4890 -1236
rect 4770 -1316 4813 -1282
rect 4847 -1316 4890 -1282
rect 4770 -1349 4890 -1316
rect 4920 -1122 5040 -1049
rect 4920 -1156 4963 -1122
rect 4997 -1156 5040 -1122
rect 4920 -1202 5040 -1156
rect 4920 -1236 4963 -1202
rect 4997 -1236 5040 -1202
rect 4920 -1282 5040 -1236
rect 4920 -1316 4963 -1282
rect 4997 -1316 5040 -1282
rect 4920 -1349 5040 -1316
rect 5390 -1122 5510 -1049
rect 5390 -1156 5433 -1122
rect 5467 -1156 5510 -1122
rect 5390 -1202 5510 -1156
rect 5390 -1236 5433 -1202
rect 5467 -1236 5510 -1202
rect 5390 -1282 5510 -1236
rect 5390 -1316 5433 -1282
rect 5467 -1316 5510 -1282
rect 5390 -1349 5510 -1316
rect 5540 -1122 5660 -1049
rect 5540 -1156 5583 -1122
rect 5617 -1156 5660 -1122
rect 5540 -1202 5660 -1156
rect 5540 -1236 5583 -1202
rect 5617 -1236 5660 -1202
rect 5540 -1282 5660 -1236
rect 5540 -1316 5583 -1282
rect 5617 -1316 5660 -1282
rect 5540 -1349 5660 -1316
rect 5690 -1122 5810 -1049
rect 5690 -1156 5733 -1122
rect 5767 -1156 5810 -1122
rect 5690 -1202 5810 -1156
rect 5690 -1236 5733 -1202
rect 5767 -1236 5810 -1202
rect 5690 -1282 5810 -1236
rect 5690 -1316 5733 -1282
rect 5767 -1316 5810 -1282
rect 5690 -1349 5810 -1316
rect 5870 -1122 5990 -1049
rect 5870 -1156 5913 -1122
rect 5947 -1156 5990 -1122
rect 5870 -1202 5990 -1156
rect 5870 -1236 5913 -1202
rect 5947 -1236 5990 -1202
rect 5870 -1282 5990 -1236
rect 5870 -1316 5913 -1282
rect 5947 -1316 5990 -1282
rect 5870 -1349 5990 -1316
rect 6020 -1122 6140 -1049
rect 6020 -1156 6063 -1122
rect 6097 -1156 6140 -1122
rect 6020 -1202 6140 -1156
rect 6020 -1236 6063 -1202
rect 6097 -1236 6140 -1202
rect 6020 -1282 6140 -1236
rect 6020 -1316 6063 -1282
rect 6097 -1316 6140 -1282
rect 6020 -1349 6140 -1316
rect 6170 -1122 6290 -1049
rect 6170 -1156 6213 -1122
rect 6247 -1156 6290 -1122
rect 6170 -1202 6290 -1156
rect 6170 -1236 6213 -1202
rect 6247 -1236 6290 -1202
rect 6170 -1282 6290 -1236
rect 6170 -1316 6213 -1282
rect 6247 -1316 6290 -1282
rect 6170 -1349 6290 -1316
rect 6320 -1122 6440 -1049
rect 6320 -1156 6363 -1122
rect 6397 -1156 6440 -1122
rect 6320 -1202 6440 -1156
rect 6320 -1236 6363 -1202
rect 6397 -1236 6440 -1202
rect 6320 -1282 6440 -1236
rect 6320 -1316 6363 -1282
rect 6397 -1316 6440 -1282
rect 6320 -1349 6440 -1316
rect 6470 -1122 6590 -1049
rect 6470 -1156 6513 -1122
rect 6547 -1156 6590 -1122
rect 6470 -1202 6590 -1156
rect 6470 -1236 6513 -1202
rect 6547 -1236 6590 -1202
rect 6470 -1282 6590 -1236
rect 6470 -1316 6513 -1282
rect 6547 -1316 6590 -1282
rect 6470 -1349 6590 -1316
rect 6650 -1122 6770 -1049
rect 6650 -1156 6693 -1122
rect 6727 -1156 6770 -1122
rect 6650 -1202 6770 -1156
rect 6650 -1236 6693 -1202
rect 6727 -1236 6770 -1202
rect 6650 -1282 6770 -1236
rect 6650 -1316 6693 -1282
rect 6727 -1316 6770 -1282
rect 6650 -1349 6770 -1316
rect 6800 -1349 6920 -1049
rect 6950 -1122 7070 -1049
rect 6950 -1156 6993 -1122
rect 7027 -1156 7070 -1122
rect 6950 -1202 7070 -1156
rect 6950 -1236 6993 -1202
rect 7027 -1236 7070 -1202
rect 6950 -1282 7070 -1236
rect 6950 -1316 6993 -1282
rect 7027 -1316 7070 -1282
rect 6950 -1349 7070 -1316
rect 1020 -1762 1140 -1729
rect 1020 -1796 1063 -1762
rect 1097 -1796 1140 -1762
rect 1020 -1842 1140 -1796
rect 1020 -1876 1063 -1842
rect 1097 -1876 1140 -1842
rect 1020 -1922 1140 -1876
rect 1020 -1956 1063 -1922
rect 1097 -1956 1140 -1922
rect 1020 -2029 1140 -1956
rect 1170 -2029 1290 -1729
rect 1320 -1762 1440 -1729
rect 1320 -1796 1363 -1762
rect 1397 -1796 1440 -1762
rect 1320 -1842 1440 -1796
rect 1320 -1876 1363 -1842
rect 1397 -1876 1440 -1842
rect 1320 -1922 1440 -1876
rect 1320 -1956 1363 -1922
rect 1397 -1956 1440 -1922
rect 1320 -2029 1440 -1956
rect 1470 -2029 1590 -1729
rect 1620 -1762 1740 -1729
rect 1620 -1796 1663 -1762
rect 1697 -1796 1740 -1762
rect 1620 -1842 1740 -1796
rect 1620 -1876 1663 -1842
rect 1697 -1876 1740 -1842
rect 1620 -1922 1740 -1876
rect 1620 -1956 1663 -1922
rect 1697 -1956 1740 -1922
rect 1620 -2029 1740 -1956
rect 1800 -1762 1920 -1729
rect 1800 -1796 1843 -1762
rect 1877 -1796 1920 -1762
rect 1800 -1842 1920 -1796
rect 1800 -1876 1843 -1842
rect 1877 -1876 1920 -1842
rect 1800 -1922 1920 -1876
rect 1800 -1956 1843 -1922
rect 1877 -1956 1920 -1922
rect 1800 -2029 1920 -1956
rect 1950 -1762 2070 -1729
rect 1950 -1796 1993 -1762
rect 2027 -1796 2070 -1762
rect 1950 -1842 2070 -1796
rect 1950 -1876 1993 -1842
rect 2027 -1876 2070 -1842
rect 1950 -1922 2070 -1876
rect 1950 -1956 1993 -1922
rect 2027 -1956 2070 -1922
rect 1950 -2029 2070 -1956
rect 2100 -1762 2220 -1729
rect 2100 -1796 2143 -1762
rect 2177 -1796 2220 -1762
rect 2100 -1842 2220 -1796
rect 2100 -1876 2143 -1842
rect 2177 -1876 2220 -1842
rect 2100 -1922 2220 -1876
rect 2100 -1956 2143 -1922
rect 2177 -1956 2220 -1922
rect 2100 -2029 2220 -1956
rect 2250 -1762 2370 -1729
rect 2250 -1796 2293 -1762
rect 2327 -1796 2370 -1762
rect 2250 -1842 2370 -1796
rect 2250 -1876 2293 -1842
rect 2327 -1876 2370 -1842
rect 2250 -1922 2370 -1876
rect 2250 -1956 2293 -1922
rect 2327 -1956 2370 -1922
rect 2250 -2029 2370 -1956
rect 2400 -1762 2520 -1729
rect 2400 -1796 2443 -1762
rect 2477 -1796 2520 -1762
rect 2400 -1842 2520 -1796
rect 2400 -1876 2443 -1842
rect 2477 -1876 2520 -1842
rect 2400 -1922 2520 -1876
rect 2400 -1956 2443 -1922
rect 2477 -1956 2520 -1922
rect 2400 -2029 2520 -1956
rect 2580 -1762 2700 -1729
rect 2580 -1796 2623 -1762
rect 2657 -1796 2700 -1762
rect 2580 -1842 2700 -1796
rect 2580 -1876 2623 -1842
rect 2657 -1876 2700 -1842
rect 2580 -1922 2700 -1876
rect 2580 -1956 2623 -1922
rect 2657 -1956 2700 -1922
rect 2580 -2029 2700 -1956
rect 2730 -2029 2850 -1729
rect 2880 -1762 3000 -1729
rect 2880 -1796 2923 -1762
rect 2957 -1796 3000 -1762
rect 2880 -1842 3000 -1796
rect 2880 -1876 2923 -1842
rect 2957 -1876 3000 -1842
rect 2880 -1922 3000 -1876
rect 2880 -1956 2923 -1922
rect 2957 -1956 3000 -1922
rect 2880 -2029 3000 -1956
rect 3030 -2029 3150 -1729
rect 3180 -1762 3300 -1729
rect 3180 -1796 3223 -1762
rect 3257 -1796 3300 -1762
rect 3180 -1842 3300 -1796
rect 3180 -1876 3223 -1842
rect 3257 -1876 3300 -1842
rect 3180 -1922 3300 -1876
rect 3180 -1956 3223 -1922
rect 3257 -1956 3300 -1922
rect 3180 -2029 3300 -1956
rect 3660 -1762 3780 -1729
rect 3660 -1796 3703 -1762
rect 3737 -1796 3780 -1762
rect 3660 -1842 3780 -1796
rect 3660 -1876 3703 -1842
rect 3737 -1876 3780 -1842
rect 3660 -1922 3780 -1876
rect 3660 -1956 3703 -1922
rect 3737 -1956 3780 -1922
rect 3660 -2029 3780 -1956
rect 3810 -1762 3930 -1729
rect 3810 -1796 3853 -1762
rect 3887 -1796 3930 -1762
rect 3810 -1842 3930 -1796
rect 3810 -1876 3853 -1842
rect 3887 -1876 3930 -1842
rect 3810 -1922 3930 -1876
rect 3810 -1956 3853 -1922
rect 3887 -1956 3930 -1922
rect 3810 -2029 3930 -1956
rect 3990 -1762 4110 -1729
rect 3990 -1796 4033 -1762
rect 4067 -1796 4110 -1762
rect 3990 -1842 4110 -1796
rect 3990 -1876 4033 -1842
rect 4067 -1876 4110 -1842
rect 3990 -1922 4110 -1876
rect 3990 -1956 4033 -1922
rect 4067 -1956 4110 -1922
rect 3990 -2029 4110 -1956
rect 4140 -1762 4260 -1729
rect 4140 -1796 4183 -1762
rect 4217 -1796 4260 -1762
rect 4140 -1842 4260 -1796
rect 4140 -1876 4183 -1842
rect 4217 -1876 4260 -1842
rect 4140 -1922 4260 -1876
rect 4140 -1956 4183 -1922
rect 4217 -1956 4260 -1922
rect 4140 -2029 4260 -1956
rect 4290 -1762 4410 -1729
rect 4290 -1796 4333 -1762
rect 4367 -1796 4410 -1762
rect 4290 -1842 4410 -1796
rect 4290 -1876 4333 -1842
rect 4367 -1876 4410 -1842
rect 4290 -1922 4410 -1876
rect 4290 -1956 4333 -1922
rect 4367 -1956 4410 -1922
rect 4290 -2029 4410 -1956
rect 4440 -1762 4560 -1729
rect 4440 -1796 4483 -1762
rect 4517 -1796 4560 -1762
rect 4440 -1842 4560 -1796
rect 4440 -1876 4483 -1842
rect 4517 -1876 4560 -1842
rect 4440 -1922 4560 -1876
rect 4440 -1956 4483 -1922
rect 4517 -1956 4560 -1922
rect 4440 -2029 4560 -1956
rect 4590 -1762 4710 -1729
rect 4590 -1796 4633 -1762
rect 4667 -1796 4710 -1762
rect 4590 -1842 4710 -1796
rect 4590 -1876 4633 -1842
rect 4667 -1876 4710 -1842
rect 4590 -1922 4710 -1876
rect 4590 -1956 4633 -1922
rect 4667 -1956 4710 -1922
rect 4590 -2029 4710 -1956
rect 4770 -1762 4890 -1729
rect 4770 -1796 4813 -1762
rect 4847 -1796 4890 -1762
rect 4770 -1842 4890 -1796
rect 4770 -1876 4813 -1842
rect 4847 -1876 4890 -1842
rect 4770 -1922 4890 -1876
rect 4770 -1956 4813 -1922
rect 4847 -1956 4890 -1922
rect 4770 -2029 4890 -1956
rect 4920 -1762 5040 -1729
rect 4920 -1796 4963 -1762
rect 4997 -1796 5040 -1762
rect 4920 -1842 5040 -1796
rect 4920 -1876 4963 -1842
rect 4997 -1876 5040 -1842
rect 4920 -1922 5040 -1876
rect 4920 -1956 4963 -1922
rect 4997 -1956 5040 -1922
rect 4920 -2029 5040 -1956
rect 5390 -1762 5510 -1729
rect 5390 -1796 5433 -1762
rect 5467 -1796 5510 -1762
rect 5390 -1842 5510 -1796
rect 5390 -1876 5433 -1842
rect 5467 -1876 5510 -1842
rect 5390 -1922 5510 -1876
rect 5390 -1956 5433 -1922
rect 5467 -1956 5510 -1922
rect 5390 -2029 5510 -1956
rect 5540 -1762 5660 -1729
rect 5540 -1796 5583 -1762
rect 5617 -1796 5660 -1762
rect 5540 -1842 5660 -1796
rect 5540 -1876 5583 -1842
rect 5617 -1876 5660 -1842
rect 5540 -1922 5660 -1876
rect 5540 -1956 5583 -1922
rect 5617 -1956 5660 -1922
rect 5540 -2029 5660 -1956
rect 5690 -1762 5810 -1729
rect 5690 -1796 5733 -1762
rect 5767 -1796 5810 -1762
rect 5690 -1842 5810 -1796
rect 5690 -1876 5733 -1842
rect 5767 -1876 5810 -1842
rect 5690 -1922 5810 -1876
rect 5690 -1956 5733 -1922
rect 5767 -1956 5810 -1922
rect 5690 -2029 5810 -1956
rect 5870 -1762 5990 -1729
rect 5870 -1796 5913 -1762
rect 5947 -1796 5990 -1762
rect 5870 -1842 5990 -1796
rect 5870 -1876 5913 -1842
rect 5947 -1876 5990 -1842
rect 5870 -1922 5990 -1876
rect 5870 -1956 5913 -1922
rect 5947 -1956 5990 -1922
rect 5870 -2029 5990 -1956
rect 6020 -1762 6140 -1729
rect 6020 -1796 6063 -1762
rect 6097 -1796 6140 -1762
rect 6020 -1842 6140 -1796
rect 6020 -1876 6063 -1842
rect 6097 -1876 6140 -1842
rect 6020 -1922 6140 -1876
rect 6020 -1956 6063 -1922
rect 6097 -1956 6140 -1922
rect 6020 -2029 6140 -1956
rect 6170 -1762 6290 -1729
rect 6170 -1796 6213 -1762
rect 6247 -1796 6290 -1762
rect 6170 -1842 6290 -1796
rect 6170 -1876 6213 -1842
rect 6247 -1876 6290 -1842
rect 6170 -1922 6290 -1876
rect 6170 -1956 6213 -1922
rect 6247 -1956 6290 -1922
rect 6170 -2029 6290 -1956
rect 6320 -1762 6440 -1729
rect 6320 -1796 6363 -1762
rect 6397 -1796 6440 -1762
rect 6320 -1842 6440 -1796
rect 6320 -1876 6363 -1842
rect 6397 -1876 6440 -1842
rect 6320 -1922 6440 -1876
rect 6320 -1956 6363 -1922
rect 6397 -1956 6440 -1922
rect 6320 -2029 6440 -1956
rect 6470 -1762 6590 -1729
rect 6470 -1796 6513 -1762
rect 6547 -1796 6590 -1762
rect 6470 -1842 6590 -1796
rect 6470 -1876 6513 -1842
rect 6547 -1876 6590 -1842
rect 6470 -1922 6590 -1876
rect 6470 -1956 6513 -1922
rect 6547 -1956 6590 -1922
rect 6470 -2029 6590 -1956
rect 6650 -1762 6770 -1729
rect 6650 -1796 6693 -1762
rect 6727 -1796 6770 -1762
rect 6650 -1842 6770 -1796
rect 6650 -1876 6693 -1842
rect 6727 -1876 6770 -1842
rect 6650 -1922 6770 -1876
rect 6650 -1956 6693 -1922
rect 6727 -1956 6770 -1922
rect 6650 -2029 6770 -1956
rect 6800 -2029 6920 -1729
rect 6950 -1762 7070 -1729
rect 6950 -1796 6993 -1762
rect 7027 -1796 7070 -1762
rect 6950 -1842 7070 -1796
rect 6950 -1876 6993 -1842
rect 7027 -1876 7070 -1842
rect 6950 -1922 7070 -1876
rect 6950 -1956 6993 -1922
rect 7027 -1956 7070 -1922
rect 6950 -2029 7070 -1956
rect 1171 -3942 1291 -3869
rect 1171 -3976 1214 -3942
rect 1248 -3976 1291 -3942
rect 1171 -4022 1291 -3976
rect 1171 -4056 1214 -4022
rect 1248 -4056 1291 -4022
rect 1171 -4102 1291 -4056
rect 1171 -4136 1214 -4102
rect 1248 -4136 1291 -4102
rect 1171 -4169 1291 -4136
rect 1321 -3942 1441 -3869
rect 1321 -3976 1364 -3942
rect 1398 -3976 1441 -3942
rect 1321 -4022 1441 -3976
rect 1321 -4056 1364 -4022
rect 1398 -4056 1441 -4022
rect 1321 -4102 1441 -4056
rect 1321 -4136 1364 -4102
rect 1398 -4136 1441 -4102
rect 1321 -4169 1441 -4136
rect 1471 -3942 1591 -3869
rect 1471 -3976 1514 -3942
rect 1548 -3976 1591 -3942
rect 1471 -4022 1591 -3976
rect 1471 -4056 1514 -4022
rect 1548 -4056 1591 -4022
rect 1471 -4102 1591 -4056
rect 1471 -4136 1514 -4102
rect 1548 -4136 1591 -4102
rect 1471 -4169 1591 -4136
rect 1621 -3942 1741 -3869
rect 1621 -3976 1664 -3942
rect 1698 -3976 1741 -3942
rect 1621 -4022 1741 -3976
rect 1621 -4056 1664 -4022
rect 1698 -4056 1741 -4022
rect 1621 -4102 1741 -4056
rect 1621 -4136 1664 -4102
rect 1698 -4136 1741 -4102
rect 1621 -4169 1741 -4136
rect 1801 -3942 1921 -3869
rect 1801 -3976 1844 -3942
rect 1878 -3976 1921 -3942
rect 1801 -4022 1921 -3976
rect 1801 -4056 1844 -4022
rect 1878 -4056 1921 -4022
rect 1801 -4102 1921 -4056
rect 1801 -4136 1844 -4102
rect 1878 -4136 1921 -4102
rect 1801 -4169 1921 -4136
rect 1951 -3942 2071 -3869
rect 1951 -3976 1994 -3942
rect 2028 -3976 2071 -3942
rect 1951 -4022 2071 -3976
rect 1951 -4056 1994 -4022
rect 2028 -4056 2071 -4022
rect 1951 -4102 2071 -4056
rect 1951 -4136 1994 -4102
rect 2028 -4136 2071 -4102
rect 1951 -4169 2071 -4136
rect 2101 -3942 2221 -3869
rect 2101 -3976 2144 -3942
rect 2178 -3976 2221 -3942
rect 2101 -4022 2221 -3976
rect 2101 -4056 2144 -4022
rect 2178 -4056 2221 -4022
rect 2101 -4102 2221 -4056
rect 2101 -4136 2144 -4102
rect 2178 -4136 2221 -4102
rect 2101 -4169 2221 -4136
rect 2251 -3942 2371 -3869
rect 2251 -3976 2294 -3942
rect 2328 -3976 2371 -3942
rect 2251 -4022 2371 -3976
rect 2251 -4056 2294 -4022
rect 2328 -4056 2371 -4022
rect 2251 -4102 2371 -4056
rect 2251 -4136 2294 -4102
rect 2328 -4136 2371 -4102
rect 2251 -4169 2371 -4136
rect 2401 -3942 2521 -3869
rect 2401 -3976 2444 -3942
rect 2478 -3976 2521 -3942
rect 2401 -4022 2521 -3976
rect 2401 -4056 2444 -4022
rect 2478 -4056 2521 -4022
rect 2401 -4102 2521 -4056
rect 2401 -4136 2444 -4102
rect 2478 -4136 2521 -4102
rect 2401 -4169 2521 -4136
rect 2581 -3942 2701 -3869
rect 2581 -3976 2624 -3942
rect 2658 -3976 2701 -3942
rect 2581 -4022 2701 -3976
rect 2581 -4056 2624 -4022
rect 2658 -4056 2701 -4022
rect 2581 -4102 2701 -4056
rect 2581 -4136 2624 -4102
rect 2658 -4136 2701 -4102
rect 2581 -4169 2701 -4136
rect 2731 -4169 2851 -3869
rect 2881 -4169 3001 -3869
rect 3031 -3942 3151 -3869
rect 3031 -3976 3074 -3942
rect 3108 -3976 3151 -3942
rect 3031 -4022 3151 -3976
rect 3031 -4056 3074 -4022
rect 3108 -4056 3151 -4022
rect 3031 -4102 3151 -4056
rect 3031 -4136 3074 -4102
rect 3108 -4136 3151 -4102
rect 3031 -4169 3151 -4136
rect 3521 -3942 3641 -3869
rect 3521 -3976 3564 -3942
rect 3598 -3976 3641 -3942
rect 3521 -4022 3641 -3976
rect 3521 -4056 3564 -4022
rect 3598 -4056 3641 -4022
rect 3521 -4102 3641 -4056
rect 3521 -4136 3564 -4102
rect 3598 -4136 3641 -4102
rect 3521 -4169 3641 -4136
rect 3671 -3942 3791 -3869
rect 3671 -3976 3714 -3942
rect 3748 -3976 3791 -3942
rect 3671 -4022 3791 -3976
rect 3671 -4056 3714 -4022
rect 3748 -4056 3791 -4022
rect 3671 -4102 3791 -4056
rect 3671 -4136 3714 -4102
rect 3748 -4136 3791 -4102
rect 3671 -4169 3791 -4136
rect 3851 -3942 3971 -3869
rect 3851 -3976 3894 -3942
rect 3928 -3976 3971 -3942
rect 3851 -4022 3971 -3976
rect 3851 -4056 3894 -4022
rect 3928 -4056 3971 -4022
rect 3851 -4102 3971 -4056
rect 3851 -4136 3894 -4102
rect 3928 -4136 3971 -4102
rect 3851 -4169 3971 -4136
rect 4001 -3942 4121 -3869
rect 4001 -3976 4044 -3942
rect 4078 -3976 4121 -3942
rect 4001 -4022 4121 -3976
rect 4001 -4056 4044 -4022
rect 4078 -4056 4121 -4022
rect 4001 -4102 4121 -4056
rect 4001 -4136 4044 -4102
rect 4078 -4136 4121 -4102
rect 4001 -4169 4121 -4136
rect 4151 -3942 4271 -3869
rect 4151 -3976 4194 -3942
rect 4228 -3976 4271 -3942
rect 4151 -4022 4271 -3976
rect 4151 -4056 4194 -4022
rect 4228 -4056 4271 -4022
rect 4151 -4102 4271 -4056
rect 4151 -4136 4194 -4102
rect 4228 -4136 4271 -4102
rect 4151 -4169 4271 -4136
rect 4301 -3942 4421 -3869
rect 4301 -3976 4344 -3942
rect 4378 -3976 4421 -3942
rect 4301 -4022 4421 -3976
rect 4301 -4056 4344 -4022
rect 4378 -4056 4421 -4022
rect 4301 -4102 4421 -4056
rect 4301 -4136 4344 -4102
rect 4378 -4136 4421 -4102
rect 4301 -4169 4421 -4136
rect 4451 -3942 4571 -3869
rect 4451 -3976 4494 -3942
rect 4528 -3976 4571 -3942
rect 4451 -4022 4571 -3976
rect 4451 -4056 4494 -4022
rect 4528 -4056 4571 -4022
rect 4451 -4102 4571 -4056
rect 4451 -4136 4494 -4102
rect 4528 -4136 4571 -4102
rect 4451 -4169 4571 -4136
rect 4631 -3942 4751 -3869
rect 4631 -3976 4674 -3942
rect 4708 -3976 4751 -3942
rect 4631 -4022 4751 -3976
rect 4631 -4056 4674 -4022
rect 4708 -4056 4751 -4022
rect 4631 -4102 4751 -4056
rect 4631 -4136 4674 -4102
rect 4708 -4136 4751 -4102
rect 4631 -4169 4751 -4136
rect 4781 -3942 4901 -3869
rect 4781 -3976 4824 -3942
rect 4858 -3976 4901 -3942
rect 4781 -4022 4901 -3976
rect 4781 -4056 4824 -4022
rect 4858 -4056 4901 -4022
rect 4781 -4102 4901 -4056
rect 4781 -4136 4824 -4102
rect 4858 -4136 4901 -4102
rect 4781 -4169 4901 -4136
rect 5261 -3943 5381 -3870
rect 5261 -3977 5304 -3943
rect 5338 -3977 5381 -3943
rect 5261 -4023 5381 -3977
rect 5261 -4057 5304 -4023
rect 5338 -4057 5381 -4023
rect 5261 -4103 5381 -4057
rect 5261 -4137 5304 -4103
rect 5338 -4137 5381 -4103
rect 5261 -4170 5381 -4137
rect 5411 -3943 5531 -3870
rect 5411 -3977 5454 -3943
rect 5488 -3977 5531 -3943
rect 5411 -4023 5531 -3977
rect 5411 -4057 5454 -4023
rect 5488 -4057 5531 -4023
rect 5411 -4103 5531 -4057
rect 5411 -4137 5454 -4103
rect 5488 -4137 5531 -4103
rect 5411 -4170 5531 -4137
rect 5561 -3943 5681 -3870
rect 5561 -3977 5604 -3943
rect 5638 -3977 5681 -3943
rect 5561 -4023 5681 -3977
rect 5561 -4057 5604 -4023
rect 5638 -4057 5681 -4023
rect 5561 -4103 5681 -4057
rect 5561 -4137 5604 -4103
rect 5638 -4137 5681 -4103
rect 5561 -4170 5681 -4137
rect 5711 -3943 5831 -3870
rect 5711 -3977 5754 -3943
rect 5788 -3977 5831 -3943
rect 5711 -4023 5831 -3977
rect 5711 -4057 5754 -4023
rect 5788 -4057 5831 -4023
rect 5711 -4103 5831 -4057
rect 5711 -4137 5754 -4103
rect 5788 -4137 5831 -4103
rect 5711 -4170 5831 -4137
rect 5891 -3943 6011 -3870
rect 5891 -3977 5934 -3943
rect 5968 -3977 6011 -3943
rect 5891 -4023 6011 -3977
rect 5891 -4057 5934 -4023
rect 5968 -4057 6011 -4023
rect 5891 -4103 6011 -4057
rect 5891 -4137 5934 -4103
rect 5968 -4137 6011 -4103
rect 5891 -4170 6011 -4137
rect 6041 -3943 6161 -3870
rect 6041 -3977 6084 -3943
rect 6118 -3977 6161 -3943
rect 6041 -4023 6161 -3977
rect 6041 -4057 6084 -4023
rect 6118 -4057 6161 -4023
rect 6041 -4103 6161 -4057
rect 6041 -4137 6084 -4103
rect 6118 -4137 6161 -4103
rect 6041 -4170 6161 -4137
rect 6191 -3943 6311 -3870
rect 6191 -3977 6234 -3943
rect 6268 -3977 6311 -3943
rect 6191 -4023 6311 -3977
rect 6191 -4057 6234 -4023
rect 6268 -4057 6311 -4023
rect 6191 -4103 6311 -4057
rect 6191 -4137 6234 -4103
rect 6268 -4137 6311 -4103
rect 6191 -4170 6311 -4137
rect 6341 -3943 6461 -3870
rect 6341 -3977 6384 -3943
rect 6418 -3977 6461 -3943
rect 6341 -4023 6461 -3977
rect 6341 -4057 6384 -4023
rect 6418 -4057 6461 -4023
rect 6341 -4103 6461 -4057
rect 6341 -4137 6384 -4103
rect 6418 -4137 6461 -4103
rect 6341 -4170 6461 -4137
rect 6491 -3943 6611 -3870
rect 6491 -3977 6534 -3943
rect 6568 -3977 6611 -3943
rect 6491 -4023 6611 -3977
rect 6491 -4057 6534 -4023
rect 6568 -4057 6611 -4023
rect 6491 -4103 6611 -4057
rect 6491 -4137 6534 -4103
rect 6568 -4137 6611 -4103
rect 6491 -4170 6611 -4137
rect 6671 -3943 6791 -3870
rect 6671 -3977 6714 -3943
rect 6748 -3977 6791 -3943
rect 6671 -4023 6791 -3977
rect 6671 -4057 6714 -4023
rect 6748 -4057 6791 -4023
rect 6671 -4103 6791 -4057
rect 6671 -4137 6714 -4103
rect 6748 -4137 6791 -4103
rect 6671 -4170 6791 -4137
rect 6821 -4170 6941 -3870
rect 6971 -4170 7091 -3870
rect 7121 -3943 7241 -3870
rect 7121 -3977 7164 -3943
rect 7198 -3977 7241 -3943
rect 7121 -4023 7241 -3977
rect 7121 -4057 7164 -4023
rect 7198 -4057 7241 -4023
rect 7121 -4103 7241 -4057
rect 7121 -4137 7164 -4103
rect 7198 -4137 7241 -4103
rect 7121 -4170 7241 -4137
rect 1060 -4662 1180 -4629
rect 1060 -4696 1103 -4662
rect 1137 -4696 1180 -4662
rect 1060 -4742 1180 -4696
rect 1060 -4776 1103 -4742
rect 1137 -4776 1180 -4742
rect 1060 -4822 1180 -4776
rect 1060 -4856 1103 -4822
rect 1137 -4856 1180 -4822
rect 1060 -4929 1180 -4856
rect 1210 -4662 1330 -4629
rect 1210 -4696 1253 -4662
rect 1287 -4696 1330 -4662
rect 1210 -4742 1330 -4696
rect 1210 -4776 1253 -4742
rect 1287 -4776 1330 -4742
rect 1210 -4822 1330 -4776
rect 1210 -4856 1253 -4822
rect 1287 -4856 1330 -4822
rect 1210 -4929 1330 -4856
rect 1360 -4662 1480 -4629
rect 1360 -4696 1403 -4662
rect 1437 -4696 1480 -4662
rect 1360 -4742 1480 -4696
rect 1360 -4776 1403 -4742
rect 1437 -4776 1480 -4742
rect 1360 -4822 1480 -4776
rect 1360 -4856 1403 -4822
rect 1437 -4856 1480 -4822
rect 1360 -4929 1480 -4856
rect 1510 -4662 1630 -4629
rect 1510 -4696 1553 -4662
rect 1587 -4696 1630 -4662
rect 1510 -4742 1630 -4696
rect 1510 -4776 1553 -4742
rect 1587 -4776 1630 -4742
rect 1510 -4822 1630 -4776
rect 1510 -4856 1553 -4822
rect 1587 -4856 1630 -4822
rect 1510 -4929 1630 -4856
rect 1660 -4662 1780 -4629
rect 1660 -4696 1703 -4662
rect 1737 -4696 1780 -4662
rect 1660 -4742 1780 -4696
rect 1660 -4776 1703 -4742
rect 1737 -4776 1780 -4742
rect 1660 -4822 1780 -4776
rect 1660 -4856 1703 -4822
rect 1737 -4856 1780 -4822
rect 1660 -4929 1780 -4856
rect 1840 -4662 1960 -4629
rect 1840 -4696 1883 -4662
rect 1917 -4696 1960 -4662
rect 1840 -4742 1960 -4696
rect 1840 -4776 1883 -4742
rect 1917 -4776 1960 -4742
rect 1840 -4822 1960 -4776
rect 1840 -4856 1883 -4822
rect 1917 -4856 1960 -4822
rect 1840 -4929 1960 -4856
rect 1990 -4662 2110 -4629
rect 1990 -4696 2033 -4662
rect 2067 -4696 2110 -4662
rect 1990 -4742 2110 -4696
rect 1990 -4776 2033 -4742
rect 2067 -4776 2110 -4742
rect 1990 -4822 2110 -4776
rect 1990 -4856 2033 -4822
rect 2067 -4856 2110 -4822
rect 1990 -4929 2110 -4856
rect 2140 -4662 2260 -4629
rect 2140 -4696 2183 -4662
rect 2217 -4696 2260 -4662
rect 2140 -4742 2260 -4696
rect 2140 -4776 2183 -4742
rect 2217 -4776 2260 -4742
rect 2140 -4822 2260 -4776
rect 2140 -4856 2183 -4822
rect 2217 -4856 2260 -4822
rect 2140 -4929 2260 -4856
rect 2290 -4662 2410 -4629
rect 2290 -4696 2333 -4662
rect 2367 -4696 2410 -4662
rect 2290 -4742 2410 -4696
rect 2290 -4776 2333 -4742
rect 2367 -4776 2410 -4742
rect 2290 -4822 2410 -4776
rect 2290 -4856 2333 -4822
rect 2367 -4856 2410 -4822
rect 2290 -4929 2410 -4856
rect 2440 -4662 2560 -4629
rect 2440 -4696 2483 -4662
rect 2517 -4696 2560 -4662
rect 2440 -4742 2560 -4696
rect 2440 -4776 2483 -4742
rect 2517 -4776 2560 -4742
rect 2440 -4822 2560 -4776
rect 2440 -4856 2483 -4822
rect 2517 -4856 2560 -4822
rect 2440 -4929 2560 -4856
rect 2620 -4662 2740 -4629
rect 2620 -4696 2663 -4662
rect 2697 -4696 2740 -4662
rect 2620 -4742 2740 -4696
rect 2620 -4776 2663 -4742
rect 2697 -4776 2740 -4742
rect 2620 -4822 2740 -4776
rect 2620 -4856 2663 -4822
rect 2697 -4856 2740 -4822
rect 2620 -4929 2740 -4856
rect 2770 -4929 2890 -4629
rect 2920 -4929 3040 -4629
rect 3070 -4929 3190 -4629
rect 3220 -4662 3340 -4629
rect 3220 -4696 3263 -4662
rect 3297 -4696 3340 -4662
rect 3220 -4742 3340 -4696
rect 3220 -4776 3263 -4742
rect 3297 -4776 3340 -4742
rect 3220 -4822 3340 -4776
rect 3220 -4856 3263 -4822
rect 3297 -4856 3340 -4822
rect 3220 -4929 3340 -4856
rect 3721 -4663 3841 -4630
rect 3721 -4697 3764 -4663
rect 3798 -4697 3841 -4663
rect 3721 -4743 3841 -4697
rect 3721 -4777 3764 -4743
rect 3798 -4777 3841 -4743
rect 3721 -4823 3841 -4777
rect 3721 -4857 3764 -4823
rect 3798 -4857 3841 -4823
rect 3721 -4930 3841 -4857
rect 3871 -4663 3991 -4630
rect 3871 -4697 3914 -4663
rect 3948 -4697 3991 -4663
rect 3871 -4743 3991 -4697
rect 3871 -4777 3914 -4743
rect 3948 -4777 3991 -4743
rect 3871 -4823 3991 -4777
rect 3871 -4857 3914 -4823
rect 3948 -4857 3991 -4823
rect 3871 -4930 3991 -4857
rect 4051 -4663 4171 -4630
rect 4051 -4697 4094 -4663
rect 4128 -4697 4171 -4663
rect 4051 -4743 4171 -4697
rect 4051 -4777 4094 -4743
rect 4128 -4777 4171 -4743
rect 4051 -4823 4171 -4777
rect 4051 -4857 4094 -4823
rect 4128 -4857 4171 -4823
rect 4051 -4930 4171 -4857
rect 4201 -4663 4321 -4630
rect 4201 -4697 4244 -4663
rect 4278 -4697 4321 -4663
rect 4201 -4743 4321 -4697
rect 4201 -4777 4244 -4743
rect 4278 -4777 4321 -4743
rect 4201 -4823 4321 -4777
rect 4201 -4857 4244 -4823
rect 4278 -4857 4321 -4823
rect 4201 -4930 4321 -4857
rect 4351 -4663 4471 -4630
rect 4351 -4697 4394 -4663
rect 4428 -4697 4471 -4663
rect 4351 -4743 4471 -4697
rect 4351 -4777 4394 -4743
rect 4428 -4777 4471 -4743
rect 4351 -4823 4471 -4777
rect 4351 -4857 4394 -4823
rect 4428 -4857 4471 -4823
rect 4351 -4930 4471 -4857
rect 4501 -4663 4621 -4630
rect 4501 -4697 4544 -4663
rect 4578 -4697 4621 -4663
rect 4501 -4743 4621 -4697
rect 4501 -4777 4544 -4743
rect 4578 -4777 4621 -4743
rect 4501 -4823 4621 -4777
rect 4501 -4857 4544 -4823
rect 4578 -4857 4621 -4823
rect 4501 -4930 4621 -4857
rect 4651 -4663 4771 -4630
rect 4651 -4697 4694 -4663
rect 4728 -4697 4771 -4663
rect 4651 -4743 4771 -4697
rect 4651 -4777 4694 -4743
rect 4728 -4777 4771 -4743
rect 4651 -4823 4771 -4777
rect 4651 -4857 4694 -4823
rect 4728 -4857 4771 -4823
rect 4651 -4930 4771 -4857
rect 4831 -4663 4951 -4630
rect 4831 -4697 4874 -4663
rect 4908 -4697 4951 -4663
rect 4831 -4743 4951 -4697
rect 4831 -4777 4874 -4743
rect 4908 -4777 4951 -4743
rect 4831 -4823 4951 -4777
rect 4831 -4857 4874 -4823
rect 4908 -4857 4951 -4823
rect 4831 -4930 4951 -4857
rect 4981 -4663 5101 -4630
rect 4981 -4697 5024 -4663
rect 5058 -4697 5101 -4663
rect 4981 -4743 5101 -4697
rect 4981 -4777 5024 -4743
rect 5058 -4777 5101 -4743
rect 4981 -4823 5101 -4777
rect 4981 -4857 5024 -4823
rect 5058 -4857 5101 -4823
rect 4981 -4930 5101 -4857
rect 5480 -4663 5600 -4630
rect 5480 -4697 5523 -4663
rect 5557 -4697 5600 -4663
rect 5480 -4743 5600 -4697
rect 5480 -4777 5523 -4743
rect 5557 -4777 5600 -4743
rect 5480 -4823 5600 -4777
rect 5480 -4857 5523 -4823
rect 5557 -4857 5600 -4823
rect 5480 -4930 5600 -4857
rect 5630 -4663 5750 -4630
rect 5630 -4697 5673 -4663
rect 5707 -4697 5750 -4663
rect 5630 -4743 5750 -4697
rect 5630 -4777 5673 -4743
rect 5707 -4777 5750 -4743
rect 5630 -4823 5750 -4777
rect 5630 -4857 5673 -4823
rect 5707 -4857 5750 -4823
rect 5630 -4930 5750 -4857
rect 5780 -4663 5900 -4630
rect 5780 -4697 5823 -4663
rect 5857 -4697 5900 -4663
rect 5780 -4743 5900 -4697
rect 5780 -4777 5823 -4743
rect 5857 -4777 5900 -4743
rect 5780 -4823 5900 -4777
rect 5780 -4857 5823 -4823
rect 5857 -4857 5900 -4823
rect 5780 -4930 5900 -4857
rect 5930 -4663 6050 -4630
rect 5930 -4697 5973 -4663
rect 6007 -4697 6050 -4663
rect 5930 -4743 6050 -4697
rect 5930 -4777 5973 -4743
rect 6007 -4777 6050 -4743
rect 5930 -4823 6050 -4777
rect 5930 -4857 5973 -4823
rect 6007 -4857 6050 -4823
rect 5930 -4930 6050 -4857
rect 6110 -4663 6230 -4630
rect 6110 -4697 6153 -4663
rect 6187 -4697 6230 -4663
rect 6110 -4743 6230 -4697
rect 6110 -4777 6153 -4743
rect 6187 -4777 6230 -4743
rect 6110 -4823 6230 -4777
rect 6110 -4857 6153 -4823
rect 6187 -4857 6230 -4823
rect 6110 -4930 6230 -4857
rect 6260 -4663 6380 -4630
rect 6260 -4697 6303 -4663
rect 6337 -4697 6380 -4663
rect 6260 -4743 6380 -4697
rect 6260 -4777 6303 -4743
rect 6337 -4777 6380 -4743
rect 6260 -4823 6380 -4777
rect 6260 -4857 6303 -4823
rect 6337 -4857 6380 -4823
rect 6260 -4930 6380 -4857
rect 6410 -4663 6530 -4630
rect 6410 -4697 6453 -4663
rect 6487 -4697 6530 -4663
rect 6410 -4743 6530 -4697
rect 6410 -4777 6453 -4743
rect 6487 -4777 6530 -4743
rect 6410 -4823 6530 -4777
rect 6410 -4857 6453 -4823
rect 6487 -4857 6530 -4823
rect 6410 -4930 6530 -4857
rect 6560 -4663 6680 -4630
rect 6560 -4697 6603 -4663
rect 6637 -4697 6680 -4663
rect 6560 -4743 6680 -4697
rect 6560 -4777 6603 -4743
rect 6637 -4777 6680 -4743
rect 6560 -4823 6680 -4777
rect 6560 -4857 6603 -4823
rect 6637 -4857 6680 -4823
rect 6560 -4930 6680 -4857
rect 6710 -4663 6830 -4630
rect 6710 -4697 6753 -4663
rect 6787 -4697 6830 -4663
rect 6710 -4743 6830 -4697
rect 6710 -4777 6753 -4743
rect 6787 -4777 6830 -4743
rect 6710 -4823 6830 -4777
rect 6710 -4857 6753 -4823
rect 6787 -4857 6830 -4823
rect 6710 -4930 6830 -4857
rect 6890 -4663 7010 -4630
rect 6890 -4697 6933 -4663
rect 6967 -4697 7010 -4663
rect 6890 -4743 7010 -4697
rect 6890 -4777 6933 -4743
rect 6967 -4777 7010 -4743
rect 6890 -4823 7010 -4777
rect 6890 -4857 6933 -4823
rect 6967 -4857 7010 -4823
rect 6890 -4930 7010 -4857
rect 7040 -4930 7160 -4630
rect 7190 -4930 7310 -4630
rect 7340 -4663 7460 -4630
rect 7340 -4697 7383 -4663
rect 7417 -4697 7460 -4663
rect 7340 -4743 7460 -4697
rect 7340 -4777 7383 -4743
rect 7417 -4777 7460 -4743
rect 7340 -4823 7460 -4777
rect 7340 -4857 7383 -4823
rect 7417 -4857 7460 -4823
rect 7340 -4930 7460 -4857
rect 1060 -6843 1180 -6770
rect 1060 -6877 1103 -6843
rect 1137 -6877 1180 -6843
rect 1060 -6923 1180 -6877
rect 1060 -6957 1103 -6923
rect 1137 -6957 1180 -6923
rect 1060 -7003 1180 -6957
rect 1060 -7037 1103 -7003
rect 1137 -7037 1180 -7003
rect 1060 -7070 1180 -7037
rect 1210 -7070 1330 -6770
rect 1360 -6843 1480 -6770
rect 1360 -6877 1403 -6843
rect 1437 -6877 1480 -6843
rect 1360 -6923 1480 -6877
rect 1360 -6957 1403 -6923
rect 1437 -6957 1480 -6923
rect 1360 -7003 1480 -6957
rect 1360 -7037 1403 -7003
rect 1437 -7037 1480 -7003
rect 1360 -7070 1480 -7037
rect 1510 -7070 1630 -6770
rect 1660 -6843 1780 -6770
rect 1660 -6877 1703 -6843
rect 1737 -6877 1780 -6843
rect 1660 -6923 1780 -6877
rect 1660 -6957 1703 -6923
rect 1737 -6957 1780 -6923
rect 1660 -7003 1780 -6957
rect 1660 -7037 1703 -7003
rect 1737 -7037 1780 -7003
rect 1660 -7070 1780 -7037
rect 1840 -6843 1960 -6770
rect 1840 -6877 1883 -6843
rect 1917 -6877 1960 -6843
rect 1840 -6923 1960 -6877
rect 1840 -6957 1883 -6923
rect 1917 -6957 1960 -6923
rect 1840 -7003 1960 -6957
rect 1840 -7037 1883 -7003
rect 1917 -7037 1960 -7003
rect 1840 -7070 1960 -7037
rect 1990 -6843 2110 -6770
rect 1990 -6877 2033 -6843
rect 2067 -6877 2110 -6843
rect 1990 -6923 2110 -6877
rect 1990 -6957 2033 -6923
rect 2067 -6957 2110 -6923
rect 1990 -7003 2110 -6957
rect 1990 -7037 2033 -7003
rect 2067 -7037 2110 -7003
rect 1990 -7070 2110 -7037
rect 2140 -6843 2260 -6770
rect 2140 -6877 2183 -6843
rect 2217 -6877 2260 -6843
rect 2140 -6923 2260 -6877
rect 2140 -6957 2183 -6923
rect 2217 -6957 2260 -6923
rect 2140 -7003 2260 -6957
rect 2140 -7037 2183 -7003
rect 2217 -7037 2260 -7003
rect 2140 -7070 2260 -7037
rect 2290 -6843 2410 -6770
rect 2290 -6877 2333 -6843
rect 2367 -6877 2410 -6843
rect 2290 -6923 2410 -6877
rect 2290 -6957 2333 -6923
rect 2367 -6957 2410 -6923
rect 2290 -7003 2410 -6957
rect 2290 -7037 2333 -7003
rect 2367 -7037 2410 -7003
rect 2290 -7070 2410 -7037
rect 2440 -6843 2560 -6770
rect 2440 -6877 2483 -6843
rect 2517 -6877 2560 -6843
rect 2440 -6923 2560 -6877
rect 2440 -6957 2483 -6923
rect 2517 -6957 2560 -6923
rect 2440 -7003 2560 -6957
rect 2440 -7037 2483 -7003
rect 2517 -7037 2560 -7003
rect 2440 -7070 2560 -7037
rect 2620 -6843 2740 -6770
rect 2620 -6877 2663 -6843
rect 2697 -6877 2740 -6843
rect 2620 -6923 2740 -6877
rect 2620 -6957 2663 -6923
rect 2697 -6957 2740 -6923
rect 2620 -7003 2740 -6957
rect 2620 -7037 2663 -7003
rect 2697 -7037 2740 -7003
rect 2620 -7070 2740 -7037
rect 2770 -7070 2890 -6770
rect 2920 -6843 3040 -6770
rect 2920 -6877 2963 -6843
rect 2997 -6877 3040 -6843
rect 2920 -6923 3040 -6877
rect 2920 -6957 2963 -6923
rect 2997 -6957 3040 -6923
rect 2920 -7003 3040 -6957
rect 2920 -7037 2963 -7003
rect 2997 -7037 3040 -7003
rect 2920 -7070 3040 -7037
rect 3070 -7070 3190 -6770
rect 3220 -6843 3340 -6770
rect 3220 -6877 3263 -6843
rect 3297 -6877 3340 -6843
rect 3220 -6923 3340 -6877
rect 3220 -6957 3263 -6923
rect 3297 -6957 3340 -6923
rect 3220 -7003 3340 -6957
rect 3220 -7037 3263 -7003
rect 3297 -7037 3340 -7003
rect 3220 -7070 3340 -7037
rect 3720 -6843 3840 -6770
rect 3720 -6877 3763 -6843
rect 3797 -6877 3840 -6843
rect 3720 -6923 3840 -6877
rect 3720 -6957 3763 -6923
rect 3797 -6957 3840 -6923
rect 3720 -7003 3840 -6957
rect 3720 -7037 3763 -7003
rect 3797 -7037 3840 -7003
rect 3720 -7070 3840 -7037
rect 3870 -6843 3990 -6770
rect 3870 -6877 3913 -6843
rect 3947 -6877 3990 -6843
rect 3870 -6923 3990 -6877
rect 3870 -6957 3913 -6923
rect 3947 -6957 3990 -6923
rect 3870 -7003 3990 -6957
rect 3870 -7037 3913 -7003
rect 3947 -7037 3990 -7003
rect 3870 -7070 3990 -7037
rect 4050 -6843 4170 -6770
rect 4050 -6877 4093 -6843
rect 4127 -6877 4170 -6843
rect 4050 -6923 4170 -6877
rect 4050 -6957 4093 -6923
rect 4127 -6957 4170 -6923
rect 4050 -7003 4170 -6957
rect 4050 -7037 4093 -7003
rect 4127 -7037 4170 -7003
rect 4050 -7070 4170 -7037
rect 4200 -6843 4320 -6770
rect 4200 -6877 4243 -6843
rect 4277 -6877 4320 -6843
rect 4200 -6923 4320 -6877
rect 4200 -6957 4243 -6923
rect 4277 -6957 4320 -6923
rect 4200 -7003 4320 -6957
rect 4200 -7037 4243 -7003
rect 4277 -7037 4320 -7003
rect 4200 -7070 4320 -7037
rect 4350 -6843 4470 -6770
rect 4350 -6877 4393 -6843
rect 4427 -6877 4470 -6843
rect 4350 -6923 4470 -6877
rect 4350 -6957 4393 -6923
rect 4427 -6957 4470 -6923
rect 4350 -7003 4470 -6957
rect 4350 -7037 4393 -7003
rect 4427 -7037 4470 -7003
rect 4350 -7070 4470 -7037
rect 4500 -6843 4620 -6770
rect 4500 -6877 4543 -6843
rect 4577 -6877 4620 -6843
rect 4500 -6923 4620 -6877
rect 4500 -6957 4543 -6923
rect 4577 -6957 4620 -6923
rect 4500 -7003 4620 -6957
rect 4500 -7037 4543 -7003
rect 4577 -7037 4620 -7003
rect 4500 -7070 4620 -7037
rect 4650 -6843 4770 -6770
rect 4650 -6877 4693 -6843
rect 4727 -6877 4770 -6843
rect 4650 -6923 4770 -6877
rect 4650 -6957 4693 -6923
rect 4727 -6957 4770 -6923
rect 4650 -7003 4770 -6957
rect 4650 -7037 4693 -7003
rect 4727 -7037 4770 -7003
rect 4650 -7070 4770 -7037
rect 4830 -6843 4950 -6770
rect 4830 -6877 4873 -6843
rect 4907 -6877 4950 -6843
rect 4830 -6923 4950 -6877
rect 4830 -6957 4873 -6923
rect 4907 -6957 4950 -6923
rect 4830 -7003 4950 -6957
rect 4830 -7037 4873 -7003
rect 4907 -7037 4950 -7003
rect 4830 -7070 4950 -7037
rect 4980 -6843 5100 -6770
rect 4980 -6877 5023 -6843
rect 5057 -6877 5100 -6843
rect 4980 -6923 5100 -6877
rect 4980 -6957 5023 -6923
rect 5057 -6957 5100 -6923
rect 4980 -7003 5100 -6957
rect 4980 -7037 5023 -7003
rect 5057 -7037 5100 -7003
rect 4980 -7070 5100 -7037
rect 5449 -6843 5569 -6770
rect 5449 -6877 5492 -6843
rect 5526 -6877 5569 -6843
rect 5449 -6923 5569 -6877
rect 5449 -6957 5492 -6923
rect 5526 -6957 5569 -6923
rect 5449 -7003 5569 -6957
rect 5449 -7037 5492 -7003
rect 5526 -7037 5569 -7003
rect 5449 -7070 5569 -7037
rect 5599 -6843 5719 -6770
rect 5599 -6877 5642 -6843
rect 5676 -6877 5719 -6843
rect 5599 -6923 5719 -6877
rect 5599 -6957 5642 -6923
rect 5676 -6957 5719 -6923
rect 5599 -7003 5719 -6957
rect 5599 -7037 5642 -7003
rect 5676 -7037 5719 -7003
rect 5599 -7070 5719 -7037
rect 5749 -6843 5869 -6770
rect 5749 -6877 5792 -6843
rect 5826 -6877 5869 -6843
rect 5749 -6923 5869 -6877
rect 5749 -6957 5792 -6923
rect 5826 -6957 5869 -6923
rect 5749 -7003 5869 -6957
rect 5749 -7037 5792 -7003
rect 5826 -7037 5869 -7003
rect 5749 -7070 5869 -7037
rect 5929 -6843 6049 -6770
rect 5929 -6877 5972 -6843
rect 6006 -6877 6049 -6843
rect 5929 -6923 6049 -6877
rect 5929 -6957 5972 -6923
rect 6006 -6957 6049 -6923
rect 5929 -7003 6049 -6957
rect 5929 -7037 5972 -7003
rect 6006 -7037 6049 -7003
rect 5929 -7070 6049 -7037
rect 6079 -6843 6199 -6770
rect 6079 -6877 6122 -6843
rect 6156 -6877 6199 -6843
rect 6079 -6923 6199 -6877
rect 6079 -6957 6122 -6923
rect 6156 -6957 6199 -6923
rect 6079 -7003 6199 -6957
rect 6079 -7037 6122 -7003
rect 6156 -7037 6199 -7003
rect 6079 -7070 6199 -7037
rect 6229 -6843 6349 -6770
rect 6229 -6877 6272 -6843
rect 6306 -6877 6349 -6843
rect 6229 -6923 6349 -6877
rect 6229 -6957 6272 -6923
rect 6306 -6957 6349 -6923
rect 6229 -7003 6349 -6957
rect 6229 -7037 6272 -7003
rect 6306 -7037 6349 -7003
rect 6229 -7070 6349 -7037
rect 6379 -6843 6499 -6770
rect 6379 -6877 6422 -6843
rect 6456 -6877 6499 -6843
rect 6379 -6923 6499 -6877
rect 6379 -6957 6422 -6923
rect 6456 -6957 6499 -6923
rect 6379 -7003 6499 -6957
rect 6379 -7037 6422 -7003
rect 6456 -7037 6499 -7003
rect 6379 -7070 6499 -7037
rect 6529 -6843 6649 -6770
rect 6529 -6877 6572 -6843
rect 6606 -6877 6649 -6843
rect 6529 -6923 6649 -6877
rect 6529 -6957 6572 -6923
rect 6606 -6957 6649 -6923
rect 6529 -7003 6649 -6957
rect 6529 -7037 6572 -7003
rect 6606 -7037 6649 -7003
rect 6529 -7070 6649 -7037
rect 6709 -6843 6829 -6770
rect 6709 -6877 6752 -6843
rect 6786 -6877 6829 -6843
rect 6709 -6923 6829 -6877
rect 6709 -6957 6752 -6923
rect 6786 -6957 6829 -6923
rect 6709 -7003 6829 -6957
rect 6709 -7037 6752 -7003
rect 6786 -7037 6829 -7003
rect 6709 -7070 6829 -7037
rect 6859 -7070 6979 -6770
rect 7009 -6843 7129 -6770
rect 7009 -6877 7052 -6843
rect 7086 -6877 7129 -6843
rect 7009 -6923 7129 -6877
rect 7009 -6957 7052 -6923
rect 7086 -6957 7129 -6923
rect 7009 -7003 7129 -6957
rect 7009 -7037 7052 -7003
rect 7086 -7037 7129 -7003
rect 7009 -7070 7129 -7037
rect 1060 -7483 1180 -7450
rect 1060 -7517 1103 -7483
rect 1137 -7517 1180 -7483
rect 1060 -7563 1180 -7517
rect 1060 -7597 1103 -7563
rect 1137 -7597 1180 -7563
rect 1060 -7643 1180 -7597
rect 1060 -7677 1103 -7643
rect 1137 -7677 1180 -7643
rect 1060 -7750 1180 -7677
rect 1210 -7750 1330 -7450
rect 1360 -7483 1480 -7450
rect 1360 -7517 1403 -7483
rect 1437 -7517 1480 -7483
rect 1360 -7563 1480 -7517
rect 1360 -7597 1403 -7563
rect 1437 -7597 1480 -7563
rect 1360 -7643 1480 -7597
rect 1360 -7677 1403 -7643
rect 1437 -7677 1480 -7643
rect 1360 -7750 1480 -7677
rect 1510 -7750 1630 -7450
rect 1660 -7483 1780 -7450
rect 1660 -7517 1703 -7483
rect 1737 -7517 1780 -7483
rect 1660 -7563 1780 -7517
rect 1660 -7597 1703 -7563
rect 1737 -7597 1780 -7563
rect 1660 -7643 1780 -7597
rect 1660 -7677 1703 -7643
rect 1737 -7677 1780 -7643
rect 1660 -7750 1780 -7677
rect 1840 -7483 1960 -7450
rect 1840 -7517 1883 -7483
rect 1917 -7517 1960 -7483
rect 1840 -7563 1960 -7517
rect 1840 -7597 1883 -7563
rect 1917 -7597 1960 -7563
rect 1840 -7643 1960 -7597
rect 1840 -7677 1883 -7643
rect 1917 -7677 1960 -7643
rect 1840 -7750 1960 -7677
rect 1990 -7483 2110 -7450
rect 1990 -7517 2033 -7483
rect 2067 -7517 2110 -7483
rect 1990 -7563 2110 -7517
rect 1990 -7597 2033 -7563
rect 2067 -7597 2110 -7563
rect 1990 -7643 2110 -7597
rect 1990 -7677 2033 -7643
rect 2067 -7677 2110 -7643
rect 1990 -7750 2110 -7677
rect 2140 -7483 2260 -7450
rect 2140 -7517 2183 -7483
rect 2217 -7517 2260 -7483
rect 2140 -7563 2260 -7517
rect 2140 -7597 2183 -7563
rect 2217 -7597 2260 -7563
rect 2140 -7643 2260 -7597
rect 2140 -7677 2183 -7643
rect 2217 -7677 2260 -7643
rect 2140 -7750 2260 -7677
rect 2290 -7483 2410 -7450
rect 2290 -7517 2333 -7483
rect 2367 -7517 2410 -7483
rect 2290 -7563 2410 -7517
rect 2290 -7597 2333 -7563
rect 2367 -7597 2410 -7563
rect 2290 -7643 2410 -7597
rect 2290 -7677 2333 -7643
rect 2367 -7677 2410 -7643
rect 2290 -7750 2410 -7677
rect 2440 -7483 2560 -7450
rect 2440 -7517 2483 -7483
rect 2517 -7517 2560 -7483
rect 2440 -7563 2560 -7517
rect 2440 -7597 2483 -7563
rect 2517 -7597 2560 -7563
rect 2440 -7643 2560 -7597
rect 2440 -7677 2483 -7643
rect 2517 -7677 2560 -7643
rect 2440 -7750 2560 -7677
rect 2620 -7483 2740 -7450
rect 2620 -7517 2663 -7483
rect 2697 -7517 2740 -7483
rect 2620 -7563 2740 -7517
rect 2620 -7597 2663 -7563
rect 2697 -7597 2740 -7563
rect 2620 -7643 2740 -7597
rect 2620 -7677 2663 -7643
rect 2697 -7677 2740 -7643
rect 2620 -7750 2740 -7677
rect 2770 -7750 2890 -7450
rect 2920 -7483 3040 -7450
rect 2920 -7517 2963 -7483
rect 2997 -7517 3040 -7483
rect 2920 -7563 3040 -7517
rect 2920 -7597 2963 -7563
rect 2997 -7597 3040 -7563
rect 2920 -7643 3040 -7597
rect 2920 -7677 2963 -7643
rect 2997 -7677 3040 -7643
rect 2920 -7750 3040 -7677
rect 3070 -7750 3190 -7450
rect 3220 -7483 3340 -7450
rect 3220 -7517 3263 -7483
rect 3297 -7517 3340 -7483
rect 3220 -7563 3340 -7517
rect 3220 -7597 3263 -7563
rect 3297 -7597 3340 -7563
rect 3220 -7643 3340 -7597
rect 3220 -7677 3263 -7643
rect 3297 -7677 3340 -7643
rect 3220 -7750 3340 -7677
rect 3720 -7483 3840 -7450
rect 3720 -7517 3763 -7483
rect 3797 -7517 3840 -7483
rect 3720 -7563 3840 -7517
rect 3720 -7597 3763 -7563
rect 3797 -7597 3840 -7563
rect 3720 -7643 3840 -7597
rect 3720 -7677 3763 -7643
rect 3797 -7677 3840 -7643
rect 3720 -7750 3840 -7677
rect 3870 -7483 3990 -7450
rect 3870 -7517 3913 -7483
rect 3947 -7517 3990 -7483
rect 3870 -7563 3990 -7517
rect 3870 -7597 3913 -7563
rect 3947 -7597 3990 -7563
rect 3870 -7643 3990 -7597
rect 3870 -7677 3913 -7643
rect 3947 -7677 3990 -7643
rect 3870 -7750 3990 -7677
rect 4050 -7483 4170 -7450
rect 4050 -7517 4093 -7483
rect 4127 -7517 4170 -7483
rect 4050 -7563 4170 -7517
rect 4050 -7597 4093 -7563
rect 4127 -7597 4170 -7563
rect 4050 -7643 4170 -7597
rect 4050 -7677 4093 -7643
rect 4127 -7677 4170 -7643
rect 4050 -7750 4170 -7677
rect 4200 -7483 4320 -7450
rect 4200 -7517 4243 -7483
rect 4277 -7517 4320 -7483
rect 4200 -7563 4320 -7517
rect 4200 -7597 4243 -7563
rect 4277 -7597 4320 -7563
rect 4200 -7643 4320 -7597
rect 4200 -7677 4243 -7643
rect 4277 -7677 4320 -7643
rect 4200 -7750 4320 -7677
rect 4350 -7483 4470 -7450
rect 4350 -7517 4393 -7483
rect 4427 -7517 4470 -7483
rect 4350 -7563 4470 -7517
rect 4350 -7597 4393 -7563
rect 4427 -7597 4470 -7563
rect 4350 -7643 4470 -7597
rect 4350 -7677 4393 -7643
rect 4427 -7677 4470 -7643
rect 4350 -7750 4470 -7677
rect 4500 -7483 4620 -7450
rect 4500 -7517 4543 -7483
rect 4577 -7517 4620 -7483
rect 4500 -7563 4620 -7517
rect 4500 -7597 4543 -7563
rect 4577 -7597 4620 -7563
rect 4500 -7643 4620 -7597
rect 4500 -7677 4543 -7643
rect 4577 -7677 4620 -7643
rect 4500 -7750 4620 -7677
rect 4650 -7483 4770 -7450
rect 4650 -7517 4693 -7483
rect 4727 -7517 4770 -7483
rect 4650 -7563 4770 -7517
rect 4650 -7597 4693 -7563
rect 4727 -7597 4770 -7563
rect 4650 -7643 4770 -7597
rect 4650 -7677 4693 -7643
rect 4727 -7677 4770 -7643
rect 4650 -7750 4770 -7677
rect 4830 -7483 4950 -7450
rect 4830 -7517 4873 -7483
rect 4907 -7517 4950 -7483
rect 4830 -7563 4950 -7517
rect 4830 -7597 4873 -7563
rect 4907 -7597 4950 -7563
rect 4830 -7643 4950 -7597
rect 4830 -7677 4873 -7643
rect 4907 -7677 4950 -7643
rect 4830 -7750 4950 -7677
rect 4980 -7483 5100 -7450
rect 4980 -7517 5023 -7483
rect 5057 -7517 5100 -7483
rect 4980 -7563 5100 -7517
rect 4980 -7597 5023 -7563
rect 5057 -7597 5100 -7563
rect 4980 -7643 5100 -7597
rect 4980 -7677 5023 -7643
rect 5057 -7677 5100 -7643
rect 4980 -7750 5100 -7677
rect 5449 -7483 5569 -7450
rect 5449 -7517 5492 -7483
rect 5526 -7517 5569 -7483
rect 5449 -7563 5569 -7517
rect 5449 -7597 5492 -7563
rect 5526 -7597 5569 -7563
rect 5449 -7643 5569 -7597
rect 5449 -7677 5492 -7643
rect 5526 -7677 5569 -7643
rect 5449 -7750 5569 -7677
rect 5599 -7483 5719 -7450
rect 5599 -7517 5642 -7483
rect 5676 -7517 5719 -7483
rect 5599 -7563 5719 -7517
rect 5599 -7597 5642 -7563
rect 5676 -7597 5719 -7563
rect 5599 -7643 5719 -7597
rect 5599 -7677 5642 -7643
rect 5676 -7677 5719 -7643
rect 5599 -7750 5719 -7677
rect 5749 -7483 5869 -7450
rect 5749 -7517 5792 -7483
rect 5826 -7517 5869 -7483
rect 5749 -7563 5869 -7517
rect 5749 -7597 5792 -7563
rect 5826 -7597 5869 -7563
rect 5749 -7643 5869 -7597
rect 5749 -7677 5792 -7643
rect 5826 -7677 5869 -7643
rect 5749 -7750 5869 -7677
rect 5929 -7483 6049 -7450
rect 5929 -7517 5972 -7483
rect 6006 -7517 6049 -7483
rect 5929 -7563 6049 -7517
rect 5929 -7597 5972 -7563
rect 6006 -7597 6049 -7563
rect 5929 -7643 6049 -7597
rect 5929 -7677 5972 -7643
rect 6006 -7677 6049 -7643
rect 5929 -7750 6049 -7677
rect 6079 -7483 6199 -7450
rect 6079 -7517 6122 -7483
rect 6156 -7517 6199 -7483
rect 6079 -7563 6199 -7517
rect 6079 -7597 6122 -7563
rect 6156 -7597 6199 -7563
rect 6079 -7643 6199 -7597
rect 6079 -7677 6122 -7643
rect 6156 -7677 6199 -7643
rect 6079 -7750 6199 -7677
rect 6229 -7483 6349 -7450
rect 6229 -7517 6272 -7483
rect 6306 -7517 6349 -7483
rect 6229 -7563 6349 -7517
rect 6229 -7597 6272 -7563
rect 6306 -7597 6349 -7563
rect 6229 -7643 6349 -7597
rect 6229 -7677 6272 -7643
rect 6306 -7677 6349 -7643
rect 6229 -7750 6349 -7677
rect 6379 -7483 6499 -7450
rect 6379 -7517 6422 -7483
rect 6456 -7517 6499 -7483
rect 6379 -7563 6499 -7517
rect 6379 -7597 6422 -7563
rect 6456 -7597 6499 -7563
rect 6379 -7643 6499 -7597
rect 6379 -7677 6422 -7643
rect 6456 -7677 6499 -7643
rect 6379 -7750 6499 -7677
rect 6529 -7483 6649 -7450
rect 6529 -7517 6572 -7483
rect 6606 -7517 6649 -7483
rect 6529 -7563 6649 -7517
rect 6529 -7597 6572 -7563
rect 6606 -7597 6649 -7563
rect 6529 -7643 6649 -7597
rect 6529 -7677 6572 -7643
rect 6606 -7677 6649 -7643
rect 6529 -7750 6649 -7677
rect 6709 -7483 6829 -7450
rect 6709 -7517 6752 -7483
rect 6786 -7517 6829 -7483
rect 6709 -7563 6829 -7517
rect 6709 -7597 6752 -7563
rect 6786 -7597 6829 -7563
rect 6709 -7643 6829 -7597
rect 6709 -7677 6752 -7643
rect 6786 -7677 6829 -7643
rect 6709 -7750 6829 -7677
rect 6859 -7750 6979 -7450
rect 7009 -7483 7129 -7450
rect 7009 -7517 7052 -7483
rect 7086 -7517 7129 -7483
rect 7009 -7563 7129 -7517
rect 7009 -7597 7052 -7563
rect 7086 -7597 7129 -7563
rect 7009 -7643 7129 -7597
rect 7009 -7677 7052 -7643
rect 7086 -7677 7129 -7643
rect 7009 -7750 7129 -7677
rect 1020 -9663 1140 -9590
rect 1020 -9697 1063 -9663
rect 1097 -9697 1140 -9663
rect 1020 -9743 1140 -9697
rect 1020 -9777 1063 -9743
rect 1097 -9777 1140 -9743
rect 1020 -9823 1140 -9777
rect 1020 -9857 1063 -9823
rect 1097 -9857 1140 -9823
rect 1020 -9890 1140 -9857
rect 1170 -9890 1290 -9590
rect 1320 -9663 1440 -9590
rect 1320 -9697 1363 -9663
rect 1397 -9697 1440 -9663
rect 1320 -9743 1440 -9697
rect 1320 -9777 1363 -9743
rect 1397 -9777 1440 -9743
rect 1320 -9823 1440 -9777
rect 1320 -9857 1363 -9823
rect 1397 -9857 1440 -9823
rect 1320 -9890 1440 -9857
rect 1470 -9890 1590 -9590
rect 1620 -9663 1740 -9590
rect 1620 -9697 1663 -9663
rect 1697 -9697 1740 -9663
rect 1620 -9743 1740 -9697
rect 1620 -9777 1663 -9743
rect 1697 -9777 1740 -9743
rect 1620 -9823 1740 -9777
rect 1620 -9857 1663 -9823
rect 1697 -9857 1740 -9823
rect 1620 -9890 1740 -9857
rect 1800 -9663 1920 -9590
rect 1800 -9697 1843 -9663
rect 1877 -9697 1920 -9663
rect 1800 -9743 1920 -9697
rect 1800 -9777 1843 -9743
rect 1877 -9777 1920 -9743
rect 1800 -9823 1920 -9777
rect 1800 -9857 1843 -9823
rect 1877 -9857 1920 -9823
rect 1800 -9890 1920 -9857
rect 1950 -9663 2070 -9590
rect 1950 -9697 1993 -9663
rect 2027 -9697 2070 -9663
rect 1950 -9743 2070 -9697
rect 1950 -9777 1993 -9743
rect 2027 -9777 2070 -9743
rect 1950 -9823 2070 -9777
rect 1950 -9857 1993 -9823
rect 2027 -9857 2070 -9823
rect 1950 -9890 2070 -9857
rect 2100 -9663 2220 -9590
rect 2100 -9697 2143 -9663
rect 2177 -9697 2220 -9663
rect 2100 -9743 2220 -9697
rect 2100 -9777 2143 -9743
rect 2177 -9777 2220 -9743
rect 2100 -9823 2220 -9777
rect 2100 -9857 2143 -9823
rect 2177 -9857 2220 -9823
rect 2100 -9890 2220 -9857
rect 2250 -9663 2370 -9590
rect 2250 -9697 2293 -9663
rect 2327 -9697 2370 -9663
rect 2250 -9743 2370 -9697
rect 2250 -9777 2293 -9743
rect 2327 -9777 2370 -9743
rect 2250 -9823 2370 -9777
rect 2250 -9857 2293 -9823
rect 2327 -9857 2370 -9823
rect 2250 -9890 2370 -9857
rect 2400 -9663 2520 -9590
rect 2400 -9697 2443 -9663
rect 2477 -9697 2520 -9663
rect 2400 -9743 2520 -9697
rect 2400 -9777 2443 -9743
rect 2477 -9777 2520 -9743
rect 2400 -9823 2520 -9777
rect 2400 -9857 2443 -9823
rect 2477 -9857 2520 -9823
rect 2400 -9890 2520 -9857
rect 2580 -9663 2700 -9590
rect 2580 -9697 2623 -9663
rect 2657 -9697 2700 -9663
rect 2580 -9743 2700 -9697
rect 2580 -9777 2623 -9743
rect 2657 -9777 2700 -9743
rect 2580 -9823 2700 -9777
rect 2580 -9857 2623 -9823
rect 2657 -9857 2700 -9823
rect 2580 -9890 2700 -9857
rect 2730 -9890 2850 -9590
rect 2880 -9663 3000 -9590
rect 2880 -9697 2923 -9663
rect 2957 -9697 3000 -9663
rect 2880 -9743 3000 -9697
rect 2880 -9777 2923 -9743
rect 2957 -9777 3000 -9743
rect 2880 -9823 3000 -9777
rect 2880 -9857 2923 -9823
rect 2957 -9857 3000 -9823
rect 2880 -9890 3000 -9857
rect 3030 -9890 3150 -9590
rect 3180 -9663 3300 -9590
rect 3180 -9697 3223 -9663
rect 3257 -9697 3300 -9663
rect 3180 -9743 3300 -9697
rect 3180 -9777 3223 -9743
rect 3257 -9777 3300 -9743
rect 3180 -9823 3300 -9777
rect 3180 -9857 3223 -9823
rect 3257 -9857 3300 -9823
rect 3180 -9890 3300 -9857
rect 3660 -9663 3780 -9590
rect 3660 -9697 3703 -9663
rect 3737 -9697 3780 -9663
rect 3660 -9743 3780 -9697
rect 3660 -9777 3703 -9743
rect 3737 -9777 3780 -9743
rect 3660 -9823 3780 -9777
rect 3660 -9857 3703 -9823
rect 3737 -9857 3780 -9823
rect 3660 -9890 3780 -9857
rect 3810 -9663 3930 -9590
rect 3810 -9697 3853 -9663
rect 3887 -9697 3930 -9663
rect 3810 -9743 3930 -9697
rect 3810 -9777 3853 -9743
rect 3887 -9777 3930 -9743
rect 3810 -9823 3930 -9777
rect 3810 -9857 3853 -9823
rect 3887 -9857 3930 -9823
rect 3810 -9890 3930 -9857
rect 3990 -9663 4110 -9590
rect 3990 -9697 4033 -9663
rect 4067 -9697 4110 -9663
rect 3990 -9743 4110 -9697
rect 3990 -9777 4033 -9743
rect 4067 -9777 4110 -9743
rect 3990 -9823 4110 -9777
rect 3990 -9857 4033 -9823
rect 4067 -9857 4110 -9823
rect 3990 -9890 4110 -9857
rect 4140 -9663 4260 -9590
rect 4140 -9697 4183 -9663
rect 4217 -9697 4260 -9663
rect 4140 -9743 4260 -9697
rect 4140 -9777 4183 -9743
rect 4217 -9777 4260 -9743
rect 4140 -9823 4260 -9777
rect 4140 -9857 4183 -9823
rect 4217 -9857 4260 -9823
rect 4140 -9890 4260 -9857
rect 4290 -9663 4410 -9590
rect 4290 -9697 4333 -9663
rect 4367 -9697 4410 -9663
rect 4290 -9743 4410 -9697
rect 4290 -9777 4333 -9743
rect 4367 -9777 4410 -9743
rect 4290 -9823 4410 -9777
rect 4290 -9857 4333 -9823
rect 4367 -9857 4410 -9823
rect 4290 -9890 4410 -9857
rect 4440 -9663 4560 -9590
rect 4440 -9697 4483 -9663
rect 4517 -9697 4560 -9663
rect 4440 -9743 4560 -9697
rect 4440 -9777 4483 -9743
rect 4517 -9777 4560 -9743
rect 4440 -9823 4560 -9777
rect 4440 -9857 4483 -9823
rect 4517 -9857 4560 -9823
rect 4440 -9890 4560 -9857
rect 4590 -9663 4710 -9590
rect 4590 -9697 4633 -9663
rect 4667 -9697 4710 -9663
rect 4590 -9743 4710 -9697
rect 4590 -9777 4633 -9743
rect 4667 -9777 4710 -9743
rect 4590 -9823 4710 -9777
rect 4590 -9857 4633 -9823
rect 4667 -9857 4710 -9823
rect 4590 -9890 4710 -9857
rect 4770 -9663 4890 -9590
rect 4770 -9697 4813 -9663
rect 4847 -9697 4890 -9663
rect 4770 -9743 4890 -9697
rect 4770 -9777 4813 -9743
rect 4847 -9777 4890 -9743
rect 4770 -9823 4890 -9777
rect 4770 -9857 4813 -9823
rect 4847 -9857 4890 -9823
rect 4770 -9890 4890 -9857
rect 4920 -9663 5040 -9590
rect 4920 -9697 4963 -9663
rect 4997 -9697 5040 -9663
rect 4920 -9743 5040 -9697
rect 4920 -9777 4963 -9743
rect 4997 -9777 5040 -9743
rect 4920 -9823 5040 -9777
rect 4920 -9857 4963 -9823
rect 4997 -9857 5040 -9823
rect 4920 -9890 5040 -9857
rect 5390 -9663 5510 -9590
rect 5390 -9697 5433 -9663
rect 5467 -9697 5510 -9663
rect 5390 -9743 5510 -9697
rect 5390 -9777 5433 -9743
rect 5467 -9777 5510 -9743
rect 5390 -9823 5510 -9777
rect 5390 -9857 5433 -9823
rect 5467 -9857 5510 -9823
rect 5390 -9890 5510 -9857
rect 5540 -9663 5660 -9590
rect 5540 -9697 5583 -9663
rect 5617 -9697 5660 -9663
rect 5540 -9743 5660 -9697
rect 5540 -9777 5583 -9743
rect 5617 -9777 5660 -9743
rect 5540 -9823 5660 -9777
rect 5540 -9857 5583 -9823
rect 5617 -9857 5660 -9823
rect 5540 -9890 5660 -9857
rect 5690 -9663 5810 -9590
rect 5690 -9697 5733 -9663
rect 5767 -9697 5810 -9663
rect 5690 -9743 5810 -9697
rect 5690 -9777 5733 -9743
rect 5767 -9777 5810 -9743
rect 5690 -9823 5810 -9777
rect 5690 -9857 5733 -9823
rect 5767 -9857 5810 -9823
rect 5690 -9890 5810 -9857
rect 5870 -9663 5990 -9590
rect 5870 -9697 5913 -9663
rect 5947 -9697 5990 -9663
rect 5870 -9743 5990 -9697
rect 5870 -9777 5913 -9743
rect 5947 -9777 5990 -9743
rect 5870 -9823 5990 -9777
rect 5870 -9857 5913 -9823
rect 5947 -9857 5990 -9823
rect 5870 -9890 5990 -9857
rect 6020 -9663 6140 -9590
rect 6020 -9697 6063 -9663
rect 6097 -9697 6140 -9663
rect 6020 -9743 6140 -9697
rect 6020 -9777 6063 -9743
rect 6097 -9777 6140 -9743
rect 6020 -9823 6140 -9777
rect 6020 -9857 6063 -9823
rect 6097 -9857 6140 -9823
rect 6020 -9890 6140 -9857
rect 6170 -9663 6290 -9590
rect 6170 -9697 6213 -9663
rect 6247 -9697 6290 -9663
rect 6170 -9743 6290 -9697
rect 6170 -9777 6213 -9743
rect 6247 -9777 6290 -9743
rect 6170 -9823 6290 -9777
rect 6170 -9857 6213 -9823
rect 6247 -9857 6290 -9823
rect 6170 -9890 6290 -9857
rect 6320 -9663 6440 -9590
rect 6320 -9697 6363 -9663
rect 6397 -9697 6440 -9663
rect 6320 -9743 6440 -9697
rect 6320 -9777 6363 -9743
rect 6397 -9777 6440 -9743
rect 6320 -9823 6440 -9777
rect 6320 -9857 6363 -9823
rect 6397 -9857 6440 -9823
rect 6320 -9890 6440 -9857
rect 6470 -9663 6590 -9590
rect 6470 -9697 6513 -9663
rect 6547 -9697 6590 -9663
rect 6470 -9743 6590 -9697
rect 6470 -9777 6513 -9743
rect 6547 -9777 6590 -9743
rect 6470 -9823 6590 -9777
rect 6470 -9857 6513 -9823
rect 6547 -9857 6590 -9823
rect 6470 -9890 6590 -9857
rect 6650 -9663 6770 -9590
rect 6650 -9697 6693 -9663
rect 6727 -9697 6770 -9663
rect 6650 -9743 6770 -9697
rect 6650 -9777 6693 -9743
rect 6727 -9777 6770 -9743
rect 6650 -9823 6770 -9777
rect 6650 -9857 6693 -9823
rect 6727 -9857 6770 -9823
rect 6650 -9890 6770 -9857
rect 6800 -9890 6920 -9590
rect 6950 -9663 7070 -9590
rect 6950 -9697 6993 -9663
rect 7027 -9697 7070 -9663
rect 6950 -9743 7070 -9697
rect 6950 -9777 6993 -9743
rect 7027 -9777 7070 -9743
rect 6950 -9823 7070 -9777
rect 6950 -9857 6993 -9823
rect 7027 -9857 7070 -9823
rect 6950 -9890 7070 -9857
rect 1020 -10303 1140 -10270
rect 1020 -10337 1063 -10303
rect 1097 -10337 1140 -10303
rect 1020 -10383 1140 -10337
rect 1020 -10417 1063 -10383
rect 1097 -10417 1140 -10383
rect 1020 -10463 1140 -10417
rect 1020 -10497 1063 -10463
rect 1097 -10497 1140 -10463
rect 1020 -10570 1140 -10497
rect 1170 -10570 1290 -10270
rect 1320 -10303 1440 -10270
rect 1320 -10337 1363 -10303
rect 1397 -10337 1440 -10303
rect 1320 -10383 1440 -10337
rect 1320 -10417 1363 -10383
rect 1397 -10417 1440 -10383
rect 1320 -10463 1440 -10417
rect 1320 -10497 1363 -10463
rect 1397 -10497 1440 -10463
rect 1320 -10570 1440 -10497
rect 1470 -10570 1590 -10270
rect 1620 -10303 1740 -10270
rect 1620 -10337 1663 -10303
rect 1697 -10337 1740 -10303
rect 1620 -10383 1740 -10337
rect 1620 -10417 1663 -10383
rect 1697 -10417 1740 -10383
rect 1620 -10463 1740 -10417
rect 1620 -10497 1663 -10463
rect 1697 -10497 1740 -10463
rect 1620 -10570 1740 -10497
rect 1800 -10303 1920 -10270
rect 1800 -10337 1843 -10303
rect 1877 -10337 1920 -10303
rect 1800 -10383 1920 -10337
rect 1800 -10417 1843 -10383
rect 1877 -10417 1920 -10383
rect 1800 -10463 1920 -10417
rect 1800 -10497 1843 -10463
rect 1877 -10497 1920 -10463
rect 1800 -10570 1920 -10497
rect 1950 -10303 2070 -10270
rect 1950 -10337 1993 -10303
rect 2027 -10337 2070 -10303
rect 1950 -10383 2070 -10337
rect 1950 -10417 1993 -10383
rect 2027 -10417 2070 -10383
rect 1950 -10463 2070 -10417
rect 1950 -10497 1993 -10463
rect 2027 -10497 2070 -10463
rect 1950 -10570 2070 -10497
rect 2100 -10303 2220 -10270
rect 2100 -10337 2143 -10303
rect 2177 -10337 2220 -10303
rect 2100 -10383 2220 -10337
rect 2100 -10417 2143 -10383
rect 2177 -10417 2220 -10383
rect 2100 -10463 2220 -10417
rect 2100 -10497 2143 -10463
rect 2177 -10497 2220 -10463
rect 2100 -10570 2220 -10497
rect 2250 -10303 2370 -10270
rect 2250 -10337 2293 -10303
rect 2327 -10337 2370 -10303
rect 2250 -10383 2370 -10337
rect 2250 -10417 2293 -10383
rect 2327 -10417 2370 -10383
rect 2250 -10463 2370 -10417
rect 2250 -10497 2293 -10463
rect 2327 -10497 2370 -10463
rect 2250 -10570 2370 -10497
rect 2400 -10303 2520 -10270
rect 2400 -10337 2443 -10303
rect 2477 -10337 2520 -10303
rect 2400 -10383 2520 -10337
rect 2400 -10417 2443 -10383
rect 2477 -10417 2520 -10383
rect 2400 -10463 2520 -10417
rect 2400 -10497 2443 -10463
rect 2477 -10497 2520 -10463
rect 2400 -10570 2520 -10497
rect 2580 -10303 2700 -10270
rect 2580 -10337 2623 -10303
rect 2657 -10337 2700 -10303
rect 2580 -10383 2700 -10337
rect 2580 -10417 2623 -10383
rect 2657 -10417 2700 -10383
rect 2580 -10463 2700 -10417
rect 2580 -10497 2623 -10463
rect 2657 -10497 2700 -10463
rect 2580 -10570 2700 -10497
rect 2730 -10570 2850 -10270
rect 2880 -10303 3000 -10270
rect 2880 -10337 2923 -10303
rect 2957 -10337 3000 -10303
rect 2880 -10383 3000 -10337
rect 2880 -10417 2923 -10383
rect 2957 -10417 3000 -10383
rect 2880 -10463 3000 -10417
rect 2880 -10497 2923 -10463
rect 2957 -10497 3000 -10463
rect 2880 -10570 3000 -10497
rect 3030 -10570 3150 -10270
rect 3180 -10303 3300 -10270
rect 3180 -10337 3223 -10303
rect 3257 -10337 3300 -10303
rect 3180 -10383 3300 -10337
rect 3180 -10417 3223 -10383
rect 3257 -10417 3300 -10383
rect 3180 -10463 3300 -10417
rect 3180 -10497 3223 -10463
rect 3257 -10497 3300 -10463
rect 3180 -10570 3300 -10497
rect 3660 -10303 3780 -10270
rect 3660 -10337 3703 -10303
rect 3737 -10337 3780 -10303
rect 3660 -10383 3780 -10337
rect 3660 -10417 3703 -10383
rect 3737 -10417 3780 -10383
rect 3660 -10463 3780 -10417
rect 3660 -10497 3703 -10463
rect 3737 -10497 3780 -10463
rect 3660 -10570 3780 -10497
rect 3810 -10303 3930 -10270
rect 3810 -10337 3853 -10303
rect 3887 -10337 3930 -10303
rect 3810 -10383 3930 -10337
rect 3810 -10417 3853 -10383
rect 3887 -10417 3930 -10383
rect 3810 -10463 3930 -10417
rect 3810 -10497 3853 -10463
rect 3887 -10497 3930 -10463
rect 3810 -10570 3930 -10497
rect 3990 -10303 4110 -10270
rect 3990 -10337 4033 -10303
rect 4067 -10337 4110 -10303
rect 3990 -10383 4110 -10337
rect 3990 -10417 4033 -10383
rect 4067 -10417 4110 -10383
rect 3990 -10463 4110 -10417
rect 3990 -10497 4033 -10463
rect 4067 -10497 4110 -10463
rect 3990 -10570 4110 -10497
rect 4140 -10303 4260 -10270
rect 4140 -10337 4183 -10303
rect 4217 -10337 4260 -10303
rect 4140 -10383 4260 -10337
rect 4140 -10417 4183 -10383
rect 4217 -10417 4260 -10383
rect 4140 -10463 4260 -10417
rect 4140 -10497 4183 -10463
rect 4217 -10497 4260 -10463
rect 4140 -10570 4260 -10497
rect 4290 -10303 4410 -10270
rect 4290 -10337 4333 -10303
rect 4367 -10337 4410 -10303
rect 4290 -10383 4410 -10337
rect 4290 -10417 4333 -10383
rect 4367 -10417 4410 -10383
rect 4290 -10463 4410 -10417
rect 4290 -10497 4333 -10463
rect 4367 -10497 4410 -10463
rect 4290 -10570 4410 -10497
rect 4440 -10303 4560 -10270
rect 4440 -10337 4483 -10303
rect 4517 -10337 4560 -10303
rect 4440 -10383 4560 -10337
rect 4440 -10417 4483 -10383
rect 4517 -10417 4560 -10383
rect 4440 -10463 4560 -10417
rect 4440 -10497 4483 -10463
rect 4517 -10497 4560 -10463
rect 4440 -10570 4560 -10497
rect 4590 -10303 4710 -10270
rect 4590 -10337 4633 -10303
rect 4667 -10337 4710 -10303
rect 4590 -10383 4710 -10337
rect 4590 -10417 4633 -10383
rect 4667 -10417 4710 -10383
rect 4590 -10463 4710 -10417
rect 4590 -10497 4633 -10463
rect 4667 -10497 4710 -10463
rect 4590 -10570 4710 -10497
rect 4770 -10303 4890 -10270
rect 4770 -10337 4813 -10303
rect 4847 -10337 4890 -10303
rect 4770 -10383 4890 -10337
rect 4770 -10417 4813 -10383
rect 4847 -10417 4890 -10383
rect 4770 -10463 4890 -10417
rect 4770 -10497 4813 -10463
rect 4847 -10497 4890 -10463
rect 4770 -10570 4890 -10497
rect 4920 -10303 5040 -10270
rect 4920 -10337 4963 -10303
rect 4997 -10337 5040 -10303
rect 4920 -10383 5040 -10337
rect 4920 -10417 4963 -10383
rect 4997 -10417 5040 -10383
rect 4920 -10463 5040 -10417
rect 4920 -10497 4963 -10463
rect 4997 -10497 5040 -10463
rect 4920 -10570 5040 -10497
rect 5390 -10303 5510 -10270
rect 5390 -10337 5433 -10303
rect 5467 -10337 5510 -10303
rect 5390 -10383 5510 -10337
rect 5390 -10417 5433 -10383
rect 5467 -10417 5510 -10383
rect 5390 -10463 5510 -10417
rect 5390 -10497 5433 -10463
rect 5467 -10497 5510 -10463
rect 5390 -10570 5510 -10497
rect 5540 -10303 5660 -10270
rect 5540 -10337 5583 -10303
rect 5617 -10337 5660 -10303
rect 5540 -10383 5660 -10337
rect 5540 -10417 5583 -10383
rect 5617 -10417 5660 -10383
rect 5540 -10463 5660 -10417
rect 5540 -10497 5583 -10463
rect 5617 -10497 5660 -10463
rect 5540 -10570 5660 -10497
rect 5690 -10303 5810 -10270
rect 5690 -10337 5733 -10303
rect 5767 -10337 5810 -10303
rect 5690 -10383 5810 -10337
rect 5690 -10417 5733 -10383
rect 5767 -10417 5810 -10383
rect 5690 -10463 5810 -10417
rect 5690 -10497 5733 -10463
rect 5767 -10497 5810 -10463
rect 5690 -10570 5810 -10497
rect 5870 -10303 5990 -10270
rect 5870 -10337 5913 -10303
rect 5947 -10337 5990 -10303
rect 5870 -10383 5990 -10337
rect 5870 -10417 5913 -10383
rect 5947 -10417 5990 -10383
rect 5870 -10463 5990 -10417
rect 5870 -10497 5913 -10463
rect 5947 -10497 5990 -10463
rect 5870 -10570 5990 -10497
rect 6020 -10303 6140 -10270
rect 6020 -10337 6063 -10303
rect 6097 -10337 6140 -10303
rect 6020 -10383 6140 -10337
rect 6020 -10417 6063 -10383
rect 6097 -10417 6140 -10383
rect 6020 -10463 6140 -10417
rect 6020 -10497 6063 -10463
rect 6097 -10497 6140 -10463
rect 6020 -10570 6140 -10497
rect 6170 -10303 6290 -10270
rect 6170 -10337 6213 -10303
rect 6247 -10337 6290 -10303
rect 6170 -10383 6290 -10337
rect 6170 -10417 6213 -10383
rect 6247 -10417 6290 -10383
rect 6170 -10463 6290 -10417
rect 6170 -10497 6213 -10463
rect 6247 -10497 6290 -10463
rect 6170 -10570 6290 -10497
rect 6320 -10303 6440 -10270
rect 6320 -10337 6363 -10303
rect 6397 -10337 6440 -10303
rect 6320 -10383 6440 -10337
rect 6320 -10417 6363 -10383
rect 6397 -10417 6440 -10383
rect 6320 -10463 6440 -10417
rect 6320 -10497 6363 -10463
rect 6397 -10497 6440 -10463
rect 6320 -10570 6440 -10497
rect 6470 -10303 6590 -10270
rect 6470 -10337 6513 -10303
rect 6547 -10337 6590 -10303
rect 6470 -10383 6590 -10337
rect 6470 -10417 6513 -10383
rect 6547 -10417 6590 -10383
rect 6470 -10463 6590 -10417
rect 6470 -10497 6513 -10463
rect 6547 -10497 6590 -10463
rect 6470 -10570 6590 -10497
rect 6650 -10303 6770 -10270
rect 6650 -10337 6693 -10303
rect 6727 -10337 6770 -10303
rect 6650 -10383 6770 -10337
rect 6650 -10417 6693 -10383
rect 6727 -10417 6770 -10383
rect 6650 -10463 6770 -10417
rect 6650 -10497 6693 -10463
rect 6727 -10497 6770 -10463
rect 6650 -10570 6770 -10497
rect 6800 -10570 6920 -10270
rect 6950 -10303 7070 -10270
rect 6950 -10337 6993 -10303
rect 7027 -10337 7070 -10303
rect 6950 -10383 7070 -10337
rect 6950 -10417 6993 -10383
rect 7027 -10417 7070 -10383
rect 6950 -10463 7070 -10417
rect 6950 -10497 6993 -10463
rect 7027 -10497 7070 -10463
rect 6950 -10570 7070 -10497
rect 1171 -12483 1291 -12410
rect 1171 -12517 1214 -12483
rect 1248 -12517 1291 -12483
rect 1171 -12563 1291 -12517
rect 1171 -12597 1214 -12563
rect 1248 -12597 1291 -12563
rect 1171 -12643 1291 -12597
rect 1171 -12677 1214 -12643
rect 1248 -12677 1291 -12643
rect 1171 -12710 1291 -12677
rect 1321 -12483 1441 -12410
rect 1321 -12517 1364 -12483
rect 1398 -12517 1441 -12483
rect 1321 -12563 1441 -12517
rect 1321 -12597 1364 -12563
rect 1398 -12597 1441 -12563
rect 1321 -12643 1441 -12597
rect 1321 -12677 1364 -12643
rect 1398 -12677 1441 -12643
rect 1321 -12710 1441 -12677
rect 1471 -12483 1591 -12410
rect 1471 -12517 1514 -12483
rect 1548 -12517 1591 -12483
rect 1471 -12563 1591 -12517
rect 1471 -12597 1514 -12563
rect 1548 -12597 1591 -12563
rect 1471 -12643 1591 -12597
rect 1471 -12677 1514 -12643
rect 1548 -12677 1591 -12643
rect 1471 -12710 1591 -12677
rect 1621 -12483 1741 -12410
rect 1621 -12517 1664 -12483
rect 1698 -12517 1741 -12483
rect 1621 -12563 1741 -12517
rect 1621 -12597 1664 -12563
rect 1698 -12597 1741 -12563
rect 1621 -12643 1741 -12597
rect 1621 -12677 1664 -12643
rect 1698 -12677 1741 -12643
rect 1621 -12710 1741 -12677
rect 1801 -12483 1921 -12410
rect 1801 -12517 1844 -12483
rect 1878 -12517 1921 -12483
rect 1801 -12563 1921 -12517
rect 1801 -12597 1844 -12563
rect 1878 -12597 1921 -12563
rect 1801 -12643 1921 -12597
rect 1801 -12677 1844 -12643
rect 1878 -12677 1921 -12643
rect 1801 -12710 1921 -12677
rect 1951 -12483 2071 -12410
rect 1951 -12517 1994 -12483
rect 2028 -12517 2071 -12483
rect 1951 -12563 2071 -12517
rect 1951 -12597 1994 -12563
rect 2028 -12597 2071 -12563
rect 1951 -12643 2071 -12597
rect 1951 -12677 1994 -12643
rect 2028 -12677 2071 -12643
rect 1951 -12710 2071 -12677
rect 2101 -12483 2221 -12410
rect 2101 -12517 2144 -12483
rect 2178 -12517 2221 -12483
rect 2101 -12563 2221 -12517
rect 2101 -12597 2144 -12563
rect 2178 -12597 2221 -12563
rect 2101 -12643 2221 -12597
rect 2101 -12677 2144 -12643
rect 2178 -12677 2221 -12643
rect 2101 -12710 2221 -12677
rect 2251 -12483 2371 -12410
rect 2251 -12517 2294 -12483
rect 2328 -12517 2371 -12483
rect 2251 -12563 2371 -12517
rect 2251 -12597 2294 -12563
rect 2328 -12597 2371 -12563
rect 2251 -12643 2371 -12597
rect 2251 -12677 2294 -12643
rect 2328 -12677 2371 -12643
rect 2251 -12710 2371 -12677
rect 2401 -12483 2521 -12410
rect 2401 -12517 2444 -12483
rect 2478 -12517 2521 -12483
rect 2401 -12563 2521 -12517
rect 2401 -12597 2444 -12563
rect 2478 -12597 2521 -12563
rect 2401 -12643 2521 -12597
rect 2401 -12677 2444 -12643
rect 2478 -12677 2521 -12643
rect 2401 -12710 2521 -12677
rect 2581 -12483 2701 -12410
rect 2581 -12517 2624 -12483
rect 2658 -12517 2701 -12483
rect 2581 -12563 2701 -12517
rect 2581 -12597 2624 -12563
rect 2658 -12597 2701 -12563
rect 2581 -12643 2701 -12597
rect 2581 -12677 2624 -12643
rect 2658 -12677 2701 -12643
rect 2581 -12710 2701 -12677
rect 2731 -12710 2851 -12410
rect 2881 -12710 3001 -12410
rect 3031 -12483 3151 -12410
rect 3031 -12517 3074 -12483
rect 3108 -12517 3151 -12483
rect 3031 -12563 3151 -12517
rect 3031 -12597 3074 -12563
rect 3108 -12597 3151 -12563
rect 3031 -12643 3151 -12597
rect 3031 -12677 3074 -12643
rect 3108 -12677 3151 -12643
rect 3031 -12710 3151 -12677
rect 3521 -12483 3641 -12410
rect 3521 -12517 3564 -12483
rect 3598 -12517 3641 -12483
rect 3521 -12563 3641 -12517
rect 3521 -12597 3564 -12563
rect 3598 -12597 3641 -12563
rect 3521 -12643 3641 -12597
rect 3521 -12677 3564 -12643
rect 3598 -12677 3641 -12643
rect 3521 -12710 3641 -12677
rect 3671 -12483 3791 -12410
rect 3671 -12517 3714 -12483
rect 3748 -12517 3791 -12483
rect 3671 -12563 3791 -12517
rect 3671 -12597 3714 -12563
rect 3748 -12597 3791 -12563
rect 3671 -12643 3791 -12597
rect 3671 -12677 3714 -12643
rect 3748 -12677 3791 -12643
rect 3671 -12710 3791 -12677
rect 3851 -12483 3971 -12410
rect 3851 -12517 3894 -12483
rect 3928 -12517 3971 -12483
rect 3851 -12563 3971 -12517
rect 3851 -12597 3894 -12563
rect 3928 -12597 3971 -12563
rect 3851 -12643 3971 -12597
rect 3851 -12677 3894 -12643
rect 3928 -12677 3971 -12643
rect 3851 -12710 3971 -12677
rect 4001 -12483 4121 -12410
rect 4001 -12517 4044 -12483
rect 4078 -12517 4121 -12483
rect 4001 -12563 4121 -12517
rect 4001 -12597 4044 -12563
rect 4078 -12597 4121 -12563
rect 4001 -12643 4121 -12597
rect 4001 -12677 4044 -12643
rect 4078 -12677 4121 -12643
rect 4001 -12710 4121 -12677
rect 4151 -12483 4271 -12410
rect 4151 -12517 4194 -12483
rect 4228 -12517 4271 -12483
rect 4151 -12563 4271 -12517
rect 4151 -12597 4194 -12563
rect 4228 -12597 4271 -12563
rect 4151 -12643 4271 -12597
rect 4151 -12677 4194 -12643
rect 4228 -12677 4271 -12643
rect 4151 -12710 4271 -12677
rect 4301 -12483 4421 -12410
rect 4301 -12517 4344 -12483
rect 4378 -12517 4421 -12483
rect 4301 -12563 4421 -12517
rect 4301 -12597 4344 -12563
rect 4378 -12597 4421 -12563
rect 4301 -12643 4421 -12597
rect 4301 -12677 4344 -12643
rect 4378 -12677 4421 -12643
rect 4301 -12710 4421 -12677
rect 4451 -12483 4571 -12410
rect 4451 -12517 4494 -12483
rect 4528 -12517 4571 -12483
rect 4451 -12563 4571 -12517
rect 4451 -12597 4494 -12563
rect 4528 -12597 4571 -12563
rect 4451 -12643 4571 -12597
rect 4451 -12677 4494 -12643
rect 4528 -12677 4571 -12643
rect 4451 -12710 4571 -12677
rect 4631 -12483 4751 -12410
rect 4631 -12517 4674 -12483
rect 4708 -12517 4751 -12483
rect 4631 -12563 4751 -12517
rect 4631 -12597 4674 -12563
rect 4708 -12597 4751 -12563
rect 4631 -12643 4751 -12597
rect 4631 -12677 4674 -12643
rect 4708 -12677 4751 -12643
rect 4631 -12710 4751 -12677
rect 4781 -12483 4901 -12410
rect 4781 -12517 4824 -12483
rect 4858 -12517 4901 -12483
rect 4781 -12563 4901 -12517
rect 4781 -12597 4824 -12563
rect 4858 -12597 4901 -12563
rect 4781 -12643 4901 -12597
rect 4781 -12677 4824 -12643
rect 4858 -12677 4901 -12643
rect 4781 -12710 4901 -12677
rect 5261 -12484 5381 -12411
rect 5261 -12518 5304 -12484
rect 5338 -12518 5381 -12484
rect 5261 -12564 5381 -12518
rect 5261 -12598 5304 -12564
rect 5338 -12598 5381 -12564
rect 5261 -12644 5381 -12598
rect 5261 -12678 5304 -12644
rect 5338 -12678 5381 -12644
rect 5261 -12711 5381 -12678
rect 5411 -12484 5531 -12411
rect 5411 -12518 5454 -12484
rect 5488 -12518 5531 -12484
rect 5411 -12564 5531 -12518
rect 5411 -12598 5454 -12564
rect 5488 -12598 5531 -12564
rect 5411 -12644 5531 -12598
rect 5411 -12678 5454 -12644
rect 5488 -12678 5531 -12644
rect 5411 -12711 5531 -12678
rect 5561 -12484 5681 -12411
rect 5561 -12518 5604 -12484
rect 5638 -12518 5681 -12484
rect 5561 -12564 5681 -12518
rect 5561 -12598 5604 -12564
rect 5638 -12598 5681 -12564
rect 5561 -12644 5681 -12598
rect 5561 -12678 5604 -12644
rect 5638 -12678 5681 -12644
rect 5561 -12711 5681 -12678
rect 5711 -12484 5831 -12411
rect 5711 -12518 5754 -12484
rect 5788 -12518 5831 -12484
rect 5711 -12564 5831 -12518
rect 5711 -12598 5754 -12564
rect 5788 -12598 5831 -12564
rect 5711 -12644 5831 -12598
rect 5711 -12678 5754 -12644
rect 5788 -12678 5831 -12644
rect 5711 -12711 5831 -12678
rect 5891 -12484 6011 -12411
rect 5891 -12518 5934 -12484
rect 5968 -12518 6011 -12484
rect 5891 -12564 6011 -12518
rect 5891 -12598 5934 -12564
rect 5968 -12598 6011 -12564
rect 5891 -12644 6011 -12598
rect 5891 -12678 5934 -12644
rect 5968 -12678 6011 -12644
rect 5891 -12711 6011 -12678
rect 6041 -12484 6161 -12411
rect 6041 -12518 6084 -12484
rect 6118 -12518 6161 -12484
rect 6041 -12564 6161 -12518
rect 6041 -12598 6084 -12564
rect 6118 -12598 6161 -12564
rect 6041 -12644 6161 -12598
rect 6041 -12678 6084 -12644
rect 6118 -12678 6161 -12644
rect 6041 -12711 6161 -12678
rect 6191 -12484 6311 -12411
rect 6191 -12518 6234 -12484
rect 6268 -12518 6311 -12484
rect 6191 -12564 6311 -12518
rect 6191 -12598 6234 -12564
rect 6268 -12598 6311 -12564
rect 6191 -12644 6311 -12598
rect 6191 -12678 6234 -12644
rect 6268 -12678 6311 -12644
rect 6191 -12711 6311 -12678
rect 6341 -12484 6461 -12411
rect 6341 -12518 6384 -12484
rect 6418 -12518 6461 -12484
rect 6341 -12564 6461 -12518
rect 6341 -12598 6384 -12564
rect 6418 -12598 6461 -12564
rect 6341 -12644 6461 -12598
rect 6341 -12678 6384 -12644
rect 6418 -12678 6461 -12644
rect 6341 -12711 6461 -12678
rect 6491 -12484 6611 -12411
rect 6491 -12518 6534 -12484
rect 6568 -12518 6611 -12484
rect 6491 -12564 6611 -12518
rect 6491 -12598 6534 -12564
rect 6568 -12598 6611 -12564
rect 6491 -12644 6611 -12598
rect 6491 -12678 6534 -12644
rect 6568 -12678 6611 -12644
rect 6491 -12711 6611 -12678
rect 6671 -12484 6791 -12411
rect 6671 -12518 6714 -12484
rect 6748 -12518 6791 -12484
rect 6671 -12564 6791 -12518
rect 6671 -12598 6714 -12564
rect 6748 -12598 6791 -12564
rect 6671 -12644 6791 -12598
rect 6671 -12678 6714 -12644
rect 6748 -12678 6791 -12644
rect 6671 -12711 6791 -12678
rect 6821 -12711 6941 -12411
rect 6971 -12711 7091 -12411
rect 7121 -12484 7241 -12411
rect 7121 -12518 7164 -12484
rect 7198 -12518 7241 -12484
rect 7121 -12564 7241 -12518
rect 7121 -12598 7164 -12564
rect 7198 -12598 7241 -12564
rect 7121 -12644 7241 -12598
rect 7121 -12678 7164 -12644
rect 7198 -12678 7241 -12644
rect 7121 -12711 7241 -12678
<< pdiff >>
rect 1800 2258 1920 2331
rect 1800 2224 1843 2258
rect 1877 2224 1920 2258
rect 1800 2178 1920 2224
rect 1800 2144 1843 2178
rect 1877 2144 1920 2178
rect 1800 2098 1920 2144
rect 1800 2064 1843 2098
rect 1877 2064 1920 2098
rect 1800 2031 1920 2064
rect 1950 2258 2070 2331
rect 1950 2224 1993 2258
rect 2027 2224 2070 2258
rect 1950 2178 2070 2224
rect 1950 2144 1993 2178
rect 2027 2144 2070 2178
rect 1950 2098 2070 2144
rect 1950 2064 1993 2098
rect 2027 2064 2070 2098
rect 1950 2031 2070 2064
rect 2100 2258 2220 2331
rect 2100 2224 2143 2258
rect 2177 2224 2220 2258
rect 2100 2178 2220 2224
rect 2100 2144 2143 2178
rect 2177 2144 2220 2178
rect 2100 2098 2220 2144
rect 2100 2064 2143 2098
rect 2177 2064 2220 2098
rect 2100 2031 2220 2064
rect 2250 2258 2370 2331
rect 2250 2224 2293 2258
rect 2327 2224 2370 2258
rect 2250 2178 2370 2224
rect 2250 2144 2293 2178
rect 2327 2144 2370 2178
rect 2250 2098 2370 2144
rect 2250 2064 2293 2098
rect 2327 2064 2370 2098
rect 2250 2031 2370 2064
rect 2400 2258 2520 2331
rect 2400 2224 2443 2258
rect 2477 2224 2520 2258
rect 2400 2178 2520 2224
rect 2400 2144 2443 2178
rect 2477 2144 2520 2178
rect 2400 2098 2520 2144
rect 2400 2064 2443 2098
rect 2477 2064 2520 2098
rect 2400 2031 2520 2064
rect 4120 2258 4240 2331
rect 4120 2224 4163 2258
rect 4197 2224 4240 2258
rect 4120 2178 4240 2224
rect 4120 2144 4163 2178
rect 4197 2144 4240 2178
rect 4120 2098 4240 2144
rect 4120 2064 4163 2098
rect 4197 2064 4240 2098
rect 4120 2031 4240 2064
rect 4270 2258 4390 2331
rect 4270 2224 4313 2258
rect 4347 2224 4390 2258
rect 4270 2178 4390 2224
rect 4270 2144 4313 2178
rect 4347 2144 4390 2178
rect 4270 2098 4390 2144
rect 4270 2064 4313 2098
rect 4347 2064 4390 2098
rect 4270 2031 4390 2064
rect 4420 2258 4540 2331
rect 4420 2224 4463 2258
rect 4497 2224 4540 2258
rect 4420 2178 4540 2224
rect 4420 2144 4463 2178
rect 4497 2144 4540 2178
rect 4420 2098 4540 2144
rect 4420 2064 4463 2098
rect 4497 2064 4540 2098
rect 4420 2031 4540 2064
rect 4570 2258 4690 2331
rect 4570 2224 4613 2258
rect 4647 2224 4690 2258
rect 4570 2178 4690 2224
rect 4570 2144 4613 2178
rect 4647 2144 4690 2178
rect 4570 2098 4690 2144
rect 4570 2064 4613 2098
rect 4647 2064 4690 2098
rect 4570 2031 4690 2064
rect 4720 2258 4840 2331
rect 4720 2224 4763 2258
rect 4797 2224 4840 2258
rect 6140 2258 6260 2331
rect 4720 2178 4840 2224
rect 4720 2144 4763 2178
rect 4797 2144 4840 2178
rect 4720 2098 4840 2144
rect 6140 2224 6183 2258
rect 6217 2224 6260 2258
rect 6140 2178 6260 2224
rect 4720 2064 4763 2098
rect 4797 2064 4840 2098
rect 4720 2031 4840 2064
rect 6140 2144 6183 2178
rect 6217 2144 6260 2178
rect 6140 2098 6260 2144
rect 6140 2064 6183 2098
rect 6217 2064 6260 2098
rect 6140 2031 6260 2064
rect 6290 2258 6410 2331
rect 6290 2224 6333 2258
rect 6367 2224 6410 2258
rect 6290 2178 6410 2224
rect 6290 2144 6333 2178
rect 6367 2144 6410 2178
rect 6290 2098 6410 2144
rect 6290 2064 6333 2098
rect 6367 2064 6410 2098
rect 6290 2031 6410 2064
rect 6440 2258 6560 2331
rect 6440 2224 6483 2258
rect 6517 2224 6560 2258
rect 6440 2178 6560 2224
rect 6440 2144 6483 2178
rect 6517 2144 6560 2178
rect 6440 2098 6560 2144
rect 6440 2064 6483 2098
rect 6517 2064 6560 2098
rect 6440 2031 6560 2064
rect 6590 2258 6710 2331
rect 6590 2224 6633 2258
rect 6667 2224 6710 2258
rect 6590 2178 6710 2224
rect 6590 2144 6633 2178
rect 6667 2144 6710 2178
rect 6590 2098 6710 2144
rect 6590 2064 6633 2098
rect 6667 2064 6710 2098
rect 6590 2031 6710 2064
rect 6740 2258 6860 2331
rect 6740 2224 6783 2258
rect 6817 2224 6860 2258
rect 6740 2178 6860 2224
rect 6740 2144 6783 2178
rect 6817 2144 6860 2178
rect 6740 2098 6860 2144
rect 6740 2064 6783 2098
rect 6817 2064 6860 2098
rect 6740 2031 6860 2064
rect 1800 498 1920 531
rect 1800 464 1843 498
rect 1877 464 1920 498
rect 1800 418 1920 464
rect 1800 384 1843 418
rect 1877 384 1920 418
rect 1800 338 1920 384
rect 1800 304 1843 338
rect 1877 304 1920 338
rect 1800 231 1920 304
rect 1950 498 2070 531
rect 1950 464 1993 498
rect 2027 464 2070 498
rect 1950 418 2070 464
rect 1950 384 1993 418
rect 2027 384 2070 418
rect 1950 338 2070 384
rect 1950 304 1993 338
rect 2027 304 2070 338
rect 1950 231 2070 304
rect 2100 498 2220 531
rect 2100 464 2143 498
rect 2177 464 2220 498
rect 2100 418 2220 464
rect 2100 384 2143 418
rect 2177 384 2220 418
rect 2100 338 2220 384
rect 2100 304 2143 338
rect 2177 304 2220 338
rect 2100 231 2220 304
rect 2250 498 2370 531
rect 2250 464 2293 498
rect 2327 464 2370 498
rect 2250 418 2370 464
rect 2250 384 2293 418
rect 2327 384 2370 418
rect 2250 338 2370 384
rect 2250 304 2293 338
rect 2327 304 2370 338
rect 2250 231 2370 304
rect 2400 498 2520 531
rect 2400 464 2443 498
rect 2477 464 2520 498
rect 2400 418 2520 464
rect 2400 384 2443 418
rect 2477 384 2520 418
rect 2400 338 2520 384
rect 2400 304 2443 338
rect 2477 304 2520 338
rect 2400 231 2520 304
rect 4120 498 4240 531
rect 4120 464 4163 498
rect 4197 464 4240 498
rect 4120 418 4240 464
rect 4120 384 4163 418
rect 4197 384 4240 418
rect 4120 338 4240 384
rect 4120 304 4163 338
rect 4197 304 4240 338
rect 4120 231 4240 304
rect 4270 498 4390 531
rect 4270 464 4313 498
rect 4347 464 4390 498
rect 4270 418 4390 464
rect 4270 384 4313 418
rect 4347 384 4390 418
rect 4270 338 4390 384
rect 4270 304 4313 338
rect 4347 304 4390 338
rect 4270 231 4390 304
rect 4420 498 4540 531
rect 4420 464 4463 498
rect 4497 464 4540 498
rect 4420 418 4540 464
rect 4420 384 4463 418
rect 4497 384 4540 418
rect 4420 338 4540 384
rect 4420 304 4463 338
rect 4497 304 4540 338
rect 4420 231 4540 304
rect 4570 498 4690 531
rect 4570 464 4613 498
rect 4647 464 4690 498
rect 4570 418 4690 464
rect 4570 384 4613 418
rect 4647 384 4690 418
rect 4570 338 4690 384
rect 4570 304 4613 338
rect 4647 304 4690 338
rect 4570 231 4690 304
rect 4720 498 4840 531
rect 4720 464 4763 498
rect 4797 464 4840 498
rect 4720 418 4840 464
rect 4720 384 4763 418
rect 4797 384 4840 418
rect 4720 338 4840 384
rect 6140 498 6260 531
rect 6140 464 6183 498
rect 6217 464 6260 498
rect 4720 304 4763 338
rect 4797 304 4840 338
rect 4720 231 4840 304
rect 6140 418 6260 464
rect 6140 384 6183 418
rect 6217 384 6260 418
rect 6140 338 6260 384
rect 6140 304 6183 338
rect 6217 304 6260 338
rect 6140 231 6260 304
rect 6290 498 6410 531
rect 6290 464 6333 498
rect 6367 464 6410 498
rect 6290 418 6410 464
rect 6290 384 6333 418
rect 6367 384 6410 418
rect 6290 338 6410 384
rect 6290 304 6333 338
rect 6367 304 6410 338
rect 6290 231 6410 304
rect 6440 498 6560 531
rect 6440 464 6483 498
rect 6517 464 6560 498
rect 6440 418 6560 464
rect 6440 384 6483 418
rect 6517 384 6560 418
rect 6440 338 6560 384
rect 6440 304 6483 338
rect 6517 304 6560 338
rect 6440 231 6560 304
rect 6590 498 6710 531
rect 6590 464 6633 498
rect 6667 464 6710 498
rect 6590 418 6710 464
rect 6590 384 6633 418
rect 6667 384 6710 418
rect 6590 338 6710 384
rect 6590 304 6633 338
rect 6667 304 6710 338
rect 6590 231 6710 304
rect 6740 498 6860 531
rect 6740 464 6783 498
rect 6817 464 6860 498
rect 6740 418 6860 464
rect 6740 384 6783 418
rect 6817 384 6860 418
rect 6740 338 6860 384
rect 6740 304 6783 338
rect 6817 304 6860 338
rect 6740 231 6860 304
rect 1800 -562 1920 -489
rect 1800 -596 1843 -562
rect 1877 -596 1920 -562
rect 1800 -642 1920 -596
rect 1800 -676 1843 -642
rect 1877 -676 1920 -642
rect 1800 -722 1920 -676
rect 1800 -756 1843 -722
rect 1877 -756 1920 -722
rect 1800 -789 1920 -756
rect 1950 -562 2070 -489
rect 1950 -596 1993 -562
rect 2027 -596 2070 -562
rect 1950 -642 2070 -596
rect 1950 -676 1993 -642
rect 2027 -676 2070 -642
rect 1950 -722 2070 -676
rect 1950 -756 1993 -722
rect 2027 -756 2070 -722
rect 1950 -789 2070 -756
rect 2100 -562 2220 -489
rect 2100 -596 2143 -562
rect 2177 -596 2220 -562
rect 2100 -642 2220 -596
rect 2100 -676 2143 -642
rect 2177 -676 2220 -642
rect 2100 -722 2220 -676
rect 2100 -756 2143 -722
rect 2177 -756 2220 -722
rect 2100 -789 2220 -756
rect 2250 -562 2370 -489
rect 2250 -596 2293 -562
rect 2327 -596 2370 -562
rect 2250 -642 2370 -596
rect 2250 -676 2293 -642
rect 2327 -676 2370 -642
rect 2250 -722 2370 -676
rect 2250 -756 2293 -722
rect 2327 -756 2370 -722
rect 2250 -789 2370 -756
rect 2400 -562 2520 -489
rect 2400 -596 2443 -562
rect 2477 -596 2520 -562
rect 2400 -642 2520 -596
rect 2400 -676 2443 -642
rect 2477 -676 2520 -642
rect 2400 -722 2520 -676
rect 2400 -756 2443 -722
rect 2477 -756 2520 -722
rect 2400 -789 2520 -756
rect 3990 -562 4110 -489
rect 3990 -596 4033 -562
rect 4067 -596 4110 -562
rect 3990 -642 4110 -596
rect 3990 -676 4033 -642
rect 4067 -676 4110 -642
rect 3990 -722 4110 -676
rect 3990 -756 4033 -722
rect 4067 -756 4110 -722
rect 3990 -789 4110 -756
rect 4140 -562 4260 -489
rect 4140 -596 4183 -562
rect 4217 -596 4260 -562
rect 4140 -642 4260 -596
rect 4140 -676 4183 -642
rect 4217 -676 4260 -642
rect 4140 -722 4260 -676
rect 4140 -756 4183 -722
rect 4217 -756 4260 -722
rect 4140 -789 4260 -756
rect 4290 -562 4410 -489
rect 4290 -596 4333 -562
rect 4367 -596 4410 -562
rect 4290 -642 4410 -596
rect 4290 -676 4333 -642
rect 4367 -676 4410 -642
rect 4290 -722 4410 -676
rect 4290 -756 4333 -722
rect 4367 -756 4410 -722
rect 4290 -789 4410 -756
rect 4440 -562 4560 -489
rect 4440 -596 4483 -562
rect 4517 -596 4560 -562
rect 4440 -642 4560 -596
rect 4440 -676 4483 -642
rect 4517 -676 4560 -642
rect 4440 -722 4560 -676
rect 4440 -756 4483 -722
rect 4517 -756 4560 -722
rect 4440 -789 4560 -756
rect 4590 -562 4710 -489
rect 4590 -596 4633 -562
rect 4667 -596 4710 -562
rect 4590 -642 4710 -596
rect 4590 -676 4633 -642
rect 4667 -676 4710 -642
rect 4590 -722 4710 -676
rect 5870 -562 5990 -489
rect 5870 -596 5913 -562
rect 5947 -596 5990 -562
rect 5870 -642 5990 -596
rect 5870 -676 5913 -642
rect 5947 -676 5990 -642
rect 4590 -756 4633 -722
rect 4667 -756 4710 -722
rect 4590 -789 4710 -756
rect 5870 -722 5990 -676
rect 5870 -756 5913 -722
rect 5947 -756 5990 -722
rect 5870 -789 5990 -756
rect 6020 -562 6140 -489
rect 6020 -596 6063 -562
rect 6097 -596 6140 -562
rect 6020 -642 6140 -596
rect 6020 -676 6063 -642
rect 6097 -676 6140 -642
rect 6020 -722 6140 -676
rect 6020 -756 6063 -722
rect 6097 -756 6140 -722
rect 6020 -789 6140 -756
rect 6170 -562 6290 -489
rect 6170 -596 6213 -562
rect 6247 -596 6290 -562
rect 6170 -642 6290 -596
rect 6170 -676 6213 -642
rect 6247 -676 6290 -642
rect 6170 -722 6290 -676
rect 6170 -756 6213 -722
rect 6247 -756 6290 -722
rect 6170 -789 6290 -756
rect 6320 -562 6440 -489
rect 6320 -596 6363 -562
rect 6397 -596 6440 -562
rect 6320 -642 6440 -596
rect 6320 -676 6363 -642
rect 6397 -676 6440 -642
rect 6320 -722 6440 -676
rect 6320 -756 6363 -722
rect 6397 -756 6440 -722
rect 6320 -789 6440 -756
rect 6470 -562 6590 -489
rect 6470 -596 6513 -562
rect 6547 -596 6590 -562
rect 6470 -642 6590 -596
rect 6470 -676 6513 -642
rect 6547 -676 6590 -642
rect 6470 -722 6590 -676
rect 6470 -756 6513 -722
rect 6547 -756 6590 -722
rect 6470 -789 6590 -756
rect 1800 -2322 1920 -2289
rect 1800 -2356 1843 -2322
rect 1877 -2356 1920 -2322
rect 1800 -2402 1920 -2356
rect 1800 -2436 1843 -2402
rect 1877 -2436 1920 -2402
rect 1800 -2482 1920 -2436
rect 1800 -2516 1843 -2482
rect 1877 -2516 1920 -2482
rect 1800 -2589 1920 -2516
rect 1950 -2322 2070 -2289
rect 1950 -2356 1993 -2322
rect 2027 -2356 2070 -2322
rect 1950 -2402 2070 -2356
rect 1950 -2436 1993 -2402
rect 2027 -2436 2070 -2402
rect 1950 -2482 2070 -2436
rect 1950 -2516 1993 -2482
rect 2027 -2516 2070 -2482
rect 1950 -2589 2070 -2516
rect 2100 -2322 2220 -2289
rect 2100 -2356 2143 -2322
rect 2177 -2356 2220 -2322
rect 2100 -2402 2220 -2356
rect 2100 -2436 2143 -2402
rect 2177 -2436 2220 -2402
rect 2100 -2482 2220 -2436
rect 2100 -2516 2143 -2482
rect 2177 -2516 2220 -2482
rect 2100 -2589 2220 -2516
rect 2250 -2322 2370 -2289
rect 2250 -2356 2293 -2322
rect 2327 -2356 2370 -2322
rect 2250 -2402 2370 -2356
rect 2250 -2436 2293 -2402
rect 2327 -2436 2370 -2402
rect 2250 -2482 2370 -2436
rect 2250 -2516 2293 -2482
rect 2327 -2516 2370 -2482
rect 2250 -2589 2370 -2516
rect 2400 -2322 2520 -2289
rect 2400 -2356 2443 -2322
rect 2477 -2356 2520 -2322
rect 2400 -2402 2520 -2356
rect 2400 -2436 2443 -2402
rect 2477 -2436 2520 -2402
rect 2400 -2482 2520 -2436
rect 2400 -2516 2443 -2482
rect 2477 -2516 2520 -2482
rect 2400 -2589 2520 -2516
rect 3990 -2322 4110 -2289
rect 3990 -2356 4033 -2322
rect 4067 -2356 4110 -2322
rect 3990 -2402 4110 -2356
rect 3990 -2436 4033 -2402
rect 4067 -2436 4110 -2402
rect 3990 -2482 4110 -2436
rect 3990 -2516 4033 -2482
rect 4067 -2516 4110 -2482
rect 3990 -2589 4110 -2516
rect 4140 -2322 4260 -2289
rect 4140 -2356 4183 -2322
rect 4217 -2356 4260 -2322
rect 4140 -2402 4260 -2356
rect 4140 -2436 4183 -2402
rect 4217 -2436 4260 -2402
rect 4140 -2482 4260 -2436
rect 4140 -2516 4183 -2482
rect 4217 -2516 4260 -2482
rect 4140 -2589 4260 -2516
rect 4290 -2322 4410 -2289
rect 4290 -2356 4333 -2322
rect 4367 -2356 4410 -2322
rect 4290 -2402 4410 -2356
rect 4290 -2436 4333 -2402
rect 4367 -2436 4410 -2402
rect 4290 -2482 4410 -2436
rect 4290 -2516 4333 -2482
rect 4367 -2516 4410 -2482
rect 4290 -2589 4410 -2516
rect 4440 -2322 4560 -2289
rect 4440 -2356 4483 -2322
rect 4517 -2356 4560 -2322
rect 4440 -2402 4560 -2356
rect 4440 -2436 4483 -2402
rect 4517 -2436 4560 -2402
rect 4440 -2482 4560 -2436
rect 4440 -2516 4483 -2482
rect 4517 -2516 4560 -2482
rect 4440 -2589 4560 -2516
rect 4590 -2322 4710 -2289
rect 4590 -2356 4633 -2322
rect 4667 -2356 4710 -2322
rect 4590 -2402 4710 -2356
rect 5870 -2322 5990 -2289
rect 5870 -2356 5913 -2322
rect 5947 -2356 5990 -2322
rect 4590 -2436 4633 -2402
rect 4667 -2436 4710 -2402
rect 4590 -2482 4710 -2436
rect 4590 -2516 4633 -2482
rect 4667 -2516 4710 -2482
rect 4590 -2589 4710 -2516
rect 5870 -2402 5990 -2356
rect 5870 -2436 5913 -2402
rect 5947 -2436 5990 -2402
rect 5870 -2482 5990 -2436
rect 5870 -2516 5913 -2482
rect 5947 -2516 5990 -2482
rect 5870 -2589 5990 -2516
rect 6020 -2322 6140 -2289
rect 6020 -2356 6063 -2322
rect 6097 -2356 6140 -2322
rect 6020 -2402 6140 -2356
rect 6020 -2436 6063 -2402
rect 6097 -2436 6140 -2402
rect 6020 -2482 6140 -2436
rect 6020 -2516 6063 -2482
rect 6097 -2516 6140 -2482
rect 6020 -2589 6140 -2516
rect 6170 -2322 6290 -2289
rect 6170 -2356 6213 -2322
rect 6247 -2356 6290 -2322
rect 6170 -2402 6290 -2356
rect 6170 -2436 6213 -2402
rect 6247 -2436 6290 -2402
rect 6170 -2482 6290 -2436
rect 6170 -2516 6213 -2482
rect 6247 -2516 6290 -2482
rect 6170 -2589 6290 -2516
rect 6320 -2322 6440 -2289
rect 6320 -2356 6363 -2322
rect 6397 -2356 6440 -2322
rect 6320 -2402 6440 -2356
rect 6320 -2436 6363 -2402
rect 6397 -2436 6440 -2402
rect 6320 -2482 6440 -2436
rect 6320 -2516 6363 -2482
rect 6397 -2516 6440 -2482
rect 6320 -2589 6440 -2516
rect 6470 -2322 6590 -2289
rect 6470 -2356 6513 -2322
rect 6547 -2356 6590 -2322
rect 6470 -2402 6590 -2356
rect 6470 -2436 6513 -2402
rect 6547 -2436 6590 -2402
rect 6470 -2482 6590 -2436
rect 6470 -2516 6513 -2482
rect 6547 -2516 6590 -2482
rect 6470 -2589 6590 -2516
rect 1801 -3382 1921 -3309
rect 1801 -3416 1844 -3382
rect 1878 -3416 1921 -3382
rect 1801 -3462 1921 -3416
rect 1801 -3496 1844 -3462
rect 1878 -3496 1921 -3462
rect 1801 -3542 1921 -3496
rect 1801 -3576 1844 -3542
rect 1878 -3576 1921 -3542
rect 1801 -3609 1921 -3576
rect 1951 -3382 2071 -3309
rect 1951 -3416 1994 -3382
rect 2028 -3416 2071 -3382
rect 1951 -3462 2071 -3416
rect 1951 -3496 1994 -3462
rect 2028 -3496 2071 -3462
rect 1951 -3542 2071 -3496
rect 1951 -3576 1994 -3542
rect 2028 -3576 2071 -3542
rect 1951 -3609 2071 -3576
rect 2101 -3382 2221 -3309
rect 2101 -3416 2144 -3382
rect 2178 -3416 2221 -3382
rect 2101 -3462 2221 -3416
rect 2101 -3496 2144 -3462
rect 2178 -3496 2221 -3462
rect 2101 -3542 2221 -3496
rect 2101 -3576 2144 -3542
rect 2178 -3576 2221 -3542
rect 2101 -3609 2221 -3576
rect 2251 -3382 2371 -3309
rect 2251 -3416 2294 -3382
rect 2328 -3416 2371 -3382
rect 2251 -3462 2371 -3416
rect 2251 -3496 2294 -3462
rect 2328 -3496 2371 -3462
rect 2251 -3542 2371 -3496
rect 2251 -3576 2294 -3542
rect 2328 -3576 2371 -3542
rect 2251 -3609 2371 -3576
rect 2401 -3382 2521 -3309
rect 2401 -3416 2444 -3382
rect 2478 -3416 2521 -3382
rect 2401 -3462 2521 -3416
rect 2401 -3496 2444 -3462
rect 2478 -3496 2521 -3462
rect 2401 -3542 2521 -3496
rect 2401 -3576 2444 -3542
rect 2478 -3576 2521 -3542
rect 2401 -3609 2521 -3576
rect 3851 -3382 3971 -3309
rect 3851 -3416 3894 -3382
rect 3928 -3416 3971 -3382
rect 3851 -3462 3971 -3416
rect 3851 -3496 3894 -3462
rect 3928 -3496 3971 -3462
rect 3851 -3542 3971 -3496
rect 3851 -3576 3894 -3542
rect 3928 -3576 3971 -3542
rect 3851 -3609 3971 -3576
rect 4001 -3382 4121 -3309
rect 4001 -3416 4044 -3382
rect 4078 -3416 4121 -3382
rect 4001 -3462 4121 -3416
rect 4001 -3496 4044 -3462
rect 4078 -3496 4121 -3462
rect 4001 -3542 4121 -3496
rect 4001 -3576 4044 -3542
rect 4078 -3576 4121 -3542
rect 4001 -3609 4121 -3576
rect 4151 -3382 4271 -3309
rect 4151 -3416 4194 -3382
rect 4228 -3416 4271 -3382
rect 4151 -3462 4271 -3416
rect 4151 -3496 4194 -3462
rect 4228 -3496 4271 -3462
rect 4151 -3542 4271 -3496
rect 4151 -3576 4194 -3542
rect 4228 -3576 4271 -3542
rect 4151 -3609 4271 -3576
rect 4301 -3382 4421 -3309
rect 4301 -3416 4344 -3382
rect 4378 -3416 4421 -3382
rect 4301 -3462 4421 -3416
rect 4301 -3496 4344 -3462
rect 4378 -3496 4421 -3462
rect 4301 -3542 4421 -3496
rect 4301 -3576 4344 -3542
rect 4378 -3576 4421 -3542
rect 4301 -3609 4421 -3576
rect 4451 -3382 4571 -3309
rect 4451 -3416 4494 -3382
rect 4528 -3416 4571 -3382
rect 4451 -3462 4571 -3416
rect 4451 -3496 4494 -3462
rect 4528 -3496 4571 -3462
rect 4451 -3542 4571 -3496
rect 4451 -3576 4494 -3542
rect 4528 -3576 4571 -3542
rect 4451 -3609 4571 -3576
rect 5891 -3383 6011 -3310
rect 5891 -3417 5934 -3383
rect 5968 -3417 6011 -3383
rect 5891 -3463 6011 -3417
rect 5891 -3497 5934 -3463
rect 5968 -3497 6011 -3463
rect 5891 -3543 6011 -3497
rect 5891 -3577 5934 -3543
rect 5968 -3577 6011 -3543
rect 5891 -3610 6011 -3577
rect 6041 -3383 6161 -3310
rect 6041 -3417 6084 -3383
rect 6118 -3417 6161 -3383
rect 6041 -3463 6161 -3417
rect 6041 -3497 6084 -3463
rect 6118 -3497 6161 -3463
rect 6041 -3543 6161 -3497
rect 6041 -3577 6084 -3543
rect 6118 -3577 6161 -3543
rect 6041 -3610 6161 -3577
rect 6191 -3383 6311 -3310
rect 6191 -3417 6234 -3383
rect 6268 -3417 6311 -3383
rect 6191 -3463 6311 -3417
rect 6191 -3497 6234 -3463
rect 6268 -3497 6311 -3463
rect 6191 -3543 6311 -3497
rect 6191 -3577 6234 -3543
rect 6268 -3577 6311 -3543
rect 6191 -3610 6311 -3577
rect 6341 -3383 6461 -3310
rect 6341 -3417 6384 -3383
rect 6418 -3417 6461 -3383
rect 6341 -3463 6461 -3417
rect 6341 -3497 6384 -3463
rect 6418 -3497 6461 -3463
rect 6341 -3543 6461 -3497
rect 6341 -3577 6384 -3543
rect 6418 -3577 6461 -3543
rect 6341 -3610 6461 -3577
rect 6491 -3383 6611 -3310
rect 6491 -3417 6534 -3383
rect 6568 -3417 6611 -3383
rect 6491 -3463 6611 -3417
rect 6491 -3497 6534 -3463
rect 6568 -3497 6611 -3463
rect 6491 -3543 6611 -3497
rect 6491 -3577 6534 -3543
rect 6568 -3577 6611 -3543
rect 6491 -3610 6611 -3577
rect 4051 -5223 4171 -5190
rect 4051 -5257 4094 -5223
rect 4128 -5257 4171 -5223
rect 4051 -5303 4171 -5257
rect 4051 -5337 4094 -5303
rect 4128 -5337 4171 -5303
rect 4051 -5383 4171 -5337
rect 4051 -5417 4094 -5383
rect 4128 -5417 4171 -5383
rect 4051 -5490 4171 -5417
rect 4201 -5223 4321 -5190
rect 4201 -5257 4244 -5223
rect 4278 -5257 4321 -5223
rect 4201 -5303 4321 -5257
rect 4201 -5337 4244 -5303
rect 4278 -5337 4321 -5303
rect 4201 -5383 4321 -5337
rect 4201 -5417 4244 -5383
rect 4278 -5417 4321 -5383
rect 4201 -5490 4321 -5417
rect 4351 -5223 4471 -5190
rect 4351 -5257 4394 -5223
rect 4428 -5257 4471 -5223
rect 4351 -5303 4471 -5257
rect 4351 -5337 4394 -5303
rect 4428 -5337 4471 -5303
rect 4351 -5383 4471 -5337
rect 4351 -5417 4394 -5383
rect 4428 -5417 4471 -5383
rect 4351 -5490 4471 -5417
rect 4501 -5223 4621 -5190
rect 4501 -5257 4544 -5223
rect 4578 -5257 4621 -5223
rect 4501 -5303 4621 -5257
rect 4501 -5337 4544 -5303
rect 4578 -5337 4621 -5303
rect 4501 -5383 4621 -5337
rect 4501 -5417 4544 -5383
rect 4578 -5417 4621 -5383
rect 4501 -5490 4621 -5417
rect 4651 -5223 4771 -5190
rect 4651 -5257 4694 -5223
rect 4728 -5257 4771 -5223
rect 4651 -5303 4771 -5257
rect 4651 -5337 4694 -5303
rect 4728 -5337 4771 -5303
rect 4651 -5383 4771 -5337
rect 4651 -5417 4694 -5383
rect 4728 -5417 4771 -5383
rect 4651 -5490 4771 -5417
rect 6110 -5223 6230 -5190
rect 6110 -5257 6153 -5223
rect 6187 -5257 6230 -5223
rect 6110 -5303 6230 -5257
rect 6110 -5337 6153 -5303
rect 6187 -5337 6230 -5303
rect 6110 -5383 6230 -5337
rect 6110 -5417 6153 -5383
rect 6187 -5417 6230 -5383
rect 1840 -5542 1960 -5509
rect 1840 -5576 1883 -5542
rect 1917 -5576 1960 -5542
rect 1840 -5622 1960 -5576
rect 1840 -5656 1883 -5622
rect 1917 -5656 1960 -5622
rect 1840 -5702 1960 -5656
rect 1840 -5736 1883 -5702
rect 1917 -5736 1960 -5702
rect 1840 -5809 1960 -5736
rect 1990 -5542 2110 -5509
rect 1990 -5576 2033 -5542
rect 2067 -5576 2110 -5542
rect 1990 -5622 2110 -5576
rect 1990 -5656 2033 -5622
rect 2067 -5656 2110 -5622
rect 1990 -5702 2110 -5656
rect 1990 -5736 2033 -5702
rect 2067 -5736 2110 -5702
rect 1990 -5809 2110 -5736
rect 2140 -5542 2260 -5509
rect 2140 -5576 2183 -5542
rect 2217 -5576 2260 -5542
rect 2140 -5622 2260 -5576
rect 2140 -5656 2183 -5622
rect 2217 -5656 2260 -5622
rect 2140 -5702 2260 -5656
rect 2140 -5736 2183 -5702
rect 2217 -5736 2260 -5702
rect 2140 -5809 2260 -5736
rect 2290 -5542 2410 -5509
rect 2290 -5576 2333 -5542
rect 2367 -5576 2410 -5542
rect 2290 -5622 2410 -5576
rect 2290 -5656 2333 -5622
rect 2367 -5656 2410 -5622
rect 2290 -5702 2410 -5656
rect 2290 -5736 2333 -5702
rect 2367 -5736 2410 -5702
rect 2290 -5809 2410 -5736
rect 2440 -5542 2560 -5509
rect 2440 -5576 2483 -5542
rect 2517 -5576 2560 -5542
rect 6110 -5490 6230 -5417
rect 6260 -5223 6380 -5190
rect 6260 -5257 6303 -5223
rect 6337 -5257 6380 -5223
rect 6260 -5303 6380 -5257
rect 6260 -5337 6303 -5303
rect 6337 -5337 6380 -5303
rect 6260 -5383 6380 -5337
rect 6260 -5417 6303 -5383
rect 6337 -5417 6380 -5383
rect 6260 -5490 6380 -5417
rect 6410 -5223 6530 -5190
rect 6410 -5257 6453 -5223
rect 6487 -5257 6530 -5223
rect 6410 -5303 6530 -5257
rect 6410 -5337 6453 -5303
rect 6487 -5337 6530 -5303
rect 6410 -5383 6530 -5337
rect 6410 -5417 6453 -5383
rect 6487 -5417 6530 -5383
rect 6410 -5490 6530 -5417
rect 6560 -5223 6680 -5190
rect 6560 -5257 6603 -5223
rect 6637 -5257 6680 -5223
rect 6560 -5303 6680 -5257
rect 6560 -5337 6603 -5303
rect 6637 -5337 6680 -5303
rect 6560 -5383 6680 -5337
rect 6560 -5417 6603 -5383
rect 6637 -5417 6680 -5383
rect 6560 -5490 6680 -5417
rect 6710 -5223 6830 -5190
rect 6710 -5257 6753 -5223
rect 6787 -5257 6830 -5223
rect 6710 -5303 6830 -5257
rect 6710 -5337 6753 -5303
rect 6787 -5337 6830 -5303
rect 6710 -5383 6830 -5337
rect 6710 -5417 6753 -5383
rect 6787 -5417 6830 -5383
rect 6710 -5490 6830 -5417
rect 2440 -5622 2560 -5576
rect 2440 -5656 2483 -5622
rect 2517 -5656 2560 -5622
rect 2440 -5702 2560 -5656
rect 2440 -5736 2483 -5702
rect 2517 -5736 2560 -5702
rect 2440 -5809 2560 -5736
rect 1840 -6283 1960 -6210
rect 1840 -6317 1883 -6283
rect 1917 -6317 1960 -6283
rect 1840 -6363 1960 -6317
rect 1840 -6397 1883 -6363
rect 1917 -6397 1960 -6363
rect 1840 -6443 1960 -6397
rect 1840 -6477 1883 -6443
rect 1917 -6477 1960 -6443
rect 1840 -6510 1960 -6477
rect 1990 -6283 2110 -6210
rect 1990 -6317 2033 -6283
rect 2067 -6317 2110 -6283
rect 1990 -6363 2110 -6317
rect 1990 -6397 2033 -6363
rect 2067 -6397 2110 -6363
rect 1990 -6443 2110 -6397
rect 1990 -6477 2033 -6443
rect 2067 -6477 2110 -6443
rect 1990 -6510 2110 -6477
rect 2140 -6283 2260 -6210
rect 2140 -6317 2183 -6283
rect 2217 -6317 2260 -6283
rect 2140 -6363 2260 -6317
rect 2140 -6397 2183 -6363
rect 2217 -6397 2260 -6363
rect 2140 -6443 2260 -6397
rect 2140 -6477 2183 -6443
rect 2217 -6477 2260 -6443
rect 2140 -6510 2260 -6477
rect 2290 -6283 2410 -6210
rect 2290 -6317 2333 -6283
rect 2367 -6317 2410 -6283
rect 2290 -6363 2410 -6317
rect 2290 -6397 2333 -6363
rect 2367 -6397 2410 -6363
rect 2290 -6443 2410 -6397
rect 2290 -6477 2333 -6443
rect 2367 -6477 2410 -6443
rect 2290 -6510 2410 -6477
rect 2440 -6283 2560 -6210
rect 2440 -6317 2483 -6283
rect 2517 -6317 2560 -6283
rect 2440 -6363 2560 -6317
rect 2440 -6397 2483 -6363
rect 2517 -6397 2560 -6363
rect 2440 -6443 2560 -6397
rect 2440 -6477 2483 -6443
rect 2517 -6477 2560 -6443
rect 2440 -6510 2560 -6477
rect 4050 -6283 4170 -6210
rect 4050 -6317 4093 -6283
rect 4127 -6317 4170 -6283
rect 4050 -6363 4170 -6317
rect 4050 -6397 4093 -6363
rect 4127 -6397 4170 -6363
rect 4050 -6443 4170 -6397
rect 4050 -6477 4093 -6443
rect 4127 -6477 4170 -6443
rect 4050 -6510 4170 -6477
rect 4200 -6283 4320 -6210
rect 4200 -6317 4243 -6283
rect 4277 -6317 4320 -6283
rect 4200 -6363 4320 -6317
rect 4200 -6397 4243 -6363
rect 4277 -6397 4320 -6363
rect 4200 -6443 4320 -6397
rect 4200 -6477 4243 -6443
rect 4277 -6477 4320 -6443
rect 4200 -6510 4320 -6477
rect 4350 -6283 4470 -6210
rect 4350 -6317 4393 -6283
rect 4427 -6317 4470 -6283
rect 4350 -6363 4470 -6317
rect 4350 -6397 4393 -6363
rect 4427 -6397 4470 -6363
rect 4350 -6443 4470 -6397
rect 4350 -6477 4393 -6443
rect 4427 -6477 4470 -6443
rect 4350 -6510 4470 -6477
rect 4500 -6283 4620 -6210
rect 4500 -6317 4543 -6283
rect 4577 -6317 4620 -6283
rect 4500 -6363 4620 -6317
rect 4500 -6397 4543 -6363
rect 4577 -6397 4620 -6363
rect 4500 -6443 4620 -6397
rect 4500 -6477 4543 -6443
rect 4577 -6477 4620 -6443
rect 4500 -6510 4620 -6477
rect 4650 -6283 4770 -6210
rect 4650 -6317 4693 -6283
rect 4727 -6317 4770 -6283
rect 4650 -6363 4770 -6317
rect 4650 -6397 4693 -6363
rect 4727 -6397 4770 -6363
rect 4650 -6443 4770 -6397
rect 5929 -6283 6049 -6210
rect 5929 -6317 5972 -6283
rect 6006 -6317 6049 -6283
rect 5929 -6363 6049 -6317
rect 5929 -6397 5972 -6363
rect 6006 -6397 6049 -6363
rect 4650 -6477 4693 -6443
rect 4727 -6477 4770 -6443
rect 4650 -6510 4770 -6477
rect 5929 -6443 6049 -6397
rect 5929 -6477 5972 -6443
rect 6006 -6477 6049 -6443
rect 5929 -6510 6049 -6477
rect 6079 -6283 6199 -6210
rect 6079 -6317 6122 -6283
rect 6156 -6317 6199 -6283
rect 6079 -6363 6199 -6317
rect 6079 -6397 6122 -6363
rect 6156 -6397 6199 -6363
rect 6079 -6443 6199 -6397
rect 6079 -6477 6122 -6443
rect 6156 -6477 6199 -6443
rect 6079 -6510 6199 -6477
rect 6229 -6283 6349 -6210
rect 6229 -6317 6272 -6283
rect 6306 -6317 6349 -6283
rect 6229 -6363 6349 -6317
rect 6229 -6397 6272 -6363
rect 6306 -6397 6349 -6363
rect 6229 -6443 6349 -6397
rect 6229 -6477 6272 -6443
rect 6306 -6477 6349 -6443
rect 6229 -6510 6349 -6477
rect 6379 -6283 6499 -6210
rect 6379 -6317 6422 -6283
rect 6456 -6317 6499 -6283
rect 6379 -6363 6499 -6317
rect 6379 -6397 6422 -6363
rect 6456 -6397 6499 -6363
rect 6379 -6443 6499 -6397
rect 6379 -6477 6422 -6443
rect 6456 -6477 6499 -6443
rect 6379 -6510 6499 -6477
rect 6529 -6283 6649 -6210
rect 6529 -6317 6572 -6283
rect 6606 -6317 6649 -6283
rect 6529 -6363 6649 -6317
rect 6529 -6397 6572 -6363
rect 6606 -6397 6649 -6363
rect 6529 -6443 6649 -6397
rect 6529 -6477 6572 -6443
rect 6606 -6477 6649 -6443
rect 6529 -6510 6649 -6477
rect 1840 -8043 1960 -8010
rect 1840 -8077 1883 -8043
rect 1917 -8077 1960 -8043
rect 1840 -8123 1960 -8077
rect 1840 -8157 1883 -8123
rect 1917 -8157 1960 -8123
rect 1840 -8203 1960 -8157
rect 1840 -8237 1883 -8203
rect 1917 -8237 1960 -8203
rect 1840 -8310 1960 -8237
rect 1990 -8043 2110 -8010
rect 1990 -8077 2033 -8043
rect 2067 -8077 2110 -8043
rect 1990 -8123 2110 -8077
rect 1990 -8157 2033 -8123
rect 2067 -8157 2110 -8123
rect 1990 -8203 2110 -8157
rect 1990 -8237 2033 -8203
rect 2067 -8237 2110 -8203
rect 1990 -8310 2110 -8237
rect 2140 -8043 2260 -8010
rect 2140 -8077 2183 -8043
rect 2217 -8077 2260 -8043
rect 2140 -8123 2260 -8077
rect 2140 -8157 2183 -8123
rect 2217 -8157 2260 -8123
rect 2140 -8203 2260 -8157
rect 2140 -8237 2183 -8203
rect 2217 -8237 2260 -8203
rect 2140 -8310 2260 -8237
rect 2290 -8043 2410 -8010
rect 2290 -8077 2333 -8043
rect 2367 -8077 2410 -8043
rect 2290 -8123 2410 -8077
rect 2290 -8157 2333 -8123
rect 2367 -8157 2410 -8123
rect 2290 -8203 2410 -8157
rect 2290 -8237 2333 -8203
rect 2367 -8237 2410 -8203
rect 2290 -8310 2410 -8237
rect 2440 -8043 2560 -8010
rect 2440 -8077 2483 -8043
rect 2517 -8077 2560 -8043
rect 2440 -8123 2560 -8077
rect 2440 -8157 2483 -8123
rect 2517 -8157 2560 -8123
rect 2440 -8203 2560 -8157
rect 2440 -8237 2483 -8203
rect 2517 -8237 2560 -8203
rect 2440 -8310 2560 -8237
rect 4050 -8043 4170 -8010
rect 4050 -8077 4093 -8043
rect 4127 -8077 4170 -8043
rect 4050 -8123 4170 -8077
rect 4050 -8157 4093 -8123
rect 4127 -8157 4170 -8123
rect 4050 -8203 4170 -8157
rect 4050 -8237 4093 -8203
rect 4127 -8237 4170 -8203
rect 4050 -8310 4170 -8237
rect 4200 -8043 4320 -8010
rect 4200 -8077 4243 -8043
rect 4277 -8077 4320 -8043
rect 4200 -8123 4320 -8077
rect 4200 -8157 4243 -8123
rect 4277 -8157 4320 -8123
rect 4200 -8203 4320 -8157
rect 4200 -8237 4243 -8203
rect 4277 -8237 4320 -8203
rect 4200 -8310 4320 -8237
rect 4350 -8043 4470 -8010
rect 4350 -8077 4393 -8043
rect 4427 -8077 4470 -8043
rect 4350 -8123 4470 -8077
rect 4350 -8157 4393 -8123
rect 4427 -8157 4470 -8123
rect 4350 -8203 4470 -8157
rect 4350 -8237 4393 -8203
rect 4427 -8237 4470 -8203
rect 4350 -8310 4470 -8237
rect 4500 -8043 4620 -8010
rect 4500 -8077 4543 -8043
rect 4577 -8077 4620 -8043
rect 4500 -8123 4620 -8077
rect 4500 -8157 4543 -8123
rect 4577 -8157 4620 -8123
rect 4500 -8203 4620 -8157
rect 4500 -8237 4543 -8203
rect 4577 -8237 4620 -8203
rect 4500 -8310 4620 -8237
rect 4650 -8043 4770 -8010
rect 4650 -8077 4693 -8043
rect 4727 -8077 4770 -8043
rect 4650 -8123 4770 -8077
rect 5929 -8043 6049 -8010
rect 5929 -8077 5972 -8043
rect 6006 -8077 6049 -8043
rect 4650 -8157 4693 -8123
rect 4727 -8157 4770 -8123
rect 4650 -8203 4770 -8157
rect 4650 -8237 4693 -8203
rect 4727 -8237 4770 -8203
rect 4650 -8310 4770 -8237
rect 5929 -8123 6049 -8077
rect 5929 -8157 5972 -8123
rect 6006 -8157 6049 -8123
rect 5929 -8203 6049 -8157
rect 5929 -8237 5972 -8203
rect 6006 -8237 6049 -8203
rect 5929 -8310 6049 -8237
rect 6079 -8043 6199 -8010
rect 6079 -8077 6122 -8043
rect 6156 -8077 6199 -8043
rect 6079 -8123 6199 -8077
rect 6079 -8157 6122 -8123
rect 6156 -8157 6199 -8123
rect 6079 -8203 6199 -8157
rect 6079 -8237 6122 -8203
rect 6156 -8237 6199 -8203
rect 6079 -8310 6199 -8237
rect 6229 -8043 6349 -8010
rect 6229 -8077 6272 -8043
rect 6306 -8077 6349 -8043
rect 6229 -8123 6349 -8077
rect 6229 -8157 6272 -8123
rect 6306 -8157 6349 -8123
rect 6229 -8203 6349 -8157
rect 6229 -8237 6272 -8203
rect 6306 -8237 6349 -8203
rect 6229 -8310 6349 -8237
rect 6379 -8043 6499 -8010
rect 6379 -8077 6422 -8043
rect 6456 -8077 6499 -8043
rect 6379 -8123 6499 -8077
rect 6379 -8157 6422 -8123
rect 6456 -8157 6499 -8123
rect 6379 -8203 6499 -8157
rect 6379 -8237 6422 -8203
rect 6456 -8237 6499 -8203
rect 6379 -8310 6499 -8237
rect 6529 -8043 6649 -8010
rect 6529 -8077 6572 -8043
rect 6606 -8077 6649 -8043
rect 6529 -8123 6649 -8077
rect 6529 -8157 6572 -8123
rect 6606 -8157 6649 -8123
rect 6529 -8203 6649 -8157
rect 6529 -8237 6572 -8203
rect 6606 -8237 6649 -8203
rect 6529 -8310 6649 -8237
rect 1800 -9103 1920 -9030
rect 1800 -9137 1843 -9103
rect 1877 -9137 1920 -9103
rect 1800 -9183 1920 -9137
rect 1800 -9217 1843 -9183
rect 1877 -9217 1920 -9183
rect 1800 -9263 1920 -9217
rect 1800 -9297 1843 -9263
rect 1877 -9297 1920 -9263
rect 1800 -9330 1920 -9297
rect 1950 -9103 2070 -9030
rect 1950 -9137 1993 -9103
rect 2027 -9137 2070 -9103
rect 1950 -9183 2070 -9137
rect 1950 -9217 1993 -9183
rect 2027 -9217 2070 -9183
rect 1950 -9263 2070 -9217
rect 1950 -9297 1993 -9263
rect 2027 -9297 2070 -9263
rect 1950 -9330 2070 -9297
rect 2100 -9103 2220 -9030
rect 2100 -9137 2143 -9103
rect 2177 -9137 2220 -9103
rect 2100 -9183 2220 -9137
rect 2100 -9217 2143 -9183
rect 2177 -9217 2220 -9183
rect 2100 -9263 2220 -9217
rect 2100 -9297 2143 -9263
rect 2177 -9297 2220 -9263
rect 2100 -9330 2220 -9297
rect 2250 -9103 2370 -9030
rect 2250 -9137 2293 -9103
rect 2327 -9137 2370 -9103
rect 2250 -9183 2370 -9137
rect 2250 -9217 2293 -9183
rect 2327 -9217 2370 -9183
rect 2250 -9263 2370 -9217
rect 2250 -9297 2293 -9263
rect 2327 -9297 2370 -9263
rect 2250 -9330 2370 -9297
rect 2400 -9103 2520 -9030
rect 2400 -9137 2443 -9103
rect 2477 -9137 2520 -9103
rect 2400 -9183 2520 -9137
rect 2400 -9217 2443 -9183
rect 2477 -9217 2520 -9183
rect 2400 -9263 2520 -9217
rect 2400 -9297 2443 -9263
rect 2477 -9297 2520 -9263
rect 2400 -9330 2520 -9297
rect 3990 -9103 4110 -9030
rect 3990 -9137 4033 -9103
rect 4067 -9137 4110 -9103
rect 3990 -9183 4110 -9137
rect 3990 -9217 4033 -9183
rect 4067 -9217 4110 -9183
rect 3990 -9263 4110 -9217
rect 3990 -9297 4033 -9263
rect 4067 -9297 4110 -9263
rect 3990 -9330 4110 -9297
rect 4140 -9103 4260 -9030
rect 4140 -9137 4183 -9103
rect 4217 -9137 4260 -9103
rect 4140 -9183 4260 -9137
rect 4140 -9217 4183 -9183
rect 4217 -9217 4260 -9183
rect 4140 -9263 4260 -9217
rect 4140 -9297 4183 -9263
rect 4217 -9297 4260 -9263
rect 4140 -9330 4260 -9297
rect 4290 -9103 4410 -9030
rect 4290 -9137 4333 -9103
rect 4367 -9137 4410 -9103
rect 4290 -9183 4410 -9137
rect 4290 -9217 4333 -9183
rect 4367 -9217 4410 -9183
rect 4290 -9263 4410 -9217
rect 4290 -9297 4333 -9263
rect 4367 -9297 4410 -9263
rect 4290 -9330 4410 -9297
rect 4440 -9103 4560 -9030
rect 4440 -9137 4483 -9103
rect 4517 -9137 4560 -9103
rect 4440 -9183 4560 -9137
rect 4440 -9217 4483 -9183
rect 4517 -9217 4560 -9183
rect 4440 -9263 4560 -9217
rect 4440 -9297 4483 -9263
rect 4517 -9297 4560 -9263
rect 4440 -9330 4560 -9297
rect 4590 -9103 4710 -9030
rect 4590 -9137 4633 -9103
rect 4667 -9137 4710 -9103
rect 4590 -9183 4710 -9137
rect 4590 -9217 4633 -9183
rect 4667 -9217 4710 -9183
rect 4590 -9263 4710 -9217
rect 5870 -9103 5990 -9030
rect 5870 -9137 5913 -9103
rect 5947 -9137 5990 -9103
rect 5870 -9183 5990 -9137
rect 5870 -9217 5913 -9183
rect 5947 -9217 5990 -9183
rect 4590 -9297 4633 -9263
rect 4667 -9297 4710 -9263
rect 4590 -9330 4710 -9297
rect 5870 -9263 5990 -9217
rect 5870 -9297 5913 -9263
rect 5947 -9297 5990 -9263
rect 5870 -9330 5990 -9297
rect 6020 -9103 6140 -9030
rect 6020 -9137 6063 -9103
rect 6097 -9137 6140 -9103
rect 6020 -9183 6140 -9137
rect 6020 -9217 6063 -9183
rect 6097 -9217 6140 -9183
rect 6020 -9263 6140 -9217
rect 6020 -9297 6063 -9263
rect 6097 -9297 6140 -9263
rect 6020 -9330 6140 -9297
rect 6170 -9103 6290 -9030
rect 6170 -9137 6213 -9103
rect 6247 -9137 6290 -9103
rect 6170 -9183 6290 -9137
rect 6170 -9217 6213 -9183
rect 6247 -9217 6290 -9183
rect 6170 -9263 6290 -9217
rect 6170 -9297 6213 -9263
rect 6247 -9297 6290 -9263
rect 6170 -9330 6290 -9297
rect 6320 -9103 6440 -9030
rect 6320 -9137 6363 -9103
rect 6397 -9137 6440 -9103
rect 6320 -9183 6440 -9137
rect 6320 -9217 6363 -9183
rect 6397 -9217 6440 -9183
rect 6320 -9263 6440 -9217
rect 6320 -9297 6363 -9263
rect 6397 -9297 6440 -9263
rect 6320 -9330 6440 -9297
rect 6470 -9103 6590 -9030
rect 6470 -9137 6513 -9103
rect 6547 -9137 6590 -9103
rect 6470 -9183 6590 -9137
rect 6470 -9217 6513 -9183
rect 6547 -9217 6590 -9183
rect 6470 -9263 6590 -9217
rect 6470 -9297 6513 -9263
rect 6547 -9297 6590 -9263
rect 6470 -9330 6590 -9297
rect 1800 -10863 1920 -10830
rect 1800 -10897 1843 -10863
rect 1877 -10897 1920 -10863
rect 1800 -10943 1920 -10897
rect 1800 -10977 1843 -10943
rect 1877 -10977 1920 -10943
rect 1800 -11023 1920 -10977
rect 1800 -11057 1843 -11023
rect 1877 -11057 1920 -11023
rect 1800 -11130 1920 -11057
rect 1950 -10863 2070 -10830
rect 1950 -10897 1993 -10863
rect 2027 -10897 2070 -10863
rect 1950 -10943 2070 -10897
rect 1950 -10977 1993 -10943
rect 2027 -10977 2070 -10943
rect 1950 -11023 2070 -10977
rect 1950 -11057 1993 -11023
rect 2027 -11057 2070 -11023
rect 1950 -11130 2070 -11057
rect 2100 -10863 2220 -10830
rect 2100 -10897 2143 -10863
rect 2177 -10897 2220 -10863
rect 2100 -10943 2220 -10897
rect 2100 -10977 2143 -10943
rect 2177 -10977 2220 -10943
rect 2100 -11023 2220 -10977
rect 2100 -11057 2143 -11023
rect 2177 -11057 2220 -11023
rect 2100 -11130 2220 -11057
rect 2250 -10863 2370 -10830
rect 2250 -10897 2293 -10863
rect 2327 -10897 2370 -10863
rect 2250 -10943 2370 -10897
rect 2250 -10977 2293 -10943
rect 2327 -10977 2370 -10943
rect 2250 -11023 2370 -10977
rect 2250 -11057 2293 -11023
rect 2327 -11057 2370 -11023
rect 2250 -11130 2370 -11057
rect 2400 -10863 2520 -10830
rect 2400 -10897 2443 -10863
rect 2477 -10897 2520 -10863
rect 2400 -10943 2520 -10897
rect 2400 -10977 2443 -10943
rect 2477 -10977 2520 -10943
rect 2400 -11023 2520 -10977
rect 2400 -11057 2443 -11023
rect 2477 -11057 2520 -11023
rect 2400 -11130 2520 -11057
rect 3990 -10863 4110 -10830
rect 3990 -10897 4033 -10863
rect 4067 -10897 4110 -10863
rect 3990 -10943 4110 -10897
rect 3990 -10977 4033 -10943
rect 4067 -10977 4110 -10943
rect 3990 -11023 4110 -10977
rect 3990 -11057 4033 -11023
rect 4067 -11057 4110 -11023
rect 3990 -11130 4110 -11057
rect 4140 -10863 4260 -10830
rect 4140 -10897 4183 -10863
rect 4217 -10897 4260 -10863
rect 4140 -10943 4260 -10897
rect 4140 -10977 4183 -10943
rect 4217 -10977 4260 -10943
rect 4140 -11023 4260 -10977
rect 4140 -11057 4183 -11023
rect 4217 -11057 4260 -11023
rect 4140 -11130 4260 -11057
rect 4290 -10863 4410 -10830
rect 4290 -10897 4333 -10863
rect 4367 -10897 4410 -10863
rect 4290 -10943 4410 -10897
rect 4290 -10977 4333 -10943
rect 4367 -10977 4410 -10943
rect 4290 -11023 4410 -10977
rect 4290 -11057 4333 -11023
rect 4367 -11057 4410 -11023
rect 4290 -11130 4410 -11057
rect 4440 -10863 4560 -10830
rect 4440 -10897 4483 -10863
rect 4517 -10897 4560 -10863
rect 4440 -10943 4560 -10897
rect 4440 -10977 4483 -10943
rect 4517 -10977 4560 -10943
rect 4440 -11023 4560 -10977
rect 4440 -11057 4483 -11023
rect 4517 -11057 4560 -11023
rect 4440 -11130 4560 -11057
rect 4590 -10863 4710 -10830
rect 4590 -10897 4633 -10863
rect 4667 -10897 4710 -10863
rect 4590 -10943 4710 -10897
rect 5870 -10863 5990 -10830
rect 5870 -10897 5913 -10863
rect 5947 -10897 5990 -10863
rect 4590 -10977 4633 -10943
rect 4667 -10977 4710 -10943
rect 4590 -11023 4710 -10977
rect 4590 -11057 4633 -11023
rect 4667 -11057 4710 -11023
rect 4590 -11130 4710 -11057
rect 5870 -10943 5990 -10897
rect 5870 -10977 5913 -10943
rect 5947 -10977 5990 -10943
rect 5870 -11023 5990 -10977
rect 5870 -11057 5913 -11023
rect 5947 -11057 5990 -11023
rect 5870 -11130 5990 -11057
rect 6020 -10863 6140 -10830
rect 6020 -10897 6063 -10863
rect 6097 -10897 6140 -10863
rect 6020 -10943 6140 -10897
rect 6020 -10977 6063 -10943
rect 6097 -10977 6140 -10943
rect 6020 -11023 6140 -10977
rect 6020 -11057 6063 -11023
rect 6097 -11057 6140 -11023
rect 6020 -11130 6140 -11057
rect 6170 -10863 6290 -10830
rect 6170 -10897 6213 -10863
rect 6247 -10897 6290 -10863
rect 6170 -10943 6290 -10897
rect 6170 -10977 6213 -10943
rect 6247 -10977 6290 -10943
rect 6170 -11023 6290 -10977
rect 6170 -11057 6213 -11023
rect 6247 -11057 6290 -11023
rect 6170 -11130 6290 -11057
rect 6320 -10863 6440 -10830
rect 6320 -10897 6363 -10863
rect 6397 -10897 6440 -10863
rect 6320 -10943 6440 -10897
rect 6320 -10977 6363 -10943
rect 6397 -10977 6440 -10943
rect 6320 -11023 6440 -10977
rect 6320 -11057 6363 -11023
rect 6397 -11057 6440 -11023
rect 6320 -11130 6440 -11057
rect 6470 -10863 6590 -10830
rect 6470 -10897 6513 -10863
rect 6547 -10897 6590 -10863
rect 6470 -10943 6590 -10897
rect 6470 -10977 6513 -10943
rect 6547 -10977 6590 -10943
rect 6470 -11023 6590 -10977
rect 6470 -11057 6513 -11023
rect 6547 -11057 6590 -11023
rect 6470 -11130 6590 -11057
rect 1801 -11923 1921 -11850
rect 1801 -11957 1844 -11923
rect 1878 -11957 1921 -11923
rect 1801 -12003 1921 -11957
rect 1801 -12037 1844 -12003
rect 1878 -12037 1921 -12003
rect 1801 -12083 1921 -12037
rect 1801 -12117 1844 -12083
rect 1878 -12117 1921 -12083
rect 1801 -12150 1921 -12117
rect 1951 -11923 2071 -11850
rect 1951 -11957 1994 -11923
rect 2028 -11957 2071 -11923
rect 1951 -12003 2071 -11957
rect 1951 -12037 1994 -12003
rect 2028 -12037 2071 -12003
rect 1951 -12083 2071 -12037
rect 1951 -12117 1994 -12083
rect 2028 -12117 2071 -12083
rect 1951 -12150 2071 -12117
rect 2101 -11923 2221 -11850
rect 2101 -11957 2144 -11923
rect 2178 -11957 2221 -11923
rect 2101 -12003 2221 -11957
rect 2101 -12037 2144 -12003
rect 2178 -12037 2221 -12003
rect 2101 -12083 2221 -12037
rect 2101 -12117 2144 -12083
rect 2178 -12117 2221 -12083
rect 2101 -12150 2221 -12117
rect 2251 -11923 2371 -11850
rect 2251 -11957 2294 -11923
rect 2328 -11957 2371 -11923
rect 2251 -12003 2371 -11957
rect 2251 -12037 2294 -12003
rect 2328 -12037 2371 -12003
rect 2251 -12083 2371 -12037
rect 2251 -12117 2294 -12083
rect 2328 -12117 2371 -12083
rect 2251 -12150 2371 -12117
rect 2401 -11923 2521 -11850
rect 2401 -11957 2444 -11923
rect 2478 -11957 2521 -11923
rect 2401 -12003 2521 -11957
rect 2401 -12037 2444 -12003
rect 2478 -12037 2521 -12003
rect 2401 -12083 2521 -12037
rect 2401 -12117 2444 -12083
rect 2478 -12117 2521 -12083
rect 2401 -12150 2521 -12117
rect 3851 -11923 3971 -11850
rect 3851 -11957 3894 -11923
rect 3928 -11957 3971 -11923
rect 3851 -12003 3971 -11957
rect 3851 -12037 3894 -12003
rect 3928 -12037 3971 -12003
rect 3851 -12083 3971 -12037
rect 3851 -12117 3894 -12083
rect 3928 -12117 3971 -12083
rect 3851 -12150 3971 -12117
rect 4001 -11923 4121 -11850
rect 4001 -11957 4044 -11923
rect 4078 -11957 4121 -11923
rect 4001 -12003 4121 -11957
rect 4001 -12037 4044 -12003
rect 4078 -12037 4121 -12003
rect 4001 -12083 4121 -12037
rect 4001 -12117 4044 -12083
rect 4078 -12117 4121 -12083
rect 4001 -12150 4121 -12117
rect 4151 -11923 4271 -11850
rect 4151 -11957 4194 -11923
rect 4228 -11957 4271 -11923
rect 4151 -12003 4271 -11957
rect 4151 -12037 4194 -12003
rect 4228 -12037 4271 -12003
rect 4151 -12083 4271 -12037
rect 4151 -12117 4194 -12083
rect 4228 -12117 4271 -12083
rect 4151 -12150 4271 -12117
rect 4301 -11923 4421 -11850
rect 4301 -11957 4344 -11923
rect 4378 -11957 4421 -11923
rect 4301 -12003 4421 -11957
rect 4301 -12037 4344 -12003
rect 4378 -12037 4421 -12003
rect 4301 -12083 4421 -12037
rect 4301 -12117 4344 -12083
rect 4378 -12117 4421 -12083
rect 4301 -12150 4421 -12117
rect 4451 -11923 4571 -11850
rect 4451 -11957 4494 -11923
rect 4528 -11957 4571 -11923
rect 4451 -12003 4571 -11957
rect 4451 -12037 4494 -12003
rect 4528 -12037 4571 -12003
rect 4451 -12083 4571 -12037
rect 4451 -12117 4494 -12083
rect 4528 -12117 4571 -12083
rect 4451 -12150 4571 -12117
rect 5891 -11924 6011 -11851
rect 5891 -11958 5934 -11924
rect 5968 -11958 6011 -11924
rect 5891 -12004 6011 -11958
rect 5891 -12038 5934 -12004
rect 5968 -12038 6011 -12004
rect 5891 -12084 6011 -12038
rect 5891 -12118 5934 -12084
rect 5968 -12118 6011 -12084
rect 5891 -12151 6011 -12118
rect 6041 -11924 6161 -11851
rect 6041 -11958 6084 -11924
rect 6118 -11958 6161 -11924
rect 6041 -12004 6161 -11958
rect 6041 -12038 6084 -12004
rect 6118 -12038 6161 -12004
rect 6041 -12084 6161 -12038
rect 6041 -12118 6084 -12084
rect 6118 -12118 6161 -12084
rect 6041 -12151 6161 -12118
rect 6191 -11924 6311 -11851
rect 6191 -11958 6234 -11924
rect 6268 -11958 6311 -11924
rect 6191 -12004 6311 -11958
rect 6191 -12038 6234 -12004
rect 6268 -12038 6311 -12004
rect 6191 -12084 6311 -12038
rect 6191 -12118 6234 -12084
rect 6268 -12118 6311 -12084
rect 6191 -12151 6311 -12118
rect 6341 -11924 6461 -11851
rect 6341 -11958 6384 -11924
rect 6418 -11958 6461 -11924
rect 6341 -12004 6461 -11958
rect 6341 -12038 6384 -12004
rect 6418 -12038 6461 -12004
rect 6341 -12084 6461 -12038
rect 6341 -12118 6384 -12084
rect 6418 -12118 6461 -12084
rect 6341 -12151 6461 -12118
rect 6491 -11924 6611 -11851
rect 6491 -11958 6534 -11924
rect 6568 -11958 6611 -11924
rect 6491 -12004 6611 -11958
rect 6491 -12038 6534 -12004
rect 6568 -12038 6611 -12004
rect 6491 -12084 6611 -12038
rect 6491 -12118 6534 -12084
rect 6568 -12118 6611 -12084
rect 6491 -12151 6611 -12118
<< ndiffc >>
rect 1063 1664 1097 1698
rect 1063 1584 1097 1618
rect 1063 1504 1097 1538
rect 1363 1664 1397 1698
rect 1363 1584 1397 1618
rect 1363 1504 1397 1538
rect 1663 1664 1697 1698
rect 1663 1584 1697 1618
rect 1663 1504 1697 1538
rect 1843 1664 1877 1698
rect 1843 1584 1877 1618
rect 1843 1504 1877 1538
rect 1993 1664 2027 1698
rect 1993 1584 2027 1618
rect 1993 1504 2027 1538
rect 2143 1664 2177 1698
rect 2143 1584 2177 1618
rect 2143 1504 2177 1538
rect 2293 1664 2327 1698
rect 2293 1584 2327 1618
rect 2293 1504 2327 1538
rect 2443 1664 2477 1698
rect 2443 1584 2477 1618
rect 2443 1504 2477 1538
rect 2623 1664 2657 1698
rect 2623 1584 2657 1618
rect 2623 1504 2657 1538
rect 2923 1664 2957 1698
rect 2923 1584 2957 1618
rect 2923 1504 2957 1538
rect 3223 1664 3257 1698
rect 3223 1584 3257 1618
rect 3223 1504 3257 1538
rect 3683 1664 3717 1698
rect 3683 1584 3717 1618
rect 3683 1504 3717 1538
rect 3983 1664 4017 1698
rect 3983 1584 4017 1618
rect 3983 1504 4017 1538
rect 4163 1664 4197 1698
rect 4163 1584 4197 1618
rect 4163 1504 4197 1538
rect 4313 1664 4347 1698
rect 4313 1584 4347 1618
rect 4313 1504 4347 1538
rect 4463 1664 4497 1698
rect 4463 1584 4497 1618
rect 4463 1504 4497 1538
rect 4613 1664 4647 1698
rect 4613 1584 4647 1618
rect 4613 1504 4647 1538
rect 4763 1664 4797 1698
rect 4763 1584 4797 1618
rect 4763 1504 4797 1538
rect 4943 1664 4977 1698
rect 4943 1584 4977 1618
rect 4943 1504 4977 1538
rect 5093 1664 5127 1698
rect 5093 1584 5127 1618
rect 5093 1504 5127 1538
rect 5243 1664 5277 1698
rect 5243 1584 5277 1618
rect 5243 1504 5277 1538
rect 5703 1664 5737 1698
rect 5703 1584 5737 1618
rect 5703 1504 5737 1538
rect 5853 1664 5887 1698
rect 5853 1584 5887 1618
rect 5853 1504 5887 1538
rect 6003 1664 6037 1698
rect 6003 1584 6037 1618
rect 6003 1504 6037 1538
rect 6183 1664 6217 1698
rect 6183 1584 6217 1618
rect 6183 1504 6217 1538
rect 6333 1664 6367 1698
rect 6333 1584 6367 1618
rect 6333 1504 6367 1538
rect 6483 1664 6517 1698
rect 6483 1584 6517 1618
rect 6483 1504 6517 1538
rect 6633 1664 6667 1698
rect 6633 1584 6667 1618
rect 6633 1504 6667 1538
rect 6783 1664 6817 1698
rect 6783 1584 6817 1618
rect 6783 1504 6817 1538
rect 6963 1664 6997 1698
rect 6963 1584 6997 1618
rect 6963 1504 6997 1538
rect 7263 1664 7297 1698
rect 7263 1584 7297 1618
rect 7263 1504 7297 1538
rect 1363 1024 1397 1058
rect 1363 944 1397 978
rect 1363 864 1397 898
rect 1513 1024 1547 1058
rect 1513 944 1547 978
rect 1513 864 1547 898
rect 1663 1024 1697 1058
rect 1663 944 1697 978
rect 1663 864 1697 898
rect 1843 1024 1877 1058
rect 1843 944 1877 978
rect 1843 864 1877 898
rect 1993 1024 2027 1058
rect 1993 944 2027 978
rect 1993 864 2027 898
rect 2143 1024 2177 1058
rect 2143 944 2177 978
rect 2143 864 2177 898
rect 2293 1024 2327 1058
rect 2293 944 2327 978
rect 2293 864 2327 898
rect 2443 1024 2477 1058
rect 2443 944 2477 978
rect 2443 864 2477 898
rect 2623 1024 2657 1058
rect 2623 944 2657 978
rect 2623 864 2657 898
rect 2923 1024 2957 1058
rect 2923 944 2957 978
rect 2923 864 2957 898
rect 3683 1024 3717 1058
rect 3683 944 3717 978
rect 3683 864 3717 898
rect 3833 1024 3867 1058
rect 3833 944 3867 978
rect 3833 864 3867 898
rect 3983 1024 4017 1058
rect 3983 944 4017 978
rect 3983 864 4017 898
rect 4163 1024 4197 1058
rect 4163 944 4197 978
rect 4163 864 4197 898
rect 4313 1024 4347 1058
rect 4313 944 4347 978
rect 4313 864 4347 898
rect 4463 1024 4497 1058
rect 4463 944 4497 978
rect 4463 864 4497 898
rect 4613 1024 4647 1058
rect 4613 944 4647 978
rect 4613 864 4647 898
rect 4763 1024 4797 1058
rect 4763 944 4797 978
rect 4763 864 4797 898
rect 4943 1024 4977 1058
rect 4943 944 4977 978
rect 4943 864 4977 898
rect 5243 1024 5277 1058
rect 5243 944 5277 978
rect 5243 864 5277 898
rect 5703 1024 5737 1058
rect 5703 944 5737 978
rect 5703 864 5737 898
rect 5853 1024 5887 1058
rect 5853 944 5887 978
rect 5853 864 5887 898
rect 6003 1024 6037 1058
rect 6003 944 6037 978
rect 6003 864 6037 898
rect 6183 1024 6217 1058
rect 6183 944 6217 978
rect 6183 864 6217 898
rect 6333 1024 6367 1058
rect 6333 944 6367 978
rect 6333 864 6367 898
rect 6483 1024 6517 1058
rect 6483 944 6517 978
rect 6483 864 6517 898
rect 6633 1024 6667 1058
rect 6633 944 6667 978
rect 6633 864 6667 898
rect 6783 1024 6817 1058
rect 6783 944 6817 978
rect 6783 864 6817 898
rect 6963 1024 6997 1058
rect 6963 944 6997 978
rect 6963 864 6997 898
rect 7263 1024 7297 1058
rect 7263 944 7297 978
rect 7263 864 7297 898
rect 1063 -1156 1097 -1122
rect 1063 -1236 1097 -1202
rect 1063 -1316 1097 -1282
rect 1363 -1156 1397 -1122
rect 1363 -1236 1397 -1202
rect 1363 -1316 1397 -1282
rect 1663 -1156 1697 -1122
rect 1663 -1236 1697 -1202
rect 1663 -1316 1697 -1282
rect 1843 -1156 1877 -1122
rect 1843 -1236 1877 -1202
rect 1843 -1316 1877 -1282
rect 1993 -1156 2027 -1122
rect 1993 -1236 2027 -1202
rect 1993 -1316 2027 -1282
rect 2143 -1156 2177 -1122
rect 2143 -1236 2177 -1202
rect 2143 -1316 2177 -1282
rect 2293 -1156 2327 -1122
rect 2293 -1236 2327 -1202
rect 2293 -1316 2327 -1282
rect 2443 -1156 2477 -1122
rect 2443 -1236 2477 -1202
rect 2443 -1316 2477 -1282
rect 2623 -1156 2657 -1122
rect 2623 -1236 2657 -1202
rect 2623 -1316 2657 -1282
rect 2923 -1156 2957 -1122
rect 2923 -1236 2957 -1202
rect 2923 -1316 2957 -1282
rect 3223 -1156 3257 -1122
rect 3223 -1236 3257 -1202
rect 3223 -1316 3257 -1282
rect 3703 -1156 3737 -1122
rect 3703 -1236 3737 -1202
rect 3703 -1316 3737 -1282
rect 3853 -1156 3887 -1122
rect 3853 -1236 3887 -1202
rect 3853 -1316 3887 -1282
rect 4033 -1156 4067 -1122
rect 4033 -1236 4067 -1202
rect 4033 -1316 4067 -1282
rect 4183 -1156 4217 -1122
rect 4183 -1236 4217 -1202
rect 4183 -1316 4217 -1282
rect 4333 -1156 4367 -1122
rect 4333 -1236 4367 -1202
rect 4333 -1316 4367 -1282
rect 4483 -1156 4517 -1122
rect 4483 -1236 4517 -1202
rect 4483 -1316 4517 -1282
rect 4633 -1156 4667 -1122
rect 4633 -1236 4667 -1202
rect 4633 -1316 4667 -1282
rect 4813 -1156 4847 -1122
rect 4813 -1236 4847 -1202
rect 4813 -1316 4847 -1282
rect 4963 -1156 4997 -1122
rect 4963 -1236 4997 -1202
rect 4963 -1316 4997 -1282
rect 5433 -1156 5467 -1122
rect 5433 -1236 5467 -1202
rect 5433 -1316 5467 -1282
rect 5583 -1156 5617 -1122
rect 5583 -1236 5617 -1202
rect 5583 -1316 5617 -1282
rect 5733 -1156 5767 -1122
rect 5733 -1236 5767 -1202
rect 5733 -1316 5767 -1282
rect 5913 -1156 5947 -1122
rect 5913 -1236 5947 -1202
rect 5913 -1316 5947 -1282
rect 6063 -1156 6097 -1122
rect 6063 -1236 6097 -1202
rect 6063 -1316 6097 -1282
rect 6213 -1156 6247 -1122
rect 6213 -1236 6247 -1202
rect 6213 -1316 6247 -1282
rect 6363 -1156 6397 -1122
rect 6363 -1236 6397 -1202
rect 6363 -1316 6397 -1282
rect 6513 -1156 6547 -1122
rect 6513 -1236 6547 -1202
rect 6513 -1316 6547 -1282
rect 6693 -1156 6727 -1122
rect 6693 -1236 6727 -1202
rect 6693 -1316 6727 -1282
rect 6993 -1156 7027 -1122
rect 6993 -1236 7027 -1202
rect 6993 -1316 7027 -1282
rect 1063 -1796 1097 -1762
rect 1063 -1876 1097 -1842
rect 1063 -1956 1097 -1922
rect 1363 -1796 1397 -1762
rect 1363 -1876 1397 -1842
rect 1363 -1956 1397 -1922
rect 1663 -1796 1697 -1762
rect 1663 -1876 1697 -1842
rect 1663 -1956 1697 -1922
rect 1843 -1796 1877 -1762
rect 1843 -1876 1877 -1842
rect 1843 -1956 1877 -1922
rect 1993 -1796 2027 -1762
rect 1993 -1876 2027 -1842
rect 1993 -1956 2027 -1922
rect 2143 -1796 2177 -1762
rect 2143 -1876 2177 -1842
rect 2143 -1956 2177 -1922
rect 2293 -1796 2327 -1762
rect 2293 -1876 2327 -1842
rect 2293 -1956 2327 -1922
rect 2443 -1796 2477 -1762
rect 2443 -1876 2477 -1842
rect 2443 -1956 2477 -1922
rect 2623 -1796 2657 -1762
rect 2623 -1876 2657 -1842
rect 2623 -1956 2657 -1922
rect 2923 -1796 2957 -1762
rect 2923 -1876 2957 -1842
rect 2923 -1956 2957 -1922
rect 3223 -1796 3257 -1762
rect 3223 -1876 3257 -1842
rect 3223 -1956 3257 -1922
rect 3703 -1796 3737 -1762
rect 3703 -1876 3737 -1842
rect 3703 -1956 3737 -1922
rect 3853 -1796 3887 -1762
rect 3853 -1876 3887 -1842
rect 3853 -1956 3887 -1922
rect 4033 -1796 4067 -1762
rect 4033 -1876 4067 -1842
rect 4033 -1956 4067 -1922
rect 4183 -1796 4217 -1762
rect 4183 -1876 4217 -1842
rect 4183 -1956 4217 -1922
rect 4333 -1796 4367 -1762
rect 4333 -1876 4367 -1842
rect 4333 -1956 4367 -1922
rect 4483 -1796 4517 -1762
rect 4483 -1876 4517 -1842
rect 4483 -1956 4517 -1922
rect 4633 -1796 4667 -1762
rect 4633 -1876 4667 -1842
rect 4633 -1956 4667 -1922
rect 4813 -1796 4847 -1762
rect 4813 -1876 4847 -1842
rect 4813 -1956 4847 -1922
rect 4963 -1796 4997 -1762
rect 4963 -1876 4997 -1842
rect 4963 -1956 4997 -1922
rect 5433 -1796 5467 -1762
rect 5433 -1876 5467 -1842
rect 5433 -1956 5467 -1922
rect 5583 -1796 5617 -1762
rect 5583 -1876 5617 -1842
rect 5583 -1956 5617 -1922
rect 5733 -1796 5767 -1762
rect 5733 -1876 5767 -1842
rect 5733 -1956 5767 -1922
rect 5913 -1796 5947 -1762
rect 5913 -1876 5947 -1842
rect 5913 -1956 5947 -1922
rect 6063 -1796 6097 -1762
rect 6063 -1876 6097 -1842
rect 6063 -1956 6097 -1922
rect 6213 -1796 6247 -1762
rect 6213 -1876 6247 -1842
rect 6213 -1956 6247 -1922
rect 6363 -1796 6397 -1762
rect 6363 -1876 6397 -1842
rect 6363 -1956 6397 -1922
rect 6513 -1796 6547 -1762
rect 6513 -1876 6547 -1842
rect 6513 -1956 6547 -1922
rect 6693 -1796 6727 -1762
rect 6693 -1876 6727 -1842
rect 6693 -1956 6727 -1922
rect 6993 -1796 7027 -1762
rect 6993 -1876 7027 -1842
rect 6993 -1956 7027 -1922
rect 1214 -3976 1248 -3942
rect 1214 -4056 1248 -4022
rect 1214 -4136 1248 -4102
rect 1364 -3976 1398 -3942
rect 1364 -4056 1398 -4022
rect 1364 -4136 1398 -4102
rect 1514 -3976 1548 -3942
rect 1514 -4056 1548 -4022
rect 1514 -4136 1548 -4102
rect 1664 -3976 1698 -3942
rect 1664 -4056 1698 -4022
rect 1664 -4136 1698 -4102
rect 1844 -3976 1878 -3942
rect 1844 -4056 1878 -4022
rect 1844 -4136 1878 -4102
rect 1994 -3976 2028 -3942
rect 1994 -4056 2028 -4022
rect 1994 -4136 2028 -4102
rect 2144 -3976 2178 -3942
rect 2144 -4056 2178 -4022
rect 2144 -4136 2178 -4102
rect 2294 -3976 2328 -3942
rect 2294 -4056 2328 -4022
rect 2294 -4136 2328 -4102
rect 2444 -3976 2478 -3942
rect 2444 -4056 2478 -4022
rect 2444 -4136 2478 -4102
rect 2624 -3976 2658 -3942
rect 2624 -4056 2658 -4022
rect 2624 -4136 2658 -4102
rect 3074 -3976 3108 -3942
rect 3074 -4056 3108 -4022
rect 3074 -4136 3108 -4102
rect 3564 -3976 3598 -3942
rect 3564 -4056 3598 -4022
rect 3564 -4136 3598 -4102
rect 3714 -3976 3748 -3942
rect 3714 -4056 3748 -4022
rect 3714 -4136 3748 -4102
rect 3894 -3976 3928 -3942
rect 3894 -4056 3928 -4022
rect 3894 -4136 3928 -4102
rect 4044 -3976 4078 -3942
rect 4044 -4056 4078 -4022
rect 4044 -4136 4078 -4102
rect 4194 -3976 4228 -3942
rect 4194 -4056 4228 -4022
rect 4194 -4136 4228 -4102
rect 4344 -3976 4378 -3942
rect 4344 -4056 4378 -4022
rect 4344 -4136 4378 -4102
rect 4494 -3976 4528 -3942
rect 4494 -4056 4528 -4022
rect 4494 -4136 4528 -4102
rect 4674 -3976 4708 -3942
rect 4674 -4056 4708 -4022
rect 4674 -4136 4708 -4102
rect 4824 -3976 4858 -3942
rect 4824 -4056 4858 -4022
rect 4824 -4136 4858 -4102
rect 5304 -3977 5338 -3943
rect 5304 -4057 5338 -4023
rect 5304 -4137 5338 -4103
rect 5454 -3977 5488 -3943
rect 5454 -4057 5488 -4023
rect 5454 -4137 5488 -4103
rect 5604 -3977 5638 -3943
rect 5604 -4057 5638 -4023
rect 5604 -4137 5638 -4103
rect 5754 -3977 5788 -3943
rect 5754 -4057 5788 -4023
rect 5754 -4137 5788 -4103
rect 5934 -3977 5968 -3943
rect 5934 -4057 5968 -4023
rect 5934 -4137 5968 -4103
rect 6084 -3977 6118 -3943
rect 6084 -4057 6118 -4023
rect 6084 -4137 6118 -4103
rect 6234 -3977 6268 -3943
rect 6234 -4057 6268 -4023
rect 6234 -4137 6268 -4103
rect 6384 -3977 6418 -3943
rect 6384 -4057 6418 -4023
rect 6384 -4137 6418 -4103
rect 6534 -3977 6568 -3943
rect 6534 -4057 6568 -4023
rect 6534 -4137 6568 -4103
rect 6714 -3977 6748 -3943
rect 6714 -4057 6748 -4023
rect 6714 -4137 6748 -4103
rect 7164 -3977 7198 -3943
rect 7164 -4057 7198 -4023
rect 7164 -4137 7198 -4103
rect 1103 -4696 1137 -4662
rect 1103 -4776 1137 -4742
rect 1103 -4856 1137 -4822
rect 1253 -4696 1287 -4662
rect 1253 -4776 1287 -4742
rect 1253 -4856 1287 -4822
rect 1403 -4696 1437 -4662
rect 1403 -4776 1437 -4742
rect 1403 -4856 1437 -4822
rect 1553 -4696 1587 -4662
rect 1553 -4776 1587 -4742
rect 1553 -4856 1587 -4822
rect 1703 -4696 1737 -4662
rect 1703 -4776 1737 -4742
rect 1703 -4856 1737 -4822
rect 1883 -4696 1917 -4662
rect 1883 -4776 1917 -4742
rect 1883 -4856 1917 -4822
rect 2033 -4696 2067 -4662
rect 2033 -4776 2067 -4742
rect 2033 -4856 2067 -4822
rect 2183 -4696 2217 -4662
rect 2183 -4776 2217 -4742
rect 2183 -4856 2217 -4822
rect 2333 -4696 2367 -4662
rect 2333 -4776 2367 -4742
rect 2333 -4856 2367 -4822
rect 2483 -4696 2517 -4662
rect 2483 -4776 2517 -4742
rect 2483 -4856 2517 -4822
rect 2663 -4696 2697 -4662
rect 2663 -4776 2697 -4742
rect 2663 -4856 2697 -4822
rect 3263 -4696 3297 -4662
rect 3263 -4776 3297 -4742
rect 3263 -4856 3297 -4822
rect 3764 -4697 3798 -4663
rect 3764 -4777 3798 -4743
rect 3764 -4857 3798 -4823
rect 3914 -4697 3948 -4663
rect 3914 -4777 3948 -4743
rect 3914 -4857 3948 -4823
rect 4094 -4697 4128 -4663
rect 4094 -4777 4128 -4743
rect 4094 -4857 4128 -4823
rect 4244 -4697 4278 -4663
rect 4244 -4777 4278 -4743
rect 4244 -4857 4278 -4823
rect 4394 -4697 4428 -4663
rect 4394 -4777 4428 -4743
rect 4394 -4857 4428 -4823
rect 4544 -4697 4578 -4663
rect 4544 -4777 4578 -4743
rect 4544 -4857 4578 -4823
rect 4694 -4697 4728 -4663
rect 4694 -4777 4728 -4743
rect 4694 -4857 4728 -4823
rect 4874 -4697 4908 -4663
rect 4874 -4777 4908 -4743
rect 4874 -4857 4908 -4823
rect 5024 -4697 5058 -4663
rect 5024 -4777 5058 -4743
rect 5024 -4857 5058 -4823
rect 5523 -4697 5557 -4663
rect 5523 -4777 5557 -4743
rect 5523 -4857 5557 -4823
rect 5673 -4697 5707 -4663
rect 5673 -4777 5707 -4743
rect 5673 -4857 5707 -4823
rect 5823 -4697 5857 -4663
rect 5823 -4777 5857 -4743
rect 5823 -4857 5857 -4823
rect 5973 -4697 6007 -4663
rect 5973 -4777 6007 -4743
rect 5973 -4857 6007 -4823
rect 6153 -4697 6187 -4663
rect 6153 -4777 6187 -4743
rect 6153 -4857 6187 -4823
rect 6303 -4697 6337 -4663
rect 6303 -4777 6337 -4743
rect 6303 -4857 6337 -4823
rect 6453 -4697 6487 -4663
rect 6453 -4777 6487 -4743
rect 6453 -4857 6487 -4823
rect 6603 -4697 6637 -4663
rect 6603 -4777 6637 -4743
rect 6603 -4857 6637 -4823
rect 6753 -4697 6787 -4663
rect 6753 -4777 6787 -4743
rect 6753 -4857 6787 -4823
rect 6933 -4697 6967 -4663
rect 6933 -4777 6967 -4743
rect 6933 -4857 6967 -4823
rect 7383 -4697 7417 -4663
rect 7383 -4777 7417 -4743
rect 7383 -4857 7417 -4823
rect 1103 -6877 1137 -6843
rect 1103 -6957 1137 -6923
rect 1103 -7037 1137 -7003
rect 1403 -6877 1437 -6843
rect 1403 -6957 1437 -6923
rect 1403 -7037 1437 -7003
rect 1703 -6877 1737 -6843
rect 1703 -6957 1737 -6923
rect 1703 -7037 1737 -7003
rect 1883 -6877 1917 -6843
rect 1883 -6957 1917 -6923
rect 1883 -7037 1917 -7003
rect 2033 -6877 2067 -6843
rect 2033 -6957 2067 -6923
rect 2033 -7037 2067 -7003
rect 2183 -6877 2217 -6843
rect 2183 -6957 2217 -6923
rect 2183 -7037 2217 -7003
rect 2333 -6877 2367 -6843
rect 2333 -6957 2367 -6923
rect 2333 -7037 2367 -7003
rect 2483 -6877 2517 -6843
rect 2483 -6957 2517 -6923
rect 2483 -7037 2517 -7003
rect 2663 -6877 2697 -6843
rect 2663 -6957 2697 -6923
rect 2663 -7037 2697 -7003
rect 2963 -6877 2997 -6843
rect 2963 -6957 2997 -6923
rect 2963 -7037 2997 -7003
rect 3263 -6877 3297 -6843
rect 3263 -6957 3297 -6923
rect 3263 -7037 3297 -7003
rect 3763 -6877 3797 -6843
rect 3763 -6957 3797 -6923
rect 3763 -7037 3797 -7003
rect 3913 -6877 3947 -6843
rect 3913 -6957 3947 -6923
rect 3913 -7037 3947 -7003
rect 4093 -6877 4127 -6843
rect 4093 -6957 4127 -6923
rect 4093 -7037 4127 -7003
rect 4243 -6877 4277 -6843
rect 4243 -6957 4277 -6923
rect 4243 -7037 4277 -7003
rect 4393 -6877 4427 -6843
rect 4393 -6957 4427 -6923
rect 4393 -7037 4427 -7003
rect 4543 -6877 4577 -6843
rect 4543 -6957 4577 -6923
rect 4543 -7037 4577 -7003
rect 4693 -6877 4727 -6843
rect 4693 -6957 4727 -6923
rect 4693 -7037 4727 -7003
rect 4873 -6877 4907 -6843
rect 4873 -6957 4907 -6923
rect 4873 -7037 4907 -7003
rect 5023 -6877 5057 -6843
rect 5023 -6957 5057 -6923
rect 5023 -7037 5057 -7003
rect 5492 -6877 5526 -6843
rect 5492 -6957 5526 -6923
rect 5492 -7037 5526 -7003
rect 5642 -6877 5676 -6843
rect 5642 -6957 5676 -6923
rect 5642 -7037 5676 -7003
rect 5792 -6877 5826 -6843
rect 5792 -6957 5826 -6923
rect 5792 -7037 5826 -7003
rect 5972 -6877 6006 -6843
rect 5972 -6957 6006 -6923
rect 5972 -7037 6006 -7003
rect 6122 -6877 6156 -6843
rect 6122 -6957 6156 -6923
rect 6122 -7037 6156 -7003
rect 6272 -6877 6306 -6843
rect 6272 -6957 6306 -6923
rect 6272 -7037 6306 -7003
rect 6422 -6877 6456 -6843
rect 6422 -6957 6456 -6923
rect 6422 -7037 6456 -7003
rect 6572 -6877 6606 -6843
rect 6572 -6957 6606 -6923
rect 6572 -7037 6606 -7003
rect 6752 -6877 6786 -6843
rect 6752 -6957 6786 -6923
rect 6752 -7037 6786 -7003
rect 7052 -6877 7086 -6843
rect 7052 -6957 7086 -6923
rect 7052 -7037 7086 -7003
rect 1103 -7517 1137 -7483
rect 1103 -7597 1137 -7563
rect 1103 -7677 1137 -7643
rect 1403 -7517 1437 -7483
rect 1403 -7597 1437 -7563
rect 1403 -7677 1437 -7643
rect 1703 -7517 1737 -7483
rect 1703 -7597 1737 -7563
rect 1703 -7677 1737 -7643
rect 1883 -7517 1917 -7483
rect 1883 -7597 1917 -7563
rect 1883 -7677 1917 -7643
rect 2033 -7517 2067 -7483
rect 2033 -7597 2067 -7563
rect 2033 -7677 2067 -7643
rect 2183 -7517 2217 -7483
rect 2183 -7597 2217 -7563
rect 2183 -7677 2217 -7643
rect 2333 -7517 2367 -7483
rect 2333 -7597 2367 -7563
rect 2333 -7677 2367 -7643
rect 2483 -7517 2517 -7483
rect 2483 -7597 2517 -7563
rect 2483 -7677 2517 -7643
rect 2663 -7517 2697 -7483
rect 2663 -7597 2697 -7563
rect 2663 -7677 2697 -7643
rect 2963 -7517 2997 -7483
rect 2963 -7597 2997 -7563
rect 2963 -7677 2997 -7643
rect 3263 -7517 3297 -7483
rect 3263 -7597 3297 -7563
rect 3263 -7677 3297 -7643
rect 3763 -7517 3797 -7483
rect 3763 -7597 3797 -7563
rect 3763 -7677 3797 -7643
rect 3913 -7517 3947 -7483
rect 3913 -7597 3947 -7563
rect 3913 -7677 3947 -7643
rect 4093 -7517 4127 -7483
rect 4093 -7597 4127 -7563
rect 4093 -7677 4127 -7643
rect 4243 -7517 4277 -7483
rect 4243 -7597 4277 -7563
rect 4243 -7677 4277 -7643
rect 4393 -7517 4427 -7483
rect 4393 -7597 4427 -7563
rect 4393 -7677 4427 -7643
rect 4543 -7517 4577 -7483
rect 4543 -7597 4577 -7563
rect 4543 -7677 4577 -7643
rect 4693 -7517 4727 -7483
rect 4693 -7597 4727 -7563
rect 4693 -7677 4727 -7643
rect 4873 -7517 4907 -7483
rect 4873 -7597 4907 -7563
rect 4873 -7677 4907 -7643
rect 5023 -7517 5057 -7483
rect 5023 -7597 5057 -7563
rect 5023 -7677 5057 -7643
rect 5492 -7517 5526 -7483
rect 5492 -7597 5526 -7563
rect 5492 -7677 5526 -7643
rect 5642 -7517 5676 -7483
rect 5642 -7597 5676 -7563
rect 5642 -7677 5676 -7643
rect 5792 -7517 5826 -7483
rect 5792 -7597 5826 -7563
rect 5792 -7677 5826 -7643
rect 5972 -7517 6006 -7483
rect 5972 -7597 6006 -7563
rect 5972 -7677 6006 -7643
rect 6122 -7517 6156 -7483
rect 6122 -7597 6156 -7563
rect 6122 -7677 6156 -7643
rect 6272 -7517 6306 -7483
rect 6272 -7597 6306 -7563
rect 6272 -7677 6306 -7643
rect 6422 -7517 6456 -7483
rect 6422 -7597 6456 -7563
rect 6422 -7677 6456 -7643
rect 6572 -7517 6606 -7483
rect 6572 -7597 6606 -7563
rect 6572 -7677 6606 -7643
rect 6752 -7517 6786 -7483
rect 6752 -7597 6786 -7563
rect 6752 -7677 6786 -7643
rect 7052 -7517 7086 -7483
rect 7052 -7597 7086 -7563
rect 7052 -7677 7086 -7643
rect 1063 -9697 1097 -9663
rect 1063 -9777 1097 -9743
rect 1063 -9857 1097 -9823
rect 1363 -9697 1397 -9663
rect 1363 -9777 1397 -9743
rect 1363 -9857 1397 -9823
rect 1663 -9697 1697 -9663
rect 1663 -9777 1697 -9743
rect 1663 -9857 1697 -9823
rect 1843 -9697 1877 -9663
rect 1843 -9777 1877 -9743
rect 1843 -9857 1877 -9823
rect 1993 -9697 2027 -9663
rect 1993 -9777 2027 -9743
rect 1993 -9857 2027 -9823
rect 2143 -9697 2177 -9663
rect 2143 -9777 2177 -9743
rect 2143 -9857 2177 -9823
rect 2293 -9697 2327 -9663
rect 2293 -9777 2327 -9743
rect 2293 -9857 2327 -9823
rect 2443 -9697 2477 -9663
rect 2443 -9777 2477 -9743
rect 2443 -9857 2477 -9823
rect 2623 -9697 2657 -9663
rect 2623 -9777 2657 -9743
rect 2623 -9857 2657 -9823
rect 2923 -9697 2957 -9663
rect 2923 -9777 2957 -9743
rect 2923 -9857 2957 -9823
rect 3223 -9697 3257 -9663
rect 3223 -9777 3257 -9743
rect 3223 -9857 3257 -9823
rect 3703 -9697 3737 -9663
rect 3703 -9777 3737 -9743
rect 3703 -9857 3737 -9823
rect 3853 -9697 3887 -9663
rect 3853 -9777 3887 -9743
rect 3853 -9857 3887 -9823
rect 4033 -9697 4067 -9663
rect 4033 -9777 4067 -9743
rect 4033 -9857 4067 -9823
rect 4183 -9697 4217 -9663
rect 4183 -9777 4217 -9743
rect 4183 -9857 4217 -9823
rect 4333 -9697 4367 -9663
rect 4333 -9777 4367 -9743
rect 4333 -9857 4367 -9823
rect 4483 -9697 4517 -9663
rect 4483 -9777 4517 -9743
rect 4483 -9857 4517 -9823
rect 4633 -9697 4667 -9663
rect 4633 -9777 4667 -9743
rect 4633 -9857 4667 -9823
rect 4813 -9697 4847 -9663
rect 4813 -9777 4847 -9743
rect 4813 -9857 4847 -9823
rect 4963 -9697 4997 -9663
rect 4963 -9777 4997 -9743
rect 4963 -9857 4997 -9823
rect 5433 -9697 5467 -9663
rect 5433 -9777 5467 -9743
rect 5433 -9857 5467 -9823
rect 5583 -9697 5617 -9663
rect 5583 -9777 5617 -9743
rect 5583 -9857 5617 -9823
rect 5733 -9697 5767 -9663
rect 5733 -9777 5767 -9743
rect 5733 -9857 5767 -9823
rect 5913 -9697 5947 -9663
rect 5913 -9777 5947 -9743
rect 5913 -9857 5947 -9823
rect 6063 -9697 6097 -9663
rect 6063 -9777 6097 -9743
rect 6063 -9857 6097 -9823
rect 6213 -9697 6247 -9663
rect 6213 -9777 6247 -9743
rect 6213 -9857 6247 -9823
rect 6363 -9697 6397 -9663
rect 6363 -9777 6397 -9743
rect 6363 -9857 6397 -9823
rect 6513 -9697 6547 -9663
rect 6513 -9777 6547 -9743
rect 6513 -9857 6547 -9823
rect 6693 -9697 6727 -9663
rect 6693 -9777 6727 -9743
rect 6693 -9857 6727 -9823
rect 6993 -9697 7027 -9663
rect 6993 -9777 7027 -9743
rect 6993 -9857 7027 -9823
rect 1063 -10337 1097 -10303
rect 1063 -10417 1097 -10383
rect 1063 -10497 1097 -10463
rect 1363 -10337 1397 -10303
rect 1363 -10417 1397 -10383
rect 1363 -10497 1397 -10463
rect 1663 -10337 1697 -10303
rect 1663 -10417 1697 -10383
rect 1663 -10497 1697 -10463
rect 1843 -10337 1877 -10303
rect 1843 -10417 1877 -10383
rect 1843 -10497 1877 -10463
rect 1993 -10337 2027 -10303
rect 1993 -10417 2027 -10383
rect 1993 -10497 2027 -10463
rect 2143 -10337 2177 -10303
rect 2143 -10417 2177 -10383
rect 2143 -10497 2177 -10463
rect 2293 -10337 2327 -10303
rect 2293 -10417 2327 -10383
rect 2293 -10497 2327 -10463
rect 2443 -10337 2477 -10303
rect 2443 -10417 2477 -10383
rect 2443 -10497 2477 -10463
rect 2623 -10337 2657 -10303
rect 2623 -10417 2657 -10383
rect 2623 -10497 2657 -10463
rect 2923 -10337 2957 -10303
rect 2923 -10417 2957 -10383
rect 2923 -10497 2957 -10463
rect 3223 -10337 3257 -10303
rect 3223 -10417 3257 -10383
rect 3223 -10497 3257 -10463
rect 3703 -10337 3737 -10303
rect 3703 -10417 3737 -10383
rect 3703 -10497 3737 -10463
rect 3853 -10337 3887 -10303
rect 3853 -10417 3887 -10383
rect 3853 -10497 3887 -10463
rect 4033 -10337 4067 -10303
rect 4033 -10417 4067 -10383
rect 4033 -10497 4067 -10463
rect 4183 -10337 4217 -10303
rect 4183 -10417 4217 -10383
rect 4183 -10497 4217 -10463
rect 4333 -10337 4367 -10303
rect 4333 -10417 4367 -10383
rect 4333 -10497 4367 -10463
rect 4483 -10337 4517 -10303
rect 4483 -10417 4517 -10383
rect 4483 -10497 4517 -10463
rect 4633 -10337 4667 -10303
rect 4633 -10417 4667 -10383
rect 4633 -10497 4667 -10463
rect 4813 -10337 4847 -10303
rect 4813 -10417 4847 -10383
rect 4813 -10497 4847 -10463
rect 4963 -10337 4997 -10303
rect 4963 -10417 4997 -10383
rect 4963 -10497 4997 -10463
rect 5433 -10337 5467 -10303
rect 5433 -10417 5467 -10383
rect 5433 -10497 5467 -10463
rect 5583 -10337 5617 -10303
rect 5583 -10417 5617 -10383
rect 5583 -10497 5617 -10463
rect 5733 -10337 5767 -10303
rect 5733 -10417 5767 -10383
rect 5733 -10497 5767 -10463
rect 5913 -10337 5947 -10303
rect 5913 -10417 5947 -10383
rect 5913 -10497 5947 -10463
rect 6063 -10337 6097 -10303
rect 6063 -10417 6097 -10383
rect 6063 -10497 6097 -10463
rect 6213 -10337 6247 -10303
rect 6213 -10417 6247 -10383
rect 6213 -10497 6247 -10463
rect 6363 -10337 6397 -10303
rect 6363 -10417 6397 -10383
rect 6363 -10497 6397 -10463
rect 6513 -10337 6547 -10303
rect 6513 -10417 6547 -10383
rect 6513 -10497 6547 -10463
rect 6693 -10337 6727 -10303
rect 6693 -10417 6727 -10383
rect 6693 -10497 6727 -10463
rect 6993 -10337 7027 -10303
rect 6993 -10417 7027 -10383
rect 6993 -10497 7027 -10463
rect 1214 -12517 1248 -12483
rect 1214 -12597 1248 -12563
rect 1214 -12677 1248 -12643
rect 1364 -12517 1398 -12483
rect 1364 -12597 1398 -12563
rect 1364 -12677 1398 -12643
rect 1514 -12517 1548 -12483
rect 1514 -12597 1548 -12563
rect 1514 -12677 1548 -12643
rect 1664 -12517 1698 -12483
rect 1664 -12597 1698 -12563
rect 1664 -12677 1698 -12643
rect 1844 -12517 1878 -12483
rect 1844 -12597 1878 -12563
rect 1844 -12677 1878 -12643
rect 1994 -12517 2028 -12483
rect 1994 -12597 2028 -12563
rect 1994 -12677 2028 -12643
rect 2144 -12517 2178 -12483
rect 2144 -12597 2178 -12563
rect 2144 -12677 2178 -12643
rect 2294 -12517 2328 -12483
rect 2294 -12597 2328 -12563
rect 2294 -12677 2328 -12643
rect 2444 -12517 2478 -12483
rect 2444 -12597 2478 -12563
rect 2444 -12677 2478 -12643
rect 2624 -12517 2658 -12483
rect 2624 -12597 2658 -12563
rect 2624 -12677 2658 -12643
rect 3074 -12517 3108 -12483
rect 3074 -12597 3108 -12563
rect 3074 -12677 3108 -12643
rect 3564 -12517 3598 -12483
rect 3564 -12597 3598 -12563
rect 3564 -12677 3598 -12643
rect 3714 -12517 3748 -12483
rect 3714 -12597 3748 -12563
rect 3714 -12677 3748 -12643
rect 3894 -12517 3928 -12483
rect 3894 -12597 3928 -12563
rect 3894 -12677 3928 -12643
rect 4044 -12517 4078 -12483
rect 4044 -12597 4078 -12563
rect 4044 -12677 4078 -12643
rect 4194 -12517 4228 -12483
rect 4194 -12597 4228 -12563
rect 4194 -12677 4228 -12643
rect 4344 -12517 4378 -12483
rect 4344 -12597 4378 -12563
rect 4344 -12677 4378 -12643
rect 4494 -12517 4528 -12483
rect 4494 -12597 4528 -12563
rect 4494 -12677 4528 -12643
rect 4674 -12517 4708 -12483
rect 4674 -12597 4708 -12563
rect 4674 -12677 4708 -12643
rect 4824 -12517 4858 -12483
rect 4824 -12597 4858 -12563
rect 4824 -12677 4858 -12643
rect 5304 -12518 5338 -12484
rect 5304 -12598 5338 -12564
rect 5304 -12678 5338 -12644
rect 5454 -12518 5488 -12484
rect 5454 -12598 5488 -12564
rect 5454 -12678 5488 -12644
rect 5604 -12518 5638 -12484
rect 5604 -12598 5638 -12564
rect 5604 -12678 5638 -12644
rect 5754 -12518 5788 -12484
rect 5754 -12598 5788 -12564
rect 5754 -12678 5788 -12644
rect 5934 -12518 5968 -12484
rect 5934 -12598 5968 -12564
rect 5934 -12678 5968 -12644
rect 6084 -12518 6118 -12484
rect 6084 -12598 6118 -12564
rect 6084 -12678 6118 -12644
rect 6234 -12518 6268 -12484
rect 6234 -12598 6268 -12564
rect 6234 -12678 6268 -12644
rect 6384 -12518 6418 -12484
rect 6384 -12598 6418 -12564
rect 6384 -12678 6418 -12644
rect 6534 -12518 6568 -12484
rect 6534 -12598 6568 -12564
rect 6534 -12678 6568 -12644
rect 6714 -12518 6748 -12484
rect 6714 -12598 6748 -12564
rect 6714 -12678 6748 -12644
rect 7164 -12518 7198 -12484
rect 7164 -12598 7198 -12564
rect 7164 -12678 7198 -12644
<< pdiffc >>
rect 1843 2224 1877 2258
rect 1843 2144 1877 2178
rect 1843 2064 1877 2098
rect 1993 2224 2027 2258
rect 1993 2144 2027 2178
rect 1993 2064 2027 2098
rect 2143 2224 2177 2258
rect 2143 2144 2177 2178
rect 2143 2064 2177 2098
rect 2293 2224 2327 2258
rect 2293 2144 2327 2178
rect 2293 2064 2327 2098
rect 2443 2224 2477 2258
rect 2443 2144 2477 2178
rect 2443 2064 2477 2098
rect 4163 2224 4197 2258
rect 4163 2144 4197 2178
rect 4163 2064 4197 2098
rect 4313 2224 4347 2258
rect 4313 2144 4347 2178
rect 4313 2064 4347 2098
rect 4463 2224 4497 2258
rect 4463 2144 4497 2178
rect 4463 2064 4497 2098
rect 4613 2224 4647 2258
rect 4613 2144 4647 2178
rect 4613 2064 4647 2098
rect 4763 2224 4797 2258
rect 4763 2144 4797 2178
rect 6183 2224 6217 2258
rect 4763 2064 4797 2098
rect 6183 2144 6217 2178
rect 6183 2064 6217 2098
rect 6333 2224 6367 2258
rect 6333 2144 6367 2178
rect 6333 2064 6367 2098
rect 6483 2224 6517 2258
rect 6483 2144 6517 2178
rect 6483 2064 6517 2098
rect 6633 2224 6667 2258
rect 6633 2144 6667 2178
rect 6633 2064 6667 2098
rect 6783 2224 6817 2258
rect 6783 2144 6817 2178
rect 6783 2064 6817 2098
rect 1843 464 1877 498
rect 1843 384 1877 418
rect 1843 304 1877 338
rect 1993 464 2027 498
rect 1993 384 2027 418
rect 1993 304 2027 338
rect 2143 464 2177 498
rect 2143 384 2177 418
rect 2143 304 2177 338
rect 2293 464 2327 498
rect 2293 384 2327 418
rect 2293 304 2327 338
rect 2443 464 2477 498
rect 2443 384 2477 418
rect 2443 304 2477 338
rect 4163 464 4197 498
rect 4163 384 4197 418
rect 4163 304 4197 338
rect 4313 464 4347 498
rect 4313 384 4347 418
rect 4313 304 4347 338
rect 4463 464 4497 498
rect 4463 384 4497 418
rect 4463 304 4497 338
rect 4613 464 4647 498
rect 4613 384 4647 418
rect 4613 304 4647 338
rect 4763 464 4797 498
rect 4763 384 4797 418
rect 6183 464 6217 498
rect 4763 304 4797 338
rect 6183 384 6217 418
rect 6183 304 6217 338
rect 6333 464 6367 498
rect 6333 384 6367 418
rect 6333 304 6367 338
rect 6483 464 6517 498
rect 6483 384 6517 418
rect 6483 304 6517 338
rect 6633 464 6667 498
rect 6633 384 6667 418
rect 6633 304 6667 338
rect 6783 464 6817 498
rect 6783 384 6817 418
rect 6783 304 6817 338
rect 1843 -596 1877 -562
rect 1843 -676 1877 -642
rect 1843 -756 1877 -722
rect 1993 -596 2027 -562
rect 1993 -676 2027 -642
rect 1993 -756 2027 -722
rect 2143 -596 2177 -562
rect 2143 -676 2177 -642
rect 2143 -756 2177 -722
rect 2293 -596 2327 -562
rect 2293 -676 2327 -642
rect 2293 -756 2327 -722
rect 2443 -596 2477 -562
rect 2443 -676 2477 -642
rect 2443 -756 2477 -722
rect 4033 -596 4067 -562
rect 4033 -676 4067 -642
rect 4033 -756 4067 -722
rect 4183 -596 4217 -562
rect 4183 -676 4217 -642
rect 4183 -756 4217 -722
rect 4333 -596 4367 -562
rect 4333 -676 4367 -642
rect 4333 -756 4367 -722
rect 4483 -596 4517 -562
rect 4483 -676 4517 -642
rect 4483 -756 4517 -722
rect 4633 -596 4667 -562
rect 4633 -676 4667 -642
rect 5913 -596 5947 -562
rect 5913 -676 5947 -642
rect 4633 -756 4667 -722
rect 5913 -756 5947 -722
rect 6063 -596 6097 -562
rect 6063 -676 6097 -642
rect 6063 -756 6097 -722
rect 6213 -596 6247 -562
rect 6213 -676 6247 -642
rect 6213 -756 6247 -722
rect 6363 -596 6397 -562
rect 6363 -676 6397 -642
rect 6363 -756 6397 -722
rect 6513 -596 6547 -562
rect 6513 -676 6547 -642
rect 6513 -756 6547 -722
rect 1843 -2356 1877 -2322
rect 1843 -2436 1877 -2402
rect 1843 -2516 1877 -2482
rect 1993 -2356 2027 -2322
rect 1993 -2436 2027 -2402
rect 1993 -2516 2027 -2482
rect 2143 -2356 2177 -2322
rect 2143 -2436 2177 -2402
rect 2143 -2516 2177 -2482
rect 2293 -2356 2327 -2322
rect 2293 -2436 2327 -2402
rect 2293 -2516 2327 -2482
rect 2443 -2356 2477 -2322
rect 2443 -2436 2477 -2402
rect 2443 -2516 2477 -2482
rect 4033 -2356 4067 -2322
rect 4033 -2436 4067 -2402
rect 4033 -2516 4067 -2482
rect 4183 -2356 4217 -2322
rect 4183 -2436 4217 -2402
rect 4183 -2516 4217 -2482
rect 4333 -2356 4367 -2322
rect 4333 -2436 4367 -2402
rect 4333 -2516 4367 -2482
rect 4483 -2356 4517 -2322
rect 4483 -2436 4517 -2402
rect 4483 -2516 4517 -2482
rect 4633 -2356 4667 -2322
rect 5913 -2356 5947 -2322
rect 4633 -2436 4667 -2402
rect 4633 -2516 4667 -2482
rect 5913 -2436 5947 -2402
rect 5913 -2516 5947 -2482
rect 6063 -2356 6097 -2322
rect 6063 -2436 6097 -2402
rect 6063 -2516 6097 -2482
rect 6213 -2356 6247 -2322
rect 6213 -2436 6247 -2402
rect 6213 -2516 6247 -2482
rect 6363 -2356 6397 -2322
rect 6363 -2436 6397 -2402
rect 6363 -2516 6397 -2482
rect 6513 -2356 6547 -2322
rect 6513 -2436 6547 -2402
rect 6513 -2516 6547 -2482
rect 1844 -3416 1878 -3382
rect 1844 -3496 1878 -3462
rect 1844 -3576 1878 -3542
rect 1994 -3416 2028 -3382
rect 1994 -3496 2028 -3462
rect 1994 -3576 2028 -3542
rect 2144 -3416 2178 -3382
rect 2144 -3496 2178 -3462
rect 2144 -3576 2178 -3542
rect 2294 -3416 2328 -3382
rect 2294 -3496 2328 -3462
rect 2294 -3576 2328 -3542
rect 2444 -3416 2478 -3382
rect 2444 -3496 2478 -3462
rect 2444 -3576 2478 -3542
rect 3894 -3416 3928 -3382
rect 3894 -3496 3928 -3462
rect 3894 -3576 3928 -3542
rect 4044 -3416 4078 -3382
rect 4044 -3496 4078 -3462
rect 4044 -3576 4078 -3542
rect 4194 -3416 4228 -3382
rect 4194 -3496 4228 -3462
rect 4194 -3576 4228 -3542
rect 4344 -3416 4378 -3382
rect 4344 -3496 4378 -3462
rect 4344 -3576 4378 -3542
rect 4494 -3416 4528 -3382
rect 4494 -3496 4528 -3462
rect 4494 -3576 4528 -3542
rect 5934 -3417 5968 -3383
rect 5934 -3497 5968 -3463
rect 5934 -3577 5968 -3543
rect 6084 -3417 6118 -3383
rect 6084 -3497 6118 -3463
rect 6084 -3577 6118 -3543
rect 6234 -3417 6268 -3383
rect 6234 -3497 6268 -3463
rect 6234 -3577 6268 -3543
rect 6384 -3417 6418 -3383
rect 6384 -3497 6418 -3463
rect 6384 -3577 6418 -3543
rect 6534 -3417 6568 -3383
rect 6534 -3497 6568 -3463
rect 6534 -3577 6568 -3543
rect 4094 -5257 4128 -5223
rect 4094 -5337 4128 -5303
rect 4094 -5417 4128 -5383
rect 4244 -5257 4278 -5223
rect 4244 -5337 4278 -5303
rect 4244 -5417 4278 -5383
rect 4394 -5257 4428 -5223
rect 4394 -5337 4428 -5303
rect 4394 -5417 4428 -5383
rect 4544 -5257 4578 -5223
rect 4544 -5337 4578 -5303
rect 4544 -5417 4578 -5383
rect 4694 -5257 4728 -5223
rect 4694 -5337 4728 -5303
rect 4694 -5417 4728 -5383
rect 6153 -5257 6187 -5223
rect 6153 -5337 6187 -5303
rect 6153 -5417 6187 -5383
rect 1883 -5576 1917 -5542
rect 1883 -5656 1917 -5622
rect 1883 -5736 1917 -5702
rect 2033 -5576 2067 -5542
rect 2033 -5656 2067 -5622
rect 2033 -5736 2067 -5702
rect 2183 -5576 2217 -5542
rect 2183 -5656 2217 -5622
rect 2183 -5736 2217 -5702
rect 2333 -5576 2367 -5542
rect 2333 -5656 2367 -5622
rect 2333 -5736 2367 -5702
rect 2483 -5576 2517 -5542
rect 6303 -5257 6337 -5223
rect 6303 -5337 6337 -5303
rect 6303 -5417 6337 -5383
rect 6453 -5257 6487 -5223
rect 6453 -5337 6487 -5303
rect 6453 -5417 6487 -5383
rect 6603 -5257 6637 -5223
rect 6603 -5337 6637 -5303
rect 6603 -5417 6637 -5383
rect 6753 -5257 6787 -5223
rect 6753 -5337 6787 -5303
rect 6753 -5417 6787 -5383
rect 2483 -5656 2517 -5622
rect 2483 -5736 2517 -5702
rect 1883 -6317 1917 -6283
rect 1883 -6397 1917 -6363
rect 1883 -6477 1917 -6443
rect 2033 -6317 2067 -6283
rect 2033 -6397 2067 -6363
rect 2033 -6477 2067 -6443
rect 2183 -6317 2217 -6283
rect 2183 -6397 2217 -6363
rect 2183 -6477 2217 -6443
rect 2333 -6317 2367 -6283
rect 2333 -6397 2367 -6363
rect 2333 -6477 2367 -6443
rect 2483 -6317 2517 -6283
rect 2483 -6397 2517 -6363
rect 2483 -6477 2517 -6443
rect 4093 -6317 4127 -6283
rect 4093 -6397 4127 -6363
rect 4093 -6477 4127 -6443
rect 4243 -6317 4277 -6283
rect 4243 -6397 4277 -6363
rect 4243 -6477 4277 -6443
rect 4393 -6317 4427 -6283
rect 4393 -6397 4427 -6363
rect 4393 -6477 4427 -6443
rect 4543 -6317 4577 -6283
rect 4543 -6397 4577 -6363
rect 4543 -6477 4577 -6443
rect 4693 -6317 4727 -6283
rect 4693 -6397 4727 -6363
rect 5972 -6317 6006 -6283
rect 5972 -6397 6006 -6363
rect 4693 -6477 4727 -6443
rect 5972 -6477 6006 -6443
rect 6122 -6317 6156 -6283
rect 6122 -6397 6156 -6363
rect 6122 -6477 6156 -6443
rect 6272 -6317 6306 -6283
rect 6272 -6397 6306 -6363
rect 6272 -6477 6306 -6443
rect 6422 -6317 6456 -6283
rect 6422 -6397 6456 -6363
rect 6422 -6477 6456 -6443
rect 6572 -6317 6606 -6283
rect 6572 -6397 6606 -6363
rect 6572 -6477 6606 -6443
rect 1883 -8077 1917 -8043
rect 1883 -8157 1917 -8123
rect 1883 -8237 1917 -8203
rect 2033 -8077 2067 -8043
rect 2033 -8157 2067 -8123
rect 2033 -8237 2067 -8203
rect 2183 -8077 2217 -8043
rect 2183 -8157 2217 -8123
rect 2183 -8237 2217 -8203
rect 2333 -8077 2367 -8043
rect 2333 -8157 2367 -8123
rect 2333 -8237 2367 -8203
rect 2483 -8077 2517 -8043
rect 2483 -8157 2517 -8123
rect 2483 -8237 2517 -8203
rect 4093 -8077 4127 -8043
rect 4093 -8157 4127 -8123
rect 4093 -8237 4127 -8203
rect 4243 -8077 4277 -8043
rect 4243 -8157 4277 -8123
rect 4243 -8237 4277 -8203
rect 4393 -8077 4427 -8043
rect 4393 -8157 4427 -8123
rect 4393 -8237 4427 -8203
rect 4543 -8077 4577 -8043
rect 4543 -8157 4577 -8123
rect 4543 -8237 4577 -8203
rect 4693 -8077 4727 -8043
rect 5972 -8077 6006 -8043
rect 4693 -8157 4727 -8123
rect 4693 -8237 4727 -8203
rect 5972 -8157 6006 -8123
rect 5972 -8237 6006 -8203
rect 6122 -8077 6156 -8043
rect 6122 -8157 6156 -8123
rect 6122 -8237 6156 -8203
rect 6272 -8077 6306 -8043
rect 6272 -8157 6306 -8123
rect 6272 -8237 6306 -8203
rect 6422 -8077 6456 -8043
rect 6422 -8157 6456 -8123
rect 6422 -8237 6456 -8203
rect 6572 -8077 6606 -8043
rect 6572 -8157 6606 -8123
rect 6572 -8237 6606 -8203
rect 1843 -9137 1877 -9103
rect 1843 -9217 1877 -9183
rect 1843 -9297 1877 -9263
rect 1993 -9137 2027 -9103
rect 1993 -9217 2027 -9183
rect 1993 -9297 2027 -9263
rect 2143 -9137 2177 -9103
rect 2143 -9217 2177 -9183
rect 2143 -9297 2177 -9263
rect 2293 -9137 2327 -9103
rect 2293 -9217 2327 -9183
rect 2293 -9297 2327 -9263
rect 2443 -9137 2477 -9103
rect 2443 -9217 2477 -9183
rect 2443 -9297 2477 -9263
rect 4033 -9137 4067 -9103
rect 4033 -9217 4067 -9183
rect 4033 -9297 4067 -9263
rect 4183 -9137 4217 -9103
rect 4183 -9217 4217 -9183
rect 4183 -9297 4217 -9263
rect 4333 -9137 4367 -9103
rect 4333 -9217 4367 -9183
rect 4333 -9297 4367 -9263
rect 4483 -9137 4517 -9103
rect 4483 -9217 4517 -9183
rect 4483 -9297 4517 -9263
rect 4633 -9137 4667 -9103
rect 4633 -9217 4667 -9183
rect 5913 -9137 5947 -9103
rect 5913 -9217 5947 -9183
rect 4633 -9297 4667 -9263
rect 5913 -9297 5947 -9263
rect 6063 -9137 6097 -9103
rect 6063 -9217 6097 -9183
rect 6063 -9297 6097 -9263
rect 6213 -9137 6247 -9103
rect 6213 -9217 6247 -9183
rect 6213 -9297 6247 -9263
rect 6363 -9137 6397 -9103
rect 6363 -9217 6397 -9183
rect 6363 -9297 6397 -9263
rect 6513 -9137 6547 -9103
rect 6513 -9217 6547 -9183
rect 6513 -9297 6547 -9263
rect 1843 -10897 1877 -10863
rect 1843 -10977 1877 -10943
rect 1843 -11057 1877 -11023
rect 1993 -10897 2027 -10863
rect 1993 -10977 2027 -10943
rect 1993 -11057 2027 -11023
rect 2143 -10897 2177 -10863
rect 2143 -10977 2177 -10943
rect 2143 -11057 2177 -11023
rect 2293 -10897 2327 -10863
rect 2293 -10977 2327 -10943
rect 2293 -11057 2327 -11023
rect 2443 -10897 2477 -10863
rect 2443 -10977 2477 -10943
rect 2443 -11057 2477 -11023
rect 4033 -10897 4067 -10863
rect 4033 -10977 4067 -10943
rect 4033 -11057 4067 -11023
rect 4183 -10897 4217 -10863
rect 4183 -10977 4217 -10943
rect 4183 -11057 4217 -11023
rect 4333 -10897 4367 -10863
rect 4333 -10977 4367 -10943
rect 4333 -11057 4367 -11023
rect 4483 -10897 4517 -10863
rect 4483 -10977 4517 -10943
rect 4483 -11057 4517 -11023
rect 4633 -10897 4667 -10863
rect 5913 -10897 5947 -10863
rect 4633 -10977 4667 -10943
rect 4633 -11057 4667 -11023
rect 5913 -10977 5947 -10943
rect 5913 -11057 5947 -11023
rect 6063 -10897 6097 -10863
rect 6063 -10977 6097 -10943
rect 6063 -11057 6097 -11023
rect 6213 -10897 6247 -10863
rect 6213 -10977 6247 -10943
rect 6213 -11057 6247 -11023
rect 6363 -10897 6397 -10863
rect 6363 -10977 6397 -10943
rect 6363 -11057 6397 -11023
rect 6513 -10897 6547 -10863
rect 6513 -10977 6547 -10943
rect 6513 -11057 6547 -11023
rect 1844 -11957 1878 -11923
rect 1844 -12037 1878 -12003
rect 1844 -12117 1878 -12083
rect 1994 -11957 2028 -11923
rect 1994 -12037 2028 -12003
rect 1994 -12117 2028 -12083
rect 2144 -11957 2178 -11923
rect 2144 -12037 2178 -12003
rect 2144 -12117 2178 -12083
rect 2294 -11957 2328 -11923
rect 2294 -12037 2328 -12003
rect 2294 -12117 2328 -12083
rect 2444 -11957 2478 -11923
rect 2444 -12037 2478 -12003
rect 2444 -12117 2478 -12083
rect 3894 -11957 3928 -11923
rect 3894 -12037 3928 -12003
rect 3894 -12117 3928 -12083
rect 4044 -11957 4078 -11923
rect 4044 -12037 4078 -12003
rect 4044 -12117 4078 -12083
rect 4194 -11957 4228 -11923
rect 4194 -12037 4228 -12003
rect 4194 -12117 4228 -12083
rect 4344 -11957 4378 -11923
rect 4344 -12037 4378 -12003
rect 4344 -12117 4378 -12083
rect 4494 -11957 4528 -11923
rect 4494 -12037 4528 -12003
rect 4494 -12117 4528 -12083
rect 5934 -11958 5968 -11924
rect 5934 -12038 5968 -12004
rect 5934 -12118 5968 -12084
rect 6084 -11958 6118 -11924
rect 6084 -12038 6118 -12004
rect 6084 -12118 6118 -12084
rect 6234 -11958 6268 -11924
rect 6234 -12038 6268 -12004
rect 6234 -12118 6268 -12084
rect 6384 -11958 6418 -11924
rect 6384 -12038 6418 -12004
rect 6384 -12118 6418 -12084
rect 6534 -11958 6568 -11924
rect 6534 -12038 6568 -12004
rect 6534 -12118 6568 -12084
<< psubdiff >>
rect 1020 1298 3300 1331
rect 1020 1264 1103 1298
rect 1137 1264 1183 1298
rect 1217 1264 1263 1298
rect 1297 1264 1343 1298
rect 1377 1264 1423 1298
rect 1457 1264 1503 1298
rect 1537 1264 1583 1298
rect 1617 1264 1663 1298
rect 1697 1264 1743 1298
rect 1777 1264 1823 1298
rect 1857 1264 1903 1298
rect 1937 1264 1983 1298
rect 2017 1264 2063 1298
rect 2097 1264 2143 1298
rect 2177 1264 2223 1298
rect 2257 1264 2303 1298
rect 2337 1264 2383 1298
rect 2417 1264 2463 1298
rect 2497 1264 2543 1298
rect 2577 1264 2623 1298
rect 2657 1264 2703 1298
rect 2737 1264 2783 1298
rect 2817 1264 2863 1298
rect 2897 1264 2943 1298
rect 2977 1264 3023 1298
rect 3057 1264 3103 1298
rect 3137 1264 3183 1298
rect 3217 1264 3300 1298
rect 1020 1231 3300 1264
rect 3640 1298 5320 1331
rect 3640 1264 3663 1298
rect 3697 1264 3743 1298
rect 3777 1264 3823 1298
rect 3857 1264 3903 1298
rect 3937 1264 3983 1298
rect 4017 1264 4063 1298
rect 4097 1264 4143 1298
rect 4177 1264 4223 1298
rect 4257 1264 4303 1298
rect 4337 1264 4383 1298
rect 4417 1264 4463 1298
rect 4497 1264 4543 1298
rect 4577 1264 4623 1298
rect 4657 1264 4703 1298
rect 4737 1264 4783 1298
rect 4817 1264 4863 1298
rect 4897 1264 4943 1298
rect 4977 1264 5023 1298
rect 5057 1264 5103 1298
rect 5137 1264 5183 1298
rect 5217 1264 5263 1298
rect 5297 1264 5320 1298
rect 3640 1231 5320 1264
rect 5660 1298 7340 1331
rect 5660 1264 5683 1298
rect 5717 1264 5763 1298
rect 5797 1264 5843 1298
rect 5877 1264 5923 1298
rect 5957 1264 6003 1298
rect 6037 1264 6083 1298
rect 6117 1264 6163 1298
rect 6197 1264 6243 1298
rect 6277 1264 6323 1298
rect 6357 1264 6403 1298
rect 6437 1264 6483 1298
rect 6517 1264 6563 1298
rect 6597 1264 6643 1298
rect 6677 1264 6723 1298
rect 6757 1264 6803 1298
rect 6837 1264 6883 1298
rect 6917 1264 6963 1298
rect 6997 1264 7043 1298
rect 7077 1264 7123 1298
rect 7157 1264 7203 1298
rect 7237 1264 7283 1298
rect 7317 1264 7340 1298
rect 5660 1231 7340 1264
rect 1020 -1522 3300 -1489
rect 1020 -1556 1103 -1522
rect 1137 -1556 1183 -1522
rect 1217 -1556 1263 -1522
rect 1297 -1556 1343 -1522
rect 1377 -1556 1423 -1522
rect 1457 -1556 1503 -1522
rect 1537 -1556 1583 -1522
rect 1617 -1556 1663 -1522
rect 1697 -1556 1743 -1522
rect 1777 -1556 1823 -1522
rect 1857 -1556 1903 -1522
rect 1937 -1556 1983 -1522
rect 2017 -1556 2063 -1522
rect 2097 -1556 2143 -1522
rect 2177 -1556 2223 -1522
rect 2257 -1556 2303 -1522
rect 2337 -1556 2383 -1522
rect 2417 -1556 2463 -1522
rect 2497 -1556 2543 -1522
rect 2577 -1556 2623 -1522
rect 2657 -1556 2703 -1522
rect 2737 -1556 2783 -1522
rect 2817 -1556 2863 -1522
rect 2897 -1556 2943 -1522
rect 2977 -1556 3023 -1522
rect 3057 -1556 3103 -1522
rect 3137 -1556 3183 -1522
rect 3217 -1556 3300 -1522
rect 1020 -1589 3300 -1556
rect 3660 -1522 5040 -1489
rect 3660 -1556 3693 -1522
rect 3727 -1556 3773 -1522
rect 3807 -1556 3853 -1522
rect 3887 -1556 3933 -1522
rect 3967 -1556 4013 -1522
rect 4047 -1556 4093 -1522
rect 4127 -1556 4173 -1522
rect 4207 -1556 4253 -1522
rect 4287 -1556 4333 -1522
rect 4367 -1556 4413 -1522
rect 4447 -1556 4493 -1522
rect 4527 -1556 4573 -1522
rect 4607 -1556 4653 -1522
rect 4687 -1556 4733 -1522
rect 4767 -1556 4813 -1522
rect 4847 -1556 4893 -1522
rect 4927 -1556 4973 -1522
rect 5007 -1556 5040 -1522
rect 3660 -1589 5040 -1556
rect 5390 -1522 7070 -1489
rect 5390 -1556 5413 -1522
rect 5447 -1556 5493 -1522
rect 5527 -1556 5573 -1522
rect 5607 -1556 5653 -1522
rect 5687 -1556 5733 -1522
rect 5767 -1556 5813 -1522
rect 5847 -1556 5893 -1522
rect 5927 -1556 5973 -1522
rect 6007 -1556 6053 -1522
rect 6087 -1556 6133 -1522
rect 6167 -1556 6213 -1522
rect 6247 -1556 6293 -1522
rect 6327 -1556 6373 -1522
rect 6407 -1556 6453 -1522
rect 6487 -1556 6533 -1522
rect 6567 -1556 6613 -1522
rect 6647 -1556 6693 -1522
rect 6727 -1556 6773 -1522
rect 6807 -1556 6853 -1522
rect 6887 -1556 6933 -1522
rect 6967 -1556 7013 -1522
rect 7047 -1556 7070 -1522
rect 5390 -1589 7070 -1556
rect 1161 -4342 3161 -4309
rect 1161 -4376 1184 -4342
rect 1218 -4376 1264 -4342
rect 1298 -4376 1344 -4342
rect 1378 -4376 1424 -4342
rect 1458 -4376 1504 -4342
rect 1538 -4376 1584 -4342
rect 1618 -4376 1664 -4342
rect 1698 -4376 1744 -4342
rect 1778 -4376 1824 -4342
rect 1858 -4376 1904 -4342
rect 1938 -4376 1984 -4342
rect 2018 -4376 2064 -4342
rect 2098 -4376 2144 -4342
rect 2178 -4376 2224 -4342
rect 2258 -4376 2304 -4342
rect 2338 -4376 2384 -4342
rect 2418 -4376 2464 -4342
rect 2498 -4376 2544 -4342
rect 2578 -4376 2624 -4342
rect 2658 -4376 2704 -4342
rect 2738 -4376 2784 -4342
rect 2818 -4376 2864 -4342
rect 2898 -4376 2944 -4342
rect 2978 -4376 3024 -4342
rect 3058 -4376 3104 -4342
rect 3138 -4376 3161 -4342
rect 1161 -4389 3161 -4376
rect 3521 -4342 4901 -4309
rect 3521 -4376 3554 -4342
rect 3588 -4376 3634 -4342
rect 3668 -4376 3714 -4342
rect 3748 -4376 3794 -4342
rect 3828 -4376 3874 -4342
rect 3908 -4376 3954 -4342
rect 3988 -4376 4034 -4342
rect 4068 -4376 4114 -4342
rect 4148 -4376 4194 -4342
rect 4228 -4376 4274 -4342
rect 4308 -4376 4354 -4342
rect 4388 -4376 4434 -4342
rect 4468 -4376 4514 -4342
rect 4548 -4376 4594 -4342
rect 4628 -4376 4674 -4342
rect 4708 -4376 4754 -4342
rect 4788 -4376 4834 -4342
rect 4868 -4376 4901 -4342
rect 1040 -4422 3360 -4389
rect 3521 -4390 4901 -4376
rect 5251 -4343 7251 -4310
rect 5251 -4377 5274 -4343
rect 5308 -4377 5354 -4343
rect 5388 -4377 5434 -4343
rect 5468 -4377 5514 -4343
rect 5548 -4377 5594 -4343
rect 5628 -4377 5674 -4343
rect 5708 -4377 5754 -4343
rect 5788 -4377 5834 -4343
rect 5868 -4377 5914 -4343
rect 5948 -4377 5994 -4343
rect 6028 -4377 6074 -4343
rect 6108 -4377 6154 -4343
rect 6188 -4377 6234 -4343
rect 6268 -4377 6314 -4343
rect 6348 -4377 6394 -4343
rect 6428 -4377 6474 -4343
rect 6508 -4377 6554 -4343
rect 6588 -4377 6634 -4343
rect 6668 -4377 6714 -4343
rect 6748 -4377 6794 -4343
rect 6828 -4377 6874 -4343
rect 6908 -4377 6954 -4343
rect 6988 -4377 7034 -4343
rect 7068 -4377 7114 -4343
rect 7148 -4377 7194 -4343
rect 7228 -4377 7251 -4343
rect 5251 -4390 7251 -4377
rect 3521 -4409 5101 -4390
rect 1040 -4456 1063 -4422
rect 1097 -4456 1143 -4422
rect 1177 -4456 1223 -4422
rect 1257 -4456 1303 -4422
rect 1337 -4456 1383 -4422
rect 1417 -4456 1463 -4422
rect 1497 -4456 1543 -4422
rect 1577 -4456 1623 -4422
rect 1657 -4456 1703 -4422
rect 1737 -4456 1783 -4422
rect 1817 -4456 1863 -4422
rect 1897 -4456 1943 -4422
rect 1977 -4456 2023 -4422
rect 2057 -4456 2103 -4422
rect 2137 -4456 2183 -4422
rect 2217 -4456 2263 -4422
rect 2297 -4456 2343 -4422
rect 2377 -4456 2423 -4422
rect 2457 -4456 2503 -4422
rect 2537 -4456 2583 -4422
rect 2617 -4456 2663 -4422
rect 2697 -4456 2743 -4422
rect 2777 -4456 2823 -4422
rect 2857 -4456 2903 -4422
rect 2937 -4456 2983 -4422
rect 3017 -4456 3063 -4422
rect 3097 -4456 3143 -4422
rect 3177 -4456 3223 -4422
rect 3257 -4456 3303 -4422
rect 3337 -4456 3360 -4422
rect 1040 -4489 3360 -4456
rect 3721 -4423 5101 -4409
rect 5251 -4410 7470 -4390
rect 3721 -4457 3754 -4423
rect 3788 -4457 3834 -4423
rect 3868 -4457 3914 -4423
rect 3948 -4457 3994 -4423
rect 4028 -4457 4074 -4423
rect 4108 -4457 4154 -4423
rect 4188 -4457 4234 -4423
rect 4268 -4457 4314 -4423
rect 4348 -4457 4394 -4423
rect 4428 -4457 4474 -4423
rect 4508 -4457 4554 -4423
rect 4588 -4457 4634 -4423
rect 4668 -4457 4714 -4423
rect 4748 -4457 4794 -4423
rect 4828 -4457 4874 -4423
rect 4908 -4457 4954 -4423
rect 4988 -4457 5034 -4423
rect 5068 -4457 5101 -4423
rect 3721 -4490 5101 -4457
rect 5470 -4423 7470 -4410
rect 5470 -4457 5493 -4423
rect 5527 -4457 5573 -4423
rect 5607 -4457 5653 -4423
rect 5687 -4457 5733 -4423
rect 5767 -4457 5813 -4423
rect 5847 -4457 5893 -4423
rect 5927 -4457 5973 -4423
rect 6007 -4457 6053 -4423
rect 6087 -4457 6133 -4423
rect 6167 -4457 6213 -4423
rect 6247 -4457 6293 -4423
rect 6327 -4457 6373 -4423
rect 6407 -4457 6453 -4423
rect 6487 -4457 6533 -4423
rect 6567 -4457 6613 -4423
rect 6647 -4457 6693 -4423
rect 6727 -4457 6773 -4423
rect 6807 -4457 6853 -4423
rect 6887 -4457 6933 -4423
rect 6967 -4457 7013 -4423
rect 7047 -4457 7093 -4423
rect 7127 -4457 7173 -4423
rect 7207 -4457 7253 -4423
rect 7287 -4457 7333 -4423
rect 7367 -4457 7413 -4423
rect 7447 -4457 7470 -4423
rect 5470 -4490 7470 -4457
rect 1060 -7243 3340 -7210
rect 1060 -7277 1143 -7243
rect 1177 -7277 1223 -7243
rect 1257 -7277 1303 -7243
rect 1337 -7277 1383 -7243
rect 1417 -7277 1463 -7243
rect 1497 -7277 1543 -7243
rect 1577 -7277 1623 -7243
rect 1657 -7277 1703 -7243
rect 1737 -7277 1783 -7243
rect 1817 -7277 1863 -7243
rect 1897 -7277 1943 -7243
rect 1977 -7277 2023 -7243
rect 2057 -7277 2103 -7243
rect 2137 -7277 2183 -7243
rect 2217 -7277 2263 -7243
rect 2297 -7277 2343 -7243
rect 2377 -7277 2423 -7243
rect 2457 -7277 2503 -7243
rect 2537 -7277 2583 -7243
rect 2617 -7277 2663 -7243
rect 2697 -7277 2743 -7243
rect 2777 -7277 2823 -7243
rect 2857 -7277 2903 -7243
rect 2937 -7277 2983 -7243
rect 3017 -7277 3063 -7243
rect 3097 -7277 3143 -7243
rect 3177 -7277 3223 -7243
rect 3257 -7277 3340 -7243
rect 1060 -7310 3340 -7277
rect 3720 -7243 5100 -7210
rect 3720 -7277 3753 -7243
rect 3787 -7277 3833 -7243
rect 3867 -7277 3913 -7243
rect 3947 -7277 3993 -7243
rect 4027 -7277 4073 -7243
rect 4107 -7277 4153 -7243
rect 4187 -7277 4233 -7243
rect 4267 -7277 4313 -7243
rect 4347 -7277 4393 -7243
rect 4427 -7277 4473 -7243
rect 4507 -7277 4553 -7243
rect 4587 -7277 4633 -7243
rect 4667 -7277 4713 -7243
rect 4747 -7277 4793 -7243
rect 4827 -7277 4873 -7243
rect 4907 -7277 4953 -7243
rect 4987 -7277 5033 -7243
rect 5067 -7277 5100 -7243
rect 3720 -7310 5100 -7277
rect 5449 -7243 7129 -7210
rect 5449 -7277 5472 -7243
rect 5506 -7277 5552 -7243
rect 5586 -7277 5632 -7243
rect 5666 -7277 5712 -7243
rect 5746 -7277 5792 -7243
rect 5826 -7277 5872 -7243
rect 5906 -7277 5952 -7243
rect 5986 -7277 6032 -7243
rect 6066 -7277 6112 -7243
rect 6146 -7277 6192 -7243
rect 6226 -7277 6272 -7243
rect 6306 -7277 6352 -7243
rect 6386 -7277 6432 -7243
rect 6466 -7277 6512 -7243
rect 6546 -7277 6592 -7243
rect 6626 -7277 6672 -7243
rect 6706 -7277 6752 -7243
rect 6786 -7277 6832 -7243
rect 6866 -7277 6912 -7243
rect 6946 -7277 6992 -7243
rect 7026 -7277 7072 -7243
rect 7106 -7277 7129 -7243
rect 5449 -7310 7129 -7277
rect 1020 -10063 3300 -10030
rect 1020 -10097 1103 -10063
rect 1137 -10097 1183 -10063
rect 1217 -10097 1263 -10063
rect 1297 -10097 1343 -10063
rect 1377 -10097 1423 -10063
rect 1457 -10097 1503 -10063
rect 1537 -10097 1583 -10063
rect 1617 -10097 1663 -10063
rect 1697 -10097 1743 -10063
rect 1777 -10097 1823 -10063
rect 1857 -10097 1903 -10063
rect 1937 -10097 1983 -10063
rect 2017 -10097 2063 -10063
rect 2097 -10097 2143 -10063
rect 2177 -10097 2223 -10063
rect 2257 -10097 2303 -10063
rect 2337 -10097 2383 -10063
rect 2417 -10097 2463 -10063
rect 2497 -10097 2543 -10063
rect 2577 -10097 2623 -10063
rect 2657 -10097 2703 -10063
rect 2737 -10097 2783 -10063
rect 2817 -10097 2863 -10063
rect 2897 -10097 2943 -10063
rect 2977 -10097 3023 -10063
rect 3057 -10097 3103 -10063
rect 3137 -10097 3183 -10063
rect 3217 -10097 3300 -10063
rect 1020 -10130 3300 -10097
rect 3660 -10063 5040 -10030
rect 3660 -10097 3693 -10063
rect 3727 -10097 3773 -10063
rect 3807 -10097 3853 -10063
rect 3887 -10097 3933 -10063
rect 3967 -10097 4013 -10063
rect 4047 -10097 4093 -10063
rect 4127 -10097 4173 -10063
rect 4207 -10097 4253 -10063
rect 4287 -10097 4333 -10063
rect 4367 -10097 4413 -10063
rect 4447 -10097 4493 -10063
rect 4527 -10097 4573 -10063
rect 4607 -10097 4653 -10063
rect 4687 -10097 4733 -10063
rect 4767 -10097 4813 -10063
rect 4847 -10097 4893 -10063
rect 4927 -10097 4973 -10063
rect 5007 -10097 5040 -10063
rect 3660 -10130 5040 -10097
rect 5390 -10063 7070 -10030
rect 5390 -10097 5413 -10063
rect 5447 -10097 5493 -10063
rect 5527 -10097 5573 -10063
rect 5607 -10097 5653 -10063
rect 5687 -10097 5733 -10063
rect 5767 -10097 5813 -10063
rect 5847 -10097 5893 -10063
rect 5927 -10097 5973 -10063
rect 6007 -10097 6053 -10063
rect 6087 -10097 6133 -10063
rect 6167 -10097 6213 -10063
rect 6247 -10097 6293 -10063
rect 6327 -10097 6373 -10063
rect 6407 -10097 6453 -10063
rect 6487 -10097 6533 -10063
rect 6567 -10097 6613 -10063
rect 6647 -10097 6693 -10063
rect 6727 -10097 6773 -10063
rect 6807 -10097 6853 -10063
rect 6887 -10097 6933 -10063
rect 6967 -10097 7013 -10063
rect 7047 -10097 7070 -10063
rect 5390 -10130 7070 -10097
rect 1161 -12883 3161 -12850
rect 1161 -12917 1184 -12883
rect 1218 -12917 1264 -12883
rect 1298 -12917 1344 -12883
rect 1378 -12917 1424 -12883
rect 1458 -12917 1504 -12883
rect 1538 -12917 1584 -12883
rect 1618 -12917 1664 -12883
rect 1698 -12917 1744 -12883
rect 1778 -12917 1824 -12883
rect 1858 -12917 1904 -12883
rect 1938 -12917 1984 -12883
rect 2018 -12917 2064 -12883
rect 2098 -12917 2144 -12883
rect 2178 -12917 2224 -12883
rect 2258 -12917 2304 -12883
rect 2338 -12917 2384 -12883
rect 2418 -12917 2464 -12883
rect 2498 -12917 2544 -12883
rect 2578 -12917 2624 -12883
rect 2658 -12917 2704 -12883
rect 2738 -12917 2784 -12883
rect 2818 -12917 2864 -12883
rect 2898 -12917 2944 -12883
rect 2978 -12917 3024 -12883
rect 3058 -12917 3104 -12883
rect 3138 -12917 3161 -12883
rect 1161 -12950 3161 -12917
rect 3521 -12883 4901 -12850
rect 3521 -12917 3554 -12883
rect 3588 -12917 3634 -12883
rect 3668 -12917 3714 -12883
rect 3748 -12917 3794 -12883
rect 3828 -12917 3874 -12883
rect 3908 -12917 3954 -12883
rect 3988 -12917 4034 -12883
rect 4068 -12917 4114 -12883
rect 4148 -12917 4194 -12883
rect 4228 -12917 4274 -12883
rect 4308 -12917 4354 -12883
rect 4388 -12917 4434 -12883
rect 4468 -12917 4514 -12883
rect 4548 -12917 4594 -12883
rect 4628 -12917 4674 -12883
rect 4708 -12917 4754 -12883
rect 4788 -12917 4834 -12883
rect 4868 -12917 4901 -12883
rect 3521 -12950 4901 -12917
rect 5251 -12884 7251 -12851
rect 5251 -12918 5274 -12884
rect 5308 -12918 5354 -12884
rect 5388 -12918 5434 -12884
rect 5468 -12918 5514 -12884
rect 5548 -12918 5594 -12884
rect 5628 -12918 5674 -12884
rect 5708 -12918 5754 -12884
rect 5788 -12918 5834 -12884
rect 5868 -12918 5914 -12884
rect 5948 -12918 5994 -12884
rect 6028 -12918 6074 -12884
rect 6108 -12918 6154 -12884
rect 6188 -12918 6234 -12884
rect 6268 -12918 6314 -12884
rect 6348 -12918 6394 -12884
rect 6428 -12918 6474 -12884
rect 6508 -12918 6554 -12884
rect 6588 -12918 6634 -12884
rect 6668 -12918 6714 -12884
rect 6748 -12918 6794 -12884
rect 6828 -12918 6874 -12884
rect 6908 -12918 6954 -12884
rect 6988 -12918 7034 -12884
rect 7068 -12918 7114 -12884
rect 7148 -12918 7194 -12884
rect 7228 -12918 7251 -12884
rect 5251 -12951 7251 -12918
<< nsubdiff >>
rect 1020 2478 3300 2511
rect 1020 2444 1103 2478
rect 1137 2444 1183 2478
rect 1217 2444 1263 2478
rect 1297 2444 1343 2478
rect 1377 2444 1423 2478
rect 1457 2444 1503 2478
rect 1537 2444 1583 2478
rect 1617 2444 1663 2478
rect 1697 2444 1743 2478
rect 1777 2444 1823 2478
rect 1857 2444 1903 2478
rect 1937 2444 1983 2478
rect 2017 2444 2063 2478
rect 2097 2444 2143 2478
rect 2177 2444 2223 2478
rect 2257 2444 2303 2478
rect 2337 2444 2383 2478
rect 2417 2444 2463 2478
rect 2497 2444 2543 2478
rect 2577 2444 2623 2478
rect 2657 2444 2703 2478
rect 2737 2444 2783 2478
rect 2817 2444 2863 2478
rect 2897 2444 2943 2478
rect 2977 2444 3023 2478
rect 3057 2444 3103 2478
rect 3137 2444 3183 2478
rect 3217 2444 3300 2478
rect 1020 2411 3300 2444
rect 3640 2478 5320 2511
rect 3640 2444 3663 2478
rect 3697 2444 3743 2478
rect 3777 2444 3823 2478
rect 3857 2444 3903 2478
rect 3937 2444 3983 2478
rect 4017 2444 4063 2478
rect 4097 2444 4143 2478
rect 4177 2444 4223 2478
rect 4257 2444 4303 2478
rect 4337 2444 4383 2478
rect 4417 2444 4463 2478
rect 4497 2444 4543 2478
rect 4577 2444 4623 2478
rect 4657 2444 4703 2478
rect 4737 2444 4783 2478
rect 4817 2444 4863 2478
rect 4897 2444 4943 2478
rect 4977 2444 5023 2478
rect 5057 2444 5103 2478
rect 5137 2444 5183 2478
rect 5217 2444 5263 2478
rect 5297 2444 5320 2478
rect 3640 2411 5320 2444
rect 5660 2478 7340 2511
rect 5660 2444 5683 2478
rect 5717 2444 5763 2478
rect 5797 2444 5843 2478
rect 5877 2444 5923 2478
rect 5957 2444 6003 2478
rect 6037 2444 6083 2478
rect 6117 2444 6163 2478
rect 6197 2444 6243 2478
rect 6277 2444 6323 2478
rect 6357 2444 6403 2478
rect 6437 2444 6483 2478
rect 6517 2444 6563 2478
rect 6597 2444 6643 2478
rect 6677 2444 6723 2478
rect 6757 2444 6803 2478
rect 6837 2444 6883 2478
rect 6917 2444 6963 2478
rect 6997 2444 7043 2478
rect 7077 2444 7123 2478
rect 7157 2444 7203 2478
rect 7237 2444 7283 2478
rect 7317 2444 7340 2478
rect 5660 2411 7340 2444
rect 1320 118 3000 151
rect 1320 84 1343 118
rect 1377 84 1423 118
rect 1457 84 1503 118
rect 1537 84 1583 118
rect 1617 84 1663 118
rect 1697 84 1743 118
rect 1777 84 1823 118
rect 1857 84 1903 118
rect 1937 84 1983 118
rect 2017 84 2063 118
rect 2097 84 2143 118
rect 2177 84 2223 118
rect 2257 84 2303 118
rect 2337 84 2383 118
rect 2417 84 2463 118
rect 2497 84 2543 118
rect 2577 84 2623 118
rect 2657 84 2703 118
rect 2737 84 2783 118
rect 2817 84 2863 118
rect 2897 84 2943 118
rect 2977 84 3000 118
rect 1320 51 3000 84
rect 3640 118 5320 151
rect 3640 84 3663 118
rect 3697 84 3743 118
rect 3777 84 3823 118
rect 3857 84 3903 118
rect 3937 84 3983 118
rect 4017 84 4063 118
rect 4097 84 4143 118
rect 4177 84 4223 118
rect 4257 84 4303 118
rect 4337 84 4383 118
rect 4417 84 4463 118
rect 4497 84 4543 118
rect 4577 84 4623 118
rect 4657 84 4703 118
rect 4737 84 4783 118
rect 4817 84 4863 118
rect 4897 84 4943 118
rect 4977 84 5023 118
rect 5057 84 5103 118
rect 5137 84 5183 118
rect 5217 84 5263 118
rect 5297 84 5320 118
rect 3640 51 5320 84
rect 5660 118 7340 151
rect 5660 84 5683 118
rect 5717 84 5763 118
rect 5797 84 5843 118
rect 5877 84 5923 118
rect 5957 84 6003 118
rect 6037 84 6083 118
rect 6117 84 6163 118
rect 6197 84 6243 118
rect 6277 84 6323 118
rect 6357 84 6403 118
rect 6437 84 6483 118
rect 6517 84 6563 118
rect 6597 84 6643 118
rect 6677 84 6723 118
rect 6757 84 6803 118
rect 6837 84 6883 118
rect 6917 84 6963 118
rect 6997 84 7043 118
rect 7077 84 7123 118
rect 7157 84 7203 118
rect 7237 84 7283 118
rect 7317 84 7340 118
rect 5660 51 7340 84
rect 1020 -342 3300 -309
rect 1020 -376 1103 -342
rect 1137 -376 1183 -342
rect 1217 -376 1263 -342
rect 1297 -376 1343 -342
rect 1377 -376 1423 -342
rect 1457 -376 1503 -342
rect 1537 -376 1583 -342
rect 1617 -376 1663 -342
rect 1697 -376 1743 -342
rect 1777 -376 1823 -342
rect 1857 -376 1903 -342
rect 1937 -376 1983 -342
rect 2017 -376 2063 -342
rect 2097 -376 2143 -342
rect 2177 -376 2223 -342
rect 2257 -376 2303 -342
rect 2337 -376 2383 -342
rect 2417 -376 2463 -342
rect 2497 -376 2543 -342
rect 2577 -376 2623 -342
rect 2657 -376 2703 -342
rect 2737 -376 2783 -342
rect 2817 -376 2863 -342
rect 2897 -376 2943 -342
rect 2977 -376 3023 -342
rect 3057 -376 3103 -342
rect 3137 -376 3183 -342
rect 3217 -376 3300 -342
rect 1020 -409 3300 -376
rect 3660 -342 5040 -309
rect 3660 -376 3693 -342
rect 3727 -376 3773 -342
rect 3807 -376 3853 -342
rect 3887 -376 3933 -342
rect 3967 -376 4013 -342
rect 4047 -376 4093 -342
rect 4127 -376 4173 -342
rect 4207 -376 4253 -342
rect 4287 -376 4333 -342
rect 4367 -376 4413 -342
rect 4447 -376 4493 -342
rect 4527 -376 4573 -342
rect 4607 -376 4653 -342
rect 4687 -376 4733 -342
rect 4767 -376 4813 -342
rect 4847 -376 4893 -342
rect 4927 -376 4973 -342
rect 5007 -376 5040 -342
rect 3660 -409 5040 -376
rect 5390 -342 7070 -309
rect 5390 -376 5413 -342
rect 5447 -376 5493 -342
rect 5527 -376 5573 -342
rect 5607 -376 5653 -342
rect 5687 -376 5733 -342
rect 5767 -376 5813 -342
rect 5847 -376 5893 -342
rect 5927 -376 5973 -342
rect 6007 -376 6053 -342
rect 6087 -376 6133 -342
rect 6167 -376 6213 -342
rect 6247 -376 6293 -342
rect 6327 -376 6373 -342
rect 6407 -376 6453 -342
rect 6487 -376 6533 -342
rect 6567 -376 6613 -342
rect 6647 -376 6693 -342
rect 6727 -376 6773 -342
rect 6807 -376 6853 -342
rect 6887 -376 6933 -342
rect 6967 -376 7013 -342
rect 7047 -376 7070 -342
rect 5390 -409 7070 -376
rect 1020 -2702 3300 -2669
rect 1020 -2736 1103 -2702
rect 1137 -2736 1183 -2702
rect 1217 -2736 1263 -2702
rect 1297 -2736 1343 -2702
rect 1377 -2736 1423 -2702
rect 1457 -2736 1503 -2702
rect 1537 -2736 1583 -2702
rect 1617 -2736 1663 -2702
rect 1697 -2736 1743 -2702
rect 1777 -2736 1823 -2702
rect 1857 -2736 1903 -2702
rect 1937 -2736 1983 -2702
rect 2017 -2736 2063 -2702
rect 2097 -2736 2143 -2702
rect 2177 -2736 2223 -2702
rect 2257 -2736 2303 -2702
rect 2337 -2736 2383 -2702
rect 2417 -2736 2463 -2702
rect 2497 -2736 2543 -2702
rect 2577 -2736 2623 -2702
rect 2657 -2736 2703 -2702
rect 2737 -2736 2783 -2702
rect 2817 -2736 2863 -2702
rect 2897 -2736 2943 -2702
rect 2977 -2736 3023 -2702
rect 3057 -2736 3103 -2702
rect 3137 -2736 3183 -2702
rect 3217 -2736 3300 -2702
rect 1020 -2769 3300 -2736
rect 3660 -2702 5040 -2669
rect 3660 -2736 3693 -2702
rect 3727 -2736 3773 -2702
rect 3807 -2736 3853 -2702
rect 3887 -2736 3933 -2702
rect 3967 -2736 4013 -2702
rect 4047 -2736 4093 -2702
rect 4127 -2736 4173 -2702
rect 4207 -2736 4253 -2702
rect 4287 -2736 4333 -2702
rect 4367 -2736 4413 -2702
rect 4447 -2736 4493 -2702
rect 4527 -2736 4573 -2702
rect 4607 -2736 4653 -2702
rect 4687 -2736 4733 -2702
rect 4767 -2736 4813 -2702
rect 4847 -2736 4893 -2702
rect 4927 -2736 4973 -2702
rect 5007 -2736 5040 -2702
rect 3660 -2769 5040 -2736
rect 5390 -2702 7070 -2669
rect 5390 -2736 5413 -2702
rect 5447 -2736 5493 -2702
rect 5527 -2736 5573 -2702
rect 5607 -2736 5653 -2702
rect 5687 -2736 5733 -2702
rect 5767 -2736 5813 -2702
rect 5847 -2736 5893 -2702
rect 5927 -2736 5973 -2702
rect 6007 -2736 6053 -2702
rect 6087 -2736 6133 -2702
rect 6167 -2736 6213 -2702
rect 6247 -2736 6293 -2702
rect 6327 -2736 6373 -2702
rect 6407 -2736 6453 -2702
rect 6487 -2736 6533 -2702
rect 6567 -2736 6613 -2702
rect 6647 -2736 6693 -2702
rect 6727 -2736 6773 -2702
rect 6807 -2736 6853 -2702
rect 6887 -2736 6933 -2702
rect 6967 -2736 7013 -2702
rect 7047 -2736 7070 -2702
rect 5390 -2769 7070 -2736
rect 1161 -3162 3161 -3129
rect 1161 -3196 1184 -3162
rect 1218 -3196 1264 -3162
rect 1298 -3196 1344 -3162
rect 1378 -3196 1424 -3162
rect 1458 -3196 1504 -3162
rect 1538 -3196 1584 -3162
rect 1618 -3196 1664 -3162
rect 1698 -3196 1744 -3162
rect 1778 -3196 1824 -3162
rect 1858 -3196 1904 -3162
rect 1938 -3196 1984 -3162
rect 2018 -3196 2064 -3162
rect 2098 -3196 2144 -3162
rect 2178 -3196 2224 -3162
rect 2258 -3196 2304 -3162
rect 2338 -3196 2384 -3162
rect 2418 -3196 2464 -3162
rect 2498 -3196 2544 -3162
rect 2578 -3196 2624 -3162
rect 2658 -3196 2704 -3162
rect 2738 -3196 2784 -3162
rect 2818 -3196 2864 -3162
rect 2898 -3196 2944 -3162
rect 2978 -3196 3024 -3162
rect 3058 -3196 3104 -3162
rect 3138 -3196 3161 -3162
rect 1161 -3229 3161 -3196
rect 3521 -3162 4901 -3129
rect 3521 -3196 3554 -3162
rect 3588 -3196 3634 -3162
rect 3668 -3196 3714 -3162
rect 3748 -3196 3794 -3162
rect 3828 -3196 3874 -3162
rect 3908 -3196 3954 -3162
rect 3988 -3196 4034 -3162
rect 4068 -3196 4114 -3162
rect 4148 -3196 4194 -3162
rect 4228 -3196 4274 -3162
rect 4308 -3196 4354 -3162
rect 4388 -3196 4434 -3162
rect 4468 -3196 4514 -3162
rect 4548 -3196 4594 -3162
rect 4628 -3196 4674 -3162
rect 4708 -3196 4754 -3162
rect 4788 -3196 4834 -3162
rect 4868 -3196 4901 -3162
rect 3521 -3229 4901 -3196
rect 5251 -3163 7251 -3130
rect 5251 -3197 5274 -3163
rect 5308 -3197 5354 -3163
rect 5388 -3197 5434 -3163
rect 5468 -3197 5514 -3163
rect 5548 -3197 5594 -3163
rect 5628 -3197 5674 -3163
rect 5708 -3197 5754 -3163
rect 5788 -3197 5834 -3163
rect 5868 -3197 5914 -3163
rect 5948 -3197 5994 -3163
rect 6028 -3197 6074 -3163
rect 6108 -3197 6154 -3163
rect 6188 -3197 6234 -3163
rect 6268 -3197 6314 -3163
rect 6348 -3197 6394 -3163
rect 6428 -3197 6474 -3163
rect 6508 -3197 6554 -3163
rect 6588 -3197 6634 -3163
rect 6668 -3197 6714 -3163
rect 6748 -3197 6794 -3163
rect 6828 -3197 6874 -3163
rect 6908 -3197 6954 -3163
rect 6988 -3197 7034 -3163
rect 7068 -3197 7114 -3163
rect 7148 -3197 7194 -3163
rect 7228 -3197 7251 -3163
rect 5251 -3230 7251 -3197
rect 3721 -5603 5101 -5570
rect 3721 -5637 3754 -5603
rect 3788 -5637 3834 -5603
rect 3868 -5637 3914 -5603
rect 3948 -5637 3994 -5603
rect 4028 -5637 4074 -5603
rect 4108 -5637 4154 -5603
rect 4188 -5637 4234 -5603
rect 4268 -5637 4314 -5603
rect 4348 -5637 4394 -5603
rect 4428 -5637 4474 -5603
rect 4508 -5637 4554 -5603
rect 4588 -5637 4634 -5603
rect 4668 -5637 4714 -5603
rect 4748 -5637 4794 -5603
rect 4828 -5637 4874 -5603
rect 4908 -5637 4954 -5603
rect 4988 -5637 5034 -5603
rect 5068 -5637 5101 -5603
rect 3721 -5670 5101 -5637
rect 5470 -5603 7470 -5570
rect 5470 -5637 5493 -5603
rect 5527 -5637 5573 -5603
rect 5607 -5637 5653 -5603
rect 5687 -5637 5733 -5603
rect 5767 -5637 5813 -5603
rect 5847 -5637 5893 -5603
rect 5927 -5637 5973 -5603
rect 6007 -5637 6053 -5603
rect 6087 -5637 6133 -5603
rect 6167 -5637 6213 -5603
rect 6247 -5637 6293 -5603
rect 6327 -5637 6373 -5603
rect 6407 -5637 6453 -5603
rect 6487 -5637 6533 -5603
rect 6567 -5637 6613 -5603
rect 6647 -5637 6693 -5603
rect 6727 -5637 6773 -5603
rect 6807 -5637 6853 -5603
rect 6887 -5637 6933 -5603
rect 6967 -5637 7013 -5603
rect 7047 -5637 7093 -5603
rect 7127 -5637 7173 -5603
rect 7207 -5637 7253 -5603
rect 7287 -5637 7333 -5603
rect 7367 -5637 7413 -5603
rect 7447 -5637 7470 -5603
rect 5470 -5670 7470 -5637
rect 1040 -5922 3360 -5889
rect 1040 -5956 1063 -5922
rect 1097 -5956 1143 -5922
rect 1177 -5956 1223 -5922
rect 1257 -5956 1303 -5922
rect 1337 -5956 1383 -5922
rect 1417 -5956 1463 -5922
rect 1497 -5956 1543 -5922
rect 1577 -5956 1623 -5922
rect 1657 -5956 1703 -5922
rect 1737 -5956 1783 -5922
rect 1817 -5956 1863 -5922
rect 1897 -5956 1943 -5922
rect 1977 -5956 2023 -5922
rect 2057 -5956 2103 -5922
rect 2137 -5956 2183 -5922
rect 2217 -5956 2263 -5922
rect 2297 -5956 2343 -5922
rect 2377 -5956 2423 -5922
rect 2457 -5956 2503 -5922
rect 2537 -5956 2583 -5922
rect 2617 -5956 2663 -5922
rect 2697 -5956 2743 -5922
rect 2777 -5956 2823 -5922
rect 2857 -5956 2903 -5922
rect 2937 -5956 2983 -5922
rect 3017 -5956 3063 -5922
rect 3097 -5956 3143 -5922
rect 3177 -5956 3223 -5922
rect 3257 -5956 3303 -5922
rect 3337 -5956 3360 -5922
rect 1040 -6063 3360 -5956
rect 1040 -6097 1063 -6063
rect 1097 -6097 1143 -6063
rect 1177 -6097 1223 -6063
rect 1257 -6097 1303 -6063
rect 1337 -6097 1383 -6063
rect 1417 -6097 1463 -6063
rect 1497 -6097 1543 -6063
rect 1577 -6097 1623 -6063
rect 1657 -6097 1703 -6063
rect 1737 -6097 1783 -6063
rect 1817 -6097 1863 -6063
rect 1897 -6097 1943 -6063
rect 1977 -6097 2023 -6063
rect 2057 -6097 2103 -6063
rect 2137 -6097 2183 -6063
rect 2217 -6097 2263 -6063
rect 2297 -6097 2343 -6063
rect 2377 -6097 2423 -6063
rect 2457 -6097 2503 -6063
rect 2537 -6097 2583 -6063
rect 2617 -6097 2663 -6063
rect 2697 -6097 2743 -6063
rect 2777 -6097 2823 -6063
rect 2857 -6097 2903 -6063
rect 2937 -6097 2983 -6063
rect 3017 -6097 3063 -6063
rect 3097 -6097 3143 -6063
rect 3177 -6097 3223 -6063
rect 3257 -6097 3303 -6063
rect 3337 -6097 3360 -6063
rect 1040 -6130 3360 -6097
rect 3720 -6063 5100 -6030
rect 3720 -6097 3753 -6063
rect 3787 -6097 3833 -6063
rect 3867 -6097 3913 -6063
rect 3947 -6097 3993 -6063
rect 4027 -6097 4073 -6063
rect 4107 -6097 4153 -6063
rect 4187 -6097 4233 -6063
rect 4267 -6097 4313 -6063
rect 4347 -6097 4393 -6063
rect 4427 -6097 4473 -6063
rect 4507 -6097 4553 -6063
rect 4587 -6097 4633 -6063
rect 4667 -6097 4713 -6063
rect 4747 -6097 4793 -6063
rect 4827 -6097 4873 -6063
rect 4907 -6097 4953 -6063
rect 4987 -6097 5033 -6063
rect 5067 -6097 5100 -6063
rect 3720 -6130 5100 -6097
rect 5449 -6063 7129 -6030
rect 5449 -6097 5472 -6063
rect 5506 -6097 5552 -6063
rect 5586 -6097 5632 -6063
rect 5666 -6097 5712 -6063
rect 5746 -6097 5792 -6063
rect 5826 -6097 5872 -6063
rect 5906 -6097 5952 -6063
rect 5986 -6097 6032 -6063
rect 6066 -6097 6112 -6063
rect 6146 -6097 6192 -6063
rect 6226 -6097 6272 -6063
rect 6306 -6097 6352 -6063
rect 6386 -6097 6432 -6063
rect 6466 -6097 6512 -6063
rect 6546 -6097 6592 -6063
rect 6626 -6097 6672 -6063
rect 6706 -6097 6752 -6063
rect 6786 -6097 6832 -6063
rect 6866 -6097 6912 -6063
rect 6946 -6097 6992 -6063
rect 7026 -6097 7072 -6063
rect 7106 -6097 7129 -6063
rect 5449 -6130 7129 -6097
rect 1060 -8423 3340 -8390
rect 1060 -8457 1143 -8423
rect 1177 -8457 1223 -8423
rect 1257 -8457 1303 -8423
rect 1337 -8457 1383 -8423
rect 1417 -8457 1463 -8423
rect 1497 -8457 1543 -8423
rect 1577 -8457 1623 -8423
rect 1657 -8457 1703 -8423
rect 1737 -8457 1783 -8423
rect 1817 -8457 1863 -8423
rect 1897 -8457 1943 -8423
rect 1977 -8457 2023 -8423
rect 2057 -8457 2103 -8423
rect 2137 -8457 2183 -8423
rect 2217 -8457 2263 -8423
rect 2297 -8457 2343 -8423
rect 2377 -8457 2423 -8423
rect 2457 -8457 2503 -8423
rect 2537 -8457 2583 -8423
rect 2617 -8457 2663 -8423
rect 2697 -8457 2743 -8423
rect 2777 -8457 2823 -8423
rect 2857 -8457 2903 -8423
rect 2937 -8457 2983 -8423
rect 3017 -8457 3063 -8423
rect 3097 -8457 3143 -8423
rect 3177 -8457 3223 -8423
rect 3257 -8457 3340 -8423
rect 1060 -8490 3340 -8457
rect 3720 -8423 5100 -8390
rect 3720 -8457 3753 -8423
rect 3787 -8457 3833 -8423
rect 3867 -8457 3913 -8423
rect 3947 -8457 3993 -8423
rect 4027 -8457 4073 -8423
rect 4107 -8457 4153 -8423
rect 4187 -8457 4233 -8423
rect 4267 -8457 4313 -8423
rect 4347 -8457 4393 -8423
rect 4427 -8457 4473 -8423
rect 4507 -8457 4553 -8423
rect 4587 -8457 4633 -8423
rect 4667 -8457 4713 -8423
rect 4747 -8457 4793 -8423
rect 4827 -8457 4873 -8423
rect 4907 -8457 4953 -8423
rect 4987 -8457 5033 -8423
rect 5067 -8457 5100 -8423
rect 3720 -8490 5100 -8457
rect 5449 -8423 7129 -8390
rect 5449 -8457 5472 -8423
rect 5506 -8457 5552 -8423
rect 5586 -8457 5632 -8423
rect 5666 -8457 5712 -8423
rect 5746 -8457 5792 -8423
rect 5826 -8457 5872 -8423
rect 5906 -8457 5952 -8423
rect 5986 -8457 6032 -8423
rect 6066 -8457 6112 -8423
rect 6146 -8457 6192 -8423
rect 6226 -8457 6272 -8423
rect 6306 -8457 6352 -8423
rect 6386 -8457 6432 -8423
rect 6466 -8457 6512 -8423
rect 6546 -8457 6592 -8423
rect 6626 -8457 6672 -8423
rect 6706 -8457 6752 -8423
rect 6786 -8457 6832 -8423
rect 6866 -8457 6912 -8423
rect 6946 -8457 6992 -8423
rect 7026 -8457 7072 -8423
rect 7106 -8457 7129 -8423
rect 5449 -8490 7129 -8457
rect 1020 -8883 3300 -8850
rect 1020 -8917 1103 -8883
rect 1137 -8917 1183 -8883
rect 1217 -8917 1263 -8883
rect 1297 -8917 1343 -8883
rect 1377 -8917 1423 -8883
rect 1457 -8917 1503 -8883
rect 1537 -8917 1583 -8883
rect 1617 -8917 1663 -8883
rect 1697 -8917 1743 -8883
rect 1777 -8917 1823 -8883
rect 1857 -8917 1903 -8883
rect 1937 -8917 1983 -8883
rect 2017 -8917 2063 -8883
rect 2097 -8917 2143 -8883
rect 2177 -8917 2223 -8883
rect 2257 -8917 2303 -8883
rect 2337 -8917 2383 -8883
rect 2417 -8917 2463 -8883
rect 2497 -8917 2543 -8883
rect 2577 -8917 2623 -8883
rect 2657 -8917 2703 -8883
rect 2737 -8917 2783 -8883
rect 2817 -8917 2863 -8883
rect 2897 -8917 2943 -8883
rect 2977 -8917 3023 -8883
rect 3057 -8917 3103 -8883
rect 3137 -8917 3183 -8883
rect 3217 -8917 3300 -8883
rect 1020 -8950 3300 -8917
rect 3660 -8883 5040 -8850
rect 3660 -8917 3693 -8883
rect 3727 -8917 3773 -8883
rect 3807 -8917 3853 -8883
rect 3887 -8917 3933 -8883
rect 3967 -8917 4013 -8883
rect 4047 -8917 4093 -8883
rect 4127 -8917 4173 -8883
rect 4207 -8917 4253 -8883
rect 4287 -8917 4333 -8883
rect 4367 -8917 4413 -8883
rect 4447 -8917 4493 -8883
rect 4527 -8917 4573 -8883
rect 4607 -8917 4653 -8883
rect 4687 -8917 4733 -8883
rect 4767 -8917 4813 -8883
rect 4847 -8917 4893 -8883
rect 4927 -8917 4973 -8883
rect 5007 -8917 5040 -8883
rect 3660 -8950 5040 -8917
rect 5390 -8883 7070 -8850
rect 5390 -8917 5413 -8883
rect 5447 -8917 5493 -8883
rect 5527 -8917 5573 -8883
rect 5607 -8917 5653 -8883
rect 5687 -8917 5733 -8883
rect 5767 -8917 5813 -8883
rect 5847 -8917 5893 -8883
rect 5927 -8917 5973 -8883
rect 6007 -8917 6053 -8883
rect 6087 -8917 6133 -8883
rect 6167 -8917 6213 -8883
rect 6247 -8917 6293 -8883
rect 6327 -8917 6373 -8883
rect 6407 -8917 6453 -8883
rect 6487 -8917 6533 -8883
rect 6567 -8917 6613 -8883
rect 6647 -8917 6693 -8883
rect 6727 -8917 6773 -8883
rect 6807 -8917 6853 -8883
rect 6887 -8917 6933 -8883
rect 6967 -8917 7013 -8883
rect 7047 -8917 7070 -8883
rect 5390 -8950 7070 -8917
rect 1020 -11243 3300 -11210
rect 1020 -11277 1103 -11243
rect 1137 -11277 1183 -11243
rect 1217 -11277 1263 -11243
rect 1297 -11277 1343 -11243
rect 1377 -11277 1423 -11243
rect 1457 -11277 1503 -11243
rect 1537 -11277 1583 -11243
rect 1617 -11277 1663 -11243
rect 1697 -11277 1743 -11243
rect 1777 -11277 1823 -11243
rect 1857 -11277 1903 -11243
rect 1937 -11277 1983 -11243
rect 2017 -11277 2063 -11243
rect 2097 -11277 2143 -11243
rect 2177 -11277 2223 -11243
rect 2257 -11277 2303 -11243
rect 2337 -11277 2383 -11243
rect 2417 -11277 2463 -11243
rect 2497 -11277 2543 -11243
rect 2577 -11277 2623 -11243
rect 2657 -11277 2703 -11243
rect 2737 -11277 2783 -11243
rect 2817 -11277 2863 -11243
rect 2897 -11277 2943 -11243
rect 2977 -11277 3023 -11243
rect 3057 -11277 3103 -11243
rect 3137 -11277 3183 -11243
rect 3217 -11277 3300 -11243
rect 1020 -11310 3300 -11277
rect 3660 -11243 5040 -11210
rect 3660 -11277 3693 -11243
rect 3727 -11277 3773 -11243
rect 3807 -11277 3853 -11243
rect 3887 -11277 3933 -11243
rect 3967 -11277 4013 -11243
rect 4047 -11277 4093 -11243
rect 4127 -11277 4173 -11243
rect 4207 -11277 4253 -11243
rect 4287 -11277 4333 -11243
rect 4367 -11277 4413 -11243
rect 4447 -11277 4493 -11243
rect 4527 -11277 4573 -11243
rect 4607 -11277 4653 -11243
rect 4687 -11277 4733 -11243
rect 4767 -11277 4813 -11243
rect 4847 -11277 4893 -11243
rect 4927 -11277 4973 -11243
rect 5007 -11277 5040 -11243
rect 3660 -11310 5040 -11277
rect 5390 -11243 7070 -11210
rect 5390 -11277 5413 -11243
rect 5447 -11277 5493 -11243
rect 5527 -11277 5573 -11243
rect 5607 -11277 5653 -11243
rect 5687 -11277 5733 -11243
rect 5767 -11277 5813 -11243
rect 5847 -11277 5893 -11243
rect 5927 -11277 5973 -11243
rect 6007 -11277 6053 -11243
rect 6087 -11277 6133 -11243
rect 6167 -11277 6213 -11243
rect 6247 -11277 6293 -11243
rect 6327 -11277 6373 -11243
rect 6407 -11277 6453 -11243
rect 6487 -11277 6533 -11243
rect 6567 -11277 6613 -11243
rect 6647 -11277 6693 -11243
rect 6727 -11277 6773 -11243
rect 6807 -11277 6853 -11243
rect 6887 -11277 6933 -11243
rect 6967 -11277 7013 -11243
rect 7047 -11277 7070 -11243
rect 5390 -11310 7070 -11277
rect 1161 -11703 3161 -11670
rect 1161 -11737 1184 -11703
rect 1218 -11737 1264 -11703
rect 1298 -11737 1344 -11703
rect 1378 -11737 1424 -11703
rect 1458 -11737 1504 -11703
rect 1538 -11737 1584 -11703
rect 1618 -11737 1664 -11703
rect 1698 -11737 1744 -11703
rect 1778 -11737 1824 -11703
rect 1858 -11737 1904 -11703
rect 1938 -11737 1984 -11703
rect 2018 -11737 2064 -11703
rect 2098 -11737 2144 -11703
rect 2178 -11737 2224 -11703
rect 2258 -11737 2304 -11703
rect 2338 -11737 2384 -11703
rect 2418 -11737 2464 -11703
rect 2498 -11737 2544 -11703
rect 2578 -11737 2624 -11703
rect 2658 -11737 2704 -11703
rect 2738 -11737 2784 -11703
rect 2818 -11737 2864 -11703
rect 2898 -11737 2944 -11703
rect 2978 -11737 3024 -11703
rect 3058 -11737 3104 -11703
rect 3138 -11737 3161 -11703
rect 1161 -11770 3161 -11737
rect 3521 -11703 4901 -11670
rect 3521 -11737 3554 -11703
rect 3588 -11737 3634 -11703
rect 3668 -11737 3714 -11703
rect 3748 -11737 3794 -11703
rect 3828 -11737 3874 -11703
rect 3908 -11737 3954 -11703
rect 3988 -11737 4034 -11703
rect 4068 -11737 4114 -11703
rect 4148 -11737 4194 -11703
rect 4228 -11737 4274 -11703
rect 4308 -11737 4354 -11703
rect 4388 -11737 4434 -11703
rect 4468 -11737 4514 -11703
rect 4548 -11737 4594 -11703
rect 4628 -11737 4674 -11703
rect 4708 -11737 4754 -11703
rect 4788 -11737 4834 -11703
rect 4868 -11737 4901 -11703
rect 3521 -11770 4901 -11737
rect 5251 -11704 7251 -11671
rect 5251 -11738 5274 -11704
rect 5308 -11738 5354 -11704
rect 5388 -11738 5434 -11704
rect 5468 -11738 5514 -11704
rect 5548 -11738 5594 -11704
rect 5628 -11738 5674 -11704
rect 5708 -11738 5754 -11704
rect 5788 -11738 5834 -11704
rect 5868 -11738 5914 -11704
rect 5948 -11738 5994 -11704
rect 6028 -11738 6074 -11704
rect 6108 -11738 6154 -11704
rect 6188 -11738 6234 -11704
rect 6268 -11738 6314 -11704
rect 6348 -11738 6394 -11704
rect 6428 -11738 6474 -11704
rect 6508 -11738 6554 -11704
rect 6588 -11738 6634 -11704
rect 6668 -11738 6714 -11704
rect 6748 -11738 6794 -11704
rect 6828 -11738 6874 -11704
rect 6908 -11738 6954 -11704
rect 6988 -11738 7034 -11704
rect 7068 -11738 7114 -11704
rect 7148 -11738 7194 -11704
rect 7228 -11738 7251 -11704
rect 5251 -11771 7251 -11738
<< psubdiffcont >>
rect 1103 1264 1137 1298
rect 1183 1264 1217 1298
rect 1263 1264 1297 1298
rect 1343 1264 1377 1298
rect 1423 1264 1457 1298
rect 1503 1264 1537 1298
rect 1583 1264 1617 1298
rect 1663 1264 1697 1298
rect 1743 1264 1777 1298
rect 1823 1264 1857 1298
rect 1903 1264 1937 1298
rect 1983 1264 2017 1298
rect 2063 1264 2097 1298
rect 2143 1264 2177 1298
rect 2223 1264 2257 1298
rect 2303 1264 2337 1298
rect 2383 1264 2417 1298
rect 2463 1264 2497 1298
rect 2543 1264 2577 1298
rect 2623 1264 2657 1298
rect 2703 1264 2737 1298
rect 2783 1264 2817 1298
rect 2863 1264 2897 1298
rect 2943 1264 2977 1298
rect 3023 1264 3057 1298
rect 3103 1264 3137 1298
rect 3183 1264 3217 1298
rect 3663 1264 3697 1298
rect 3743 1264 3777 1298
rect 3823 1264 3857 1298
rect 3903 1264 3937 1298
rect 3983 1264 4017 1298
rect 4063 1264 4097 1298
rect 4143 1264 4177 1298
rect 4223 1264 4257 1298
rect 4303 1264 4337 1298
rect 4383 1264 4417 1298
rect 4463 1264 4497 1298
rect 4543 1264 4577 1298
rect 4623 1264 4657 1298
rect 4703 1264 4737 1298
rect 4783 1264 4817 1298
rect 4863 1264 4897 1298
rect 4943 1264 4977 1298
rect 5023 1264 5057 1298
rect 5103 1264 5137 1298
rect 5183 1264 5217 1298
rect 5263 1264 5297 1298
rect 5683 1264 5717 1298
rect 5763 1264 5797 1298
rect 5843 1264 5877 1298
rect 5923 1264 5957 1298
rect 6003 1264 6037 1298
rect 6083 1264 6117 1298
rect 6163 1264 6197 1298
rect 6243 1264 6277 1298
rect 6323 1264 6357 1298
rect 6403 1264 6437 1298
rect 6483 1264 6517 1298
rect 6563 1264 6597 1298
rect 6643 1264 6677 1298
rect 6723 1264 6757 1298
rect 6803 1264 6837 1298
rect 6883 1264 6917 1298
rect 6963 1264 6997 1298
rect 7043 1264 7077 1298
rect 7123 1264 7157 1298
rect 7203 1264 7237 1298
rect 7283 1264 7317 1298
rect 1103 -1556 1137 -1522
rect 1183 -1556 1217 -1522
rect 1263 -1556 1297 -1522
rect 1343 -1556 1377 -1522
rect 1423 -1556 1457 -1522
rect 1503 -1556 1537 -1522
rect 1583 -1556 1617 -1522
rect 1663 -1556 1697 -1522
rect 1743 -1556 1777 -1522
rect 1823 -1556 1857 -1522
rect 1903 -1556 1937 -1522
rect 1983 -1556 2017 -1522
rect 2063 -1556 2097 -1522
rect 2143 -1556 2177 -1522
rect 2223 -1556 2257 -1522
rect 2303 -1556 2337 -1522
rect 2383 -1556 2417 -1522
rect 2463 -1556 2497 -1522
rect 2543 -1556 2577 -1522
rect 2623 -1556 2657 -1522
rect 2703 -1556 2737 -1522
rect 2783 -1556 2817 -1522
rect 2863 -1556 2897 -1522
rect 2943 -1556 2977 -1522
rect 3023 -1556 3057 -1522
rect 3103 -1556 3137 -1522
rect 3183 -1556 3217 -1522
rect 3693 -1556 3727 -1522
rect 3773 -1556 3807 -1522
rect 3853 -1556 3887 -1522
rect 3933 -1556 3967 -1522
rect 4013 -1556 4047 -1522
rect 4093 -1556 4127 -1522
rect 4173 -1556 4207 -1522
rect 4253 -1556 4287 -1522
rect 4333 -1556 4367 -1522
rect 4413 -1556 4447 -1522
rect 4493 -1556 4527 -1522
rect 4573 -1556 4607 -1522
rect 4653 -1556 4687 -1522
rect 4733 -1556 4767 -1522
rect 4813 -1556 4847 -1522
rect 4893 -1556 4927 -1522
rect 4973 -1556 5007 -1522
rect 5413 -1556 5447 -1522
rect 5493 -1556 5527 -1522
rect 5573 -1556 5607 -1522
rect 5653 -1556 5687 -1522
rect 5733 -1556 5767 -1522
rect 5813 -1556 5847 -1522
rect 5893 -1556 5927 -1522
rect 5973 -1556 6007 -1522
rect 6053 -1556 6087 -1522
rect 6133 -1556 6167 -1522
rect 6213 -1556 6247 -1522
rect 6293 -1556 6327 -1522
rect 6373 -1556 6407 -1522
rect 6453 -1556 6487 -1522
rect 6533 -1556 6567 -1522
rect 6613 -1556 6647 -1522
rect 6693 -1556 6727 -1522
rect 6773 -1556 6807 -1522
rect 6853 -1556 6887 -1522
rect 6933 -1556 6967 -1522
rect 7013 -1556 7047 -1522
rect 1184 -4376 1218 -4342
rect 1264 -4376 1298 -4342
rect 1344 -4376 1378 -4342
rect 1424 -4376 1458 -4342
rect 1504 -4376 1538 -4342
rect 1584 -4376 1618 -4342
rect 1664 -4376 1698 -4342
rect 1744 -4376 1778 -4342
rect 1824 -4376 1858 -4342
rect 1904 -4376 1938 -4342
rect 1984 -4376 2018 -4342
rect 2064 -4376 2098 -4342
rect 2144 -4376 2178 -4342
rect 2224 -4376 2258 -4342
rect 2304 -4376 2338 -4342
rect 2384 -4376 2418 -4342
rect 2464 -4376 2498 -4342
rect 2544 -4376 2578 -4342
rect 2624 -4376 2658 -4342
rect 2704 -4376 2738 -4342
rect 2784 -4376 2818 -4342
rect 2864 -4376 2898 -4342
rect 2944 -4376 2978 -4342
rect 3024 -4376 3058 -4342
rect 3104 -4376 3138 -4342
rect 3554 -4376 3588 -4342
rect 3634 -4376 3668 -4342
rect 3714 -4376 3748 -4342
rect 3794 -4376 3828 -4342
rect 3874 -4376 3908 -4342
rect 3954 -4376 3988 -4342
rect 4034 -4376 4068 -4342
rect 4114 -4376 4148 -4342
rect 4194 -4376 4228 -4342
rect 4274 -4376 4308 -4342
rect 4354 -4376 4388 -4342
rect 4434 -4376 4468 -4342
rect 4514 -4376 4548 -4342
rect 4594 -4376 4628 -4342
rect 4674 -4376 4708 -4342
rect 4754 -4376 4788 -4342
rect 4834 -4376 4868 -4342
rect 5274 -4377 5308 -4343
rect 5354 -4377 5388 -4343
rect 5434 -4377 5468 -4343
rect 5514 -4377 5548 -4343
rect 5594 -4377 5628 -4343
rect 5674 -4377 5708 -4343
rect 5754 -4377 5788 -4343
rect 5834 -4377 5868 -4343
rect 5914 -4377 5948 -4343
rect 5994 -4377 6028 -4343
rect 6074 -4377 6108 -4343
rect 6154 -4377 6188 -4343
rect 6234 -4377 6268 -4343
rect 6314 -4377 6348 -4343
rect 6394 -4377 6428 -4343
rect 6474 -4377 6508 -4343
rect 6554 -4377 6588 -4343
rect 6634 -4377 6668 -4343
rect 6714 -4377 6748 -4343
rect 6794 -4377 6828 -4343
rect 6874 -4377 6908 -4343
rect 6954 -4377 6988 -4343
rect 7034 -4377 7068 -4343
rect 7114 -4377 7148 -4343
rect 7194 -4377 7228 -4343
rect 1063 -4456 1097 -4422
rect 1143 -4456 1177 -4422
rect 1223 -4456 1257 -4422
rect 1303 -4456 1337 -4422
rect 1383 -4456 1417 -4422
rect 1463 -4456 1497 -4422
rect 1543 -4456 1577 -4422
rect 1623 -4456 1657 -4422
rect 1703 -4456 1737 -4422
rect 1783 -4456 1817 -4422
rect 1863 -4456 1897 -4422
rect 1943 -4456 1977 -4422
rect 2023 -4456 2057 -4422
rect 2103 -4456 2137 -4422
rect 2183 -4456 2217 -4422
rect 2263 -4456 2297 -4422
rect 2343 -4456 2377 -4422
rect 2423 -4456 2457 -4422
rect 2503 -4456 2537 -4422
rect 2583 -4456 2617 -4422
rect 2663 -4456 2697 -4422
rect 2743 -4456 2777 -4422
rect 2823 -4456 2857 -4422
rect 2903 -4456 2937 -4422
rect 2983 -4456 3017 -4422
rect 3063 -4456 3097 -4422
rect 3143 -4456 3177 -4422
rect 3223 -4456 3257 -4422
rect 3303 -4456 3337 -4422
rect 3754 -4457 3788 -4423
rect 3834 -4457 3868 -4423
rect 3914 -4457 3948 -4423
rect 3994 -4457 4028 -4423
rect 4074 -4457 4108 -4423
rect 4154 -4457 4188 -4423
rect 4234 -4457 4268 -4423
rect 4314 -4457 4348 -4423
rect 4394 -4457 4428 -4423
rect 4474 -4457 4508 -4423
rect 4554 -4457 4588 -4423
rect 4634 -4457 4668 -4423
rect 4714 -4457 4748 -4423
rect 4794 -4457 4828 -4423
rect 4874 -4457 4908 -4423
rect 4954 -4457 4988 -4423
rect 5034 -4457 5068 -4423
rect 5493 -4457 5527 -4423
rect 5573 -4457 5607 -4423
rect 5653 -4457 5687 -4423
rect 5733 -4457 5767 -4423
rect 5813 -4457 5847 -4423
rect 5893 -4457 5927 -4423
rect 5973 -4457 6007 -4423
rect 6053 -4457 6087 -4423
rect 6133 -4457 6167 -4423
rect 6213 -4457 6247 -4423
rect 6293 -4457 6327 -4423
rect 6373 -4457 6407 -4423
rect 6453 -4457 6487 -4423
rect 6533 -4457 6567 -4423
rect 6613 -4457 6647 -4423
rect 6693 -4457 6727 -4423
rect 6773 -4457 6807 -4423
rect 6853 -4457 6887 -4423
rect 6933 -4457 6967 -4423
rect 7013 -4457 7047 -4423
rect 7093 -4457 7127 -4423
rect 7173 -4457 7207 -4423
rect 7253 -4457 7287 -4423
rect 7333 -4457 7367 -4423
rect 7413 -4457 7447 -4423
rect 1143 -7277 1177 -7243
rect 1223 -7277 1257 -7243
rect 1303 -7277 1337 -7243
rect 1383 -7277 1417 -7243
rect 1463 -7277 1497 -7243
rect 1543 -7277 1577 -7243
rect 1623 -7277 1657 -7243
rect 1703 -7277 1737 -7243
rect 1783 -7277 1817 -7243
rect 1863 -7277 1897 -7243
rect 1943 -7277 1977 -7243
rect 2023 -7277 2057 -7243
rect 2103 -7277 2137 -7243
rect 2183 -7277 2217 -7243
rect 2263 -7277 2297 -7243
rect 2343 -7277 2377 -7243
rect 2423 -7277 2457 -7243
rect 2503 -7277 2537 -7243
rect 2583 -7277 2617 -7243
rect 2663 -7277 2697 -7243
rect 2743 -7277 2777 -7243
rect 2823 -7277 2857 -7243
rect 2903 -7277 2937 -7243
rect 2983 -7277 3017 -7243
rect 3063 -7277 3097 -7243
rect 3143 -7277 3177 -7243
rect 3223 -7277 3257 -7243
rect 3753 -7277 3787 -7243
rect 3833 -7277 3867 -7243
rect 3913 -7277 3947 -7243
rect 3993 -7277 4027 -7243
rect 4073 -7277 4107 -7243
rect 4153 -7277 4187 -7243
rect 4233 -7277 4267 -7243
rect 4313 -7277 4347 -7243
rect 4393 -7277 4427 -7243
rect 4473 -7277 4507 -7243
rect 4553 -7277 4587 -7243
rect 4633 -7277 4667 -7243
rect 4713 -7277 4747 -7243
rect 4793 -7277 4827 -7243
rect 4873 -7277 4907 -7243
rect 4953 -7277 4987 -7243
rect 5033 -7277 5067 -7243
rect 5472 -7277 5506 -7243
rect 5552 -7277 5586 -7243
rect 5632 -7277 5666 -7243
rect 5712 -7277 5746 -7243
rect 5792 -7277 5826 -7243
rect 5872 -7277 5906 -7243
rect 5952 -7277 5986 -7243
rect 6032 -7277 6066 -7243
rect 6112 -7277 6146 -7243
rect 6192 -7277 6226 -7243
rect 6272 -7277 6306 -7243
rect 6352 -7277 6386 -7243
rect 6432 -7277 6466 -7243
rect 6512 -7277 6546 -7243
rect 6592 -7277 6626 -7243
rect 6672 -7277 6706 -7243
rect 6752 -7277 6786 -7243
rect 6832 -7277 6866 -7243
rect 6912 -7277 6946 -7243
rect 6992 -7277 7026 -7243
rect 7072 -7277 7106 -7243
rect 1103 -10097 1137 -10063
rect 1183 -10097 1217 -10063
rect 1263 -10097 1297 -10063
rect 1343 -10097 1377 -10063
rect 1423 -10097 1457 -10063
rect 1503 -10097 1537 -10063
rect 1583 -10097 1617 -10063
rect 1663 -10097 1697 -10063
rect 1743 -10097 1777 -10063
rect 1823 -10097 1857 -10063
rect 1903 -10097 1937 -10063
rect 1983 -10097 2017 -10063
rect 2063 -10097 2097 -10063
rect 2143 -10097 2177 -10063
rect 2223 -10097 2257 -10063
rect 2303 -10097 2337 -10063
rect 2383 -10097 2417 -10063
rect 2463 -10097 2497 -10063
rect 2543 -10097 2577 -10063
rect 2623 -10097 2657 -10063
rect 2703 -10097 2737 -10063
rect 2783 -10097 2817 -10063
rect 2863 -10097 2897 -10063
rect 2943 -10097 2977 -10063
rect 3023 -10097 3057 -10063
rect 3103 -10097 3137 -10063
rect 3183 -10097 3217 -10063
rect 3693 -10097 3727 -10063
rect 3773 -10097 3807 -10063
rect 3853 -10097 3887 -10063
rect 3933 -10097 3967 -10063
rect 4013 -10097 4047 -10063
rect 4093 -10097 4127 -10063
rect 4173 -10097 4207 -10063
rect 4253 -10097 4287 -10063
rect 4333 -10097 4367 -10063
rect 4413 -10097 4447 -10063
rect 4493 -10097 4527 -10063
rect 4573 -10097 4607 -10063
rect 4653 -10097 4687 -10063
rect 4733 -10097 4767 -10063
rect 4813 -10097 4847 -10063
rect 4893 -10097 4927 -10063
rect 4973 -10097 5007 -10063
rect 5413 -10097 5447 -10063
rect 5493 -10097 5527 -10063
rect 5573 -10097 5607 -10063
rect 5653 -10097 5687 -10063
rect 5733 -10097 5767 -10063
rect 5813 -10097 5847 -10063
rect 5893 -10097 5927 -10063
rect 5973 -10097 6007 -10063
rect 6053 -10097 6087 -10063
rect 6133 -10097 6167 -10063
rect 6213 -10097 6247 -10063
rect 6293 -10097 6327 -10063
rect 6373 -10097 6407 -10063
rect 6453 -10097 6487 -10063
rect 6533 -10097 6567 -10063
rect 6613 -10097 6647 -10063
rect 6693 -10097 6727 -10063
rect 6773 -10097 6807 -10063
rect 6853 -10097 6887 -10063
rect 6933 -10097 6967 -10063
rect 7013 -10097 7047 -10063
rect 1184 -12917 1218 -12883
rect 1264 -12917 1298 -12883
rect 1344 -12917 1378 -12883
rect 1424 -12917 1458 -12883
rect 1504 -12917 1538 -12883
rect 1584 -12917 1618 -12883
rect 1664 -12917 1698 -12883
rect 1744 -12917 1778 -12883
rect 1824 -12917 1858 -12883
rect 1904 -12917 1938 -12883
rect 1984 -12917 2018 -12883
rect 2064 -12917 2098 -12883
rect 2144 -12917 2178 -12883
rect 2224 -12917 2258 -12883
rect 2304 -12917 2338 -12883
rect 2384 -12917 2418 -12883
rect 2464 -12917 2498 -12883
rect 2544 -12917 2578 -12883
rect 2624 -12917 2658 -12883
rect 2704 -12917 2738 -12883
rect 2784 -12917 2818 -12883
rect 2864 -12917 2898 -12883
rect 2944 -12917 2978 -12883
rect 3024 -12917 3058 -12883
rect 3104 -12917 3138 -12883
rect 3554 -12917 3588 -12883
rect 3634 -12917 3668 -12883
rect 3714 -12917 3748 -12883
rect 3794 -12917 3828 -12883
rect 3874 -12917 3908 -12883
rect 3954 -12917 3988 -12883
rect 4034 -12917 4068 -12883
rect 4114 -12917 4148 -12883
rect 4194 -12917 4228 -12883
rect 4274 -12917 4308 -12883
rect 4354 -12917 4388 -12883
rect 4434 -12917 4468 -12883
rect 4514 -12917 4548 -12883
rect 4594 -12917 4628 -12883
rect 4674 -12917 4708 -12883
rect 4754 -12917 4788 -12883
rect 4834 -12917 4868 -12883
rect 5274 -12918 5308 -12884
rect 5354 -12918 5388 -12884
rect 5434 -12918 5468 -12884
rect 5514 -12918 5548 -12884
rect 5594 -12918 5628 -12884
rect 5674 -12918 5708 -12884
rect 5754 -12918 5788 -12884
rect 5834 -12918 5868 -12884
rect 5914 -12918 5948 -12884
rect 5994 -12918 6028 -12884
rect 6074 -12918 6108 -12884
rect 6154 -12918 6188 -12884
rect 6234 -12918 6268 -12884
rect 6314 -12918 6348 -12884
rect 6394 -12918 6428 -12884
rect 6474 -12918 6508 -12884
rect 6554 -12918 6588 -12884
rect 6634 -12918 6668 -12884
rect 6714 -12918 6748 -12884
rect 6794 -12918 6828 -12884
rect 6874 -12918 6908 -12884
rect 6954 -12918 6988 -12884
rect 7034 -12918 7068 -12884
rect 7114 -12918 7148 -12884
rect 7194 -12918 7228 -12884
<< nsubdiffcont >>
rect 1103 2444 1137 2478
rect 1183 2444 1217 2478
rect 1263 2444 1297 2478
rect 1343 2444 1377 2478
rect 1423 2444 1457 2478
rect 1503 2444 1537 2478
rect 1583 2444 1617 2478
rect 1663 2444 1697 2478
rect 1743 2444 1777 2478
rect 1823 2444 1857 2478
rect 1903 2444 1937 2478
rect 1983 2444 2017 2478
rect 2063 2444 2097 2478
rect 2143 2444 2177 2478
rect 2223 2444 2257 2478
rect 2303 2444 2337 2478
rect 2383 2444 2417 2478
rect 2463 2444 2497 2478
rect 2543 2444 2577 2478
rect 2623 2444 2657 2478
rect 2703 2444 2737 2478
rect 2783 2444 2817 2478
rect 2863 2444 2897 2478
rect 2943 2444 2977 2478
rect 3023 2444 3057 2478
rect 3103 2444 3137 2478
rect 3183 2444 3217 2478
rect 3663 2444 3697 2478
rect 3743 2444 3777 2478
rect 3823 2444 3857 2478
rect 3903 2444 3937 2478
rect 3983 2444 4017 2478
rect 4063 2444 4097 2478
rect 4143 2444 4177 2478
rect 4223 2444 4257 2478
rect 4303 2444 4337 2478
rect 4383 2444 4417 2478
rect 4463 2444 4497 2478
rect 4543 2444 4577 2478
rect 4623 2444 4657 2478
rect 4703 2444 4737 2478
rect 4783 2444 4817 2478
rect 4863 2444 4897 2478
rect 4943 2444 4977 2478
rect 5023 2444 5057 2478
rect 5103 2444 5137 2478
rect 5183 2444 5217 2478
rect 5263 2444 5297 2478
rect 5683 2444 5717 2478
rect 5763 2444 5797 2478
rect 5843 2444 5877 2478
rect 5923 2444 5957 2478
rect 6003 2444 6037 2478
rect 6083 2444 6117 2478
rect 6163 2444 6197 2478
rect 6243 2444 6277 2478
rect 6323 2444 6357 2478
rect 6403 2444 6437 2478
rect 6483 2444 6517 2478
rect 6563 2444 6597 2478
rect 6643 2444 6677 2478
rect 6723 2444 6757 2478
rect 6803 2444 6837 2478
rect 6883 2444 6917 2478
rect 6963 2444 6997 2478
rect 7043 2444 7077 2478
rect 7123 2444 7157 2478
rect 7203 2444 7237 2478
rect 7283 2444 7317 2478
rect 1343 84 1377 118
rect 1423 84 1457 118
rect 1503 84 1537 118
rect 1583 84 1617 118
rect 1663 84 1697 118
rect 1743 84 1777 118
rect 1823 84 1857 118
rect 1903 84 1937 118
rect 1983 84 2017 118
rect 2063 84 2097 118
rect 2143 84 2177 118
rect 2223 84 2257 118
rect 2303 84 2337 118
rect 2383 84 2417 118
rect 2463 84 2497 118
rect 2543 84 2577 118
rect 2623 84 2657 118
rect 2703 84 2737 118
rect 2783 84 2817 118
rect 2863 84 2897 118
rect 2943 84 2977 118
rect 3663 84 3697 118
rect 3743 84 3777 118
rect 3823 84 3857 118
rect 3903 84 3937 118
rect 3983 84 4017 118
rect 4063 84 4097 118
rect 4143 84 4177 118
rect 4223 84 4257 118
rect 4303 84 4337 118
rect 4383 84 4417 118
rect 4463 84 4497 118
rect 4543 84 4577 118
rect 4623 84 4657 118
rect 4703 84 4737 118
rect 4783 84 4817 118
rect 4863 84 4897 118
rect 4943 84 4977 118
rect 5023 84 5057 118
rect 5103 84 5137 118
rect 5183 84 5217 118
rect 5263 84 5297 118
rect 5683 84 5717 118
rect 5763 84 5797 118
rect 5843 84 5877 118
rect 5923 84 5957 118
rect 6003 84 6037 118
rect 6083 84 6117 118
rect 6163 84 6197 118
rect 6243 84 6277 118
rect 6323 84 6357 118
rect 6403 84 6437 118
rect 6483 84 6517 118
rect 6563 84 6597 118
rect 6643 84 6677 118
rect 6723 84 6757 118
rect 6803 84 6837 118
rect 6883 84 6917 118
rect 6963 84 6997 118
rect 7043 84 7077 118
rect 7123 84 7157 118
rect 7203 84 7237 118
rect 7283 84 7317 118
rect 1103 -376 1137 -342
rect 1183 -376 1217 -342
rect 1263 -376 1297 -342
rect 1343 -376 1377 -342
rect 1423 -376 1457 -342
rect 1503 -376 1537 -342
rect 1583 -376 1617 -342
rect 1663 -376 1697 -342
rect 1743 -376 1777 -342
rect 1823 -376 1857 -342
rect 1903 -376 1937 -342
rect 1983 -376 2017 -342
rect 2063 -376 2097 -342
rect 2143 -376 2177 -342
rect 2223 -376 2257 -342
rect 2303 -376 2337 -342
rect 2383 -376 2417 -342
rect 2463 -376 2497 -342
rect 2543 -376 2577 -342
rect 2623 -376 2657 -342
rect 2703 -376 2737 -342
rect 2783 -376 2817 -342
rect 2863 -376 2897 -342
rect 2943 -376 2977 -342
rect 3023 -376 3057 -342
rect 3103 -376 3137 -342
rect 3183 -376 3217 -342
rect 3693 -376 3727 -342
rect 3773 -376 3807 -342
rect 3853 -376 3887 -342
rect 3933 -376 3967 -342
rect 4013 -376 4047 -342
rect 4093 -376 4127 -342
rect 4173 -376 4207 -342
rect 4253 -376 4287 -342
rect 4333 -376 4367 -342
rect 4413 -376 4447 -342
rect 4493 -376 4527 -342
rect 4573 -376 4607 -342
rect 4653 -376 4687 -342
rect 4733 -376 4767 -342
rect 4813 -376 4847 -342
rect 4893 -376 4927 -342
rect 4973 -376 5007 -342
rect 5413 -376 5447 -342
rect 5493 -376 5527 -342
rect 5573 -376 5607 -342
rect 5653 -376 5687 -342
rect 5733 -376 5767 -342
rect 5813 -376 5847 -342
rect 5893 -376 5927 -342
rect 5973 -376 6007 -342
rect 6053 -376 6087 -342
rect 6133 -376 6167 -342
rect 6213 -376 6247 -342
rect 6293 -376 6327 -342
rect 6373 -376 6407 -342
rect 6453 -376 6487 -342
rect 6533 -376 6567 -342
rect 6613 -376 6647 -342
rect 6693 -376 6727 -342
rect 6773 -376 6807 -342
rect 6853 -376 6887 -342
rect 6933 -376 6967 -342
rect 7013 -376 7047 -342
rect 1103 -2736 1137 -2702
rect 1183 -2736 1217 -2702
rect 1263 -2736 1297 -2702
rect 1343 -2736 1377 -2702
rect 1423 -2736 1457 -2702
rect 1503 -2736 1537 -2702
rect 1583 -2736 1617 -2702
rect 1663 -2736 1697 -2702
rect 1743 -2736 1777 -2702
rect 1823 -2736 1857 -2702
rect 1903 -2736 1937 -2702
rect 1983 -2736 2017 -2702
rect 2063 -2736 2097 -2702
rect 2143 -2736 2177 -2702
rect 2223 -2736 2257 -2702
rect 2303 -2736 2337 -2702
rect 2383 -2736 2417 -2702
rect 2463 -2736 2497 -2702
rect 2543 -2736 2577 -2702
rect 2623 -2736 2657 -2702
rect 2703 -2736 2737 -2702
rect 2783 -2736 2817 -2702
rect 2863 -2736 2897 -2702
rect 2943 -2736 2977 -2702
rect 3023 -2736 3057 -2702
rect 3103 -2736 3137 -2702
rect 3183 -2736 3217 -2702
rect 3693 -2736 3727 -2702
rect 3773 -2736 3807 -2702
rect 3853 -2736 3887 -2702
rect 3933 -2736 3967 -2702
rect 4013 -2736 4047 -2702
rect 4093 -2736 4127 -2702
rect 4173 -2736 4207 -2702
rect 4253 -2736 4287 -2702
rect 4333 -2736 4367 -2702
rect 4413 -2736 4447 -2702
rect 4493 -2736 4527 -2702
rect 4573 -2736 4607 -2702
rect 4653 -2736 4687 -2702
rect 4733 -2736 4767 -2702
rect 4813 -2736 4847 -2702
rect 4893 -2736 4927 -2702
rect 4973 -2736 5007 -2702
rect 5413 -2736 5447 -2702
rect 5493 -2736 5527 -2702
rect 5573 -2736 5607 -2702
rect 5653 -2736 5687 -2702
rect 5733 -2736 5767 -2702
rect 5813 -2736 5847 -2702
rect 5893 -2736 5927 -2702
rect 5973 -2736 6007 -2702
rect 6053 -2736 6087 -2702
rect 6133 -2736 6167 -2702
rect 6213 -2736 6247 -2702
rect 6293 -2736 6327 -2702
rect 6373 -2736 6407 -2702
rect 6453 -2736 6487 -2702
rect 6533 -2736 6567 -2702
rect 6613 -2736 6647 -2702
rect 6693 -2736 6727 -2702
rect 6773 -2736 6807 -2702
rect 6853 -2736 6887 -2702
rect 6933 -2736 6967 -2702
rect 7013 -2736 7047 -2702
rect 1184 -3196 1218 -3162
rect 1264 -3196 1298 -3162
rect 1344 -3196 1378 -3162
rect 1424 -3196 1458 -3162
rect 1504 -3196 1538 -3162
rect 1584 -3196 1618 -3162
rect 1664 -3196 1698 -3162
rect 1744 -3196 1778 -3162
rect 1824 -3196 1858 -3162
rect 1904 -3196 1938 -3162
rect 1984 -3196 2018 -3162
rect 2064 -3196 2098 -3162
rect 2144 -3196 2178 -3162
rect 2224 -3196 2258 -3162
rect 2304 -3196 2338 -3162
rect 2384 -3196 2418 -3162
rect 2464 -3196 2498 -3162
rect 2544 -3196 2578 -3162
rect 2624 -3196 2658 -3162
rect 2704 -3196 2738 -3162
rect 2784 -3196 2818 -3162
rect 2864 -3196 2898 -3162
rect 2944 -3196 2978 -3162
rect 3024 -3196 3058 -3162
rect 3104 -3196 3138 -3162
rect 3554 -3196 3588 -3162
rect 3634 -3196 3668 -3162
rect 3714 -3196 3748 -3162
rect 3794 -3196 3828 -3162
rect 3874 -3196 3908 -3162
rect 3954 -3196 3988 -3162
rect 4034 -3196 4068 -3162
rect 4114 -3196 4148 -3162
rect 4194 -3196 4228 -3162
rect 4274 -3196 4308 -3162
rect 4354 -3196 4388 -3162
rect 4434 -3196 4468 -3162
rect 4514 -3196 4548 -3162
rect 4594 -3196 4628 -3162
rect 4674 -3196 4708 -3162
rect 4754 -3196 4788 -3162
rect 4834 -3196 4868 -3162
rect 5274 -3197 5308 -3163
rect 5354 -3197 5388 -3163
rect 5434 -3197 5468 -3163
rect 5514 -3197 5548 -3163
rect 5594 -3197 5628 -3163
rect 5674 -3197 5708 -3163
rect 5754 -3197 5788 -3163
rect 5834 -3197 5868 -3163
rect 5914 -3197 5948 -3163
rect 5994 -3197 6028 -3163
rect 6074 -3197 6108 -3163
rect 6154 -3197 6188 -3163
rect 6234 -3197 6268 -3163
rect 6314 -3197 6348 -3163
rect 6394 -3197 6428 -3163
rect 6474 -3197 6508 -3163
rect 6554 -3197 6588 -3163
rect 6634 -3197 6668 -3163
rect 6714 -3197 6748 -3163
rect 6794 -3197 6828 -3163
rect 6874 -3197 6908 -3163
rect 6954 -3197 6988 -3163
rect 7034 -3197 7068 -3163
rect 7114 -3197 7148 -3163
rect 7194 -3197 7228 -3163
rect 3754 -5637 3788 -5603
rect 3834 -5637 3868 -5603
rect 3914 -5637 3948 -5603
rect 3994 -5637 4028 -5603
rect 4074 -5637 4108 -5603
rect 4154 -5637 4188 -5603
rect 4234 -5637 4268 -5603
rect 4314 -5637 4348 -5603
rect 4394 -5637 4428 -5603
rect 4474 -5637 4508 -5603
rect 4554 -5637 4588 -5603
rect 4634 -5637 4668 -5603
rect 4714 -5637 4748 -5603
rect 4794 -5637 4828 -5603
rect 4874 -5637 4908 -5603
rect 4954 -5637 4988 -5603
rect 5034 -5637 5068 -5603
rect 5493 -5637 5527 -5603
rect 5573 -5637 5607 -5603
rect 5653 -5637 5687 -5603
rect 5733 -5637 5767 -5603
rect 5813 -5637 5847 -5603
rect 5893 -5637 5927 -5603
rect 5973 -5637 6007 -5603
rect 6053 -5637 6087 -5603
rect 6133 -5637 6167 -5603
rect 6213 -5637 6247 -5603
rect 6293 -5637 6327 -5603
rect 6373 -5637 6407 -5603
rect 6453 -5637 6487 -5603
rect 6533 -5637 6567 -5603
rect 6613 -5637 6647 -5603
rect 6693 -5637 6727 -5603
rect 6773 -5637 6807 -5603
rect 6853 -5637 6887 -5603
rect 6933 -5637 6967 -5603
rect 7013 -5637 7047 -5603
rect 7093 -5637 7127 -5603
rect 7173 -5637 7207 -5603
rect 7253 -5637 7287 -5603
rect 7333 -5637 7367 -5603
rect 7413 -5637 7447 -5603
rect 1063 -5956 1097 -5922
rect 1143 -5956 1177 -5922
rect 1223 -5956 1257 -5922
rect 1303 -5956 1337 -5922
rect 1383 -5956 1417 -5922
rect 1463 -5956 1497 -5922
rect 1543 -5956 1577 -5922
rect 1623 -5956 1657 -5922
rect 1703 -5956 1737 -5922
rect 1783 -5956 1817 -5922
rect 1863 -5956 1897 -5922
rect 1943 -5956 1977 -5922
rect 2023 -5956 2057 -5922
rect 2103 -5956 2137 -5922
rect 2183 -5956 2217 -5922
rect 2263 -5956 2297 -5922
rect 2343 -5956 2377 -5922
rect 2423 -5956 2457 -5922
rect 2503 -5956 2537 -5922
rect 2583 -5956 2617 -5922
rect 2663 -5956 2697 -5922
rect 2743 -5956 2777 -5922
rect 2823 -5956 2857 -5922
rect 2903 -5956 2937 -5922
rect 2983 -5956 3017 -5922
rect 3063 -5956 3097 -5922
rect 3143 -5956 3177 -5922
rect 3223 -5956 3257 -5922
rect 3303 -5956 3337 -5922
rect 1063 -6097 1097 -6063
rect 1143 -6097 1177 -6063
rect 1223 -6097 1257 -6063
rect 1303 -6097 1337 -6063
rect 1383 -6097 1417 -6063
rect 1463 -6097 1497 -6063
rect 1543 -6097 1577 -6063
rect 1623 -6097 1657 -6063
rect 1703 -6097 1737 -6063
rect 1783 -6097 1817 -6063
rect 1863 -6097 1897 -6063
rect 1943 -6097 1977 -6063
rect 2023 -6097 2057 -6063
rect 2103 -6097 2137 -6063
rect 2183 -6097 2217 -6063
rect 2263 -6097 2297 -6063
rect 2343 -6097 2377 -6063
rect 2423 -6097 2457 -6063
rect 2503 -6097 2537 -6063
rect 2583 -6097 2617 -6063
rect 2663 -6097 2697 -6063
rect 2743 -6097 2777 -6063
rect 2823 -6097 2857 -6063
rect 2903 -6097 2937 -6063
rect 2983 -6097 3017 -6063
rect 3063 -6097 3097 -6063
rect 3143 -6097 3177 -6063
rect 3223 -6097 3257 -6063
rect 3303 -6097 3337 -6063
rect 3753 -6097 3787 -6063
rect 3833 -6097 3867 -6063
rect 3913 -6097 3947 -6063
rect 3993 -6097 4027 -6063
rect 4073 -6097 4107 -6063
rect 4153 -6097 4187 -6063
rect 4233 -6097 4267 -6063
rect 4313 -6097 4347 -6063
rect 4393 -6097 4427 -6063
rect 4473 -6097 4507 -6063
rect 4553 -6097 4587 -6063
rect 4633 -6097 4667 -6063
rect 4713 -6097 4747 -6063
rect 4793 -6097 4827 -6063
rect 4873 -6097 4907 -6063
rect 4953 -6097 4987 -6063
rect 5033 -6097 5067 -6063
rect 5472 -6097 5506 -6063
rect 5552 -6097 5586 -6063
rect 5632 -6097 5666 -6063
rect 5712 -6097 5746 -6063
rect 5792 -6097 5826 -6063
rect 5872 -6097 5906 -6063
rect 5952 -6097 5986 -6063
rect 6032 -6097 6066 -6063
rect 6112 -6097 6146 -6063
rect 6192 -6097 6226 -6063
rect 6272 -6097 6306 -6063
rect 6352 -6097 6386 -6063
rect 6432 -6097 6466 -6063
rect 6512 -6097 6546 -6063
rect 6592 -6097 6626 -6063
rect 6672 -6097 6706 -6063
rect 6752 -6097 6786 -6063
rect 6832 -6097 6866 -6063
rect 6912 -6097 6946 -6063
rect 6992 -6097 7026 -6063
rect 7072 -6097 7106 -6063
rect 1143 -8457 1177 -8423
rect 1223 -8457 1257 -8423
rect 1303 -8457 1337 -8423
rect 1383 -8457 1417 -8423
rect 1463 -8457 1497 -8423
rect 1543 -8457 1577 -8423
rect 1623 -8457 1657 -8423
rect 1703 -8457 1737 -8423
rect 1783 -8457 1817 -8423
rect 1863 -8457 1897 -8423
rect 1943 -8457 1977 -8423
rect 2023 -8457 2057 -8423
rect 2103 -8457 2137 -8423
rect 2183 -8457 2217 -8423
rect 2263 -8457 2297 -8423
rect 2343 -8457 2377 -8423
rect 2423 -8457 2457 -8423
rect 2503 -8457 2537 -8423
rect 2583 -8457 2617 -8423
rect 2663 -8457 2697 -8423
rect 2743 -8457 2777 -8423
rect 2823 -8457 2857 -8423
rect 2903 -8457 2937 -8423
rect 2983 -8457 3017 -8423
rect 3063 -8457 3097 -8423
rect 3143 -8457 3177 -8423
rect 3223 -8457 3257 -8423
rect 3753 -8457 3787 -8423
rect 3833 -8457 3867 -8423
rect 3913 -8457 3947 -8423
rect 3993 -8457 4027 -8423
rect 4073 -8457 4107 -8423
rect 4153 -8457 4187 -8423
rect 4233 -8457 4267 -8423
rect 4313 -8457 4347 -8423
rect 4393 -8457 4427 -8423
rect 4473 -8457 4507 -8423
rect 4553 -8457 4587 -8423
rect 4633 -8457 4667 -8423
rect 4713 -8457 4747 -8423
rect 4793 -8457 4827 -8423
rect 4873 -8457 4907 -8423
rect 4953 -8457 4987 -8423
rect 5033 -8457 5067 -8423
rect 5472 -8457 5506 -8423
rect 5552 -8457 5586 -8423
rect 5632 -8457 5666 -8423
rect 5712 -8457 5746 -8423
rect 5792 -8457 5826 -8423
rect 5872 -8457 5906 -8423
rect 5952 -8457 5986 -8423
rect 6032 -8457 6066 -8423
rect 6112 -8457 6146 -8423
rect 6192 -8457 6226 -8423
rect 6272 -8457 6306 -8423
rect 6352 -8457 6386 -8423
rect 6432 -8457 6466 -8423
rect 6512 -8457 6546 -8423
rect 6592 -8457 6626 -8423
rect 6672 -8457 6706 -8423
rect 6752 -8457 6786 -8423
rect 6832 -8457 6866 -8423
rect 6912 -8457 6946 -8423
rect 6992 -8457 7026 -8423
rect 7072 -8457 7106 -8423
rect 1103 -8917 1137 -8883
rect 1183 -8917 1217 -8883
rect 1263 -8917 1297 -8883
rect 1343 -8917 1377 -8883
rect 1423 -8917 1457 -8883
rect 1503 -8917 1537 -8883
rect 1583 -8917 1617 -8883
rect 1663 -8917 1697 -8883
rect 1743 -8917 1777 -8883
rect 1823 -8917 1857 -8883
rect 1903 -8917 1937 -8883
rect 1983 -8917 2017 -8883
rect 2063 -8917 2097 -8883
rect 2143 -8917 2177 -8883
rect 2223 -8917 2257 -8883
rect 2303 -8917 2337 -8883
rect 2383 -8917 2417 -8883
rect 2463 -8917 2497 -8883
rect 2543 -8917 2577 -8883
rect 2623 -8917 2657 -8883
rect 2703 -8917 2737 -8883
rect 2783 -8917 2817 -8883
rect 2863 -8917 2897 -8883
rect 2943 -8917 2977 -8883
rect 3023 -8917 3057 -8883
rect 3103 -8917 3137 -8883
rect 3183 -8917 3217 -8883
rect 3693 -8917 3727 -8883
rect 3773 -8917 3807 -8883
rect 3853 -8917 3887 -8883
rect 3933 -8917 3967 -8883
rect 4013 -8917 4047 -8883
rect 4093 -8917 4127 -8883
rect 4173 -8917 4207 -8883
rect 4253 -8917 4287 -8883
rect 4333 -8917 4367 -8883
rect 4413 -8917 4447 -8883
rect 4493 -8917 4527 -8883
rect 4573 -8917 4607 -8883
rect 4653 -8917 4687 -8883
rect 4733 -8917 4767 -8883
rect 4813 -8917 4847 -8883
rect 4893 -8917 4927 -8883
rect 4973 -8917 5007 -8883
rect 5413 -8917 5447 -8883
rect 5493 -8917 5527 -8883
rect 5573 -8917 5607 -8883
rect 5653 -8917 5687 -8883
rect 5733 -8917 5767 -8883
rect 5813 -8917 5847 -8883
rect 5893 -8917 5927 -8883
rect 5973 -8917 6007 -8883
rect 6053 -8917 6087 -8883
rect 6133 -8917 6167 -8883
rect 6213 -8917 6247 -8883
rect 6293 -8917 6327 -8883
rect 6373 -8917 6407 -8883
rect 6453 -8917 6487 -8883
rect 6533 -8917 6567 -8883
rect 6613 -8917 6647 -8883
rect 6693 -8917 6727 -8883
rect 6773 -8917 6807 -8883
rect 6853 -8917 6887 -8883
rect 6933 -8917 6967 -8883
rect 7013 -8917 7047 -8883
rect 1103 -11277 1137 -11243
rect 1183 -11277 1217 -11243
rect 1263 -11277 1297 -11243
rect 1343 -11277 1377 -11243
rect 1423 -11277 1457 -11243
rect 1503 -11277 1537 -11243
rect 1583 -11277 1617 -11243
rect 1663 -11277 1697 -11243
rect 1743 -11277 1777 -11243
rect 1823 -11277 1857 -11243
rect 1903 -11277 1937 -11243
rect 1983 -11277 2017 -11243
rect 2063 -11277 2097 -11243
rect 2143 -11277 2177 -11243
rect 2223 -11277 2257 -11243
rect 2303 -11277 2337 -11243
rect 2383 -11277 2417 -11243
rect 2463 -11277 2497 -11243
rect 2543 -11277 2577 -11243
rect 2623 -11277 2657 -11243
rect 2703 -11277 2737 -11243
rect 2783 -11277 2817 -11243
rect 2863 -11277 2897 -11243
rect 2943 -11277 2977 -11243
rect 3023 -11277 3057 -11243
rect 3103 -11277 3137 -11243
rect 3183 -11277 3217 -11243
rect 3693 -11277 3727 -11243
rect 3773 -11277 3807 -11243
rect 3853 -11277 3887 -11243
rect 3933 -11277 3967 -11243
rect 4013 -11277 4047 -11243
rect 4093 -11277 4127 -11243
rect 4173 -11277 4207 -11243
rect 4253 -11277 4287 -11243
rect 4333 -11277 4367 -11243
rect 4413 -11277 4447 -11243
rect 4493 -11277 4527 -11243
rect 4573 -11277 4607 -11243
rect 4653 -11277 4687 -11243
rect 4733 -11277 4767 -11243
rect 4813 -11277 4847 -11243
rect 4893 -11277 4927 -11243
rect 4973 -11277 5007 -11243
rect 5413 -11277 5447 -11243
rect 5493 -11277 5527 -11243
rect 5573 -11277 5607 -11243
rect 5653 -11277 5687 -11243
rect 5733 -11277 5767 -11243
rect 5813 -11277 5847 -11243
rect 5893 -11277 5927 -11243
rect 5973 -11277 6007 -11243
rect 6053 -11277 6087 -11243
rect 6133 -11277 6167 -11243
rect 6213 -11277 6247 -11243
rect 6293 -11277 6327 -11243
rect 6373 -11277 6407 -11243
rect 6453 -11277 6487 -11243
rect 6533 -11277 6567 -11243
rect 6613 -11277 6647 -11243
rect 6693 -11277 6727 -11243
rect 6773 -11277 6807 -11243
rect 6853 -11277 6887 -11243
rect 6933 -11277 6967 -11243
rect 7013 -11277 7047 -11243
rect 1184 -11737 1218 -11703
rect 1264 -11737 1298 -11703
rect 1344 -11737 1378 -11703
rect 1424 -11737 1458 -11703
rect 1504 -11737 1538 -11703
rect 1584 -11737 1618 -11703
rect 1664 -11737 1698 -11703
rect 1744 -11737 1778 -11703
rect 1824 -11737 1858 -11703
rect 1904 -11737 1938 -11703
rect 1984 -11737 2018 -11703
rect 2064 -11737 2098 -11703
rect 2144 -11737 2178 -11703
rect 2224 -11737 2258 -11703
rect 2304 -11737 2338 -11703
rect 2384 -11737 2418 -11703
rect 2464 -11737 2498 -11703
rect 2544 -11737 2578 -11703
rect 2624 -11737 2658 -11703
rect 2704 -11737 2738 -11703
rect 2784 -11737 2818 -11703
rect 2864 -11737 2898 -11703
rect 2944 -11737 2978 -11703
rect 3024 -11737 3058 -11703
rect 3104 -11737 3138 -11703
rect 3554 -11737 3588 -11703
rect 3634 -11737 3668 -11703
rect 3714 -11737 3748 -11703
rect 3794 -11737 3828 -11703
rect 3874 -11737 3908 -11703
rect 3954 -11737 3988 -11703
rect 4034 -11737 4068 -11703
rect 4114 -11737 4148 -11703
rect 4194 -11737 4228 -11703
rect 4274 -11737 4308 -11703
rect 4354 -11737 4388 -11703
rect 4434 -11737 4468 -11703
rect 4514 -11737 4548 -11703
rect 4594 -11737 4628 -11703
rect 4674 -11737 4708 -11703
rect 4754 -11737 4788 -11703
rect 4834 -11737 4868 -11703
rect 5274 -11738 5308 -11704
rect 5354 -11738 5388 -11704
rect 5434 -11738 5468 -11704
rect 5514 -11738 5548 -11704
rect 5594 -11738 5628 -11704
rect 5674 -11738 5708 -11704
rect 5754 -11738 5788 -11704
rect 5834 -11738 5868 -11704
rect 5914 -11738 5948 -11704
rect 5994 -11738 6028 -11704
rect 6074 -11738 6108 -11704
rect 6154 -11738 6188 -11704
rect 6234 -11738 6268 -11704
rect 6314 -11738 6348 -11704
rect 6394 -11738 6428 -11704
rect 6474 -11738 6508 -11704
rect 6554 -11738 6588 -11704
rect 6634 -11738 6668 -11704
rect 6714 -11738 6748 -11704
rect 6794 -11738 6828 -11704
rect 6874 -11738 6908 -11704
rect 6954 -11738 6988 -11704
rect 7034 -11738 7068 -11704
rect 7114 -11738 7148 -11704
rect 7194 -11738 7228 -11704
<< poly >>
rect 1410 2348 1490 2371
rect 1410 2314 1433 2348
rect 1467 2314 1490 2348
rect 1920 2361 2100 2391
rect 1920 2331 1950 2361
rect 2070 2331 2100 2361
rect 2220 2361 2400 2391
rect 2220 2331 2250 2361
rect 2370 2331 2400 2361
rect 2800 2348 2880 2371
rect 1410 2291 1490 2314
rect 1290 2248 1370 2271
rect 1290 2214 1313 2248
rect 1347 2214 1370 2248
rect 1290 2191 1370 2214
rect 1090 2048 1170 2071
rect 1090 2014 1113 2048
rect 1147 2014 1170 2048
rect 1090 1991 1170 2014
rect 1140 1771 1170 1991
rect 1290 1771 1320 2191
rect 1440 1771 1470 2291
rect 1540 2148 1620 2171
rect 1540 2114 1563 2148
rect 1597 2114 1620 2148
rect 1540 2091 1620 2114
rect 1590 1771 1620 2091
rect 2800 2314 2823 2348
rect 2857 2314 2880 2348
rect 4240 2361 4420 2391
rect 4240 2331 4270 2361
rect 4390 2331 4420 2361
rect 4540 2361 4720 2391
rect 4540 2331 4570 2361
rect 4690 2331 4720 2361
rect 6260 2361 6440 2391
rect 6260 2331 6290 2361
rect 6410 2331 6440 2361
rect 6560 2361 6740 2391
rect 6560 2331 6590 2361
rect 6710 2331 6740 2361
rect 2800 2291 2880 2314
rect 2700 2048 2780 2071
rect 1920 2001 1950 2031
rect 2070 1876 2100 2031
rect 2220 2001 2250 2031
rect 2370 2001 2400 2031
rect 2700 2014 2723 2048
rect 2757 2014 2780 2048
rect 2170 1978 2250 2001
rect 2170 1944 2193 1978
rect 2227 1944 2250 1978
rect 2170 1921 2250 1944
rect 2070 1853 2150 1876
rect 2070 1819 2093 1853
rect 2127 1819 2150 1853
rect 1920 1771 1950 1801
rect 2070 1796 2150 1819
rect 2070 1771 2100 1796
rect 2220 1771 2250 1921
rect 2700 1991 2780 2014
rect 2370 1771 2400 1801
rect 2700 1771 2730 1991
rect 2850 1771 2880 2291
rect 3000 2248 3080 2271
rect 3000 2214 3023 2248
rect 3057 2214 3080 2248
rect 3000 2191 3080 2214
rect 3000 1771 3030 2191
rect 3150 2148 3230 2171
rect 3150 2114 3173 2148
rect 3207 2114 3230 2148
rect 3150 2091 3230 2114
rect 3150 1771 3180 2091
rect 5170 2218 5250 2241
rect 5170 2184 5193 2218
rect 5227 2184 5250 2218
rect 5170 2161 5250 2184
rect 4970 2098 5050 2121
rect 4970 2064 4993 2098
rect 5027 2064 5050 2098
rect 4970 2041 5050 2064
rect 3860 1998 3940 2021
rect 4240 2001 4270 2031
rect 3860 1964 3883 1998
rect 3917 1964 3940 1998
rect 3860 1941 3940 1964
rect 3710 1898 3790 1921
rect 3710 1864 3733 1898
rect 3767 1864 3790 1898
rect 3710 1841 3790 1864
rect 3760 1771 3790 1841
rect 3910 1771 3940 1941
rect 4390 1876 4420 2031
rect 4540 2001 4570 2031
rect 4690 2001 4720 2031
rect 4490 1978 4570 2001
rect 4490 1944 4513 1978
rect 4547 1944 4570 1978
rect 4490 1921 4570 1944
rect 4390 1853 4470 1876
rect 4390 1819 4413 1853
rect 4447 1819 4470 1853
rect 4240 1771 4270 1801
rect 4390 1796 4470 1819
rect 4390 1771 4420 1796
rect 4540 1771 4570 1921
rect 4690 1771 4720 1801
rect 5020 1771 5050 2041
rect 5170 1771 5200 2161
rect 5880 2028 5960 2051
rect 7140 2248 7220 2271
rect 7140 2214 7163 2248
rect 7197 2214 7220 2248
rect 7140 2191 7220 2214
rect 6990 2128 7070 2151
rect 6990 2094 7013 2128
rect 7047 2094 7070 2128
rect 6990 2071 7070 2094
rect 5880 1994 5903 2028
rect 5937 1994 5960 2028
rect 6260 2001 6290 2031
rect 5880 1971 5960 1994
rect 5730 1928 5810 1951
rect 5730 1894 5753 1928
rect 5787 1894 5810 1928
rect 5730 1871 5810 1894
rect 5780 1771 5810 1871
rect 5930 1771 5960 1971
rect 6410 1876 6440 2031
rect 6560 2001 6590 2031
rect 6710 2001 6740 2031
rect 6510 1978 6590 2001
rect 6510 1944 6533 1978
rect 6567 1944 6590 1978
rect 6510 1921 6590 1944
rect 6410 1853 6490 1876
rect 6410 1819 6433 1853
rect 6467 1819 6490 1853
rect 6260 1771 6290 1801
rect 6410 1796 6490 1819
rect 6410 1771 6440 1796
rect 6560 1771 6590 1921
rect 6710 1771 6740 1801
rect 7040 1771 7070 2071
rect 7190 1771 7220 2191
rect 1140 1441 1170 1471
rect 1290 1441 1320 1471
rect 1440 1441 1470 1471
rect 1590 1441 1620 1471
rect 1920 1441 1950 1471
rect 2070 1441 2100 1471
rect 2220 1441 2250 1471
rect 2370 1441 2400 1471
rect 2700 1441 2730 1471
rect 1920 1418 2000 1441
rect 1920 1384 1943 1418
rect 1977 1384 2000 1418
rect 1920 1361 2000 1384
rect 2320 1418 2400 1441
rect 2850 1431 2880 1471
rect 3000 1431 3030 1471
rect 3150 1431 3180 1471
rect 3760 1441 3790 1471
rect 3910 1441 3940 1471
rect 4240 1441 4270 1471
rect 4390 1441 4420 1471
rect 4540 1441 4570 1471
rect 4690 1441 4720 1471
rect 5020 1441 5050 1471
rect 5170 1441 5200 1471
rect 5780 1441 5810 1471
rect 5930 1441 5960 1471
rect 6260 1441 6290 1471
rect 6410 1441 6440 1471
rect 6560 1441 6590 1471
rect 6710 1441 6740 1471
rect 7040 1441 7070 1471
rect 7190 1441 7220 1471
rect 2320 1384 2343 1418
rect 2377 1384 2400 1418
rect 2320 1361 2400 1384
rect 4240 1418 4320 1441
rect 4240 1384 4263 1418
rect 4297 1384 4320 1418
rect 4240 1361 4320 1384
rect 4640 1418 4720 1441
rect 4640 1384 4663 1418
rect 4697 1384 4720 1418
rect 4640 1361 4720 1384
rect 6260 1418 6340 1441
rect 6260 1384 6283 1418
rect 6317 1384 6340 1418
rect 6260 1361 6340 1384
rect 6660 1418 6740 1441
rect 6660 1384 6683 1418
rect 6717 1384 6740 1418
rect 6660 1361 6740 1384
rect 1920 1178 2000 1201
rect 1920 1144 1943 1178
rect 1977 1144 2000 1178
rect 1920 1121 2000 1144
rect 2320 1178 2400 1201
rect 2320 1144 2343 1178
rect 2377 1144 2400 1178
rect 2320 1121 2400 1144
rect 4240 1178 4320 1201
rect 4240 1144 4263 1178
rect 4297 1144 4320 1178
rect 4240 1121 4320 1144
rect 4640 1178 4720 1201
rect 4640 1144 4663 1178
rect 4697 1144 4720 1178
rect 4640 1121 4720 1144
rect 6260 1178 6340 1201
rect 6260 1144 6283 1178
rect 6317 1144 6340 1178
rect 6260 1121 6340 1144
rect 6660 1178 6740 1201
rect 6660 1144 6683 1178
rect 6717 1144 6740 1178
rect 6660 1121 6740 1144
rect 1440 1091 1470 1121
rect 1590 1091 1620 1121
rect 1920 1091 1950 1121
rect 2070 1091 2100 1121
rect 2220 1091 2250 1121
rect 2370 1091 2400 1121
rect 2700 1091 2730 1121
rect 2850 1091 2880 1121
rect 3760 1091 3790 1121
rect 3910 1091 3940 1121
rect 4240 1091 4270 1121
rect 4390 1091 4420 1121
rect 4540 1091 4570 1121
rect 4690 1091 4720 1121
rect 5020 1091 5050 1121
rect 5170 1091 5200 1121
rect 5780 1091 5810 1121
rect 5930 1091 5960 1121
rect 6260 1091 6290 1121
rect 6410 1091 6440 1121
rect 6560 1091 6590 1121
rect 6710 1091 6740 1121
rect 7040 1091 7070 1121
rect 7190 1091 7220 1121
rect 1440 691 1470 791
rect 1390 668 1470 691
rect 1390 634 1413 668
rect 1447 634 1470 668
rect 1390 611 1470 634
rect 1590 591 1620 791
rect 1920 761 1950 791
rect 2070 766 2100 791
rect 1540 568 1620 591
rect 1540 534 1563 568
rect 1597 534 1620 568
rect 2070 743 2150 766
rect 2070 709 2093 743
rect 2127 709 2150 743
rect 2070 686 2150 709
rect 1540 511 1620 534
rect 1920 531 1950 561
rect 2070 531 2100 686
rect 2220 641 2250 791
rect 2370 761 2400 791
rect 2170 618 2250 641
rect 2170 584 2193 618
rect 2227 584 2250 618
rect 2170 561 2250 584
rect 2220 531 2250 561
rect 2370 531 2400 561
rect 2700 491 2730 791
rect 2650 468 2730 491
rect 2650 434 2673 468
rect 2707 434 2730 468
rect 2650 411 2730 434
rect 2850 371 2880 791
rect 3760 691 3790 791
rect 3710 668 3790 691
rect 3710 634 3733 668
rect 3767 634 3790 668
rect 3710 611 3790 634
rect 3910 591 3940 791
rect 4240 761 4270 791
rect 4390 766 4420 791
rect 3860 568 3940 591
rect 3860 534 3883 568
rect 3917 534 3940 568
rect 4390 743 4470 766
rect 4390 709 4413 743
rect 4447 709 4470 743
rect 4390 686 4470 709
rect 3860 511 3940 534
rect 4240 531 4270 561
rect 4390 531 4420 686
rect 4540 641 4570 791
rect 4690 761 4720 791
rect 4490 618 4570 641
rect 4490 584 4513 618
rect 4547 584 4570 618
rect 4490 561 4570 584
rect 4540 531 4570 561
rect 4690 531 4720 561
rect 2800 348 2880 371
rect 2800 314 2823 348
rect 2857 314 2880 348
rect 2800 291 2880 314
rect 5020 491 5050 791
rect 4970 468 5050 491
rect 4970 434 4993 468
rect 5027 434 5050 468
rect 4970 411 5050 434
rect 5170 371 5200 791
rect 5780 401 5810 791
rect 5930 521 5960 791
rect 6260 761 6290 791
rect 6410 641 6440 791
rect 6560 766 6590 791
rect 6510 743 6590 766
rect 6710 761 6740 791
rect 6510 709 6533 743
rect 6567 709 6590 743
rect 6510 686 6590 709
rect 6410 618 6490 641
rect 6410 584 6433 618
rect 6467 584 6490 618
rect 6410 561 6490 584
rect 6260 531 6290 561
rect 6410 531 6440 561
rect 6560 531 6590 686
rect 7040 621 7070 791
rect 7190 721 7220 791
rect 7190 698 7270 721
rect 7190 664 7213 698
rect 7247 664 7270 698
rect 7190 641 7270 664
rect 7040 598 7120 621
rect 7040 564 7063 598
rect 7097 564 7120 598
rect 6710 531 6740 561
rect 7040 541 7120 564
rect 5930 498 6010 521
rect 5930 464 5953 498
rect 5987 464 6010 498
rect 5930 441 6010 464
rect 5120 348 5200 371
rect 5120 314 5143 348
rect 5177 314 5200 348
rect 5730 378 5810 401
rect 5730 344 5753 378
rect 5787 344 5810 378
rect 5730 321 5810 344
rect 5120 291 5200 314
rect 1920 201 1950 231
rect 2070 201 2100 231
rect 1920 171 2100 201
rect 2220 201 2250 231
rect 2370 201 2400 231
rect 2220 171 2400 201
rect 4240 201 4270 231
rect 4390 201 4420 231
rect 4240 171 4420 201
rect 4540 201 4570 231
rect 4690 201 4720 231
rect 4540 171 4720 201
rect 6260 201 6290 231
rect 6410 201 6440 231
rect 6260 171 6440 201
rect 6560 201 6590 231
rect 6710 201 6740 231
rect 6560 171 6740 201
rect 1410 -472 1490 -449
rect 1410 -506 1433 -472
rect 1467 -506 1490 -472
rect 1920 -459 2100 -429
rect 1920 -489 1950 -459
rect 2070 -489 2100 -459
rect 2220 -459 2400 -429
rect 2220 -489 2250 -459
rect 2370 -489 2400 -459
rect 2800 -472 2880 -449
rect 1410 -529 1490 -506
rect 1290 -572 1370 -549
rect 1290 -606 1313 -572
rect 1347 -606 1370 -572
rect 1290 -629 1370 -606
rect 1090 -772 1170 -749
rect 1090 -806 1113 -772
rect 1147 -806 1170 -772
rect 1090 -829 1170 -806
rect 1140 -1049 1170 -829
rect 1290 -1049 1320 -629
rect 1440 -1049 1470 -529
rect 1540 -672 1620 -649
rect 1540 -706 1563 -672
rect 1597 -706 1620 -672
rect 1540 -729 1620 -706
rect 1590 -1049 1620 -729
rect 2800 -506 2823 -472
rect 2857 -506 2880 -472
rect 4110 -459 4290 -429
rect 4110 -489 4140 -459
rect 4260 -489 4290 -459
rect 4410 -459 4590 -429
rect 4410 -489 4440 -459
rect 4560 -489 4590 -459
rect 5990 -459 6170 -429
rect 5990 -489 6020 -459
rect 6140 -489 6170 -459
rect 6290 -459 6470 -429
rect 6290 -489 6320 -459
rect 6440 -489 6470 -459
rect 2800 -529 2880 -506
rect 2700 -772 2780 -749
rect 1920 -819 1950 -789
rect 2070 -944 2100 -789
rect 2220 -819 2250 -789
rect 2370 -819 2400 -789
rect 2700 -806 2723 -772
rect 2757 -806 2780 -772
rect 2170 -842 2250 -819
rect 2170 -876 2193 -842
rect 2227 -876 2250 -842
rect 2170 -899 2250 -876
rect 2070 -967 2150 -944
rect 2070 -1001 2093 -967
rect 2127 -1001 2150 -967
rect 1920 -1049 1950 -1019
rect 2070 -1024 2150 -1001
rect 2070 -1049 2100 -1024
rect 2220 -1049 2250 -899
rect 2700 -829 2780 -806
rect 2370 -1049 2400 -1019
rect 2700 -1049 2730 -829
rect 2850 -1049 2880 -529
rect 3000 -572 3080 -549
rect 3000 -606 3023 -572
rect 3057 -606 3080 -572
rect 3000 -629 3080 -606
rect 3000 -1049 3030 -629
rect 3150 -672 3230 -649
rect 3150 -706 3173 -672
rect 3207 -706 3230 -672
rect 3150 -729 3230 -706
rect 3150 -1049 3180 -729
rect 4890 -722 4970 -699
rect 4890 -756 4913 -722
rect 4947 -756 4970 -722
rect 4890 -779 4970 -756
rect 4110 -819 4140 -789
rect 3730 -962 3810 -939
rect 3730 -996 3753 -962
rect 3787 -996 3810 -962
rect 3730 -1019 3810 -996
rect 4260 -944 4290 -789
rect 4410 -819 4440 -789
rect 4560 -819 4590 -789
rect 4360 -842 4440 -819
rect 4360 -876 4383 -842
rect 4417 -876 4440 -842
rect 4360 -899 4440 -876
rect 4260 -967 4340 -944
rect 4260 -1001 4283 -967
rect 4317 -1001 4340 -967
rect 3780 -1049 3810 -1019
rect 4110 -1049 4140 -1019
rect 4260 -1024 4340 -1001
rect 4260 -1049 4290 -1024
rect 4410 -1049 4440 -899
rect 4560 -1049 4590 -1019
rect 4890 -1049 4920 -779
rect 5610 -792 5690 -769
rect 6870 -572 6950 -549
rect 6870 -606 6893 -572
rect 6927 -606 6950 -572
rect 6870 -629 6950 -606
rect 6720 -692 6800 -669
rect 6720 -726 6743 -692
rect 6777 -726 6800 -692
rect 6720 -749 6800 -726
rect 5610 -826 5633 -792
rect 5667 -826 5690 -792
rect 5990 -819 6020 -789
rect 5610 -849 5690 -826
rect 5460 -892 5540 -869
rect 5460 -926 5483 -892
rect 5517 -926 5540 -892
rect 5460 -949 5540 -926
rect 5510 -1049 5540 -949
rect 5660 -1049 5690 -849
rect 6140 -944 6170 -789
rect 6290 -819 6320 -789
rect 6440 -819 6470 -789
rect 6240 -842 6320 -819
rect 6240 -876 6263 -842
rect 6297 -876 6320 -842
rect 6240 -899 6320 -876
rect 6140 -967 6220 -944
rect 6140 -1001 6163 -967
rect 6197 -1001 6220 -967
rect 5990 -1049 6020 -1019
rect 6140 -1024 6220 -1001
rect 6140 -1049 6170 -1024
rect 6290 -1049 6320 -899
rect 6440 -1049 6470 -1019
rect 6770 -1049 6800 -749
rect 6920 -1049 6950 -629
rect 1140 -1379 1170 -1349
rect 1290 -1379 1320 -1349
rect 1440 -1379 1470 -1349
rect 1590 -1379 1620 -1349
rect 1920 -1379 1950 -1349
rect 2070 -1379 2100 -1349
rect 2220 -1379 2250 -1349
rect 2370 -1379 2400 -1349
rect 2700 -1379 2730 -1349
rect 1920 -1402 2000 -1379
rect 1920 -1436 1943 -1402
rect 1977 -1436 2000 -1402
rect 1920 -1459 2000 -1436
rect 2320 -1402 2400 -1379
rect 2850 -1389 2880 -1349
rect 3000 -1389 3030 -1349
rect 3150 -1389 3180 -1349
rect 3780 -1379 3810 -1349
rect 4110 -1379 4140 -1349
rect 4260 -1379 4290 -1349
rect 4410 -1379 4440 -1349
rect 4560 -1379 4590 -1349
rect 4890 -1379 4920 -1349
rect 5510 -1379 5540 -1349
rect 5660 -1379 5690 -1349
rect 5990 -1379 6020 -1349
rect 6140 -1379 6170 -1349
rect 6290 -1379 6320 -1349
rect 6440 -1379 6470 -1349
rect 6770 -1379 6800 -1349
rect 6920 -1379 6950 -1349
rect 2320 -1436 2343 -1402
rect 2377 -1436 2400 -1402
rect 2320 -1459 2400 -1436
rect 4110 -1402 4190 -1379
rect 4110 -1436 4133 -1402
rect 4167 -1436 4190 -1402
rect 4110 -1459 4190 -1436
rect 4510 -1402 4590 -1379
rect 4510 -1436 4533 -1402
rect 4567 -1436 4590 -1402
rect 4510 -1459 4590 -1436
rect 5990 -1402 6070 -1379
rect 5990 -1436 6013 -1402
rect 6047 -1436 6070 -1402
rect 5990 -1459 6070 -1436
rect 6390 -1402 6470 -1379
rect 6390 -1436 6413 -1402
rect 6447 -1436 6470 -1402
rect 6390 -1459 6470 -1436
rect 1920 -1642 2000 -1619
rect 1920 -1676 1943 -1642
rect 1977 -1676 2000 -1642
rect 1920 -1699 2000 -1676
rect 2320 -1642 2400 -1619
rect 2320 -1676 2343 -1642
rect 2377 -1676 2400 -1642
rect 2320 -1699 2400 -1676
rect 4110 -1642 4190 -1619
rect 4110 -1676 4133 -1642
rect 4167 -1676 4190 -1642
rect 1140 -1729 1170 -1699
rect 1290 -1729 1320 -1699
rect 1440 -1729 1470 -1699
rect 1590 -1729 1620 -1699
rect 1920 -1729 1950 -1699
rect 2070 -1729 2100 -1699
rect 2220 -1729 2250 -1699
rect 2370 -1729 2400 -1699
rect 2700 -1729 2730 -1699
rect 2850 -1729 2880 -1689
rect 3000 -1729 3030 -1689
rect 3150 -1729 3180 -1689
rect 4110 -1699 4190 -1676
rect 4510 -1642 4590 -1619
rect 4510 -1676 4533 -1642
rect 4567 -1676 4590 -1642
rect 4510 -1699 4590 -1676
rect 5990 -1642 6070 -1619
rect 5990 -1676 6013 -1642
rect 6047 -1676 6070 -1642
rect 5990 -1699 6070 -1676
rect 6390 -1642 6470 -1619
rect 6390 -1676 6413 -1642
rect 6447 -1676 6470 -1642
rect 6390 -1699 6470 -1676
rect 3780 -1729 3810 -1699
rect 4110 -1729 4140 -1699
rect 4260 -1729 4290 -1699
rect 4410 -1729 4440 -1699
rect 4560 -1729 4590 -1699
rect 4890 -1729 4920 -1699
rect 5510 -1729 5540 -1699
rect 5660 -1729 5690 -1699
rect 5990 -1729 6020 -1699
rect 6140 -1729 6170 -1699
rect 6290 -1729 6320 -1699
rect 6440 -1729 6470 -1699
rect 6770 -1729 6800 -1699
rect 6920 -1729 6950 -1699
rect 1140 -2249 1170 -2029
rect 1090 -2272 1170 -2249
rect 1090 -2306 1113 -2272
rect 1147 -2306 1170 -2272
rect 1090 -2329 1170 -2306
rect 1290 -2449 1320 -2029
rect 1290 -2472 1370 -2449
rect 1290 -2506 1313 -2472
rect 1347 -2506 1370 -2472
rect 1290 -2529 1370 -2506
rect 1440 -2549 1470 -2029
rect 1590 -2349 1620 -2029
rect 1920 -2059 1950 -2029
rect 2070 -2054 2100 -2029
rect 2070 -2077 2150 -2054
rect 2070 -2111 2093 -2077
rect 2127 -2111 2150 -2077
rect 2070 -2134 2150 -2111
rect 1920 -2289 1950 -2259
rect 2070 -2289 2100 -2134
rect 2220 -2179 2250 -2029
rect 2370 -2059 2400 -2029
rect 2170 -2202 2250 -2179
rect 2170 -2236 2193 -2202
rect 2227 -2236 2250 -2202
rect 2170 -2259 2250 -2236
rect 2700 -2249 2730 -2029
rect 2220 -2289 2250 -2259
rect 2370 -2289 2400 -2259
rect 2700 -2272 2780 -2249
rect 1540 -2372 1620 -2349
rect 1540 -2406 1563 -2372
rect 1597 -2406 1620 -2372
rect 1540 -2429 1620 -2406
rect 1410 -2572 1490 -2549
rect 1410 -2606 1433 -2572
rect 1467 -2606 1490 -2572
rect 2700 -2306 2723 -2272
rect 2757 -2306 2780 -2272
rect 2700 -2329 2780 -2306
rect 2850 -2549 2880 -2029
rect 3000 -2449 3030 -2029
rect 3150 -2349 3180 -2029
rect 3780 -2059 3810 -2029
rect 4110 -2059 4140 -2029
rect 4260 -2054 4290 -2029
rect 3730 -2082 3810 -2059
rect 3730 -2116 3753 -2082
rect 3787 -2116 3810 -2082
rect 3730 -2139 3810 -2116
rect 4260 -2077 4340 -2054
rect 4260 -2111 4283 -2077
rect 4317 -2111 4340 -2077
rect 4260 -2134 4340 -2111
rect 4110 -2289 4140 -2259
rect 4260 -2289 4290 -2134
rect 4410 -2179 4440 -2029
rect 4560 -2059 4590 -2029
rect 4360 -2202 4440 -2179
rect 4360 -2236 4383 -2202
rect 4417 -2236 4440 -2202
rect 4360 -2259 4440 -2236
rect 4410 -2289 4440 -2259
rect 4560 -2289 4590 -2259
rect 3150 -2372 3230 -2349
rect 3150 -2406 3173 -2372
rect 3207 -2406 3230 -2372
rect 3150 -2429 3230 -2406
rect 3000 -2472 3080 -2449
rect 3000 -2506 3023 -2472
rect 3057 -2506 3080 -2472
rect 3000 -2529 3080 -2506
rect 2800 -2572 2880 -2549
rect 1410 -2629 1490 -2606
rect 1920 -2619 1950 -2589
rect 2070 -2619 2100 -2589
rect 1920 -2649 2100 -2619
rect 2220 -2619 2250 -2589
rect 2370 -2619 2400 -2589
rect 2220 -2649 2400 -2619
rect 2800 -2606 2823 -2572
rect 2857 -2606 2880 -2572
rect 4890 -2299 4920 -2029
rect 5510 -2129 5540 -2029
rect 5460 -2152 5540 -2129
rect 5460 -2186 5483 -2152
rect 5517 -2186 5540 -2152
rect 5460 -2209 5540 -2186
rect 5660 -2229 5690 -2029
rect 5990 -2059 6020 -2029
rect 6140 -2054 6170 -2029
rect 5610 -2252 5690 -2229
rect 5610 -2286 5633 -2252
rect 5667 -2286 5690 -2252
rect 6140 -2077 6220 -2054
rect 6140 -2111 6163 -2077
rect 6197 -2111 6220 -2077
rect 6140 -2134 6220 -2111
rect 4890 -2322 4970 -2299
rect 5610 -2309 5690 -2286
rect 5990 -2289 6020 -2259
rect 6140 -2289 6170 -2134
rect 6290 -2179 6320 -2029
rect 6440 -2059 6470 -2029
rect 6240 -2202 6320 -2179
rect 6240 -2236 6263 -2202
rect 6297 -2236 6320 -2202
rect 6240 -2259 6320 -2236
rect 6290 -2289 6320 -2259
rect 6440 -2289 6470 -2259
rect 4890 -2356 4913 -2322
rect 4947 -2356 4970 -2322
rect 4890 -2379 4970 -2356
rect 6770 -2329 6800 -2029
rect 6720 -2352 6800 -2329
rect 6720 -2386 6743 -2352
rect 6777 -2386 6800 -2352
rect 6720 -2409 6800 -2386
rect 6920 -2449 6950 -2029
rect 6870 -2472 6950 -2449
rect 6870 -2506 6893 -2472
rect 6927 -2506 6950 -2472
rect 6870 -2529 6950 -2506
rect 2800 -2629 2880 -2606
rect 4110 -2619 4140 -2589
rect 4260 -2619 4290 -2589
rect 4110 -2649 4290 -2619
rect 4410 -2619 4440 -2589
rect 4560 -2619 4590 -2589
rect 4410 -2649 4590 -2619
rect 5990 -2619 6020 -2589
rect 6140 -2619 6170 -2589
rect 5990 -2649 6170 -2619
rect 6290 -2619 6320 -2589
rect 6440 -2619 6470 -2589
rect 6290 -2649 6470 -2619
rect 1921 -3279 2101 -3249
rect 1921 -3309 1951 -3279
rect 2071 -3309 2101 -3279
rect 2221 -3279 2401 -3249
rect 2221 -3309 2251 -3279
rect 2371 -3309 2401 -3279
rect 2951 -3282 3031 -3259
rect 2951 -3316 2974 -3282
rect 3008 -3316 3031 -3282
rect 3971 -3279 4151 -3249
rect 3971 -3309 4001 -3279
rect 4121 -3309 4151 -3279
rect 4271 -3279 4451 -3249
rect 4271 -3309 4301 -3279
rect 4421 -3309 4451 -3279
rect 5381 -3288 5461 -3265
rect 2951 -3339 3031 -3316
rect 2801 -3402 2881 -3379
rect 2801 -3436 2824 -3402
rect 2858 -3436 2881 -3402
rect 2801 -3459 2881 -3436
rect 2671 -3522 2751 -3499
rect 2671 -3556 2694 -3522
rect 2728 -3556 2751 -3522
rect 2671 -3579 2751 -3556
rect 1921 -3639 1951 -3609
rect 1371 -3692 1471 -3669
rect 1371 -3726 1394 -3692
rect 1428 -3726 1471 -3692
rect 1371 -3749 1471 -3726
rect 1541 -3672 1621 -3649
rect 1541 -3706 1564 -3672
rect 1598 -3706 1621 -3672
rect 1541 -3729 1621 -3706
rect 1241 -3772 1321 -3749
rect 1241 -3806 1264 -3772
rect 1298 -3806 1321 -3772
rect 1241 -3829 1321 -3806
rect 1291 -3869 1321 -3829
rect 1441 -3869 1471 -3749
rect 1591 -3869 1621 -3729
rect 2071 -3764 2101 -3609
rect 2221 -3639 2251 -3609
rect 2371 -3639 2401 -3609
rect 2171 -3662 2251 -3639
rect 2171 -3696 2194 -3662
rect 2228 -3696 2251 -3662
rect 2171 -3719 2251 -3696
rect 2071 -3787 2151 -3764
rect 2071 -3821 2094 -3787
rect 2128 -3821 2151 -3787
rect 1921 -3869 1951 -3839
rect 2071 -3844 2151 -3821
rect 2071 -3869 2101 -3844
rect 2221 -3869 2251 -3719
rect 2371 -3869 2401 -3839
rect 2701 -3869 2731 -3579
rect 2851 -3869 2881 -3459
rect 3001 -3869 3031 -3339
rect 5381 -3322 5404 -3288
rect 5438 -3322 5461 -3288
rect 6011 -3280 6191 -3250
rect 6011 -3310 6041 -3280
rect 6161 -3310 6191 -3280
rect 6311 -3280 6491 -3250
rect 6311 -3310 6341 -3280
rect 6461 -3310 6491 -3280
rect 5381 -3345 5461 -3322
rect 4751 -3542 4831 -3519
rect 4751 -3576 4774 -3542
rect 4808 -3576 4831 -3542
rect 4751 -3599 4831 -3576
rect 3971 -3639 4001 -3609
rect 3591 -3782 3671 -3759
rect 3591 -3816 3614 -3782
rect 3648 -3816 3671 -3782
rect 3591 -3839 3671 -3816
rect 4121 -3764 4151 -3609
rect 4271 -3639 4301 -3609
rect 4421 -3639 4451 -3609
rect 4221 -3662 4301 -3639
rect 4221 -3696 4244 -3662
rect 4278 -3696 4301 -3662
rect 4221 -3719 4301 -3696
rect 4121 -3787 4201 -3764
rect 4121 -3821 4144 -3787
rect 4178 -3821 4201 -3787
rect 3641 -3869 3671 -3839
rect 3971 -3869 4001 -3839
rect 4121 -3844 4201 -3821
rect 4121 -3869 4151 -3844
rect 4271 -3869 4301 -3719
rect 4421 -3869 4451 -3839
rect 4751 -3869 4781 -3599
rect 5381 -3870 5411 -3345
rect 5481 -3413 5561 -3390
rect 5481 -3447 5504 -3413
rect 5538 -3447 5561 -3413
rect 5481 -3470 5561 -3447
rect 5531 -3870 5561 -3470
rect 5681 -3503 5761 -3480
rect 5681 -3537 5704 -3503
rect 5738 -3537 5761 -3503
rect 5681 -3560 5761 -3537
rect 5681 -3870 5711 -3560
rect 6011 -3640 6041 -3610
rect 6161 -3640 6191 -3610
rect 6161 -3663 6241 -3640
rect 6161 -3697 6184 -3663
rect 6218 -3697 6241 -3663
rect 6161 -3720 6241 -3697
rect 6011 -3870 6041 -3840
rect 6161 -3870 6191 -3720
rect 6311 -3765 6341 -3610
rect 6461 -3640 6491 -3610
rect 7081 -3613 7161 -3590
rect 7081 -3647 7104 -3613
rect 7138 -3647 7161 -3613
rect 7081 -3670 7161 -3647
rect 6261 -3788 6341 -3765
rect 6941 -3713 7021 -3690
rect 6941 -3747 6964 -3713
rect 6998 -3747 7021 -3713
rect 6941 -3770 7021 -3747
rect 6261 -3822 6284 -3788
rect 6318 -3822 6341 -3788
rect 6261 -3845 6341 -3822
rect 6791 -3793 6871 -3770
rect 6791 -3827 6814 -3793
rect 6848 -3827 6871 -3793
rect 6311 -3870 6341 -3845
rect 6461 -3870 6491 -3840
rect 6791 -3850 6871 -3827
rect 6791 -3870 6821 -3850
rect 6941 -3870 6971 -3770
rect 7091 -3870 7121 -3670
rect 1291 -4199 1321 -4169
rect 1441 -4199 1471 -4169
rect 1591 -4199 1621 -4169
rect 1921 -4199 1951 -4169
rect 2071 -4199 2101 -4169
rect 2221 -4199 2251 -4169
rect 2371 -4199 2401 -4169
rect 2701 -4199 2731 -4169
rect 2851 -4199 2881 -4169
rect 3001 -4199 3031 -4169
rect 3641 -4199 3671 -4169
rect 3971 -4199 4001 -4169
rect 4121 -4199 4151 -4169
rect 4271 -4199 4301 -4169
rect 4421 -4199 4451 -4169
rect 4751 -4199 4781 -4169
rect 1921 -4222 2001 -4199
rect 1921 -4256 1944 -4222
rect 1978 -4256 2001 -4222
rect 1921 -4279 2001 -4256
rect 2321 -4222 2401 -4199
rect 2321 -4256 2344 -4222
rect 2378 -4256 2401 -4222
rect 2321 -4279 2401 -4256
rect 3971 -4222 4051 -4199
rect 3971 -4256 3994 -4222
rect 4028 -4256 4051 -4222
rect 3971 -4279 4051 -4256
rect 4371 -4222 4451 -4199
rect 5381 -4200 5411 -4170
rect 5531 -4200 5561 -4170
rect 5681 -4200 5711 -4170
rect 6011 -4200 6041 -4170
rect 6161 -4200 6191 -4170
rect 6311 -4200 6341 -4170
rect 6461 -4200 6491 -4170
rect 6791 -4200 6821 -4170
rect 6941 -4200 6971 -4170
rect 7091 -4200 7121 -4170
rect 4371 -4256 4394 -4222
rect 4428 -4256 4451 -4222
rect 4371 -4279 4451 -4256
rect 6011 -4223 6091 -4200
rect 6011 -4257 6034 -4223
rect 6068 -4257 6091 -4223
rect 6011 -4280 6091 -4257
rect 6411 -4223 6491 -4200
rect 6411 -4257 6434 -4223
rect 6468 -4257 6491 -4223
rect 6411 -4280 6491 -4257
rect 1960 -4542 2040 -4519
rect 1960 -4576 1983 -4542
rect 2017 -4576 2040 -4542
rect 1960 -4599 2040 -4576
rect 2360 -4542 2440 -4519
rect 2360 -4576 2383 -4542
rect 2417 -4576 2440 -4542
rect 2360 -4599 2440 -4576
rect 4171 -4543 4251 -4520
rect 4171 -4577 4194 -4543
rect 4228 -4577 4251 -4543
rect 1180 -4629 1210 -4599
rect 1330 -4629 1360 -4599
rect 1480 -4629 1510 -4599
rect 1630 -4629 1660 -4599
rect 1960 -4629 1990 -4599
rect 2110 -4629 2140 -4599
rect 2260 -4629 2290 -4599
rect 2410 -4629 2440 -4599
rect 2740 -4629 2770 -4599
rect 2890 -4629 2920 -4599
rect 3040 -4629 3070 -4599
rect 3190 -4629 3220 -4599
rect 4171 -4600 4251 -4577
rect 4571 -4543 4651 -4520
rect 4571 -4577 4594 -4543
rect 4628 -4577 4651 -4543
rect 4571 -4600 4651 -4577
rect 6230 -4543 6310 -4520
rect 6230 -4577 6253 -4543
rect 6287 -4577 6310 -4543
rect 6230 -4600 6310 -4577
rect 6630 -4543 6710 -4520
rect 6630 -4577 6653 -4543
rect 6687 -4577 6710 -4543
rect 6630 -4600 6710 -4577
rect 3841 -4630 3871 -4600
rect 4171 -4630 4201 -4600
rect 4321 -4630 4351 -4600
rect 4471 -4630 4501 -4600
rect 4621 -4630 4651 -4600
rect 4951 -4630 4981 -4600
rect 5600 -4630 5630 -4600
rect 5750 -4630 5780 -4600
rect 5900 -4630 5930 -4600
rect 6230 -4630 6260 -4600
rect 6380 -4630 6410 -4600
rect 6530 -4630 6560 -4600
rect 6680 -4630 6710 -4600
rect 7010 -4630 7040 -4600
rect 7160 -4630 7190 -4600
rect 7310 -4630 7340 -4600
rect 1180 -5009 1210 -4929
rect 1130 -5032 1210 -5009
rect 1130 -5066 1153 -5032
rect 1187 -5066 1210 -5032
rect 1130 -5089 1210 -5066
rect 1330 -5109 1360 -4929
rect 1280 -5132 1360 -5109
rect 1280 -5166 1303 -5132
rect 1337 -5166 1360 -5132
rect 1280 -5189 1360 -5166
rect 1480 -5209 1510 -4929
rect 1430 -5232 1510 -5209
rect 1430 -5266 1453 -5232
rect 1487 -5266 1510 -5232
rect 1430 -5289 1510 -5266
rect 1630 -5309 1660 -4929
rect 1960 -4959 1990 -4929
rect 1580 -5332 1660 -5309
rect 1580 -5366 1603 -5332
rect 1637 -5366 1660 -5332
rect 1580 -5389 1660 -5366
rect 2110 -5169 2140 -4929
rect 2110 -5192 2190 -5169
rect 2110 -5226 2133 -5192
rect 2167 -5226 2190 -5192
rect 2110 -5249 2190 -5226
rect 1960 -5509 1990 -5479
rect 2110 -5509 2140 -5249
rect 2260 -5309 2290 -4929
rect 2410 -4959 2440 -4929
rect 2740 -5009 2770 -4929
rect 2890 -5009 2920 -4929
rect 3040 -5009 3070 -4929
rect 3190 -5009 3220 -4929
rect 3841 -4960 3871 -4930
rect 4171 -4960 4201 -4930
rect 4321 -4955 4351 -4930
rect 2690 -5032 2770 -5009
rect 2690 -5066 2713 -5032
rect 2747 -5066 2770 -5032
rect 2690 -5089 2770 -5066
rect 2840 -5032 2920 -5009
rect 2840 -5066 2863 -5032
rect 2897 -5066 2920 -5032
rect 2840 -5089 2920 -5066
rect 2990 -5032 3070 -5009
rect 2990 -5066 3013 -5032
rect 3047 -5066 3070 -5032
rect 2990 -5089 3070 -5066
rect 3140 -5032 3220 -5009
rect 3140 -5066 3163 -5032
rect 3197 -5066 3220 -5032
rect 3791 -4983 3871 -4960
rect 3791 -5017 3814 -4983
rect 3848 -5017 3871 -4983
rect 3791 -5040 3871 -5017
rect 4321 -4978 4401 -4955
rect 4321 -5012 4344 -4978
rect 4378 -5012 4401 -4978
rect 4321 -5035 4401 -5012
rect 3140 -5089 3220 -5066
rect 4171 -5190 4201 -5160
rect 4321 -5190 4351 -5035
rect 4471 -5080 4501 -4930
rect 4621 -4960 4651 -4930
rect 4421 -5103 4501 -5080
rect 4421 -5137 4444 -5103
rect 4478 -5137 4501 -5103
rect 4421 -5160 4501 -5137
rect 4471 -5190 4501 -5160
rect 4621 -5190 4651 -5160
rect 2210 -5332 2290 -5309
rect 2210 -5366 2233 -5332
rect 2267 -5366 2290 -5332
rect 2210 -5389 2290 -5366
rect 2260 -5509 2290 -5389
rect 2410 -5509 2440 -5479
rect 4951 -5200 4981 -4930
rect 4951 -5223 5031 -5200
rect 4951 -5257 4974 -5223
rect 5008 -5257 5031 -5223
rect 4951 -5280 5031 -5257
rect 5600 -5455 5630 -4930
rect 5750 -5330 5780 -4930
rect 5900 -5240 5930 -4930
rect 6230 -4960 6260 -4930
rect 6380 -5080 6410 -4930
rect 6530 -4955 6560 -4930
rect 6480 -4978 6560 -4955
rect 6680 -4960 6710 -4930
rect 7010 -4950 7040 -4930
rect 6480 -5012 6503 -4978
rect 6537 -5012 6560 -4978
rect 6480 -5035 6560 -5012
rect 7010 -4973 7090 -4950
rect 7010 -5007 7033 -4973
rect 7067 -5007 7090 -4973
rect 7010 -5030 7090 -5007
rect 7160 -5030 7190 -4930
rect 6380 -5103 6460 -5080
rect 6380 -5137 6403 -5103
rect 6437 -5137 6460 -5103
rect 6380 -5160 6460 -5137
rect 6230 -5190 6260 -5160
rect 6380 -5190 6410 -5160
rect 6530 -5190 6560 -5035
rect 7160 -5053 7240 -5030
rect 7160 -5087 7183 -5053
rect 7217 -5087 7240 -5053
rect 7160 -5110 7240 -5087
rect 7310 -5130 7340 -4930
rect 7300 -5153 7380 -5130
rect 6680 -5190 6710 -5160
rect 7300 -5187 7323 -5153
rect 7357 -5187 7380 -5153
rect 5900 -5263 5980 -5240
rect 5900 -5297 5923 -5263
rect 5957 -5297 5980 -5263
rect 5900 -5320 5980 -5297
rect 5700 -5353 5780 -5330
rect 5700 -5387 5723 -5353
rect 5757 -5387 5780 -5353
rect 5700 -5410 5780 -5387
rect 5600 -5478 5680 -5455
rect 4171 -5520 4201 -5490
rect 4321 -5520 4351 -5490
rect 4171 -5550 4351 -5520
rect 4471 -5520 4501 -5490
rect 4621 -5520 4651 -5490
rect 4471 -5550 4651 -5520
rect 5600 -5512 5623 -5478
rect 5657 -5512 5680 -5478
rect 7300 -5210 7380 -5187
rect 5600 -5535 5680 -5512
rect 6230 -5520 6260 -5490
rect 6380 -5520 6410 -5490
rect 6230 -5550 6410 -5520
rect 6530 -5520 6560 -5490
rect 6680 -5520 6710 -5490
rect 6530 -5550 6710 -5520
rect 1960 -5839 1990 -5809
rect 2110 -5839 2140 -5809
rect 1960 -5869 2140 -5839
rect 2260 -5839 2290 -5809
rect 2410 -5839 2440 -5809
rect 2260 -5869 2440 -5839
rect 1450 -6193 1530 -6170
rect 1450 -6227 1473 -6193
rect 1507 -6227 1530 -6193
rect 1960 -6180 2140 -6150
rect 1960 -6210 1990 -6180
rect 2110 -6210 2140 -6180
rect 2260 -6180 2440 -6150
rect 2260 -6210 2290 -6180
rect 2410 -6210 2440 -6180
rect 2840 -6193 2920 -6170
rect 1450 -6250 1530 -6227
rect 1330 -6293 1410 -6270
rect 1330 -6327 1353 -6293
rect 1387 -6327 1410 -6293
rect 1330 -6350 1410 -6327
rect 1130 -6493 1210 -6470
rect 1130 -6527 1153 -6493
rect 1187 -6527 1210 -6493
rect 1130 -6550 1210 -6527
rect 1180 -6770 1210 -6550
rect 1330 -6770 1360 -6350
rect 1480 -6770 1510 -6250
rect 1580 -6393 1660 -6370
rect 1580 -6427 1603 -6393
rect 1637 -6427 1660 -6393
rect 1580 -6450 1660 -6427
rect 1630 -6770 1660 -6450
rect 2840 -6227 2863 -6193
rect 2897 -6227 2920 -6193
rect 4170 -6180 4350 -6150
rect 4170 -6210 4200 -6180
rect 4320 -6210 4350 -6180
rect 4470 -6180 4650 -6150
rect 4470 -6210 4500 -6180
rect 4620 -6210 4650 -6180
rect 6049 -6180 6229 -6150
rect 6049 -6210 6079 -6180
rect 6199 -6210 6229 -6180
rect 6349 -6180 6529 -6150
rect 6349 -6210 6379 -6180
rect 6499 -6210 6529 -6180
rect 2840 -6250 2920 -6227
rect 2740 -6493 2820 -6470
rect 1960 -6540 1990 -6510
rect 2110 -6665 2140 -6510
rect 2260 -6540 2290 -6510
rect 2410 -6540 2440 -6510
rect 2740 -6527 2763 -6493
rect 2797 -6527 2820 -6493
rect 2210 -6563 2290 -6540
rect 2210 -6597 2233 -6563
rect 2267 -6597 2290 -6563
rect 2210 -6620 2290 -6597
rect 2110 -6688 2190 -6665
rect 2110 -6722 2133 -6688
rect 2167 -6722 2190 -6688
rect 1960 -6770 1990 -6740
rect 2110 -6745 2190 -6722
rect 2110 -6770 2140 -6745
rect 2260 -6770 2290 -6620
rect 2740 -6550 2820 -6527
rect 2410 -6770 2440 -6740
rect 2740 -6770 2770 -6550
rect 2890 -6770 2920 -6250
rect 3040 -6293 3120 -6270
rect 3040 -6327 3063 -6293
rect 3097 -6327 3120 -6293
rect 3040 -6350 3120 -6327
rect 3040 -6770 3070 -6350
rect 3190 -6393 3270 -6370
rect 3190 -6427 3213 -6393
rect 3247 -6427 3270 -6393
rect 3190 -6450 3270 -6427
rect 3190 -6770 3220 -6450
rect 4950 -6443 5030 -6420
rect 4950 -6477 4973 -6443
rect 5007 -6477 5030 -6443
rect 4950 -6500 5030 -6477
rect 4170 -6540 4200 -6510
rect 3790 -6683 3870 -6660
rect 3790 -6717 3813 -6683
rect 3847 -6717 3870 -6683
rect 3790 -6740 3870 -6717
rect 4320 -6665 4350 -6510
rect 4470 -6540 4500 -6510
rect 4620 -6540 4650 -6510
rect 4420 -6563 4500 -6540
rect 4420 -6597 4443 -6563
rect 4477 -6597 4500 -6563
rect 4420 -6620 4500 -6597
rect 4320 -6688 4400 -6665
rect 4320 -6722 4343 -6688
rect 4377 -6722 4400 -6688
rect 3840 -6770 3870 -6740
rect 4170 -6770 4200 -6740
rect 4320 -6745 4400 -6722
rect 4320 -6770 4350 -6745
rect 4470 -6770 4500 -6620
rect 4620 -6770 4650 -6740
rect 4950 -6770 4980 -6500
rect 5669 -6513 5749 -6490
rect 6929 -6293 7009 -6270
rect 6929 -6327 6952 -6293
rect 6986 -6327 7009 -6293
rect 6929 -6350 7009 -6327
rect 6779 -6413 6859 -6390
rect 6779 -6447 6802 -6413
rect 6836 -6447 6859 -6413
rect 6779 -6470 6859 -6447
rect 5669 -6547 5692 -6513
rect 5726 -6547 5749 -6513
rect 6049 -6540 6079 -6510
rect 5669 -6570 5749 -6547
rect 5519 -6613 5599 -6590
rect 5519 -6647 5542 -6613
rect 5576 -6647 5599 -6613
rect 5519 -6670 5599 -6647
rect 5569 -6770 5599 -6670
rect 5719 -6770 5749 -6570
rect 6199 -6665 6229 -6510
rect 6349 -6540 6379 -6510
rect 6499 -6540 6529 -6510
rect 6299 -6563 6379 -6540
rect 6299 -6597 6322 -6563
rect 6356 -6597 6379 -6563
rect 6299 -6620 6379 -6597
rect 6199 -6688 6279 -6665
rect 6199 -6722 6222 -6688
rect 6256 -6722 6279 -6688
rect 6049 -6770 6079 -6740
rect 6199 -6745 6279 -6722
rect 6199 -6770 6229 -6745
rect 6349 -6770 6379 -6620
rect 6499 -6770 6529 -6740
rect 6829 -6770 6859 -6470
rect 6979 -6770 7009 -6350
rect 1180 -7100 1210 -7070
rect 1330 -7100 1360 -7070
rect 1480 -7100 1510 -7070
rect 1630 -7100 1660 -7070
rect 1960 -7100 1990 -7070
rect 2110 -7100 2140 -7070
rect 2260 -7100 2290 -7070
rect 2410 -7100 2440 -7070
rect 2740 -7100 2770 -7070
rect 1960 -7123 2040 -7100
rect 1960 -7157 1983 -7123
rect 2017 -7157 2040 -7123
rect 1960 -7180 2040 -7157
rect 2360 -7123 2440 -7100
rect 2890 -7110 2920 -7070
rect 3040 -7110 3070 -7070
rect 3190 -7110 3220 -7070
rect 3840 -7100 3870 -7070
rect 4170 -7100 4200 -7070
rect 4320 -7100 4350 -7070
rect 4470 -7100 4500 -7070
rect 4620 -7100 4650 -7070
rect 4950 -7100 4980 -7070
rect 5569 -7100 5599 -7070
rect 5719 -7100 5749 -7070
rect 6049 -7100 6079 -7070
rect 6199 -7100 6229 -7070
rect 6349 -7100 6379 -7070
rect 6499 -7100 6529 -7070
rect 6829 -7100 6859 -7070
rect 6979 -7100 7009 -7070
rect 2360 -7157 2383 -7123
rect 2417 -7157 2440 -7123
rect 2360 -7180 2440 -7157
rect 4170 -7123 4250 -7100
rect 4170 -7157 4193 -7123
rect 4227 -7157 4250 -7123
rect 4170 -7180 4250 -7157
rect 4570 -7123 4650 -7100
rect 4570 -7157 4593 -7123
rect 4627 -7157 4650 -7123
rect 4570 -7180 4650 -7157
rect 6049 -7123 6129 -7100
rect 6049 -7157 6072 -7123
rect 6106 -7157 6129 -7123
rect 6049 -7180 6129 -7157
rect 6449 -7123 6529 -7100
rect 6449 -7157 6472 -7123
rect 6506 -7157 6529 -7123
rect 6449 -7180 6529 -7157
rect 1960 -7363 2040 -7340
rect 1960 -7397 1983 -7363
rect 2017 -7397 2040 -7363
rect 1960 -7420 2040 -7397
rect 2360 -7363 2440 -7340
rect 2360 -7397 2383 -7363
rect 2417 -7397 2440 -7363
rect 2360 -7420 2440 -7397
rect 4170 -7363 4250 -7340
rect 4170 -7397 4193 -7363
rect 4227 -7397 4250 -7363
rect 1180 -7450 1210 -7420
rect 1330 -7450 1360 -7420
rect 1480 -7450 1510 -7420
rect 1630 -7450 1660 -7420
rect 1960 -7450 1990 -7420
rect 2110 -7450 2140 -7420
rect 2260 -7450 2290 -7420
rect 2410 -7450 2440 -7420
rect 2740 -7450 2770 -7420
rect 2890 -7450 2920 -7410
rect 3040 -7450 3070 -7410
rect 3190 -7450 3220 -7410
rect 4170 -7420 4250 -7397
rect 4570 -7363 4650 -7340
rect 4570 -7397 4593 -7363
rect 4627 -7397 4650 -7363
rect 4570 -7420 4650 -7397
rect 6049 -7363 6129 -7340
rect 6049 -7397 6072 -7363
rect 6106 -7397 6129 -7363
rect 6049 -7420 6129 -7397
rect 6449 -7363 6529 -7340
rect 6449 -7397 6472 -7363
rect 6506 -7397 6529 -7363
rect 6449 -7420 6529 -7397
rect 3840 -7450 3870 -7420
rect 4170 -7450 4200 -7420
rect 4320 -7450 4350 -7420
rect 4470 -7450 4500 -7420
rect 4620 -7450 4650 -7420
rect 4950 -7450 4980 -7420
rect 5569 -7450 5599 -7420
rect 5719 -7450 5749 -7420
rect 6049 -7450 6079 -7420
rect 6199 -7450 6229 -7420
rect 6349 -7450 6379 -7420
rect 6499 -7450 6529 -7420
rect 6829 -7450 6859 -7420
rect 6979 -7450 7009 -7420
rect 1180 -7970 1210 -7750
rect 1130 -7993 1210 -7970
rect 1130 -8027 1153 -7993
rect 1187 -8027 1210 -7993
rect 1130 -8050 1210 -8027
rect 1330 -8170 1360 -7750
rect 1330 -8193 1410 -8170
rect 1330 -8227 1353 -8193
rect 1387 -8227 1410 -8193
rect 1330 -8250 1410 -8227
rect 1480 -8270 1510 -7750
rect 1630 -8070 1660 -7750
rect 1960 -7780 1990 -7750
rect 2110 -7775 2140 -7750
rect 2110 -7798 2190 -7775
rect 2110 -7832 2133 -7798
rect 2167 -7832 2190 -7798
rect 2110 -7855 2190 -7832
rect 1960 -8010 1990 -7980
rect 2110 -8010 2140 -7855
rect 2260 -7900 2290 -7750
rect 2410 -7780 2440 -7750
rect 2210 -7923 2290 -7900
rect 2210 -7957 2233 -7923
rect 2267 -7957 2290 -7923
rect 2210 -7980 2290 -7957
rect 2740 -7970 2770 -7750
rect 2260 -8010 2290 -7980
rect 2410 -8010 2440 -7980
rect 2740 -7993 2820 -7970
rect 1580 -8093 1660 -8070
rect 1580 -8127 1603 -8093
rect 1637 -8127 1660 -8093
rect 1580 -8150 1660 -8127
rect 1450 -8293 1530 -8270
rect 1450 -8327 1473 -8293
rect 1507 -8327 1530 -8293
rect 2740 -8027 2763 -7993
rect 2797 -8027 2820 -7993
rect 2740 -8050 2820 -8027
rect 2890 -8270 2920 -7750
rect 3040 -8170 3070 -7750
rect 3190 -8070 3220 -7750
rect 3840 -7780 3870 -7750
rect 4170 -7780 4200 -7750
rect 4320 -7775 4350 -7750
rect 3790 -7803 3870 -7780
rect 3790 -7837 3813 -7803
rect 3847 -7837 3870 -7803
rect 3790 -7860 3870 -7837
rect 4320 -7798 4400 -7775
rect 4320 -7832 4343 -7798
rect 4377 -7832 4400 -7798
rect 4320 -7855 4400 -7832
rect 4170 -8010 4200 -7980
rect 4320 -8010 4350 -7855
rect 4470 -7900 4500 -7750
rect 4620 -7780 4650 -7750
rect 4420 -7923 4500 -7900
rect 4420 -7957 4443 -7923
rect 4477 -7957 4500 -7923
rect 4420 -7980 4500 -7957
rect 4470 -8010 4500 -7980
rect 4620 -8010 4650 -7980
rect 3190 -8093 3270 -8070
rect 3190 -8127 3213 -8093
rect 3247 -8127 3270 -8093
rect 3190 -8150 3270 -8127
rect 3040 -8193 3120 -8170
rect 3040 -8227 3063 -8193
rect 3097 -8227 3120 -8193
rect 3040 -8250 3120 -8227
rect 2840 -8293 2920 -8270
rect 1450 -8350 1530 -8327
rect 1960 -8340 1990 -8310
rect 2110 -8340 2140 -8310
rect 1960 -8370 2140 -8340
rect 2260 -8340 2290 -8310
rect 2410 -8340 2440 -8310
rect 2260 -8370 2440 -8340
rect 2840 -8327 2863 -8293
rect 2897 -8327 2920 -8293
rect 4950 -8020 4980 -7750
rect 5569 -7850 5599 -7750
rect 5519 -7873 5599 -7850
rect 5519 -7907 5542 -7873
rect 5576 -7907 5599 -7873
rect 5519 -7930 5599 -7907
rect 5719 -7950 5749 -7750
rect 6049 -7780 6079 -7750
rect 6199 -7775 6229 -7750
rect 5669 -7973 5749 -7950
rect 5669 -8007 5692 -7973
rect 5726 -8007 5749 -7973
rect 6199 -7798 6279 -7775
rect 6199 -7832 6222 -7798
rect 6256 -7832 6279 -7798
rect 6199 -7855 6279 -7832
rect 4950 -8043 5030 -8020
rect 5669 -8030 5749 -8007
rect 6049 -8010 6079 -7980
rect 6199 -8010 6229 -7855
rect 6349 -7900 6379 -7750
rect 6499 -7780 6529 -7750
rect 6299 -7923 6379 -7900
rect 6299 -7957 6322 -7923
rect 6356 -7957 6379 -7923
rect 6299 -7980 6379 -7957
rect 6349 -8010 6379 -7980
rect 6499 -8010 6529 -7980
rect 4950 -8077 4973 -8043
rect 5007 -8077 5030 -8043
rect 4950 -8100 5030 -8077
rect 6829 -8050 6859 -7750
rect 6779 -8073 6859 -8050
rect 6779 -8107 6802 -8073
rect 6836 -8107 6859 -8073
rect 6779 -8130 6859 -8107
rect 6979 -8170 7009 -7750
rect 6929 -8193 7009 -8170
rect 6929 -8227 6952 -8193
rect 6986 -8227 7009 -8193
rect 6929 -8250 7009 -8227
rect 2840 -8350 2920 -8327
rect 4170 -8340 4200 -8310
rect 4320 -8340 4350 -8310
rect 4170 -8370 4350 -8340
rect 4470 -8340 4500 -8310
rect 4620 -8340 4650 -8310
rect 4470 -8370 4650 -8340
rect 6049 -8340 6079 -8310
rect 6199 -8340 6229 -8310
rect 6049 -8370 6229 -8340
rect 6349 -8340 6379 -8310
rect 6499 -8340 6529 -8310
rect 6349 -8370 6529 -8340
rect 1410 -9013 1490 -8990
rect 1410 -9047 1433 -9013
rect 1467 -9047 1490 -9013
rect 1920 -9000 2100 -8970
rect 1920 -9030 1950 -9000
rect 2070 -9030 2100 -9000
rect 2220 -9000 2400 -8970
rect 2220 -9030 2250 -9000
rect 2370 -9030 2400 -9000
rect 2800 -9013 2880 -8990
rect 1410 -9070 1490 -9047
rect 1290 -9113 1370 -9090
rect 1290 -9147 1313 -9113
rect 1347 -9147 1370 -9113
rect 1290 -9170 1370 -9147
rect 1090 -9313 1170 -9290
rect 1090 -9347 1113 -9313
rect 1147 -9347 1170 -9313
rect 1090 -9370 1170 -9347
rect 1140 -9590 1170 -9370
rect 1290 -9590 1320 -9170
rect 1440 -9590 1470 -9070
rect 1540 -9213 1620 -9190
rect 1540 -9247 1563 -9213
rect 1597 -9247 1620 -9213
rect 1540 -9270 1620 -9247
rect 1590 -9590 1620 -9270
rect 2800 -9047 2823 -9013
rect 2857 -9047 2880 -9013
rect 4110 -9000 4290 -8970
rect 4110 -9030 4140 -9000
rect 4260 -9030 4290 -9000
rect 4410 -9000 4590 -8970
rect 4410 -9030 4440 -9000
rect 4560 -9030 4590 -9000
rect 5990 -9000 6170 -8970
rect 5990 -9030 6020 -9000
rect 6140 -9030 6170 -9000
rect 6290 -9000 6470 -8970
rect 6290 -9030 6320 -9000
rect 6440 -9030 6470 -9000
rect 2800 -9070 2880 -9047
rect 2700 -9313 2780 -9290
rect 1920 -9360 1950 -9330
rect 2070 -9485 2100 -9330
rect 2220 -9360 2250 -9330
rect 2370 -9360 2400 -9330
rect 2700 -9347 2723 -9313
rect 2757 -9347 2780 -9313
rect 2170 -9383 2250 -9360
rect 2170 -9417 2193 -9383
rect 2227 -9417 2250 -9383
rect 2170 -9440 2250 -9417
rect 2070 -9508 2150 -9485
rect 2070 -9542 2093 -9508
rect 2127 -9542 2150 -9508
rect 1920 -9590 1950 -9560
rect 2070 -9565 2150 -9542
rect 2070 -9590 2100 -9565
rect 2220 -9590 2250 -9440
rect 2700 -9370 2780 -9347
rect 2370 -9590 2400 -9560
rect 2700 -9590 2730 -9370
rect 2850 -9590 2880 -9070
rect 3000 -9113 3080 -9090
rect 3000 -9147 3023 -9113
rect 3057 -9147 3080 -9113
rect 3000 -9170 3080 -9147
rect 3000 -9590 3030 -9170
rect 3150 -9213 3230 -9190
rect 3150 -9247 3173 -9213
rect 3207 -9247 3230 -9213
rect 3150 -9270 3230 -9247
rect 3150 -9590 3180 -9270
rect 4890 -9263 4970 -9240
rect 4890 -9297 4913 -9263
rect 4947 -9297 4970 -9263
rect 4890 -9320 4970 -9297
rect 4110 -9360 4140 -9330
rect 3730 -9503 3810 -9480
rect 3730 -9537 3753 -9503
rect 3787 -9537 3810 -9503
rect 3730 -9560 3810 -9537
rect 4260 -9485 4290 -9330
rect 4410 -9360 4440 -9330
rect 4560 -9360 4590 -9330
rect 4360 -9383 4440 -9360
rect 4360 -9417 4383 -9383
rect 4417 -9417 4440 -9383
rect 4360 -9440 4440 -9417
rect 4260 -9508 4340 -9485
rect 4260 -9542 4283 -9508
rect 4317 -9542 4340 -9508
rect 3780 -9590 3810 -9560
rect 4110 -9590 4140 -9560
rect 4260 -9565 4340 -9542
rect 4260 -9590 4290 -9565
rect 4410 -9590 4440 -9440
rect 4560 -9590 4590 -9560
rect 4890 -9590 4920 -9320
rect 5610 -9333 5690 -9310
rect 6870 -9113 6950 -9090
rect 6870 -9147 6893 -9113
rect 6927 -9147 6950 -9113
rect 6870 -9170 6950 -9147
rect 6720 -9233 6800 -9210
rect 6720 -9267 6743 -9233
rect 6777 -9267 6800 -9233
rect 6720 -9290 6800 -9267
rect 5610 -9367 5633 -9333
rect 5667 -9367 5690 -9333
rect 5990 -9360 6020 -9330
rect 5610 -9390 5690 -9367
rect 5460 -9433 5540 -9410
rect 5460 -9467 5483 -9433
rect 5517 -9467 5540 -9433
rect 5460 -9490 5540 -9467
rect 5510 -9590 5540 -9490
rect 5660 -9590 5690 -9390
rect 6140 -9485 6170 -9330
rect 6290 -9360 6320 -9330
rect 6440 -9360 6470 -9330
rect 6240 -9383 6320 -9360
rect 6240 -9417 6263 -9383
rect 6297 -9417 6320 -9383
rect 6240 -9440 6320 -9417
rect 6140 -9508 6220 -9485
rect 6140 -9542 6163 -9508
rect 6197 -9542 6220 -9508
rect 5990 -9590 6020 -9560
rect 6140 -9565 6220 -9542
rect 6140 -9590 6170 -9565
rect 6290 -9590 6320 -9440
rect 6440 -9590 6470 -9560
rect 6770 -9590 6800 -9290
rect 6920 -9590 6950 -9170
rect 1140 -9920 1170 -9890
rect 1290 -9920 1320 -9890
rect 1440 -9920 1470 -9890
rect 1590 -9920 1620 -9890
rect 1920 -9920 1950 -9890
rect 2070 -9920 2100 -9890
rect 2220 -9920 2250 -9890
rect 2370 -9920 2400 -9890
rect 2700 -9920 2730 -9890
rect 1920 -9943 2000 -9920
rect 1920 -9977 1943 -9943
rect 1977 -9977 2000 -9943
rect 1920 -10000 2000 -9977
rect 2320 -9943 2400 -9920
rect 2850 -9930 2880 -9890
rect 3000 -9930 3030 -9890
rect 3150 -9930 3180 -9890
rect 3780 -9920 3810 -9890
rect 4110 -9920 4140 -9890
rect 4260 -9920 4290 -9890
rect 4410 -9920 4440 -9890
rect 4560 -9920 4590 -9890
rect 4890 -9920 4920 -9890
rect 5510 -9920 5540 -9890
rect 5660 -9920 5690 -9890
rect 5990 -9920 6020 -9890
rect 6140 -9920 6170 -9890
rect 6290 -9920 6320 -9890
rect 6440 -9920 6470 -9890
rect 6770 -9920 6800 -9890
rect 6920 -9920 6950 -9890
rect 2320 -9977 2343 -9943
rect 2377 -9977 2400 -9943
rect 2320 -10000 2400 -9977
rect 4110 -9943 4190 -9920
rect 4110 -9977 4133 -9943
rect 4167 -9977 4190 -9943
rect 4110 -10000 4190 -9977
rect 4510 -9943 4590 -9920
rect 4510 -9977 4533 -9943
rect 4567 -9977 4590 -9943
rect 4510 -10000 4590 -9977
rect 5990 -9943 6070 -9920
rect 5990 -9977 6013 -9943
rect 6047 -9977 6070 -9943
rect 5990 -10000 6070 -9977
rect 6390 -9943 6470 -9920
rect 6390 -9977 6413 -9943
rect 6447 -9977 6470 -9943
rect 6390 -10000 6470 -9977
rect 1920 -10183 2000 -10160
rect 1920 -10217 1943 -10183
rect 1977 -10217 2000 -10183
rect 1920 -10240 2000 -10217
rect 2320 -10183 2400 -10160
rect 2320 -10217 2343 -10183
rect 2377 -10217 2400 -10183
rect 2320 -10240 2400 -10217
rect 4110 -10183 4190 -10160
rect 4110 -10217 4133 -10183
rect 4167 -10217 4190 -10183
rect 1140 -10270 1170 -10240
rect 1290 -10270 1320 -10240
rect 1440 -10270 1470 -10240
rect 1590 -10270 1620 -10240
rect 1920 -10270 1950 -10240
rect 2070 -10270 2100 -10240
rect 2220 -10270 2250 -10240
rect 2370 -10270 2400 -10240
rect 2700 -10270 2730 -10240
rect 2850 -10270 2880 -10230
rect 3000 -10270 3030 -10230
rect 3150 -10270 3180 -10230
rect 4110 -10240 4190 -10217
rect 4510 -10183 4590 -10160
rect 4510 -10217 4533 -10183
rect 4567 -10217 4590 -10183
rect 4510 -10240 4590 -10217
rect 5990 -10183 6070 -10160
rect 5990 -10217 6013 -10183
rect 6047 -10217 6070 -10183
rect 5990 -10240 6070 -10217
rect 6390 -10183 6470 -10160
rect 6390 -10217 6413 -10183
rect 6447 -10217 6470 -10183
rect 6390 -10240 6470 -10217
rect 3780 -10270 3810 -10240
rect 4110 -10270 4140 -10240
rect 4260 -10270 4290 -10240
rect 4410 -10270 4440 -10240
rect 4560 -10270 4590 -10240
rect 4890 -10270 4920 -10240
rect 5510 -10270 5540 -10240
rect 5660 -10270 5690 -10240
rect 5990 -10270 6020 -10240
rect 6140 -10270 6170 -10240
rect 6290 -10270 6320 -10240
rect 6440 -10270 6470 -10240
rect 6770 -10270 6800 -10240
rect 6920 -10270 6950 -10240
rect 1140 -10790 1170 -10570
rect 1090 -10813 1170 -10790
rect 1090 -10847 1113 -10813
rect 1147 -10847 1170 -10813
rect 1090 -10870 1170 -10847
rect 1290 -10990 1320 -10570
rect 1290 -11013 1370 -10990
rect 1290 -11047 1313 -11013
rect 1347 -11047 1370 -11013
rect 1290 -11070 1370 -11047
rect 1440 -11090 1470 -10570
rect 1590 -10890 1620 -10570
rect 1920 -10600 1950 -10570
rect 2070 -10595 2100 -10570
rect 2070 -10618 2150 -10595
rect 2070 -10652 2093 -10618
rect 2127 -10652 2150 -10618
rect 2070 -10675 2150 -10652
rect 1920 -10830 1950 -10800
rect 2070 -10830 2100 -10675
rect 2220 -10720 2250 -10570
rect 2370 -10600 2400 -10570
rect 2170 -10743 2250 -10720
rect 2170 -10777 2193 -10743
rect 2227 -10777 2250 -10743
rect 2170 -10800 2250 -10777
rect 2700 -10790 2730 -10570
rect 2220 -10830 2250 -10800
rect 2370 -10830 2400 -10800
rect 2700 -10813 2780 -10790
rect 1540 -10913 1620 -10890
rect 1540 -10947 1563 -10913
rect 1597 -10947 1620 -10913
rect 1540 -10970 1620 -10947
rect 1410 -11113 1490 -11090
rect 1410 -11147 1433 -11113
rect 1467 -11147 1490 -11113
rect 2700 -10847 2723 -10813
rect 2757 -10847 2780 -10813
rect 2700 -10870 2780 -10847
rect 2850 -11090 2880 -10570
rect 3000 -10990 3030 -10570
rect 3150 -10890 3180 -10570
rect 3780 -10600 3810 -10570
rect 4110 -10600 4140 -10570
rect 4260 -10595 4290 -10570
rect 3730 -10623 3810 -10600
rect 3730 -10657 3753 -10623
rect 3787 -10657 3810 -10623
rect 3730 -10680 3810 -10657
rect 4260 -10618 4340 -10595
rect 4260 -10652 4283 -10618
rect 4317 -10652 4340 -10618
rect 4260 -10675 4340 -10652
rect 4110 -10830 4140 -10800
rect 4260 -10830 4290 -10675
rect 4410 -10720 4440 -10570
rect 4560 -10600 4590 -10570
rect 4360 -10743 4440 -10720
rect 4360 -10777 4383 -10743
rect 4417 -10777 4440 -10743
rect 4360 -10800 4440 -10777
rect 4410 -10830 4440 -10800
rect 4560 -10830 4590 -10800
rect 3150 -10913 3230 -10890
rect 3150 -10947 3173 -10913
rect 3207 -10947 3230 -10913
rect 3150 -10970 3230 -10947
rect 3000 -11013 3080 -10990
rect 3000 -11047 3023 -11013
rect 3057 -11047 3080 -11013
rect 3000 -11070 3080 -11047
rect 2800 -11113 2880 -11090
rect 1410 -11170 1490 -11147
rect 1920 -11160 1950 -11130
rect 2070 -11160 2100 -11130
rect 1920 -11190 2100 -11160
rect 2220 -11160 2250 -11130
rect 2370 -11160 2400 -11130
rect 2220 -11190 2400 -11160
rect 2800 -11147 2823 -11113
rect 2857 -11147 2880 -11113
rect 4890 -10840 4920 -10570
rect 5510 -10670 5540 -10570
rect 5460 -10693 5540 -10670
rect 5460 -10727 5483 -10693
rect 5517 -10727 5540 -10693
rect 5460 -10750 5540 -10727
rect 5660 -10770 5690 -10570
rect 5990 -10600 6020 -10570
rect 6140 -10595 6170 -10570
rect 5610 -10793 5690 -10770
rect 5610 -10827 5633 -10793
rect 5667 -10827 5690 -10793
rect 6140 -10618 6220 -10595
rect 6140 -10652 6163 -10618
rect 6197 -10652 6220 -10618
rect 6140 -10675 6220 -10652
rect 4890 -10863 4970 -10840
rect 5610 -10850 5690 -10827
rect 5990 -10830 6020 -10800
rect 6140 -10830 6170 -10675
rect 6290 -10720 6320 -10570
rect 6440 -10600 6470 -10570
rect 6240 -10743 6320 -10720
rect 6240 -10777 6263 -10743
rect 6297 -10777 6320 -10743
rect 6240 -10800 6320 -10777
rect 6290 -10830 6320 -10800
rect 6440 -10830 6470 -10800
rect 4890 -10897 4913 -10863
rect 4947 -10897 4970 -10863
rect 4890 -10920 4970 -10897
rect 6770 -10870 6800 -10570
rect 6720 -10893 6800 -10870
rect 6720 -10927 6743 -10893
rect 6777 -10927 6800 -10893
rect 6720 -10950 6800 -10927
rect 6920 -10990 6950 -10570
rect 6870 -11013 6950 -10990
rect 6870 -11047 6893 -11013
rect 6927 -11047 6950 -11013
rect 6870 -11070 6950 -11047
rect 2800 -11170 2880 -11147
rect 4110 -11160 4140 -11130
rect 4260 -11160 4290 -11130
rect 4110 -11190 4290 -11160
rect 4410 -11160 4440 -11130
rect 4560 -11160 4590 -11130
rect 4410 -11190 4590 -11160
rect 5990 -11160 6020 -11130
rect 6140 -11160 6170 -11130
rect 5990 -11190 6170 -11160
rect 6290 -11160 6320 -11130
rect 6440 -11160 6470 -11130
rect 6290 -11190 6470 -11160
rect 1921 -11820 2101 -11790
rect 1921 -11850 1951 -11820
rect 2071 -11850 2101 -11820
rect 2221 -11820 2401 -11790
rect 2221 -11850 2251 -11820
rect 2371 -11850 2401 -11820
rect 2951 -11823 3031 -11800
rect 2951 -11857 2974 -11823
rect 3008 -11857 3031 -11823
rect 3971 -11820 4151 -11790
rect 3971 -11850 4001 -11820
rect 4121 -11850 4151 -11820
rect 4271 -11820 4451 -11790
rect 4271 -11850 4301 -11820
rect 4421 -11850 4451 -11820
rect 5381 -11829 5461 -11806
rect 2951 -11880 3031 -11857
rect 2801 -11943 2881 -11920
rect 2801 -11977 2824 -11943
rect 2858 -11977 2881 -11943
rect 2801 -12000 2881 -11977
rect 2671 -12063 2751 -12040
rect 2671 -12097 2694 -12063
rect 2728 -12097 2751 -12063
rect 2671 -12120 2751 -12097
rect 1921 -12180 1951 -12150
rect 1371 -12233 1471 -12210
rect 1371 -12267 1394 -12233
rect 1428 -12267 1471 -12233
rect 1371 -12290 1471 -12267
rect 1541 -12213 1621 -12190
rect 1541 -12247 1564 -12213
rect 1598 -12247 1621 -12213
rect 1541 -12270 1621 -12247
rect 1241 -12313 1321 -12290
rect 1241 -12347 1264 -12313
rect 1298 -12347 1321 -12313
rect 1241 -12370 1321 -12347
rect 1291 -12410 1321 -12370
rect 1441 -12410 1471 -12290
rect 1591 -12410 1621 -12270
rect 2071 -12305 2101 -12150
rect 2221 -12180 2251 -12150
rect 2371 -12180 2401 -12150
rect 2171 -12203 2251 -12180
rect 2171 -12237 2194 -12203
rect 2228 -12237 2251 -12203
rect 2171 -12260 2251 -12237
rect 2071 -12328 2151 -12305
rect 2071 -12362 2094 -12328
rect 2128 -12362 2151 -12328
rect 1921 -12410 1951 -12380
rect 2071 -12385 2151 -12362
rect 2071 -12410 2101 -12385
rect 2221 -12410 2251 -12260
rect 2371 -12410 2401 -12380
rect 2701 -12410 2731 -12120
rect 2851 -12410 2881 -12000
rect 3001 -12410 3031 -11880
rect 5381 -11863 5404 -11829
rect 5438 -11863 5461 -11829
rect 6011 -11821 6191 -11791
rect 6011 -11851 6041 -11821
rect 6161 -11851 6191 -11821
rect 6311 -11821 6491 -11791
rect 6311 -11851 6341 -11821
rect 6461 -11851 6491 -11821
rect 5381 -11886 5461 -11863
rect 4751 -12083 4831 -12060
rect 4751 -12117 4774 -12083
rect 4808 -12117 4831 -12083
rect 4751 -12140 4831 -12117
rect 3971 -12180 4001 -12150
rect 3591 -12323 3671 -12300
rect 3591 -12357 3614 -12323
rect 3648 -12357 3671 -12323
rect 3591 -12380 3671 -12357
rect 4121 -12305 4151 -12150
rect 4271 -12180 4301 -12150
rect 4421 -12180 4451 -12150
rect 4221 -12203 4301 -12180
rect 4221 -12237 4244 -12203
rect 4278 -12237 4301 -12203
rect 4221 -12260 4301 -12237
rect 4121 -12328 4201 -12305
rect 4121 -12362 4144 -12328
rect 4178 -12362 4201 -12328
rect 3641 -12410 3671 -12380
rect 3971 -12410 4001 -12380
rect 4121 -12385 4201 -12362
rect 4121 -12410 4151 -12385
rect 4271 -12410 4301 -12260
rect 4421 -12410 4451 -12380
rect 4751 -12410 4781 -12140
rect 5381 -12411 5411 -11886
rect 5481 -11954 5561 -11931
rect 5481 -11988 5504 -11954
rect 5538 -11988 5561 -11954
rect 5481 -12011 5561 -11988
rect 5531 -12411 5561 -12011
rect 5681 -12044 5761 -12021
rect 5681 -12078 5704 -12044
rect 5738 -12078 5761 -12044
rect 5681 -12101 5761 -12078
rect 5681 -12411 5711 -12101
rect 6011 -12181 6041 -12151
rect 6161 -12181 6191 -12151
rect 6161 -12204 6241 -12181
rect 6161 -12238 6184 -12204
rect 6218 -12238 6241 -12204
rect 6161 -12261 6241 -12238
rect 6011 -12411 6041 -12381
rect 6161 -12411 6191 -12261
rect 6311 -12306 6341 -12151
rect 6461 -12181 6491 -12151
rect 7081 -12154 7161 -12131
rect 7081 -12188 7104 -12154
rect 7138 -12188 7161 -12154
rect 7081 -12211 7161 -12188
rect 6261 -12329 6341 -12306
rect 6941 -12254 7021 -12231
rect 6941 -12288 6964 -12254
rect 6998 -12288 7021 -12254
rect 6941 -12311 7021 -12288
rect 6261 -12363 6284 -12329
rect 6318 -12363 6341 -12329
rect 6261 -12386 6341 -12363
rect 6791 -12334 6871 -12311
rect 6791 -12368 6814 -12334
rect 6848 -12368 6871 -12334
rect 6311 -12411 6341 -12386
rect 6461 -12411 6491 -12381
rect 6791 -12391 6871 -12368
rect 6791 -12411 6821 -12391
rect 6941 -12411 6971 -12311
rect 7091 -12411 7121 -12211
rect 1291 -12740 1321 -12710
rect 1441 -12740 1471 -12710
rect 1591 -12740 1621 -12710
rect 1921 -12740 1951 -12710
rect 2071 -12740 2101 -12710
rect 2221 -12740 2251 -12710
rect 2371 -12740 2401 -12710
rect 2701 -12740 2731 -12710
rect 2851 -12740 2881 -12710
rect 3001 -12740 3031 -12710
rect 3641 -12740 3671 -12710
rect 3971 -12740 4001 -12710
rect 4121 -12740 4151 -12710
rect 4271 -12740 4301 -12710
rect 4421 -12740 4451 -12710
rect 4751 -12740 4781 -12710
rect 1921 -12763 2001 -12740
rect 1921 -12797 1944 -12763
rect 1978 -12797 2001 -12763
rect 1921 -12820 2001 -12797
rect 2321 -12763 2401 -12740
rect 2321 -12797 2344 -12763
rect 2378 -12797 2401 -12763
rect 2321 -12820 2401 -12797
rect 3971 -12763 4051 -12740
rect 3971 -12797 3994 -12763
rect 4028 -12797 4051 -12763
rect 3971 -12820 4051 -12797
rect 4371 -12763 4451 -12740
rect 5381 -12741 5411 -12711
rect 5531 -12741 5561 -12711
rect 5681 -12741 5711 -12711
rect 6011 -12741 6041 -12711
rect 6161 -12741 6191 -12711
rect 6311 -12741 6341 -12711
rect 6461 -12741 6491 -12711
rect 6791 -12741 6821 -12711
rect 6941 -12741 6971 -12711
rect 7091 -12741 7121 -12711
rect 4371 -12797 4394 -12763
rect 4428 -12797 4451 -12763
rect 4371 -12820 4451 -12797
rect 6011 -12764 6091 -12741
rect 6011 -12798 6034 -12764
rect 6068 -12798 6091 -12764
rect 6011 -12821 6091 -12798
rect 6411 -12764 6491 -12741
rect 6411 -12798 6434 -12764
rect 6468 -12798 6491 -12764
rect 6411 -12821 6491 -12798
<< polycont >>
rect 1433 2314 1467 2348
rect 1313 2214 1347 2248
rect 1113 2014 1147 2048
rect 1563 2114 1597 2148
rect 2823 2314 2857 2348
rect 2723 2014 2757 2048
rect 2193 1944 2227 1978
rect 2093 1819 2127 1853
rect 3023 2214 3057 2248
rect 3173 2114 3207 2148
rect 5193 2184 5227 2218
rect 4993 2064 5027 2098
rect 3883 1964 3917 1998
rect 3733 1864 3767 1898
rect 4513 1944 4547 1978
rect 4413 1819 4447 1853
rect 7163 2214 7197 2248
rect 7013 2094 7047 2128
rect 5903 1994 5937 2028
rect 5753 1894 5787 1928
rect 6533 1944 6567 1978
rect 6433 1819 6467 1853
rect 1943 1384 1977 1418
rect 2343 1384 2377 1418
rect 4263 1384 4297 1418
rect 4663 1384 4697 1418
rect 6283 1384 6317 1418
rect 6683 1384 6717 1418
rect 1943 1144 1977 1178
rect 2343 1144 2377 1178
rect 4263 1144 4297 1178
rect 4663 1144 4697 1178
rect 6283 1144 6317 1178
rect 6683 1144 6717 1178
rect 1413 634 1447 668
rect 1563 534 1597 568
rect 2093 709 2127 743
rect 2193 584 2227 618
rect 2673 434 2707 468
rect 3733 634 3767 668
rect 3883 534 3917 568
rect 4413 709 4447 743
rect 4513 584 4547 618
rect 2823 314 2857 348
rect 4993 434 5027 468
rect 6533 709 6567 743
rect 6433 584 6467 618
rect 7213 664 7247 698
rect 7063 564 7097 598
rect 5953 464 5987 498
rect 5143 314 5177 348
rect 5753 344 5787 378
rect 1433 -506 1467 -472
rect 1313 -606 1347 -572
rect 1113 -806 1147 -772
rect 1563 -706 1597 -672
rect 2823 -506 2857 -472
rect 2723 -806 2757 -772
rect 2193 -876 2227 -842
rect 2093 -1001 2127 -967
rect 3023 -606 3057 -572
rect 3173 -706 3207 -672
rect 4913 -756 4947 -722
rect 3753 -996 3787 -962
rect 4383 -876 4417 -842
rect 4283 -1001 4317 -967
rect 6893 -606 6927 -572
rect 6743 -726 6777 -692
rect 5633 -826 5667 -792
rect 5483 -926 5517 -892
rect 6263 -876 6297 -842
rect 6163 -1001 6197 -967
rect 1943 -1436 1977 -1402
rect 2343 -1436 2377 -1402
rect 4133 -1436 4167 -1402
rect 4533 -1436 4567 -1402
rect 6013 -1436 6047 -1402
rect 6413 -1436 6447 -1402
rect 1943 -1676 1977 -1642
rect 2343 -1676 2377 -1642
rect 4133 -1676 4167 -1642
rect 4533 -1676 4567 -1642
rect 6013 -1676 6047 -1642
rect 6413 -1676 6447 -1642
rect 1113 -2306 1147 -2272
rect 1313 -2506 1347 -2472
rect 2093 -2111 2127 -2077
rect 2193 -2236 2227 -2202
rect 1563 -2406 1597 -2372
rect 1433 -2606 1467 -2572
rect 2723 -2306 2757 -2272
rect 3753 -2116 3787 -2082
rect 4283 -2111 4317 -2077
rect 4383 -2236 4417 -2202
rect 3173 -2406 3207 -2372
rect 3023 -2506 3057 -2472
rect 2823 -2606 2857 -2572
rect 5483 -2186 5517 -2152
rect 5633 -2286 5667 -2252
rect 6163 -2111 6197 -2077
rect 6263 -2236 6297 -2202
rect 4913 -2356 4947 -2322
rect 6743 -2386 6777 -2352
rect 6893 -2506 6927 -2472
rect 2974 -3316 3008 -3282
rect 2824 -3436 2858 -3402
rect 2694 -3556 2728 -3522
rect 1394 -3726 1428 -3692
rect 1564 -3706 1598 -3672
rect 1264 -3806 1298 -3772
rect 2194 -3696 2228 -3662
rect 2094 -3821 2128 -3787
rect 5404 -3322 5438 -3288
rect 4774 -3576 4808 -3542
rect 3614 -3816 3648 -3782
rect 4244 -3696 4278 -3662
rect 4144 -3821 4178 -3787
rect 5504 -3447 5538 -3413
rect 5704 -3537 5738 -3503
rect 6184 -3697 6218 -3663
rect 7104 -3647 7138 -3613
rect 6964 -3747 6998 -3713
rect 6284 -3822 6318 -3788
rect 6814 -3827 6848 -3793
rect 1944 -4256 1978 -4222
rect 2344 -4256 2378 -4222
rect 3994 -4256 4028 -4222
rect 4394 -4256 4428 -4222
rect 6034 -4257 6068 -4223
rect 6434 -4257 6468 -4223
rect 1983 -4576 2017 -4542
rect 2383 -4576 2417 -4542
rect 4194 -4577 4228 -4543
rect 4594 -4577 4628 -4543
rect 6253 -4577 6287 -4543
rect 6653 -4577 6687 -4543
rect 1153 -5066 1187 -5032
rect 1303 -5166 1337 -5132
rect 1453 -5266 1487 -5232
rect 1603 -5366 1637 -5332
rect 2133 -5226 2167 -5192
rect 2713 -5066 2747 -5032
rect 2863 -5066 2897 -5032
rect 3013 -5066 3047 -5032
rect 3163 -5066 3197 -5032
rect 3814 -5017 3848 -4983
rect 4344 -5012 4378 -4978
rect 4444 -5137 4478 -5103
rect 2233 -5366 2267 -5332
rect 4974 -5257 5008 -5223
rect 6503 -5012 6537 -4978
rect 7033 -5007 7067 -4973
rect 6403 -5137 6437 -5103
rect 7183 -5087 7217 -5053
rect 7323 -5187 7357 -5153
rect 5923 -5297 5957 -5263
rect 5723 -5387 5757 -5353
rect 5623 -5512 5657 -5478
rect 1473 -6227 1507 -6193
rect 1353 -6327 1387 -6293
rect 1153 -6527 1187 -6493
rect 1603 -6427 1637 -6393
rect 2863 -6227 2897 -6193
rect 2763 -6527 2797 -6493
rect 2233 -6597 2267 -6563
rect 2133 -6722 2167 -6688
rect 3063 -6327 3097 -6293
rect 3213 -6427 3247 -6393
rect 4973 -6477 5007 -6443
rect 3813 -6717 3847 -6683
rect 4443 -6597 4477 -6563
rect 4343 -6722 4377 -6688
rect 6952 -6327 6986 -6293
rect 6802 -6447 6836 -6413
rect 5692 -6547 5726 -6513
rect 5542 -6647 5576 -6613
rect 6322 -6597 6356 -6563
rect 6222 -6722 6256 -6688
rect 1983 -7157 2017 -7123
rect 2383 -7157 2417 -7123
rect 4193 -7157 4227 -7123
rect 4593 -7157 4627 -7123
rect 6072 -7157 6106 -7123
rect 6472 -7157 6506 -7123
rect 1983 -7397 2017 -7363
rect 2383 -7397 2417 -7363
rect 4193 -7397 4227 -7363
rect 4593 -7397 4627 -7363
rect 6072 -7397 6106 -7363
rect 6472 -7397 6506 -7363
rect 1153 -8027 1187 -7993
rect 1353 -8227 1387 -8193
rect 2133 -7832 2167 -7798
rect 2233 -7957 2267 -7923
rect 1603 -8127 1637 -8093
rect 1473 -8327 1507 -8293
rect 2763 -8027 2797 -7993
rect 3813 -7837 3847 -7803
rect 4343 -7832 4377 -7798
rect 4443 -7957 4477 -7923
rect 3213 -8127 3247 -8093
rect 3063 -8227 3097 -8193
rect 2863 -8327 2897 -8293
rect 5542 -7907 5576 -7873
rect 5692 -8007 5726 -7973
rect 6222 -7832 6256 -7798
rect 6322 -7957 6356 -7923
rect 4973 -8077 5007 -8043
rect 6802 -8107 6836 -8073
rect 6952 -8227 6986 -8193
rect 1433 -9047 1467 -9013
rect 1313 -9147 1347 -9113
rect 1113 -9347 1147 -9313
rect 1563 -9247 1597 -9213
rect 2823 -9047 2857 -9013
rect 2723 -9347 2757 -9313
rect 2193 -9417 2227 -9383
rect 2093 -9542 2127 -9508
rect 3023 -9147 3057 -9113
rect 3173 -9247 3207 -9213
rect 4913 -9297 4947 -9263
rect 3753 -9537 3787 -9503
rect 4383 -9417 4417 -9383
rect 4283 -9542 4317 -9508
rect 6893 -9147 6927 -9113
rect 6743 -9267 6777 -9233
rect 5633 -9367 5667 -9333
rect 5483 -9467 5517 -9433
rect 6263 -9417 6297 -9383
rect 6163 -9542 6197 -9508
rect 1943 -9977 1977 -9943
rect 2343 -9977 2377 -9943
rect 4133 -9977 4167 -9943
rect 4533 -9977 4567 -9943
rect 6013 -9977 6047 -9943
rect 6413 -9977 6447 -9943
rect 1943 -10217 1977 -10183
rect 2343 -10217 2377 -10183
rect 4133 -10217 4167 -10183
rect 4533 -10217 4567 -10183
rect 6013 -10217 6047 -10183
rect 6413 -10217 6447 -10183
rect 1113 -10847 1147 -10813
rect 1313 -11047 1347 -11013
rect 2093 -10652 2127 -10618
rect 2193 -10777 2227 -10743
rect 1563 -10947 1597 -10913
rect 1433 -11147 1467 -11113
rect 2723 -10847 2757 -10813
rect 3753 -10657 3787 -10623
rect 4283 -10652 4317 -10618
rect 4383 -10777 4417 -10743
rect 3173 -10947 3207 -10913
rect 3023 -11047 3057 -11013
rect 2823 -11147 2857 -11113
rect 5483 -10727 5517 -10693
rect 5633 -10827 5667 -10793
rect 6163 -10652 6197 -10618
rect 6263 -10777 6297 -10743
rect 4913 -10897 4947 -10863
rect 6743 -10927 6777 -10893
rect 6893 -11047 6927 -11013
rect 2974 -11857 3008 -11823
rect 2824 -11977 2858 -11943
rect 2694 -12097 2728 -12063
rect 1394 -12267 1428 -12233
rect 1564 -12247 1598 -12213
rect 1264 -12347 1298 -12313
rect 2194 -12237 2228 -12203
rect 2094 -12362 2128 -12328
rect 5404 -11863 5438 -11829
rect 4774 -12117 4808 -12083
rect 3614 -12357 3648 -12323
rect 4244 -12237 4278 -12203
rect 4144 -12362 4178 -12328
rect 5504 -11988 5538 -11954
rect 5704 -12078 5738 -12044
rect 6184 -12238 6218 -12204
rect 7104 -12188 7138 -12154
rect 6964 -12288 6998 -12254
rect 6284 -12363 6318 -12329
rect 6814 -12368 6848 -12334
rect 1944 -12797 1978 -12763
rect 2344 -12797 2378 -12763
rect 3994 -12797 4028 -12763
rect 4394 -12797 4428 -12763
rect 6034 -12798 6068 -12764
rect 6434 -12798 6468 -12764
<< locali >>
rect 1020 2478 3300 2501
rect 1020 2444 1103 2478
rect 1137 2444 1183 2478
rect 1217 2444 1263 2478
rect 1297 2444 1343 2478
rect 1377 2444 1423 2478
rect 1457 2444 1503 2478
rect 1537 2444 1583 2478
rect 1617 2444 1663 2478
rect 1697 2444 1743 2478
rect 1777 2444 1823 2478
rect 1857 2444 1903 2478
rect 1937 2444 1983 2478
rect 2017 2444 2063 2478
rect 2097 2444 2143 2478
rect 2177 2444 2223 2478
rect 2257 2444 2303 2478
rect 2337 2444 2383 2478
rect 2417 2444 2463 2478
rect 2497 2444 2543 2478
rect 2577 2444 2623 2478
rect 2657 2444 2703 2478
rect 2737 2444 2783 2478
rect 2817 2444 2863 2478
rect 2897 2444 2943 2478
rect 2977 2444 3023 2478
rect 3057 2444 3103 2478
rect 3137 2444 3183 2478
rect 3217 2444 3300 2478
rect 1020 2421 3300 2444
rect 3640 2478 5320 2501
rect 3640 2444 3663 2478
rect 3697 2444 3743 2478
rect 3777 2444 3823 2478
rect 3857 2444 3903 2478
rect 3937 2444 3983 2478
rect 4017 2444 4063 2478
rect 4097 2444 4143 2478
rect 4177 2444 4223 2478
rect 4257 2444 4303 2478
rect 4337 2444 4383 2478
rect 4417 2444 4463 2478
rect 4497 2444 4543 2478
rect 4577 2444 4623 2478
rect 4657 2444 4703 2478
rect 4737 2444 4783 2478
rect 4817 2444 4863 2478
rect 4897 2444 4943 2478
rect 4977 2444 5023 2478
rect 5057 2444 5103 2478
rect 5137 2444 5183 2478
rect 5217 2444 5263 2478
rect 5297 2444 5320 2478
rect 3640 2421 5320 2444
rect 5660 2478 7340 2501
rect 5660 2444 5683 2478
rect 5717 2444 5763 2478
rect 5797 2444 5843 2478
rect 5877 2444 5923 2478
rect 5957 2444 6003 2478
rect 6037 2444 6083 2478
rect 6117 2444 6163 2478
rect 6197 2444 6243 2478
rect 6277 2444 6323 2478
rect 6357 2444 6403 2478
rect 6437 2444 6483 2478
rect 6517 2444 6563 2478
rect 6597 2444 6643 2478
rect 6677 2444 6723 2478
rect 6757 2444 6803 2478
rect 6837 2444 6883 2478
rect 6917 2444 6963 2478
rect 6997 2444 7043 2478
rect 7077 2444 7123 2478
rect 7157 2444 7203 2478
rect 7237 2444 7283 2478
rect 7317 2444 7340 2478
rect 5660 2421 7340 2444
rect 1410 2351 1490 2371
rect 1540 2351 1620 2371
rect 0 2348 1620 2351
rect 0 2328 1433 2348
rect 0 2294 23 2328
rect 57 2314 1433 2328
rect 1467 2314 1563 2348
rect 1597 2314 1620 2348
rect 57 2311 1620 2314
rect 57 2294 80 2311
rect 0 2271 80 2294
rect 1410 2291 1490 2311
rect 1540 2291 1620 2311
rect 2800 2348 2880 2371
rect 2800 2314 2823 2348
rect 2857 2314 2880 2348
rect 2800 2291 2880 2314
rect 1290 2251 1370 2271
rect 1670 2251 1750 2271
rect 114 2248 1750 2251
rect 114 2228 1313 2248
rect 114 2194 137 2228
rect 171 2214 1313 2228
rect 1347 2214 1693 2248
rect 1727 2214 1750 2248
rect 171 2211 1750 2214
rect 171 2194 194 2211
rect 114 2171 194 2194
rect 1290 2191 1370 2211
rect 1670 2191 1750 2211
rect 1820 2258 1900 2291
rect 1820 2224 1843 2258
rect 1877 2224 1900 2258
rect 1820 2178 1900 2224
rect 1540 2151 1620 2171
rect 684 2148 1620 2151
rect 684 2128 1563 2148
rect 684 2094 707 2128
rect 741 2114 1563 2128
rect 1597 2114 1620 2148
rect 741 2111 1620 2114
rect 741 2094 764 2111
rect 684 2071 764 2094
rect 1540 2091 1620 2111
rect 1820 2144 1843 2178
rect 1877 2144 1900 2178
rect 1820 2098 1900 2144
rect 1090 2051 1170 2071
rect 1670 2051 1750 2071
rect 798 2048 1750 2051
rect 798 2028 1113 2048
rect 798 1994 821 2028
rect 855 2014 1113 2028
rect 1147 2014 1693 2048
rect 1727 2014 1750 2048
rect 1820 2064 1843 2098
rect 1877 2064 1900 2098
rect 1820 2041 1900 2064
rect 1970 2258 2050 2291
rect 1970 2224 1993 2258
rect 2027 2224 2050 2258
rect 1970 2178 2050 2224
rect 1970 2144 1993 2178
rect 2027 2144 2050 2178
rect 1970 2098 2050 2144
rect 1970 2064 1993 2098
rect 2027 2064 2050 2098
rect 1970 2031 2050 2064
rect 2120 2258 2200 2291
rect 2120 2224 2143 2258
rect 2177 2224 2200 2258
rect 2120 2178 2200 2224
rect 2120 2144 2143 2178
rect 2177 2144 2200 2178
rect 2120 2098 2200 2144
rect 2120 2064 2143 2098
rect 2177 2064 2200 2098
rect 2120 2041 2200 2064
rect 2270 2258 2350 2291
rect 2270 2224 2293 2258
rect 2327 2224 2350 2258
rect 2270 2178 2350 2224
rect 2270 2144 2293 2178
rect 2327 2144 2350 2178
rect 2270 2098 2350 2144
rect 2270 2064 2293 2098
rect 2327 2064 2350 2098
rect 2270 2031 2350 2064
rect 2420 2258 2500 2291
rect 2420 2224 2443 2258
rect 2477 2224 2500 2258
rect 2420 2178 2500 2224
rect 3000 2248 3080 2271
rect 3000 2214 3023 2248
rect 3057 2214 3080 2248
rect 3000 2191 3080 2214
rect 3560 2238 3640 2261
rect 4140 2258 4220 2291
rect 3560 2204 3583 2238
rect 3617 2221 3640 2238
rect 3990 2221 4070 2241
rect 3617 2218 4070 2221
rect 3617 2204 4013 2218
rect 3560 2184 4013 2204
rect 4047 2184 4070 2218
rect 3560 2181 4070 2184
rect 2420 2144 2443 2178
rect 2477 2144 2500 2178
rect 2420 2098 2500 2144
rect 2420 2064 2443 2098
rect 2477 2064 2500 2098
rect 3150 2148 3230 2171
rect 3990 2161 4070 2181
rect 4140 2224 4163 2258
rect 4197 2224 4220 2258
rect 4140 2178 4220 2224
rect 3150 2114 3173 2148
rect 3207 2114 3230 2148
rect 4140 2144 4163 2178
rect 4197 2144 4220 2178
rect 3150 2091 3230 2114
rect 3560 2118 3640 2141
rect 3560 2084 3583 2118
rect 3617 2101 3640 2118
rect 3990 2101 4070 2121
rect 3617 2098 4070 2101
rect 3617 2084 4013 2098
rect 2420 2041 2500 2064
rect 2700 2048 2780 2071
rect 855 2011 1750 2014
rect 855 1994 878 2011
rect 798 1971 878 1994
rect 1090 1991 1170 2011
rect 1670 1991 1750 2011
rect 1990 1981 2030 2031
rect 2170 1981 2250 2001
rect 1990 1978 2250 1981
rect 1990 1944 2193 1978
rect 2227 1944 2250 1978
rect 1990 1941 2250 1944
rect 1990 1811 2030 1941
rect 2170 1921 2250 1941
rect 1060 1771 2030 1811
rect 2070 1861 2150 1876
rect 2290 1861 2330 2031
rect 2700 2014 2723 2048
rect 2757 2014 2780 2048
rect 2700 1991 2780 2014
rect 3300 2056 3380 2079
rect 3560 2064 4013 2084
rect 4047 2064 4070 2098
rect 3560 2061 4070 2064
rect 3300 2022 3323 2056
rect 3357 2022 3380 2056
rect 3990 2041 4070 2061
rect 4140 2098 4220 2144
rect 4140 2064 4163 2098
rect 4197 2064 4220 2098
rect 4140 2041 4220 2064
rect 4290 2258 4370 2291
rect 4290 2224 4313 2258
rect 4347 2224 4370 2258
rect 4290 2178 4370 2224
rect 4290 2144 4313 2178
rect 4347 2144 4370 2178
rect 4290 2098 4370 2144
rect 4290 2064 4313 2098
rect 4347 2064 4370 2098
rect 4290 2031 4370 2064
rect 4440 2258 4520 2291
rect 4440 2224 4463 2258
rect 4497 2224 4520 2258
rect 4440 2178 4520 2224
rect 4440 2144 4463 2178
rect 4497 2144 4520 2178
rect 4440 2098 4520 2144
rect 4440 2064 4463 2098
rect 4497 2064 4520 2098
rect 4440 2041 4520 2064
rect 4590 2258 4670 2291
rect 4590 2224 4613 2258
rect 4647 2224 4670 2258
rect 4590 2178 4670 2224
rect 4590 2144 4613 2178
rect 4647 2144 4670 2178
rect 4590 2098 4670 2144
rect 4590 2064 4613 2098
rect 4647 2064 4670 2098
rect 4590 2031 4670 2064
rect 4740 2258 4820 2291
rect 4740 2224 4763 2258
rect 4797 2224 4820 2258
rect 5580 2251 5660 2271
rect 6010 2251 6090 2271
rect 5580 2248 6090 2251
rect 4740 2178 4820 2224
rect 4740 2144 4763 2178
rect 4797 2144 4820 2178
rect 5170 2218 5250 2241
rect 5170 2184 5193 2218
rect 5227 2184 5250 2218
rect 5580 2214 5603 2248
rect 5637 2214 6033 2248
rect 6067 2214 6090 2248
rect 5580 2211 6090 2214
rect 5580 2191 5660 2211
rect 6010 2191 6090 2211
rect 6160 2258 6240 2291
rect 6160 2224 6183 2258
rect 6217 2224 6240 2258
rect 5170 2161 5250 2184
rect 6160 2178 6240 2224
rect 4740 2098 4820 2144
rect 6010 2131 6090 2151
rect 5472 2128 6090 2131
rect 5472 2127 6033 2128
rect 4740 2064 4763 2098
rect 4797 2064 4820 2098
rect 4740 2041 4820 2064
rect 4970 2098 5050 2121
rect 4970 2064 4993 2098
rect 5027 2064 5050 2098
rect 4970 2041 5050 2064
rect 5250 2104 6033 2127
rect 5250 2070 5273 2104
rect 5307 2094 6033 2104
rect 6067 2094 6090 2128
rect 5307 2091 6090 2094
rect 5307 2087 5472 2091
rect 5307 2070 5330 2087
rect 6010 2071 6090 2091
rect 6160 2144 6183 2178
rect 6217 2144 6240 2178
rect 6160 2098 6240 2144
rect 5250 2047 5330 2070
rect 6160 2064 6183 2098
rect 6217 2064 6240 2098
rect 5580 2031 5660 2050
rect 5880 2031 5960 2051
rect 6160 2041 6240 2064
rect 6310 2258 6390 2291
rect 6310 2224 6333 2258
rect 6367 2224 6390 2258
rect 6310 2178 6390 2224
rect 6310 2144 6333 2178
rect 6367 2144 6390 2178
rect 6310 2098 6390 2144
rect 6310 2064 6333 2098
rect 6367 2064 6390 2098
rect 6310 2031 6390 2064
rect 6460 2258 6540 2291
rect 6460 2224 6483 2258
rect 6517 2224 6540 2258
rect 6460 2178 6540 2224
rect 6460 2144 6483 2178
rect 6517 2144 6540 2178
rect 6460 2098 6540 2144
rect 6460 2064 6483 2098
rect 6517 2064 6540 2098
rect 6460 2041 6540 2064
rect 6610 2258 6690 2291
rect 6610 2224 6633 2258
rect 6667 2224 6690 2258
rect 6610 2178 6690 2224
rect 6610 2144 6633 2178
rect 6667 2144 6690 2178
rect 6610 2098 6690 2144
rect 6610 2064 6633 2098
rect 6667 2064 6690 2098
rect 6610 2031 6690 2064
rect 6760 2258 6840 2291
rect 6760 2224 6783 2258
rect 6817 2224 6840 2258
rect 6760 2178 6840 2224
rect 7140 2248 7220 2271
rect 7140 2214 7163 2248
rect 7197 2214 7220 2248
rect 7140 2191 7220 2214
rect 6760 2144 6783 2178
rect 6817 2144 6840 2178
rect 6760 2098 6840 2144
rect 6760 2064 6783 2098
rect 6817 2064 6840 2098
rect 6990 2128 7070 2151
rect 6990 2094 7013 2128
rect 7047 2094 7070 2128
rect 6990 2071 7070 2094
rect 6760 2041 6840 2064
rect 3300 1999 3380 2022
rect 2540 1968 2620 1991
rect 2540 1934 2563 1968
rect 2597 1951 2620 1968
rect 3054 1968 3134 1991
rect 3054 1951 3077 1968
rect 2597 1934 3077 1951
rect 3111 1951 3134 1968
rect 3111 1934 3300 1951
rect 2540 1911 3300 1934
rect 3340 1877 3380 1999
rect 3560 2001 3640 2021
rect 3860 2001 3940 2021
rect 3560 1998 3940 2001
rect 3560 1964 3583 1998
rect 3617 1964 3883 1998
rect 3917 1964 3940 1998
rect 3560 1961 3940 1964
rect 3560 1941 3640 1961
rect 3860 1941 3940 1961
rect 4310 1981 4350 2031
rect 4490 1981 4570 2001
rect 4310 1978 4570 1981
rect 4310 1944 4513 1978
rect 4547 1944 4570 1978
rect 4310 1941 4570 1944
rect 3710 1901 3790 1921
rect 3300 1861 3380 1877
rect 2070 1854 3380 1861
rect 2070 1853 3323 1854
rect 2070 1819 2093 1853
rect 2127 1821 3323 1853
rect 2127 1819 2150 1821
rect 2070 1796 2150 1819
rect 1060 1731 1100 1771
rect 1660 1731 1700 1771
rect 1990 1731 2030 1771
rect 2290 1731 2330 1821
rect 2620 1731 2660 1821
rect 3220 1731 3260 1821
rect 3300 1820 3323 1821
rect 3357 1820 3380 1854
rect 3560 1898 3790 1901
rect 3560 1878 3733 1898
rect 3560 1844 3583 1878
rect 3617 1864 3733 1878
rect 3767 1864 3790 1898
rect 3617 1861 3790 1864
rect 3617 1844 3640 1861
rect 3560 1821 3640 1844
rect 3710 1841 3790 1861
rect 3300 1797 3380 1820
rect 4310 1811 4350 1941
rect 4490 1921 4570 1941
rect 3980 1771 4350 1811
rect 4390 1861 4470 1876
rect 4610 1861 4650 2031
rect 5580 2028 5960 2031
rect 5580 2027 5903 2028
rect 4890 1981 4970 2001
rect 5580 1993 5603 2027
rect 5637 1994 5903 2027
rect 5937 1994 5960 2028
rect 5637 1993 5960 1994
rect 5580 1991 5960 1993
rect 4890 1978 5546 1981
rect 4890 1944 4913 1978
rect 4947 1944 5546 1978
rect 5580 1970 5660 1991
rect 5880 1971 5960 1991
rect 6330 1981 6370 2031
rect 6510 1981 6590 2001
rect 6330 1978 6590 1981
rect 4890 1941 5546 1944
rect 4890 1921 4970 1941
rect 5506 1930 5546 1941
rect 5730 1931 5810 1951
rect 5660 1930 5810 1931
rect 5506 1928 5810 1930
rect 5250 1878 5330 1901
rect 5506 1894 5753 1928
rect 5787 1894 5810 1928
rect 5506 1891 5810 1894
rect 5506 1890 5660 1891
rect 5250 1861 5273 1878
rect 4390 1853 5273 1861
rect 4390 1819 4413 1853
rect 4447 1844 5273 1853
rect 5307 1844 5330 1878
rect 5730 1871 5810 1891
rect 6330 1944 6533 1978
rect 6567 1944 6590 1978
rect 6330 1941 6590 1944
rect 4447 1821 5330 1844
rect 4447 1819 4470 1821
rect 4390 1796 4470 1819
rect 3980 1731 4020 1771
rect 4310 1731 4350 1771
rect 4610 1731 4650 1821
rect 4920 1731 4960 1821
rect 5240 1731 5280 1821
rect 6330 1811 6370 1941
rect 6510 1921 6590 1941
rect 5700 1771 6370 1811
rect 6410 1861 6490 1876
rect 6630 1861 6670 2031
rect 6910 1981 6990 2001
rect 7340 1981 7420 2001
rect 6910 1978 7420 1981
rect 6910 1944 6933 1978
rect 6967 1944 7363 1978
rect 7397 1944 7420 1978
rect 6910 1941 7420 1944
rect 6910 1921 6990 1941
rect 7340 1921 7420 1941
rect 6410 1853 7488 1861
rect 6410 1819 6433 1853
rect 6467 1821 7488 1853
rect 6467 1819 6490 1821
rect 6410 1796 6490 1819
rect 5700 1731 5740 1771
rect 6000 1731 6040 1771
rect 6331 1731 6370 1771
rect 6630 1731 6670 1821
rect 6960 1731 7000 1821
rect 1040 1698 1120 1731
rect 1040 1664 1063 1698
rect 1097 1664 1120 1698
rect 1040 1618 1120 1664
rect 1040 1584 1063 1618
rect 1097 1584 1120 1618
rect 1040 1538 1120 1584
rect 1040 1504 1063 1538
rect 1097 1504 1120 1538
rect 1040 1481 1120 1504
rect 1340 1698 1420 1731
rect 1340 1664 1363 1698
rect 1397 1664 1420 1698
rect 1340 1618 1420 1664
rect 1340 1584 1363 1618
rect 1397 1584 1420 1618
rect 1340 1538 1420 1584
rect 1340 1504 1363 1538
rect 1397 1504 1420 1538
rect 1340 1481 1420 1504
rect 1640 1698 1720 1731
rect 1640 1664 1663 1698
rect 1697 1664 1720 1698
rect 1640 1618 1720 1664
rect 1640 1584 1663 1618
rect 1697 1584 1720 1618
rect 1640 1538 1720 1584
rect 1640 1504 1663 1538
rect 1697 1504 1720 1538
rect 1640 1481 1720 1504
rect 1820 1698 1900 1731
rect 1820 1664 1843 1698
rect 1877 1664 1900 1698
rect 1820 1618 1900 1664
rect 1820 1584 1843 1618
rect 1877 1584 1900 1618
rect 1820 1538 1900 1584
rect 1820 1504 1843 1538
rect 1877 1504 1900 1538
rect 1820 1481 1900 1504
rect 1970 1698 2050 1731
rect 1970 1664 1993 1698
rect 2027 1664 2050 1698
rect 1970 1618 2050 1664
rect 1970 1584 1993 1618
rect 2027 1584 2050 1618
rect 1970 1538 2050 1584
rect 1970 1504 1993 1538
rect 2027 1504 2050 1538
rect 1970 1481 2050 1504
rect 2120 1698 2200 1731
rect 2120 1664 2143 1698
rect 2177 1664 2200 1698
rect 2120 1618 2200 1664
rect 2120 1584 2143 1618
rect 2177 1584 2200 1618
rect 2120 1538 2200 1584
rect 2120 1504 2143 1538
rect 2177 1504 2200 1538
rect 2120 1481 2200 1504
rect 2270 1698 2350 1731
rect 2270 1664 2293 1698
rect 2327 1664 2350 1698
rect 2270 1618 2350 1664
rect 2270 1584 2293 1618
rect 2327 1584 2350 1618
rect 2270 1538 2350 1584
rect 2270 1504 2293 1538
rect 2327 1504 2350 1538
rect 2270 1481 2350 1504
rect 2420 1698 2500 1731
rect 2420 1664 2443 1698
rect 2477 1664 2500 1698
rect 2420 1618 2500 1664
rect 2420 1584 2443 1618
rect 2477 1584 2500 1618
rect 2420 1538 2500 1584
rect 2420 1504 2443 1538
rect 2477 1504 2500 1538
rect 2420 1481 2500 1504
rect 2600 1698 2680 1731
rect 2600 1664 2623 1698
rect 2657 1664 2680 1698
rect 2600 1618 2680 1664
rect 2600 1584 2623 1618
rect 2657 1584 2680 1618
rect 2600 1538 2680 1584
rect 2600 1504 2623 1538
rect 2657 1504 2680 1538
rect 2600 1481 2680 1504
rect 2900 1698 2980 1731
rect 2900 1664 2923 1698
rect 2957 1664 2980 1698
rect 2900 1618 2980 1664
rect 2900 1584 2923 1618
rect 2957 1584 2980 1618
rect 2900 1538 2980 1584
rect 2900 1504 2923 1538
rect 2957 1504 2980 1538
rect 2900 1481 2980 1504
rect 3200 1698 3280 1731
rect 3200 1664 3223 1698
rect 3257 1664 3280 1698
rect 3200 1618 3280 1664
rect 3200 1584 3223 1618
rect 3257 1584 3280 1618
rect 3200 1538 3280 1584
rect 3200 1504 3223 1538
rect 3257 1504 3280 1538
rect 3200 1481 3280 1504
rect 3660 1698 3740 1731
rect 3660 1664 3683 1698
rect 3717 1664 3740 1698
rect 3660 1618 3740 1664
rect 3660 1584 3683 1618
rect 3717 1584 3740 1618
rect 3660 1538 3740 1584
rect 3660 1504 3683 1538
rect 3717 1504 3740 1538
rect 3660 1481 3740 1504
rect 3960 1698 4040 1731
rect 3960 1664 3983 1698
rect 4017 1664 4040 1698
rect 3960 1618 4040 1664
rect 3960 1584 3983 1618
rect 4017 1584 4040 1618
rect 3960 1538 4040 1584
rect 3960 1504 3983 1538
rect 4017 1504 4040 1538
rect 3960 1481 4040 1504
rect 4140 1698 4220 1731
rect 4140 1664 4163 1698
rect 4197 1664 4220 1698
rect 4140 1618 4220 1664
rect 4140 1584 4163 1618
rect 4197 1584 4220 1618
rect 4140 1538 4220 1584
rect 4140 1504 4163 1538
rect 4197 1504 4220 1538
rect 4140 1481 4220 1504
rect 4290 1698 4370 1731
rect 4290 1664 4313 1698
rect 4347 1664 4370 1698
rect 4290 1618 4370 1664
rect 4290 1584 4313 1618
rect 4347 1584 4370 1618
rect 4290 1538 4370 1584
rect 4290 1504 4313 1538
rect 4347 1504 4370 1538
rect 4290 1481 4370 1504
rect 4440 1698 4520 1731
rect 4440 1664 4463 1698
rect 4497 1664 4520 1698
rect 4440 1618 4520 1664
rect 4440 1584 4463 1618
rect 4497 1584 4520 1618
rect 4440 1538 4520 1584
rect 4440 1504 4463 1538
rect 4497 1504 4520 1538
rect 4440 1481 4520 1504
rect 4590 1698 4670 1731
rect 4590 1664 4613 1698
rect 4647 1664 4670 1698
rect 4590 1618 4670 1664
rect 4590 1584 4613 1618
rect 4647 1584 4670 1618
rect 4590 1538 4670 1584
rect 4590 1504 4613 1538
rect 4647 1504 4670 1538
rect 4590 1481 4670 1504
rect 4740 1698 4820 1731
rect 4740 1664 4763 1698
rect 4797 1664 4820 1698
rect 4740 1618 4820 1664
rect 4740 1584 4763 1618
rect 4797 1584 4820 1618
rect 4740 1538 4820 1584
rect 4740 1504 4763 1538
rect 4797 1504 4820 1538
rect 4740 1481 4820 1504
rect 4920 1698 5000 1731
rect 4920 1664 4943 1698
rect 4977 1664 5000 1698
rect 4920 1618 5000 1664
rect 4920 1584 4943 1618
rect 4977 1584 5000 1618
rect 4920 1538 5000 1584
rect 4920 1504 4943 1538
rect 4977 1504 5000 1538
rect 4920 1481 5000 1504
rect 5070 1698 5150 1731
rect 5070 1664 5093 1698
rect 5127 1664 5150 1698
rect 5070 1618 5150 1664
rect 5070 1584 5093 1618
rect 5127 1584 5150 1618
rect 5070 1538 5150 1584
rect 5070 1504 5093 1538
rect 5127 1504 5150 1538
rect 5070 1481 5150 1504
rect 5220 1698 5300 1731
rect 5220 1664 5243 1698
rect 5277 1664 5300 1698
rect 5220 1618 5300 1664
rect 5220 1584 5243 1618
rect 5277 1584 5300 1618
rect 5220 1538 5300 1584
rect 5220 1504 5243 1538
rect 5277 1504 5300 1538
rect 5220 1481 5300 1504
rect 5680 1698 5760 1731
rect 5680 1664 5703 1698
rect 5737 1664 5760 1698
rect 5680 1618 5760 1664
rect 5680 1584 5703 1618
rect 5737 1584 5760 1618
rect 5680 1538 5760 1584
rect 5680 1504 5703 1538
rect 5737 1504 5760 1538
rect 5680 1481 5760 1504
rect 5830 1698 5910 1731
rect 5830 1664 5853 1698
rect 5887 1664 5910 1698
rect 5830 1618 5910 1664
rect 5830 1584 5853 1618
rect 5887 1584 5910 1618
rect 5830 1538 5910 1584
rect 5830 1504 5853 1538
rect 5887 1504 5910 1538
rect 5830 1481 5910 1504
rect 5980 1698 6060 1731
rect 5980 1664 6003 1698
rect 6037 1664 6060 1698
rect 5980 1618 6060 1664
rect 5980 1584 6003 1618
rect 6037 1584 6060 1618
rect 5980 1538 6060 1584
rect 5980 1504 6003 1538
rect 6037 1504 6060 1538
rect 5980 1481 6060 1504
rect 6160 1698 6240 1731
rect 6160 1664 6183 1698
rect 6217 1664 6240 1698
rect 6160 1618 6240 1664
rect 6160 1584 6183 1618
rect 6217 1584 6240 1618
rect 6160 1538 6240 1584
rect 6160 1504 6183 1538
rect 6217 1504 6240 1538
rect 6160 1481 6240 1504
rect 6310 1698 6390 1731
rect 6310 1664 6333 1698
rect 6367 1664 6390 1698
rect 6310 1618 6390 1664
rect 6310 1584 6333 1618
rect 6367 1584 6390 1618
rect 6310 1538 6390 1584
rect 6310 1504 6333 1538
rect 6367 1504 6390 1538
rect 6310 1481 6390 1504
rect 6460 1698 6540 1731
rect 6460 1664 6483 1698
rect 6517 1664 6540 1698
rect 6460 1618 6540 1664
rect 6460 1584 6483 1618
rect 6517 1584 6540 1618
rect 6460 1538 6540 1584
rect 6460 1504 6483 1538
rect 6517 1504 6540 1538
rect 6460 1481 6540 1504
rect 6610 1698 6690 1731
rect 6610 1664 6633 1698
rect 6667 1664 6690 1698
rect 6610 1618 6690 1664
rect 6610 1584 6633 1618
rect 6667 1584 6690 1618
rect 6610 1538 6690 1584
rect 6610 1504 6633 1538
rect 6667 1504 6690 1538
rect 6610 1481 6690 1504
rect 6760 1698 6840 1731
rect 6760 1664 6783 1698
rect 6817 1664 6840 1698
rect 6760 1618 6840 1664
rect 6760 1584 6783 1618
rect 6817 1584 6840 1618
rect 6760 1538 6840 1584
rect 6760 1504 6783 1538
rect 6817 1504 6840 1538
rect 6760 1481 6840 1504
rect 6940 1698 7020 1731
rect 6940 1664 6963 1698
rect 6997 1664 7020 1698
rect 6940 1618 7020 1664
rect 6940 1584 6963 1618
rect 6997 1584 7020 1618
rect 6940 1538 7020 1584
rect 6940 1504 6963 1538
rect 6997 1504 7020 1538
rect 6940 1481 7020 1504
rect 7240 1698 7320 1731
rect 7240 1664 7263 1698
rect 7297 1664 7320 1698
rect 7240 1618 7320 1664
rect 7240 1584 7263 1618
rect 7297 1584 7320 1618
rect 7240 1538 7320 1584
rect 7240 1504 7263 1538
rect 7297 1504 7320 1538
rect 7240 1481 7320 1504
rect 1129 1421 1209 1441
rect 1920 1421 2000 1441
rect 2320 1421 2400 1441
rect 4240 1421 4320 1441
rect 4640 1421 4720 1441
rect 5742 1421 5822 1441
rect 6260 1421 6340 1441
rect 6660 1421 6740 1441
rect 1020 1418 4720 1421
rect 1020 1384 1152 1418
rect 1186 1384 1943 1418
rect 1977 1384 2343 1418
rect 2377 1384 4263 1418
rect 4297 1384 4663 1418
rect 4697 1384 4720 1418
rect 1020 1381 4720 1384
rect 1129 1361 1209 1381
rect 1920 1361 2000 1381
rect 2320 1361 2400 1381
rect 4240 1361 4320 1381
rect 4640 1361 4720 1381
rect 5487 1418 6740 1421
rect 5487 1384 5765 1418
rect 5799 1384 6283 1418
rect 6317 1384 6683 1418
rect 6717 1384 6740 1418
rect 5487 1381 6740 1384
rect 912 1298 3300 1321
rect 912 1264 935 1298
rect 969 1264 1103 1298
rect 1137 1264 1183 1298
rect 1217 1264 1263 1298
rect 1297 1264 1343 1298
rect 1377 1264 1423 1298
rect 1457 1264 1503 1298
rect 1537 1264 1583 1298
rect 1617 1264 1663 1298
rect 1697 1264 1743 1298
rect 1777 1264 1823 1298
rect 1857 1264 1903 1298
rect 1937 1264 1983 1298
rect 2017 1264 2063 1298
rect 2097 1264 2143 1298
rect 2177 1264 2223 1298
rect 2257 1264 2303 1298
rect 2337 1264 2383 1298
rect 2417 1264 2463 1298
rect 2497 1264 2543 1298
rect 2577 1264 2623 1298
rect 2657 1264 2703 1298
rect 2737 1264 2783 1298
rect 2817 1264 2863 1298
rect 2897 1264 2943 1298
rect 2977 1264 3023 1298
rect 3057 1264 3103 1298
rect 3137 1264 3183 1298
rect 3217 1264 3300 1298
rect 912 1241 3300 1264
rect 3640 1298 5320 1321
rect 3640 1264 3663 1298
rect 3697 1264 3743 1298
rect 3777 1264 3823 1298
rect 3857 1264 3903 1298
rect 3937 1264 3983 1298
rect 4017 1264 4063 1298
rect 4097 1264 4143 1298
rect 4177 1264 4223 1298
rect 4257 1264 4303 1298
rect 4337 1264 4383 1298
rect 4417 1264 4463 1298
rect 4497 1264 4543 1298
rect 4577 1264 4623 1298
rect 4657 1264 4703 1298
rect 4737 1264 4783 1298
rect 4817 1264 4863 1298
rect 4897 1264 4943 1298
rect 4977 1264 5023 1298
rect 5057 1264 5103 1298
rect 5137 1264 5183 1298
rect 5217 1264 5263 1298
rect 5297 1264 5320 1298
rect 3640 1241 5320 1264
rect 1128 1181 1208 1201
rect 1920 1181 2000 1201
rect 2320 1181 2400 1201
rect 4240 1181 4320 1201
rect 4640 1181 4720 1201
rect 5073 1181 5153 1202
rect 5487 1181 5527 1381
rect 5742 1361 5822 1381
rect 6260 1361 6340 1381
rect 6660 1361 6740 1381
rect 5660 1298 7340 1321
rect 5660 1264 5683 1298
rect 5717 1264 5763 1298
rect 5797 1264 5843 1298
rect 5877 1264 5923 1298
rect 5957 1264 6003 1298
rect 6037 1264 6083 1298
rect 6117 1264 6163 1298
rect 6197 1264 6243 1298
rect 6277 1264 6323 1298
rect 6357 1264 6403 1298
rect 6437 1264 6483 1298
rect 6517 1264 6563 1298
rect 6597 1264 6643 1298
rect 6677 1264 6723 1298
rect 6757 1264 6803 1298
rect 6837 1264 6883 1298
rect 6917 1264 6963 1298
rect 6997 1264 7043 1298
rect 7077 1264 7123 1298
rect 7157 1264 7203 1298
rect 7237 1264 7283 1298
rect 7317 1264 7340 1298
rect 5660 1241 7340 1264
rect 1128 1178 2400 1181
rect 1128 1144 1151 1178
rect 1185 1144 1943 1178
rect 1977 1144 2343 1178
rect 2377 1144 2400 1178
rect 1128 1141 2400 1144
rect 3640 1179 5527 1181
rect 3640 1178 5096 1179
rect 3640 1144 4263 1178
rect 4297 1144 4663 1178
rect 4697 1145 5096 1178
rect 5130 1145 5527 1179
rect 4697 1144 5527 1145
rect 3640 1141 5527 1144
rect 5922 1181 6002 1201
rect 6260 1181 6340 1201
rect 6660 1181 6740 1201
rect 5922 1178 7340 1181
rect 5922 1144 5945 1178
rect 5979 1144 6283 1178
rect 6317 1144 6683 1178
rect 6717 1144 7340 1178
rect 5922 1141 7340 1144
rect 1128 1121 1208 1141
rect 1920 1121 2000 1141
rect 2320 1121 2400 1141
rect 4240 1121 4320 1141
rect 4640 1121 4720 1141
rect 5073 1122 5153 1141
rect 5922 1121 6002 1141
rect 6260 1121 6340 1141
rect 6660 1121 6740 1141
rect 1340 1058 1420 1081
rect 1340 1024 1363 1058
rect 1397 1024 1420 1058
rect 1340 978 1420 1024
rect 1340 944 1363 978
rect 1397 944 1420 978
rect 1340 898 1420 944
rect 1340 864 1363 898
rect 1397 864 1420 898
rect 1340 831 1420 864
rect 1490 1058 1570 1081
rect 1490 1024 1513 1058
rect 1547 1024 1570 1058
rect 1490 978 1570 1024
rect 1490 944 1513 978
rect 1547 944 1570 978
rect 1490 898 1570 944
rect 1490 864 1513 898
rect 1547 864 1570 898
rect 1490 831 1570 864
rect 1640 1058 1720 1081
rect 1640 1024 1663 1058
rect 1697 1024 1720 1058
rect 1640 978 1720 1024
rect 1640 944 1663 978
rect 1697 944 1720 978
rect 1640 898 1720 944
rect 1640 864 1663 898
rect 1697 864 1720 898
rect 1640 831 1720 864
rect 1820 1058 1900 1081
rect 1820 1024 1843 1058
rect 1877 1024 1900 1058
rect 1820 978 1900 1024
rect 1820 944 1843 978
rect 1877 944 1900 978
rect 1820 898 1900 944
rect 1820 864 1843 898
rect 1877 864 1900 898
rect 1820 831 1900 864
rect 1970 1058 2050 1081
rect 1970 1024 1993 1058
rect 2027 1024 2050 1058
rect 1970 978 2050 1024
rect 1970 944 1993 978
rect 2027 944 2050 978
rect 1970 898 2050 944
rect 1970 864 1993 898
rect 2027 864 2050 898
rect 1970 831 2050 864
rect 2120 1058 2200 1081
rect 2120 1024 2143 1058
rect 2177 1024 2200 1058
rect 2120 978 2200 1024
rect 2120 944 2143 978
rect 2177 944 2200 978
rect 2120 898 2200 944
rect 2120 864 2143 898
rect 2177 864 2200 898
rect 2120 831 2200 864
rect 2270 1058 2350 1081
rect 2270 1024 2293 1058
rect 2327 1024 2350 1058
rect 2270 978 2350 1024
rect 2270 944 2293 978
rect 2327 944 2350 978
rect 2270 898 2350 944
rect 2270 864 2293 898
rect 2327 864 2350 898
rect 2270 831 2350 864
rect 2420 1058 2500 1081
rect 2420 1024 2443 1058
rect 2477 1024 2500 1058
rect 2420 978 2500 1024
rect 2420 944 2443 978
rect 2477 944 2500 978
rect 2420 898 2500 944
rect 2420 864 2443 898
rect 2477 864 2500 898
rect 2420 831 2500 864
rect 2600 1058 2680 1081
rect 2600 1024 2623 1058
rect 2657 1024 2680 1058
rect 2600 978 2680 1024
rect 2600 944 2623 978
rect 2657 944 2680 978
rect 2600 898 2680 944
rect 2600 864 2623 898
rect 2657 864 2680 898
rect 2600 831 2680 864
rect 2900 1058 2980 1081
rect 2900 1024 2923 1058
rect 2957 1024 2980 1058
rect 2900 978 2980 1024
rect 2900 944 2923 978
rect 2957 944 2980 978
rect 2900 898 2980 944
rect 2900 864 2923 898
rect 2957 864 2980 898
rect 2900 831 2980 864
rect 3660 1058 3740 1081
rect 3660 1024 3683 1058
rect 3717 1024 3740 1058
rect 3660 978 3740 1024
rect 3660 944 3683 978
rect 3717 944 3740 978
rect 3660 898 3740 944
rect 3660 864 3683 898
rect 3717 864 3740 898
rect 3660 831 3740 864
rect 3810 1058 3890 1081
rect 3810 1024 3833 1058
rect 3867 1024 3890 1058
rect 3810 978 3890 1024
rect 3810 944 3833 978
rect 3867 944 3890 978
rect 3810 898 3890 944
rect 3810 864 3833 898
rect 3867 864 3890 898
rect 3810 831 3890 864
rect 3960 1058 4040 1081
rect 3960 1024 3983 1058
rect 4017 1024 4040 1058
rect 3960 978 4040 1024
rect 3960 944 3983 978
rect 4017 944 4040 978
rect 3960 898 4040 944
rect 3960 864 3983 898
rect 4017 864 4040 898
rect 3960 831 4040 864
rect 4140 1058 4220 1081
rect 4140 1024 4163 1058
rect 4197 1024 4220 1058
rect 4140 978 4220 1024
rect 4140 944 4163 978
rect 4197 944 4220 978
rect 4140 898 4220 944
rect 4140 864 4163 898
rect 4197 864 4220 898
rect 4140 831 4220 864
rect 4290 1058 4370 1081
rect 4290 1024 4313 1058
rect 4347 1024 4370 1058
rect 4290 978 4370 1024
rect 4290 944 4313 978
rect 4347 944 4370 978
rect 4290 898 4370 944
rect 4290 864 4313 898
rect 4347 864 4370 898
rect 4290 831 4370 864
rect 4440 1058 4520 1081
rect 4440 1024 4463 1058
rect 4497 1024 4520 1058
rect 4440 978 4520 1024
rect 4440 944 4463 978
rect 4497 944 4520 978
rect 4440 898 4520 944
rect 4440 864 4463 898
rect 4497 864 4520 898
rect 4440 831 4520 864
rect 4590 1058 4670 1081
rect 4590 1024 4613 1058
rect 4647 1024 4670 1058
rect 4590 978 4670 1024
rect 4590 944 4613 978
rect 4647 944 4670 978
rect 4590 898 4670 944
rect 4590 864 4613 898
rect 4647 864 4670 898
rect 4590 831 4670 864
rect 4740 1058 4820 1081
rect 4740 1024 4763 1058
rect 4797 1024 4820 1058
rect 4740 978 4820 1024
rect 4740 944 4763 978
rect 4797 944 4820 978
rect 4740 898 4820 944
rect 4740 864 4763 898
rect 4797 864 4820 898
rect 4740 831 4820 864
rect 4920 1058 5000 1081
rect 4920 1024 4943 1058
rect 4977 1024 5000 1058
rect 4920 978 5000 1024
rect 4920 944 4943 978
rect 4977 944 5000 978
rect 4920 898 5000 944
rect 4920 864 4943 898
rect 4977 864 5000 898
rect 4920 831 5000 864
rect 5220 1058 5300 1081
rect 5220 1024 5243 1058
rect 5277 1024 5300 1058
rect 5220 978 5300 1024
rect 5220 944 5243 978
rect 5277 944 5300 978
rect 5220 898 5300 944
rect 5220 864 5243 898
rect 5277 864 5300 898
rect 5220 831 5300 864
rect 5680 1058 5760 1081
rect 5680 1024 5703 1058
rect 5737 1024 5760 1058
rect 5680 978 5760 1024
rect 5680 944 5703 978
rect 5737 944 5760 978
rect 5680 898 5760 944
rect 5680 864 5703 898
rect 5737 864 5760 898
rect 5680 831 5760 864
rect 5830 1058 5910 1081
rect 5830 1024 5853 1058
rect 5887 1024 5910 1058
rect 5830 978 5910 1024
rect 5830 944 5853 978
rect 5887 944 5910 978
rect 5830 898 5910 944
rect 5830 864 5853 898
rect 5887 864 5910 898
rect 5830 831 5910 864
rect 5980 1058 6060 1081
rect 5980 1024 6003 1058
rect 6037 1024 6060 1058
rect 5980 978 6060 1024
rect 5980 944 6003 978
rect 6037 944 6060 978
rect 5980 898 6060 944
rect 5980 864 6003 898
rect 6037 864 6060 898
rect 5980 831 6060 864
rect 6160 1058 6240 1081
rect 6160 1024 6183 1058
rect 6217 1024 6240 1058
rect 6160 978 6240 1024
rect 6160 944 6183 978
rect 6217 944 6240 978
rect 6160 898 6240 944
rect 6160 864 6183 898
rect 6217 864 6240 898
rect 6160 831 6240 864
rect 6310 1058 6390 1081
rect 6310 1024 6333 1058
rect 6367 1024 6390 1058
rect 6310 978 6390 1024
rect 6310 944 6333 978
rect 6367 944 6390 978
rect 6310 898 6390 944
rect 6310 864 6333 898
rect 6367 864 6390 898
rect 6310 831 6390 864
rect 6460 1058 6540 1081
rect 6460 1024 6483 1058
rect 6517 1024 6540 1058
rect 6460 978 6540 1024
rect 6460 944 6483 978
rect 6517 944 6540 978
rect 6460 898 6540 944
rect 6460 864 6483 898
rect 6517 864 6540 898
rect 6460 831 6540 864
rect 6610 1058 6690 1081
rect 6610 1024 6633 1058
rect 6667 1024 6690 1058
rect 6610 978 6690 1024
rect 6610 944 6633 978
rect 6667 944 6690 978
rect 6610 898 6690 944
rect 6610 864 6633 898
rect 6667 864 6690 898
rect 6610 831 6690 864
rect 6760 1058 6840 1081
rect 6760 1024 6783 1058
rect 6817 1024 6840 1058
rect 6760 978 6840 1024
rect 6760 944 6783 978
rect 6817 944 6840 978
rect 6760 898 6840 944
rect 6760 864 6783 898
rect 6817 864 6840 898
rect 6760 831 6840 864
rect 6940 1058 7020 1081
rect 6940 1024 6963 1058
rect 6997 1024 7020 1058
rect 6940 978 7020 1024
rect 6940 944 6963 978
rect 6997 944 7020 978
rect 6940 898 7020 944
rect 7240 1058 7320 1081
rect 7240 1024 7263 1058
rect 7297 1024 7320 1058
rect 7240 978 7320 1024
rect 7240 944 7263 978
rect 7297 944 7320 978
rect 6940 864 6963 898
rect 6997 864 7020 898
rect 6940 831 7020 864
rect 7090 888 7170 911
rect 7090 854 7113 888
rect 7147 854 7170 888
rect 7090 831 7170 854
rect 7240 898 7320 944
rect 7240 864 7263 898
rect 7297 864 7320 898
rect 7240 831 7320 864
rect 1360 791 1400 831
rect 1660 791 1700 831
rect 1991 791 2030 831
rect 1360 751 2030 791
rect 228 688 308 711
rect 228 654 251 688
rect 285 671 308 688
rect 1390 671 1470 691
rect 285 668 1470 671
rect 285 654 1413 668
rect 228 634 1413 654
rect 1447 634 1470 668
rect 228 631 1470 634
rect 1390 611 1470 631
rect 1990 621 2030 751
rect 2070 743 2150 766
rect 2070 709 2093 743
rect 2127 741 2150 743
rect 2290 741 2330 831
rect 2620 741 2660 831
rect 3680 791 3720 831
rect 3980 791 4020 831
rect 4311 791 4350 831
rect 3000 741 3080 761
rect 3680 751 4350 791
rect 2127 738 3080 741
rect 2127 709 3023 738
rect 2070 704 3023 709
rect 3057 704 3080 738
rect 2070 701 3080 704
rect 2070 686 2150 701
rect 2170 621 2250 641
rect 1990 618 2250 621
rect 570 574 650 597
rect 570 540 593 574
rect 627 571 650 574
rect 1540 571 1620 591
rect 627 568 1620 571
rect 627 540 1563 568
rect 570 534 1563 540
rect 1597 534 1620 568
rect 570 531 1620 534
rect 1990 584 2193 618
rect 2227 584 2250 618
rect 1990 581 2250 584
rect 1990 531 2030 581
rect 2170 561 2250 581
rect 2290 531 2330 701
rect 3000 681 3080 701
rect 3710 671 3790 691
rect 3270 668 3790 671
rect 2570 621 2650 641
rect 3270 634 3733 668
rect 3767 634 3790 668
rect 3270 631 3790 634
rect 3270 621 3310 631
rect 2570 618 3310 621
rect 2570 584 2593 618
rect 2627 584 3310 618
rect 3710 611 3790 631
rect 4310 621 4350 751
rect 4390 743 4470 766
rect 4390 709 4413 743
rect 4447 741 4470 743
rect 4610 741 4650 831
rect 4940 741 4980 831
rect 5700 761 5740 831
rect 5660 741 5740 761
rect 6020 741 6060 831
rect 6330 741 6370 831
rect 6630 791 6670 831
rect 6960 791 7000 831
rect 6510 743 6590 766
rect 6510 741 6533 743
rect 4447 709 5625 741
rect 4390 701 5625 709
rect 4390 686 4470 701
rect 4490 621 4570 641
rect 4310 618 4570 621
rect 2570 581 3310 584
rect 2570 561 2650 581
rect 3560 571 3640 591
rect 3860 571 3940 591
rect 3560 568 3940 571
rect 3560 534 3583 568
rect 3617 534 3883 568
rect 3917 534 3940 568
rect 3560 531 3940 534
rect 4310 584 4513 618
rect 4547 584 4570 618
rect 4310 581 4570 584
rect 4310 531 4350 581
rect 4490 561 4570 581
rect 4610 531 4650 701
rect 4890 621 4970 641
rect 5471 621 5551 641
rect 4890 618 5551 621
rect 4890 584 4913 618
rect 4947 584 5494 618
rect 5528 584 5551 618
rect 4890 581 5551 584
rect 4890 561 4970 581
rect 5471 561 5551 581
rect 570 517 650 531
rect 1540 511 1620 531
rect 1820 498 1900 521
rect 342 471 422 491
rect 1670 471 1750 491
rect 342 468 1750 471
rect 342 434 365 468
rect 399 434 1693 468
rect 1727 434 1750 468
rect 342 431 1750 434
rect 342 411 422 431
rect 1670 411 1750 431
rect 1820 464 1843 498
rect 1877 464 1900 498
rect 1820 418 1900 464
rect 1820 384 1843 418
rect 1877 384 1900 418
rect 456 351 536 371
rect 1670 351 1750 371
rect 456 348 1750 351
rect 456 314 479 348
rect 513 314 1693 348
rect 1727 314 1750 348
rect 456 311 1750 314
rect 456 291 536 311
rect 1670 291 1750 311
rect 1820 338 1900 384
rect 1820 304 1843 338
rect 1877 304 1900 338
rect 1820 271 1900 304
rect 1970 498 2050 531
rect 1970 464 1993 498
rect 2027 464 2050 498
rect 1970 418 2050 464
rect 1970 384 1993 418
rect 2027 384 2050 418
rect 1970 338 2050 384
rect 1970 304 1993 338
rect 2027 304 2050 338
rect 1970 271 2050 304
rect 2120 498 2200 521
rect 2120 464 2143 498
rect 2177 464 2200 498
rect 2120 418 2200 464
rect 2120 384 2143 418
rect 2177 384 2200 418
rect 2120 338 2200 384
rect 2120 304 2143 338
rect 2177 304 2200 338
rect 2120 271 2200 304
rect 2270 498 2350 531
rect 2270 464 2293 498
rect 2327 464 2350 498
rect 2270 418 2350 464
rect 2270 384 2293 418
rect 2327 384 2350 418
rect 2270 338 2350 384
rect 2270 304 2293 338
rect 2327 304 2350 338
rect 2270 271 2350 304
rect 2420 498 2500 521
rect 3560 511 3640 531
rect 3860 511 3940 531
rect 2420 464 2443 498
rect 2477 464 2500 498
rect 2420 418 2500 464
rect 2420 384 2443 418
rect 2477 384 2500 418
rect 2650 468 2730 491
rect 2650 434 2673 468
rect 2707 434 2730 468
rect 2650 411 2730 434
rect 3000 488 3080 511
rect 4140 498 4220 521
rect 3000 454 3023 488
rect 3057 471 3080 488
rect 3990 471 4070 491
rect 3057 468 4070 471
rect 3057 454 4013 468
rect 3000 434 4013 454
rect 4047 434 4070 468
rect 3000 431 4070 434
rect 3990 411 4070 431
rect 4140 464 4163 498
rect 4197 464 4220 498
rect 4140 418 4220 464
rect 2420 338 2500 384
rect 4140 384 4163 418
rect 4197 384 4220 418
rect 2420 304 2443 338
rect 2477 304 2500 338
rect 2420 271 2500 304
rect 2800 348 2880 371
rect 2800 314 2823 348
rect 2857 314 2880 348
rect 2800 291 2880 314
rect 3054 351 3134 371
rect 3990 351 4070 371
rect 3054 348 4070 351
rect 3054 314 3077 348
rect 3111 314 4013 348
rect 4047 314 4070 348
rect 3054 311 4070 314
rect 3054 291 3134 311
rect 3990 291 4070 311
rect 4140 338 4220 384
rect 4140 304 4163 338
rect 4197 304 4220 338
rect 4140 271 4220 304
rect 4290 498 4370 531
rect 4290 464 4313 498
rect 4347 464 4370 498
rect 4290 418 4370 464
rect 4290 384 4313 418
rect 4347 384 4370 418
rect 4290 338 4370 384
rect 4290 304 4313 338
rect 4347 304 4370 338
rect 4290 271 4370 304
rect 4440 498 4520 521
rect 4440 464 4463 498
rect 4497 464 4520 498
rect 4440 418 4520 464
rect 4440 384 4463 418
rect 4497 384 4520 418
rect 4440 338 4520 384
rect 4440 304 4463 338
rect 4497 304 4520 338
rect 4440 271 4520 304
rect 4590 498 4670 531
rect 4590 464 4613 498
rect 4647 464 4670 498
rect 4590 418 4670 464
rect 4590 384 4613 418
rect 4647 384 4670 418
rect 4590 338 4670 384
rect 4590 304 4613 338
rect 4647 304 4670 338
rect 4590 271 4670 304
rect 4740 498 4820 521
rect 4740 464 4763 498
rect 4797 464 4820 498
rect 5585 501 5625 701
rect 5660 738 6533 741
rect 5660 704 5683 738
rect 5717 709 6533 738
rect 6567 709 6590 743
rect 5717 704 6590 709
rect 5660 701 6590 704
rect 5660 681 5740 701
rect 5660 621 5740 641
rect 6010 621 6090 641
rect 5660 618 6090 621
rect 5660 584 5683 618
rect 5717 584 6033 618
rect 6067 584 6090 618
rect 5660 581 6090 584
rect 5660 561 5740 581
rect 6010 561 6090 581
rect 6330 531 6370 701
rect 6510 686 6590 701
rect 6630 751 7000 791
rect 6410 621 6490 641
rect 6630 621 6670 751
rect 7111 701 7151 831
rect 7060 661 7151 701
rect 7190 701 7270 721
rect 7334 701 7414 722
rect 7190 699 7414 701
rect 7190 698 7357 699
rect 7190 664 7213 698
rect 7247 665 7357 698
rect 7391 665 7414 699
rect 7247 664 7414 665
rect 7190 661 7414 664
rect 7060 621 7100 661
rect 7190 641 7270 661
rect 7334 642 7414 661
rect 6410 618 6670 621
rect 6410 584 6433 618
rect 6467 584 6670 618
rect 6410 581 6670 584
rect 6410 561 6490 581
rect 6630 531 6670 581
rect 7040 601 7120 621
rect 7040 598 7340 601
rect 7040 564 7063 598
rect 7097 564 7340 598
rect 7040 561 7340 564
rect 7040 541 7120 561
rect 5930 501 6010 521
rect 5585 498 6010 501
rect 4740 418 4820 464
rect 4740 384 4763 418
rect 4797 384 4820 418
rect 4970 468 5050 491
rect 4970 434 4993 468
rect 5027 434 5050 468
rect 5585 464 5953 498
rect 5987 464 6010 498
rect 5585 461 6010 464
rect 5930 441 6010 461
rect 6160 498 6240 521
rect 6160 464 6183 498
rect 6217 464 6240 498
rect 4970 411 5050 434
rect 6160 418 6240 464
rect 4740 338 4820 384
rect 5730 378 5810 401
rect 4740 304 4763 338
rect 4797 304 4820 338
rect 4740 271 4820 304
rect 5120 348 5200 371
rect 5120 314 5143 348
rect 5177 314 5200 348
rect 5730 344 5753 378
rect 5787 344 5810 378
rect 5730 321 5810 344
rect 6160 384 6183 418
rect 6217 384 6240 418
rect 6160 338 6240 384
rect 5120 291 5200 314
rect 6160 304 6183 338
rect 6217 304 6240 338
rect 6160 271 6240 304
rect 6310 498 6390 531
rect 6310 464 6333 498
rect 6367 464 6390 498
rect 6310 418 6390 464
rect 6310 384 6333 418
rect 6367 384 6390 418
rect 6310 338 6390 384
rect 6310 304 6333 338
rect 6367 304 6390 338
rect 6310 271 6390 304
rect 6460 498 6540 521
rect 6460 464 6483 498
rect 6517 464 6540 498
rect 6460 418 6540 464
rect 6460 384 6483 418
rect 6517 384 6540 418
rect 6460 338 6540 384
rect 6460 304 6483 338
rect 6517 304 6540 338
rect 6460 271 6540 304
rect 6610 498 6690 531
rect 6610 464 6633 498
rect 6667 464 6690 498
rect 6610 418 6690 464
rect 6610 384 6633 418
rect 6667 384 6690 418
rect 6610 338 6690 384
rect 6610 304 6633 338
rect 6667 304 6690 338
rect 6610 271 6690 304
rect 6760 498 6840 521
rect 6760 464 6783 498
rect 6817 464 6840 498
rect 6760 418 6840 464
rect 6910 501 6990 521
rect 6910 498 7340 501
rect 6910 464 6933 498
rect 6967 464 7340 498
rect 6910 461 7340 464
rect 6910 441 6990 461
rect 6760 384 6783 418
rect 6817 384 6840 418
rect 6760 338 6840 384
rect 6760 304 6783 338
rect 6817 304 6840 338
rect 6910 381 6990 401
rect 7448 381 7488 1821
rect 6910 378 7488 381
rect 6910 344 6933 378
rect 6967 344 7488 378
rect 6910 341 7488 344
rect 6910 321 6990 341
rect 6760 271 6840 304
rect 1320 118 3000 141
rect 1320 84 1343 118
rect 1377 84 1423 118
rect 1457 84 1503 118
rect 1537 84 1583 118
rect 1617 84 1663 118
rect 1697 84 1743 118
rect 1777 84 1823 118
rect 1857 84 1903 118
rect 1937 84 1983 118
rect 2017 84 2063 118
rect 2097 84 2143 118
rect 2177 84 2223 118
rect 2257 84 2303 118
rect 2337 84 2383 118
rect 2417 84 2463 118
rect 2497 84 2543 118
rect 2577 84 2623 118
rect 2657 84 2703 118
rect 2737 84 2783 118
rect 2817 84 2863 118
rect 2897 84 2943 118
rect 2977 84 3000 118
rect 1320 61 3000 84
rect 3640 118 5592 141
rect 3640 84 3663 118
rect 3697 84 3743 118
rect 3777 84 3823 118
rect 3857 84 3903 118
rect 3937 84 3983 118
rect 4017 84 4063 118
rect 4097 84 4143 118
rect 4177 84 4223 118
rect 4257 84 4303 118
rect 4337 84 4383 118
rect 4417 84 4463 118
rect 4497 84 4543 118
rect 4577 84 4623 118
rect 4657 84 4703 118
rect 4737 84 4783 118
rect 4817 84 4863 118
rect 4897 84 4943 118
rect 4977 84 5023 118
rect 5057 84 5103 118
rect 5137 84 5183 118
rect 5217 84 5263 118
rect 5297 84 5592 118
rect 3640 61 5592 84
rect 5660 118 7340 141
rect 5660 84 5683 118
rect 5717 84 5763 118
rect 5797 84 5843 118
rect 5877 84 5923 118
rect 5957 84 6003 118
rect 6037 84 6083 118
rect 6117 84 6163 118
rect 6197 84 6243 118
rect 6277 84 6323 118
rect 6357 84 6403 118
rect 6437 84 6483 118
rect 6517 84 6563 118
rect 6597 84 6643 118
rect 6677 84 6723 118
rect 6757 84 6803 118
rect 6837 84 6883 118
rect 6917 84 6963 118
rect 6997 84 7043 118
rect 7077 84 7123 118
rect 7157 84 7203 118
rect 7237 84 7283 118
rect 7317 84 7340 118
rect 5660 61 7340 84
rect 5512 -319 5592 61
rect 1020 -342 3300 -319
rect 1020 -376 1103 -342
rect 1137 -376 1183 -342
rect 1217 -376 1263 -342
rect 1297 -376 1343 -342
rect 1377 -376 1423 -342
rect 1457 -376 1503 -342
rect 1537 -376 1583 -342
rect 1617 -376 1663 -342
rect 1697 -376 1743 -342
rect 1777 -376 1823 -342
rect 1857 -376 1903 -342
rect 1937 -376 1983 -342
rect 2017 -376 2063 -342
rect 2097 -376 2143 -342
rect 2177 -376 2223 -342
rect 2257 -376 2303 -342
rect 2337 -376 2383 -342
rect 2417 -376 2463 -342
rect 2497 -376 2543 -342
rect 2577 -376 2623 -342
rect 2657 -376 2703 -342
rect 2737 -376 2783 -342
rect 2817 -376 2863 -342
rect 2897 -376 2943 -342
rect 2977 -376 3023 -342
rect 3057 -376 3103 -342
rect 3137 -376 3183 -342
rect 3217 -376 3300 -342
rect 1020 -399 3300 -376
rect 3660 -342 5040 -319
rect 3660 -376 3693 -342
rect 3727 -376 3773 -342
rect 3807 -376 3853 -342
rect 3887 -376 3933 -342
rect 3967 -376 4013 -342
rect 4047 -376 4093 -342
rect 4127 -376 4173 -342
rect 4207 -376 4253 -342
rect 4287 -376 4333 -342
rect 4367 -376 4413 -342
rect 4447 -376 4493 -342
rect 4527 -376 4573 -342
rect 4607 -376 4653 -342
rect 4687 -376 4733 -342
rect 4767 -376 4813 -342
rect 4847 -376 4893 -342
rect 4927 -376 4973 -342
rect 5007 -376 5040 -342
rect 3660 -399 5040 -376
rect 5390 -342 7070 -319
rect 5390 -376 5413 -342
rect 5447 -376 5493 -342
rect 5527 -376 5573 -342
rect 5607 -376 5653 -342
rect 5687 -376 5733 -342
rect 5767 -376 5813 -342
rect 5847 -376 5893 -342
rect 5927 -376 5973 -342
rect 6007 -376 6053 -342
rect 6087 -376 6133 -342
rect 6167 -376 6213 -342
rect 6247 -376 6293 -342
rect 6327 -376 6373 -342
rect 6407 -376 6453 -342
rect 6487 -376 6533 -342
rect 6567 -376 6613 -342
rect 6647 -376 6693 -342
rect 6727 -376 6773 -342
rect 6807 -376 6853 -342
rect 6887 -376 6933 -342
rect 6967 -376 7013 -342
rect 7047 -376 7070 -342
rect 5390 -399 7070 -376
rect 1410 -469 1490 -449
rect 1540 -469 1620 -449
rect 456 -472 1620 -469
rect 456 -492 1433 -472
rect 456 -526 479 -492
rect 513 -506 1433 -492
rect 1467 -506 1563 -472
rect 1597 -506 1620 -472
rect 513 -509 1620 -506
rect 513 -526 536 -509
rect 456 -549 536 -526
rect 1410 -529 1490 -509
rect 1540 -529 1620 -509
rect 2800 -472 2880 -449
rect 2800 -506 2823 -472
rect 2857 -506 2880 -472
rect 2800 -529 2880 -506
rect 5251 -458 5552 -435
rect 5251 -492 5274 -458
rect 5308 -460 5552 -458
rect 5308 -492 5495 -460
rect 5251 -494 5495 -492
rect 5529 -494 5552 -460
rect 5251 -515 5552 -494
rect 570 -569 650 -549
rect 1290 -569 1370 -549
rect 1670 -569 1750 -549
rect 570 -572 1750 -569
rect 570 -606 593 -572
rect 627 -606 1313 -572
rect 1347 -606 1693 -572
rect 1727 -606 1750 -572
rect 570 -609 1750 -606
rect 570 -629 650 -609
rect 1290 -629 1370 -609
rect 1670 -629 1750 -609
rect 1820 -562 1900 -529
rect 1820 -596 1843 -562
rect 1877 -596 1900 -562
rect 1820 -642 1900 -596
rect 0 -669 80 -649
rect 1540 -669 1620 -649
rect 0 -672 1620 -669
rect 0 -706 23 -672
rect 57 -706 1563 -672
rect 1597 -706 1620 -672
rect 0 -709 1620 -706
rect 0 -729 80 -709
rect 1540 -729 1620 -709
rect 1820 -676 1843 -642
rect 1877 -676 1900 -642
rect 1820 -722 1900 -676
rect 1090 -769 1170 -749
rect 1670 -769 1750 -749
rect 1020 -770 1750 -769
rect 114 -772 1750 -770
rect 114 -793 1113 -772
rect 114 -827 137 -793
rect 171 -806 1113 -793
rect 1147 -806 1693 -772
rect 1727 -806 1750 -772
rect 1820 -756 1843 -722
rect 1877 -756 1900 -722
rect 1820 -779 1900 -756
rect 1970 -562 2050 -529
rect 1970 -596 1993 -562
rect 2027 -596 2050 -562
rect 1970 -642 2050 -596
rect 1970 -676 1993 -642
rect 2027 -676 2050 -642
rect 1970 -722 2050 -676
rect 1970 -756 1993 -722
rect 2027 -756 2050 -722
rect 1970 -789 2050 -756
rect 2120 -562 2200 -529
rect 2120 -596 2143 -562
rect 2177 -596 2200 -562
rect 2120 -642 2200 -596
rect 2120 -676 2143 -642
rect 2177 -676 2200 -642
rect 2120 -722 2200 -676
rect 2120 -756 2143 -722
rect 2177 -756 2200 -722
rect 2120 -779 2200 -756
rect 2270 -562 2350 -529
rect 2270 -596 2293 -562
rect 2327 -596 2350 -562
rect 2270 -642 2350 -596
rect 2270 -676 2293 -642
rect 2327 -676 2350 -642
rect 2270 -722 2350 -676
rect 2270 -756 2293 -722
rect 2327 -756 2350 -722
rect 2270 -789 2350 -756
rect 2420 -562 2500 -529
rect 3572 -537 3652 -515
rect 5472 -517 5552 -515
rect 3299 -538 3652 -537
rect 2420 -596 2443 -562
rect 2477 -596 2500 -562
rect 2420 -642 2500 -596
rect 3000 -572 3080 -549
rect 3000 -606 3023 -572
rect 3057 -606 3080 -572
rect 3000 -629 3080 -606
rect 3299 -572 3595 -538
rect 3629 -572 3652 -538
rect 3299 -577 3652 -572
rect 2420 -676 2443 -642
rect 2477 -676 2500 -642
rect 2420 -722 2500 -676
rect 2420 -756 2443 -722
rect 2477 -756 2500 -722
rect 3150 -672 3230 -649
rect 3150 -706 3173 -672
rect 3207 -706 3230 -672
rect 3150 -729 3230 -706
rect 2420 -779 2500 -756
rect 2700 -772 2780 -749
rect 171 -809 1750 -806
rect 171 -810 1020 -809
rect 171 -827 194 -810
rect 114 -850 194 -827
rect 1090 -829 1170 -809
rect 1670 -829 1750 -809
rect 1990 -839 2030 -789
rect 2170 -839 2250 -819
rect 1990 -842 2250 -839
rect 1990 -876 2193 -842
rect 2227 -876 2250 -842
rect 1990 -879 2250 -876
rect 1990 -1009 2030 -879
rect 2170 -899 2250 -879
rect 1060 -1049 2030 -1009
rect 2070 -959 2150 -944
rect 2290 -959 2330 -789
rect 2700 -806 2723 -772
rect 2757 -806 2780 -772
rect 2700 -829 2780 -806
rect 2540 -852 2620 -829
rect 2540 -886 2563 -852
rect 2597 -869 2620 -852
rect 3299 -869 3339 -577
rect 3572 -595 3652 -577
rect 4010 -562 4090 -529
rect 4010 -596 4033 -562
rect 4067 -596 4090 -562
rect 4010 -642 4090 -596
rect 4010 -676 4033 -642
rect 4067 -676 4090 -642
rect 3860 -719 3940 -699
rect 3660 -722 3940 -719
rect 3660 -756 3883 -722
rect 3917 -756 3940 -722
rect 3660 -759 3940 -756
rect 3860 -779 3940 -759
rect 4010 -722 4090 -676
rect 4010 -756 4033 -722
rect 4067 -756 4090 -722
rect 4010 -779 4090 -756
rect 4160 -562 4240 -529
rect 4160 -596 4183 -562
rect 4217 -596 4240 -562
rect 4160 -642 4240 -596
rect 4160 -676 4183 -642
rect 4217 -676 4240 -642
rect 4160 -722 4240 -676
rect 4160 -756 4183 -722
rect 4217 -756 4240 -722
rect 4160 -789 4240 -756
rect 4310 -562 4390 -529
rect 4310 -596 4333 -562
rect 4367 -596 4390 -562
rect 4310 -642 4390 -596
rect 4310 -676 4333 -642
rect 4367 -676 4390 -642
rect 4310 -722 4390 -676
rect 4310 -756 4333 -722
rect 4367 -756 4390 -722
rect 4310 -779 4390 -756
rect 4460 -562 4540 -529
rect 4460 -596 4483 -562
rect 4517 -596 4540 -562
rect 4460 -642 4540 -596
rect 4460 -676 4483 -642
rect 4517 -676 4540 -642
rect 4460 -722 4540 -676
rect 4460 -756 4483 -722
rect 4517 -756 4540 -722
rect 4460 -789 4540 -756
rect 4610 -562 4690 -529
rect 4610 -596 4633 -562
rect 4667 -596 4690 -562
rect 4610 -642 4690 -596
rect 5310 -569 5390 -549
rect 5740 -569 5820 -549
rect 5310 -572 5820 -569
rect 5310 -606 5333 -572
rect 5367 -606 5763 -572
rect 5797 -606 5820 -572
rect 5310 -609 5820 -606
rect 5310 -629 5390 -609
rect 5740 -629 5820 -609
rect 5890 -562 5970 -529
rect 5890 -596 5913 -562
rect 5947 -596 5970 -562
rect 4610 -676 4633 -642
rect 4667 -676 4690 -642
rect 5890 -642 5970 -596
rect 4610 -722 4690 -676
rect 5162 -689 5551 -684
rect 5740 -689 5820 -669
rect 5162 -692 5820 -689
rect 4610 -756 4633 -722
rect 4667 -756 4690 -722
rect 4610 -779 4690 -756
rect 4760 -719 4840 -699
rect 4890 -719 4970 -699
rect 4760 -722 4970 -719
rect 4760 -756 4783 -722
rect 4817 -756 4913 -722
rect 4947 -756 4970 -722
rect 4760 -759 4970 -756
rect 4760 -779 4840 -759
rect 4890 -779 4970 -759
rect 5162 -724 5763 -692
rect 2597 -886 3339 -869
rect 2540 -909 3339 -886
rect 4180 -839 4220 -789
rect 4360 -839 4440 -819
rect 4180 -842 4440 -839
rect 4180 -876 4383 -842
rect 4417 -876 4440 -842
rect 4180 -879 4440 -876
rect 3300 -959 3380 -943
rect 3730 -959 3810 -939
rect 2070 -966 3380 -959
rect 2070 -967 3323 -966
rect 2070 -1001 2093 -967
rect 2127 -999 3323 -967
rect 2127 -1001 2150 -999
rect 2070 -1024 2150 -1001
rect 1060 -1089 1100 -1049
rect 1660 -1089 1700 -1049
rect 1990 -1089 2030 -1049
rect 2290 -1089 2330 -999
rect 2620 -1089 2660 -999
rect 3220 -1089 3260 -999
rect 3300 -1000 3323 -999
rect 3357 -1000 3380 -966
rect 3300 -1023 3380 -1000
rect 3606 -962 3810 -959
rect 3606 -996 3753 -962
rect 3787 -996 3810 -962
rect 3606 -999 3810 -996
rect 1040 -1122 1120 -1089
rect 1040 -1156 1063 -1122
rect 1097 -1156 1120 -1122
rect 1040 -1202 1120 -1156
rect 1040 -1236 1063 -1202
rect 1097 -1236 1120 -1202
rect 1040 -1282 1120 -1236
rect 1040 -1316 1063 -1282
rect 1097 -1316 1120 -1282
rect 1040 -1339 1120 -1316
rect 1340 -1122 1420 -1089
rect 1340 -1156 1363 -1122
rect 1397 -1156 1420 -1122
rect 1340 -1202 1420 -1156
rect 1340 -1236 1363 -1202
rect 1397 -1236 1420 -1202
rect 1340 -1282 1420 -1236
rect 1340 -1316 1363 -1282
rect 1397 -1316 1420 -1282
rect 1340 -1339 1420 -1316
rect 1640 -1122 1720 -1089
rect 1640 -1156 1663 -1122
rect 1697 -1156 1720 -1122
rect 1640 -1202 1720 -1156
rect 1640 -1236 1663 -1202
rect 1697 -1236 1720 -1202
rect 1640 -1282 1720 -1236
rect 1640 -1316 1663 -1282
rect 1697 -1316 1720 -1282
rect 1640 -1339 1720 -1316
rect 1820 -1122 1900 -1089
rect 1820 -1156 1843 -1122
rect 1877 -1156 1900 -1122
rect 1820 -1202 1900 -1156
rect 1820 -1236 1843 -1202
rect 1877 -1236 1900 -1202
rect 1820 -1282 1900 -1236
rect 1820 -1316 1843 -1282
rect 1877 -1316 1900 -1282
rect 1820 -1339 1900 -1316
rect 1970 -1122 2050 -1089
rect 1970 -1156 1993 -1122
rect 2027 -1156 2050 -1122
rect 1970 -1202 2050 -1156
rect 1970 -1236 1993 -1202
rect 2027 -1236 2050 -1202
rect 1970 -1282 2050 -1236
rect 1970 -1316 1993 -1282
rect 2027 -1316 2050 -1282
rect 1970 -1339 2050 -1316
rect 2120 -1122 2200 -1089
rect 2120 -1156 2143 -1122
rect 2177 -1156 2200 -1122
rect 2120 -1202 2200 -1156
rect 2120 -1236 2143 -1202
rect 2177 -1236 2200 -1202
rect 2120 -1282 2200 -1236
rect 2120 -1316 2143 -1282
rect 2177 -1316 2200 -1282
rect 2120 -1339 2200 -1316
rect 2270 -1122 2350 -1089
rect 2270 -1156 2293 -1122
rect 2327 -1156 2350 -1122
rect 2270 -1202 2350 -1156
rect 2270 -1236 2293 -1202
rect 2327 -1236 2350 -1202
rect 2270 -1282 2350 -1236
rect 2270 -1316 2293 -1282
rect 2327 -1316 2350 -1282
rect 2270 -1339 2350 -1316
rect 2420 -1122 2500 -1089
rect 2420 -1156 2443 -1122
rect 2477 -1156 2500 -1122
rect 2420 -1202 2500 -1156
rect 2420 -1236 2443 -1202
rect 2477 -1236 2500 -1202
rect 2420 -1282 2500 -1236
rect 2420 -1316 2443 -1282
rect 2477 -1316 2500 -1282
rect 2420 -1339 2500 -1316
rect 2600 -1122 2680 -1089
rect 2600 -1156 2623 -1122
rect 2657 -1156 2680 -1122
rect 2600 -1202 2680 -1156
rect 2600 -1236 2623 -1202
rect 2657 -1236 2680 -1202
rect 2600 -1282 2680 -1236
rect 2600 -1316 2623 -1282
rect 2657 -1316 2680 -1282
rect 2600 -1339 2680 -1316
rect 2900 -1122 2980 -1089
rect 2900 -1156 2923 -1122
rect 2957 -1156 2980 -1122
rect 2900 -1202 2980 -1156
rect 2900 -1236 2923 -1202
rect 2957 -1236 2980 -1202
rect 2900 -1282 2980 -1236
rect 2900 -1316 2923 -1282
rect 2957 -1316 2980 -1282
rect 2900 -1339 2980 -1316
rect 3200 -1122 3280 -1089
rect 3200 -1156 3223 -1122
rect 3257 -1156 3280 -1122
rect 3200 -1202 3280 -1156
rect 3200 -1236 3223 -1202
rect 3257 -1236 3280 -1202
rect 3314 -1167 3394 -1148
rect 3606 -1167 3646 -999
rect 3730 -1019 3810 -999
rect 4180 -1009 4220 -879
rect 4360 -899 4440 -879
rect 3850 -1049 4220 -1009
rect 4260 -959 4340 -944
rect 4480 -959 4520 -789
rect 4760 -839 4840 -819
rect 5048 -839 5128 -825
rect 4760 -842 5128 -839
rect 4760 -876 4783 -842
rect 4817 -848 5128 -842
rect 4817 -876 5071 -848
rect 4760 -879 5071 -876
rect 4760 -899 4840 -879
rect 5048 -882 5071 -879
rect 5105 -882 5128 -848
rect 5048 -905 5128 -882
rect 4260 -967 4520 -959
rect 4260 -1001 4283 -967
rect 4317 -999 4520 -967
rect 4317 -1001 4340 -999
rect 4260 -1024 4340 -1001
rect 4480 -1009 4520 -999
rect 5162 -1009 5202 -724
rect 5390 -726 5763 -724
rect 5797 -726 5820 -692
rect 5390 -729 5820 -726
rect 5740 -749 5820 -729
rect 5890 -676 5913 -642
rect 5947 -676 5970 -642
rect 5890 -722 5970 -676
rect 5890 -756 5913 -722
rect 5947 -756 5970 -722
rect 5310 -789 5390 -769
rect 5610 -789 5690 -769
rect 5890 -779 5970 -756
rect 6040 -562 6120 -529
rect 6040 -596 6063 -562
rect 6097 -596 6120 -562
rect 6040 -642 6120 -596
rect 6040 -676 6063 -642
rect 6097 -676 6120 -642
rect 6040 -722 6120 -676
rect 6040 -756 6063 -722
rect 6097 -756 6120 -722
rect 6040 -789 6120 -756
rect 6190 -562 6270 -529
rect 6190 -596 6213 -562
rect 6247 -596 6270 -562
rect 6190 -642 6270 -596
rect 6190 -676 6213 -642
rect 6247 -676 6270 -642
rect 6190 -722 6270 -676
rect 6190 -756 6213 -722
rect 6247 -756 6270 -722
rect 6190 -779 6270 -756
rect 6340 -562 6420 -529
rect 6340 -596 6363 -562
rect 6397 -596 6420 -562
rect 6340 -642 6420 -596
rect 6340 -676 6363 -642
rect 6397 -676 6420 -642
rect 6340 -722 6420 -676
rect 6340 -756 6363 -722
rect 6397 -756 6420 -722
rect 6340 -789 6420 -756
rect 6490 -562 6570 -529
rect 6490 -596 6513 -562
rect 6547 -596 6570 -562
rect 6490 -642 6570 -596
rect 6870 -572 6950 -549
rect 6870 -606 6893 -572
rect 6927 -606 6950 -572
rect 6870 -629 6950 -606
rect 6490 -676 6513 -642
rect 6547 -676 6570 -642
rect 6490 -722 6570 -676
rect 6490 -756 6513 -722
rect 6547 -756 6570 -722
rect 6720 -692 6800 -669
rect 6720 -726 6743 -692
rect 6777 -726 6800 -692
rect 6720 -749 6800 -726
rect 6490 -779 6570 -756
rect 5310 -792 5690 -789
rect 5310 -826 5333 -792
rect 5367 -826 5633 -792
rect 5667 -826 5690 -792
rect 5310 -829 5690 -826
rect 5310 -849 5390 -829
rect 5610 -849 5690 -829
rect 6060 -839 6100 -789
rect 6240 -839 6320 -819
rect 6060 -842 6320 -839
rect 5460 -889 5540 -869
rect 5310 -892 5540 -889
rect 5310 -912 5483 -892
rect 5310 -946 5333 -912
rect 5367 -926 5483 -912
rect 5517 -926 5540 -892
rect 5367 -929 5540 -926
rect 5367 -946 5390 -929
rect 5310 -969 5390 -946
rect 5460 -949 5540 -929
rect 6060 -876 6263 -842
rect 6297 -876 6320 -842
rect 6060 -879 6320 -876
rect 6060 -1009 6100 -879
rect 6240 -899 6320 -879
rect 4480 -1049 5202 -1009
rect 5430 -1049 6100 -1009
rect 6140 -959 6220 -944
rect 6360 -959 6400 -789
rect 6640 -839 6720 -819
rect 6640 -842 7227 -839
rect 6640 -876 6663 -842
rect 6697 -876 7227 -842
rect 6640 -879 7227 -876
rect 6640 -899 6720 -879
rect 7073 -959 7153 -939
rect 6140 -962 7153 -959
rect 6140 -967 7096 -962
rect 6140 -1001 6163 -967
rect 6197 -996 7096 -967
rect 7130 -996 7153 -962
rect 6197 -999 7153 -996
rect 6197 -1001 6220 -999
rect 6140 -1024 6220 -1001
rect 3850 -1089 3890 -1049
rect 4180 -1089 4220 -1049
rect 3314 -1170 3646 -1167
rect 3314 -1204 3337 -1170
rect 3371 -1204 3646 -1170
rect 3314 -1207 3646 -1204
rect 3680 -1122 3760 -1089
rect 3680 -1156 3703 -1122
rect 3737 -1156 3760 -1122
rect 3680 -1202 3760 -1156
rect 3314 -1228 3394 -1207
rect 3200 -1282 3280 -1236
rect 3200 -1316 3223 -1282
rect 3257 -1316 3280 -1282
rect 3200 -1339 3280 -1316
rect 3680 -1236 3703 -1202
rect 3737 -1236 3760 -1202
rect 3680 -1282 3760 -1236
rect 3680 -1316 3703 -1282
rect 3737 -1316 3760 -1282
rect 3680 -1339 3760 -1316
rect 3830 -1122 3910 -1089
rect 3830 -1156 3853 -1122
rect 3887 -1156 3910 -1122
rect 3830 -1202 3910 -1156
rect 3830 -1236 3853 -1202
rect 3887 -1236 3910 -1202
rect 3830 -1282 3910 -1236
rect 3830 -1316 3853 -1282
rect 3887 -1316 3910 -1282
rect 3830 -1339 3910 -1316
rect 4010 -1122 4090 -1089
rect 4010 -1156 4033 -1122
rect 4067 -1156 4090 -1122
rect 4010 -1202 4090 -1156
rect 4010 -1236 4033 -1202
rect 4067 -1236 4090 -1202
rect 4010 -1282 4090 -1236
rect 4010 -1316 4033 -1282
rect 4067 -1316 4090 -1282
rect 4010 -1339 4090 -1316
rect 4160 -1122 4240 -1089
rect 4160 -1156 4183 -1122
rect 4217 -1156 4240 -1122
rect 4160 -1202 4240 -1156
rect 4160 -1236 4183 -1202
rect 4217 -1236 4240 -1202
rect 4160 -1282 4240 -1236
rect 4160 -1316 4183 -1282
rect 4217 -1316 4240 -1282
rect 4160 -1339 4240 -1316
rect 4310 -1122 4390 -1089
rect 4310 -1156 4333 -1122
rect 4367 -1156 4390 -1122
rect 4310 -1202 4390 -1156
rect 4310 -1236 4333 -1202
rect 4367 -1236 4390 -1202
rect 4310 -1282 4390 -1236
rect 4310 -1316 4333 -1282
rect 4367 -1316 4390 -1282
rect 4310 -1339 4390 -1316
rect 4460 -1122 4540 -1049
rect 4810 -1089 4850 -1049
rect 5430 -1089 5470 -1049
rect 5730 -1089 5770 -1049
rect 6061 -1089 6100 -1049
rect 6360 -1089 6400 -999
rect 6690 -1089 6730 -999
rect 7073 -1019 7153 -999
rect 4460 -1156 4483 -1122
rect 4517 -1156 4540 -1122
rect 4460 -1202 4540 -1156
rect 4460 -1236 4483 -1202
rect 4517 -1236 4540 -1202
rect 4460 -1282 4540 -1236
rect 4460 -1316 4483 -1282
rect 4517 -1316 4540 -1282
rect 4460 -1339 4540 -1316
rect 4610 -1122 4690 -1089
rect 4610 -1156 4633 -1122
rect 4667 -1156 4690 -1122
rect 4610 -1202 4690 -1156
rect 4610 -1236 4633 -1202
rect 4667 -1236 4690 -1202
rect 4610 -1282 4690 -1236
rect 4610 -1316 4633 -1282
rect 4667 -1316 4690 -1282
rect 4610 -1339 4690 -1316
rect 4790 -1122 4870 -1089
rect 4790 -1156 4813 -1122
rect 4847 -1156 4870 -1122
rect 4790 -1202 4870 -1156
rect 4790 -1236 4813 -1202
rect 4847 -1236 4870 -1202
rect 4790 -1282 4870 -1236
rect 4790 -1316 4813 -1282
rect 4847 -1316 4870 -1282
rect 4790 -1339 4870 -1316
rect 4940 -1122 5020 -1089
rect 4940 -1156 4963 -1122
rect 4997 -1156 5020 -1122
rect 4940 -1202 5020 -1156
rect 4940 -1236 4963 -1202
rect 4997 -1236 5020 -1202
rect 4940 -1282 5020 -1236
rect 4940 -1316 4963 -1282
rect 4997 -1316 5020 -1282
rect 4940 -1339 5020 -1316
rect 5410 -1122 5490 -1089
rect 5410 -1156 5433 -1122
rect 5467 -1156 5490 -1122
rect 5410 -1202 5490 -1156
rect 5410 -1236 5433 -1202
rect 5467 -1236 5490 -1202
rect 5410 -1282 5490 -1236
rect 5410 -1316 5433 -1282
rect 5467 -1316 5490 -1282
rect 5410 -1339 5490 -1316
rect 5560 -1122 5640 -1089
rect 5560 -1156 5583 -1122
rect 5617 -1156 5640 -1122
rect 5560 -1202 5640 -1156
rect 5560 -1236 5583 -1202
rect 5617 -1236 5640 -1202
rect 5560 -1282 5640 -1236
rect 5560 -1316 5583 -1282
rect 5617 -1316 5640 -1282
rect 5560 -1339 5640 -1316
rect 5710 -1122 5790 -1089
rect 5710 -1156 5733 -1122
rect 5767 -1156 5790 -1122
rect 5710 -1202 5790 -1156
rect 5710 -1236 5733 -1202
rect 5767 -1236 5790 -1202
rect 5710 -1282 5790 -1236
rect 5710 -1316 5733 -1282
rect 5767 -1316 5790 -1282
rect 5710 -1339 5790 -1316
rect 5890 -1122 5970 -1089
rect 5890 -1156 5913 -1122
rect 5947 -1156 5970 -1122
rect 5890 -1202 5970 -1156
rect 5890 -1236 5913 -1202
rect 5947 -1236 5970 -1202
rect 5890 -1282 5970 -1236
rect 5890 -1316 5913 -1282
rect 5947 -1316 5970 -1282
rect 5890 -1339 5970 -1316
rect 6040 -1122 6120 -1089
rect 6040 -1156 6063 -1122
rect 6097 -1156 6120 -1122
rect 6040 -1202 6120 -1156
rect 6040 -1236 6063 -1202
rect 6097 -1236 6120 -1202
rect 6040 -1282 6120 -1236
rect 6040 -1316 6063 -1282
rect 6097 -1316 6120 -1282
rect 6040 -1339 6120 -1316
rect 6190 -1122 6270 -1089
rect 6190 -1156 6213 -1122
rect 6247 -1156 6270 -1122
rect 6190 -1202 6270 -1156
rect 6190 -1236 6213 -1202
rect 6247 -1236 6270 -1202
rect 6190 -1282 6270 -1236
rect 6190 -1316 6213 -1282
rect 6247 -1316 6270 -1282
rect 6190 -1339 6270 -1316
rect 6340 -1122 6420 -1089
rect 6340 -1156 6363 -1122
rect 6397 -1156 6420 -1122
rect 6340 -1202 6420 -1156
rect 6340 -1236 6363 -1202
rect 6397 -1236 6420 -1202
rect 6340 -1282 6420 -1236
rect 6340 -1316 6363 -1282
rect 6397 -1316 6420 -1282
rect 6340 -1339 6420 -1316
rect 6490 -1122 6570 -1089
rect 6490 -1156 6513 -1122
rect 6547 -1156 6570 -1122
rect 6490 -1202 6570 -1156
rect 6490 -1236 6513 -1202
rect 6547 -1236 6570 -1202
rect 6490 -1282 6570 -1236
rect 6490 -1316 6513 -1282
rect 6547 -1316 6570 -1282
rect 6490 -1339 6570 -1316
rect 6670 -1122 6750 -1089
rect 6670 -1156 6693 -1122
rect 6727 -1156 6750 -1122
rect 6670 -1202 6750 -1156
rect 6670 -1236 6693 -1202
rect 6727 -1236 6750 -1202
rect 6670 -1282 6750 -1236
rect 6670 -1316 6693 -1282
rect 6727 -1316 6750 -1282
rect 6670 -1339 6750 -1316
rect 6970 -1122 7050 -1089
rect 6970 -1156 6993 -1122
rect 7027 -1156 7050 -1122
rect 6970 -1202 7050 -1156
rect 6970 -1236 6993 -1202
rect 7027 -1236 7050 -1202
rect 6970 -1282 7050 -1236
rect 6970 -1316 6993 -1282
rect 7027 -1316 7050 -1282
rect 6970 -1339 7050 -1316
rect 1171 -1399 1251 -1379
rect 1920 -1399 2000 -1379
rect 2320 -1399 2400 -1379
rect 4110 -1399 4190 -1379
rect 4510 -1399 4590 -1379
rect 5398 -1399 5478 -1379
rect 5990 -1399 6070 -1379
rect 6390 -1399 6470 -1379
rect 1020 -1402 4590 -1399
rect 1020 -1436 1194 -1402
rect 1228 -1436 1943 -1402
rect 1977 -1436 2343 -1402
rect 2377 -1436 4133 -1402
rect 4167 -1436 4533 -1402
rect 4567 -1436 4590 -1402
rect 1020 -1439 4590 -1436
rect 5390 -1402 6470 -1399
rect 5390 -1436 5421 -1402
rect 5455 -1436 6013 -1402
rect 6047 -1436 6413 -1402
rect 6447 -1436 6470 -1402
rect 5390 -1439 6470 -1436
rect 1171 -1459 1251 -1439
rect 1920 -1459 2000 -1439
rect 2320 -1459 2400 -1439
rect 4110 -1459 4190 -1439
rect 4510 -1459 4590 -1439
rect 5398 -1459 5478 -1439
rect 5990 -1459 6070 -1439
rect 6390 -1459 6470 -1439
rect 912 -1522 3300 -1499
rect 912 -1556 935 -1522
rect 969 -1556 1103 -1522
rect 1137 -1556 1183 -1522
rect 1217 -1556 1263 -1522
rect 1297 -1556 1343 -1522
rect 1377 -1556 1423 -1522
rect 1457 -1556 1503 -1522
rect 1537 -1556 1583 -1522
rect 1617 -1556 1663 -1522
rect 1697 -1556 1743 -1522
rect 1777 -1556 1823 -1522
rect 1857 -1556 1903 -1522
rect 1937 -1556 1983 -1522
rect 2017 -1556 2063 -1522
rect 2097 -1556 2143 -1522
rect 2177 -1556 2223 -1522
rect 2257 -1556 2303 -1522
rect 2337 -1556 2383 -1522
rect 2417 -1556 2463 -1522
rect 2497 -1556 2543 -1522
rect 2577 -1556 2623 -1522
rect 2657 -1556 2703 -1522
rect 2737 -1556 2783 -1522
rect 2817 -1556 2863 -1522
rect 2897 -1556 2943 -1522
rect 2977 -1556 3023 -1522
rect 3057 -1556 3103 -1522
rect 3137 -1556 3183 -1522
rect 3217 -1556 3300 -1522
rect 912 -1579 3300 -1556
rect 3660 -1522 5040 -1499
rect 3660 -1556 3693 -1522
rect 3727 -1556 3773 -1522
rect 3807 -1556 3853 -1522
rect 3887 -1556 3933 -1522
rect 3967 -1556 4013 -1522
rect 4047 -1556 4093 -1522
rect 4127 -1556 4173 -1522
rect 4207 -1556 4253 -1522
rect 4287 -1556 4333 -1522
rect 4367 -1556 4413 -1522
rect 4447 -1556 4493 -1522
rect 4527 -1556 4573 -1522
rect 4607 -1556 4653 -1522
rect 4687 -1556 4733 -1522
rect 4767 -1556 4813 -1522
rect 4847 -1556 4893 -1522
rect 4927 -1556 4973 -1522
rect 5007 -1556 5040 -1522
rect 3660 -1579 5040 -1556
rect 5390 -1522 7070 -1499
rect 5390 -1556 5413 -1522
rect 5447 -1556 5493 -1522
rect 5527 -1556 5573 -1522
rect 5607 -1556 5653 -1522
rect 5687 -1556 5733 -1522
rect 5767 -1556 5813 -1522
rect 5847 -1556 5893 -1522
rect 5927 -1556 5973 -1522
rect 6007 -1556 6053 -1522
rect 6087 -1556 6133 -1522
rect 6167 -1556 6213 -1522
rect 6247 -1556 6293 -1522
rect 6327 -1556 6373 -1522
rect 6407 -1556 6453 -1522
rect 6487 -1556 6533 -1522
rect 6567 -1556 6613 -1522
rect 6647 -1556 6693 -1522
rect 6727 -1556 6773 -1522
rect 6807 -1556 6853 -1522
rect 6887 -1556 6933 -1522
rect 6967 -1556 7013 -1522
rect 7047 -1556 7070 -1522
rect 5390 -1579 7070 -1556
rect 1171 -1639 1251 -1619
rect 1920 -1639 2000 -1619
rect 2320 -1639 2400 -1619
rect 4110 -1639 4190 -1619
rect 4510 -1639 4590 -1619
rect 5398 -1639 5478 -1618
rect 5990 -1639 6070 -1619
rect 6390 -1639 6470 -1619
rect 1020 -1642 4590 -1639
rect 1020 -1676 1194 -1642
rect 1228 -1676 1943 -1642
rect 1977 -1676 2343 -1642
rect 2377 -1676 4133 -1642
rect 4167 -1676 4533 -1642
rect 4567 -1676 4590 -1642
rect 1020 -1679 4590 -1676
rect 5390 -1641 6470 -1639
rect 5390 -1675 5421 -1641
rect 5455 -1642 6470 -1641
rect 5455 -1675 6013 -1642
rect 5390 -1676 6013 -1675
rect 6047 -1676 6413 -1642
rect 6447 -1676 6470 -1642
rect 5390 -1679 6470 -1676
rect 1171 -1699 1251 -1679
rect 1920 -1699 2000 -1679
rect 2320 -1699 2400 -1679
rect 4110 -1699 4190 -1679
rect 4510 -1699 4590 -1679
rect 5398 -1698 5478 -1679
rect 5990 -1699 6070 -1679
rect 6390 -1699 6470 -1679
rect 1040 -1762 1120 -1739
rect 1040 -1796 1063 -1762
rect 1097 -1796 1120 -1762
rect 1040 -1842 1120 -1796
rect 1040 -1876 1063 -1842
rect 1097 -1876 1120 -1842
rect 1040 -1922 1120 -1876
rect 1040 -1956 1063 -1922
rect 1097 -1956 1120 -1922
rect 1040 -1989 1120 -1956
rect 1340 -1762 1420 -1739
rect 1340 -1796 1363 -1762
rect 1397 -1796 1420 -1762
rect 1340 -1842 1420 -1796
rect 1340 -1876 1363 -1842
rect 1397 -1876 1420 -1842
rect 1340 -1922 1420 -1876
rect 1340 -1956 1363 -1922
rect 1397 -1956 1420 -1922
rect 1340 -1989 1420 -1956
rect 1640 -1762 1720 -1739
rect 1640 -1796 1663 -1762
rect 1697 -1796 1720 -1762
rect 1640 -1842 1720 -1796
rect 1640 -1876 1663 -1842
rect 1697 -1876 1720 -1842
rect 1640 -1922 1720 -1876
rect 1640 -1956 1663 -1922
rect 1697 -1956 1720 -1922
rect 1640 -1989 1720 -1956
rect 1820 -1762 1900 -1739
rect 1820 -1796 1843 -1762
rect 1877 -1796 1900 -1762
rect 1820 -1842 1900 -1796
rect 1820 -1876 1843 -1842
rect 1877 -1876 1900 -1842
rect 1820 -1922 1900 -1876
rect 1820 -1956 1843 -1922
rect 1877 -1956 1900 -1922
rect 1820 -1989 1900 -1956
rect 1970 -1762 2050 -1739
rect 1970 -1796 1993 -1762
rect 2027 -1796 2050 -1762
rect 1970 -1842 2050 -1796
rect 1970 -1876 1993 -1842
rect 2027 -1876 2050 -1842
rect 1970 -1922 2050 -1876
rect 1970 -1956 1993 -1922
rect 2027 -1956 2050 -1922
rect 1970 -1989 2050 -1956
rect 2120 -1762 2200 -1739
rect 2120 -1796 2143 -1762
rect 2177 -1796 2200 -1762
rect 2120 -1842 2200 -1796
rect 2120 -1876 2143 -1842
rect 2177 -1876 2200 -1842
rect 2120 -1922 2200 -1876
rect 2120 -1956 2143 -1922
rect 2177 -1956 2200 -1922
rect 2120 -1989 2200 -1956
rect 2270 -1762 2350 -1739
rect 2270 -1796 2293 -1762
rect 2327 -1796 2350 -1762
rect 2270 -1842 2350 -1796
rect 2270 -1876 2293 -1842
rect 2327 -1876 2350 -1842
rect 2270 -1922 2350 -1876
rect 2270 -1956 2293 -1922
rect 2327 -1956 2350 -1922
rect 2270 -1989 2350 -1956
rect 2420 -1762 2500 -1739
rect 2420 -1796 2443 -1762
rect 2477 -1796 2500 -1762
rect 2420 -1842 2500 -1796
rect 2420 -1876 2443 -1842
rect 2477 -1876 2500 -1842
rect 2420 -1922 2500 -1876
rect 2420 -1956 2443 -1922
rect 2477 -1956 2500 -1922
rect 2420 -1989 2500 -1956
rect 2600 -1762 2680 -1739
rect 2600 -1796 2623 -1762
rect 2657 -1796 2680 -1762
rect 2600 -1842 2680 -1796
rect 2600 -1876 2623 -1842
rect 2657 -1876 2680 -1842
rect 2600 -1922 2680 -1876
rect 2600 -1956 2623 -1922
rect 2657 -1956 2680 -1922
rect 2600 -1989 2680 -1956
rect 2900 -1762 2980 -1739
rect 2900 -1796 2923 -1762
rect 2957 -1796 2980 -1762
rect 2900 -1842 2980 -1796
rect 2900 -1876 2923 -1842
rect 2957 -1876 2980 -1842
rect 2900 -1922 2980 -1876
rect 2900 -1956 2923 -1922
rect 2957 -1956 2980 -1922
rect 2900 -1989 2980 -1956
rect 3200 -1762 3280 -1739
rect 3200 -1796 3223 -1762
rect 3257 -1796 3280 -1762
rect 3200 -1842 3280 -1796
rect 3200 -1876 3223 -1842
rect 3257 -1876 3280 -1842
rect 3680 -1762 3760 -1739
rect 3680 -1796 3703 -1762
rect 3737 -1796 3760 -1762
rect 3680 -1842 3760 -1796
rect 3200 -1922 3280 -1876
rect 3200 -1956 3223 -1922
rect 3257 -1956 3280 -1922
rect 3314 -1862 3394 -1843
rect 3314 -1865 3646 -1862
rect 3314 -1899 3337 -1865
rect 3371 -1899 3646 -1865
rect 3314 -1902 3646 -1899
rect 3314 -1923 3394 -1902
rect 3200 -1989 3280 -1956
rect 1060 -2029 1100 -1989
rect 1660 -2029 1700 -1989
rect 1990 -2029 2030 -1989
rect 1060 -2069 2030 -2029
rect 1990 -2199 2030 -2069
rect 2070 -2077 2150 -2054
rect 2070 -2111 2093 -2077
rect 2127 -2079 2150 -2077
rect 2290 -2079 2330 -1989
rect 2620 -2079 2660 -1989
rect 3220 -2079 3260 -1989
rect 3606 -2079 3646 -1902
rect 3680 -1876 3703 -1842
rect 3737 -1876 3760 -1842
rect 3680 -1922 3760 -1876
rect 3680 -1956 3703 -1922
rect 3737 -1956 3760 -1922
rect 3680 -1989 3760 -1956
rect 3830 -1762 3910 -1739
rect 3830 -1796 3853 -1762
rect 3887 -1796 3910 -1762
rect 3830 -1842 3910 -1796
rect 3830 -1876 3853 -1842
rect 3887 -1876 3910 -1842
rect 3830 -1922 3910 -1876
rect 3830 -1956 3853 -1922
rect 3887 -1956 3910 -1922
rect 3830 -1989 3910 -1956
rect 4010 -1762 4090 -1739
rect 4010 -1796 4033 -1762
rect 4067 -1796 4090 -1762
rect 4010 -1842 4090 -1796
rect 4010 -1876 4033 -1842
rect 4067 -1876 4090 -1842
rect 4010 -1922 4090 -1876
rect 4010 -1956 4033 -1922
rect 4067 -1956 4090 -1922
rect 4010 -1989 4090 -1956
rect 4160 -1762 4240 -1739
rect 4160 -1796 4183 -1762
rect 4217 -1796 4240 -1762
rect 4160 -1842 4240 -1796
rect 4160 -1876 4183 -1842
rect 4217 -1876 4240 -1842
rect 4160 -1922 4240 -1876
rect 4160 -1956 4183 -1922
rect 4217 -1956 4240 -1922
rect 4160 -1989 4240 -1956
rect 4310 -1762 4390 -1739
rect 4310 -1796 4333 -1762
rect 4367 -1796 4390 -1762
rect 4310 -1842 4390 -1796
rect 4310 -1876 4333 -1842
rect 4367 -1876 4390 -1842
rect 4310 -1922 4390 -1876
rect 4310 -1956 4333 -1922
rect 4367 -1956 4390 -1922
rect 4310 -1989 4390 -1956
rect 4460 -1762 4540 -1739
rect 4460 -1796 4483 -1762
rect 4517 -1796 4540 -1762
rect 4460 -1842 4540 -1796
rect 4460 -1876 4483 -1842
rect 4517 -1876 4540 -1842
rect 4460 -1922 4540 -1876
rect 4460 -1956 4483 -1922
rect 4517 -1956 4540 -1922
rect 3850 -2029 3890 -1989
rect 4180 -2029 4220 -1989
rect 4460 -2029 4540 -1956
rect 4610 -1762 4690 -1739
rect 4610 -1796 4633 -1762
rect 4667 -1796 4690 -1762
rect 4610 -1842 4690 -1796
rect 4610 -1876 4633 -1842
rect 4667 -1876 4690 -1842
rect 4610 -1922 4690 -1876
rect 4610 -1956 4633 -1922
rect 4667 -1956 4690 -1922
rect 4610 -1989 4690 -1956
rect 4790 -1762 4870 -1739
rect 4790 -1796 4813 -1762
rect 4847 -1796 4870 -1762
rect 4790 -1842 4870 -1796
rect 4790 -1876 4813 -1842
rect 4847 -1876 4870 -1842
rect 4790 -1922 4870 -1876
rect 4790 -1956 4813 -1922
rect 4847 -1956 4870 -1922
rect 4790 -1989 4870 -1956
rect 4940 -1762 5020 -1739
rect 4940 -1796 4963 -1762
rect 4997 -1796 5020 -1762
rect 4940 -1842 5020 -1796
rect 4940 -1876 4963 -1842
rect 4997 -1876 5020 -1842
rect 4940 -1922 5020 -1876
rect 4940 -1956 4963 -1922
rect 4997 -1956 5020 -1922
rect 4940 -1989 5020 -1956
rect 5410 -1762 5490 -1739
rect 5410 -1796 5433 -1762
rect 5467 -1796 5490 -1762
rect 5410 -1842 5490 -1796
rect 5410 -1876 5433 -1842
rect 5467 -1876 5490 -1842
rect 5410 -1922 5490 -1876
rect 5410 -1956 5433 -1922
rect 5467 -1956 5490 -1922
rect 5410 -1989 5490 -1956
rect 5560 -1762 5640 -1739
rect 5560 -1796 5583 -1762
rect 5617 -1796 5640 -1762
rect 5560 -1842 5640 -1796
rect 5560 -1876 5583 -1842
rect 5617 -1876 5640 -1842
rect 5560 -1922 5640 -1876
rect 5560 -1956 5583 -1922
rect 5617 -1956 5640 -1922
rect 5560 -1989 5640 -1956
rect 5710 -1762 5790 -1739
rect 5710 -1796 5733 -1762
rect 5767 -1796 5790 -1762
rect 5710 -1842 5790 -1796
rect 5710 -1876 5733 -1842
rect 5767 -1876 5790 -1842
rect 5710 -1922 5790 -1876
rect 5710 -1956 5733 -1922
rect 5767 -1956 5790 -1922
rect 5710 -1989 5790 -1956
rect 5890 -1762 5970 -1739
rect 5890 -1796 5913 -1762
rect 5947 -1796 5970 -1762
rect 5890 -1842 5970 -1796
rect 5890 -1876 5913 -1842
rect 5947 -1876 5970 -1842
rect 5890 -1922 5970 -1876
rect 5890 -1956 5913 -1922
rect 5947 -1956 5970 -1922
rect 5890 -1989 5970 -1956
rect 6040 -1762 6120 -1739
rect 6040 -1796 6063 -1762
rect 6097 -1796 6120 -1762
rect 6040 -1842 6120 -1796
rect 6040 -1876 6063 -1842
rect 6097 -1876 6120 -1842
rect 6040 -1922 6120 -1876
rect 6040 -1956 6063 -1922
rect 6097 -1956 6120 -1922
rect 6040 -1989 6120 -1956
rect 6190 -1762 6270 -1739
rect 6190 -1796 6213 -1762
rect 6247 -1796 6270 -1762
rect 6190 -1842 6270 -1796
rect 6190 -1876 6213 -1842
rect 6247 -1876 6270 -1842
rect 6190 -1922 6270 -1876
rect 6190 -1956 6213 -1922
rect 6247 -1956 6270 -1922
rect 6190 -1989 6270 -1956
rect 6340 -1762 6420 -1739
rect 6340 -1796 6363 -1762
rect 6397 -1796 6420 -1762
rect 6340 -1842 6420 -1796
rect 6340 -1876 6363 -1842
rect 6397 -1876 6420 -1842
rect 6340 -1922 6420 -1876
rect 6340 -1956 6363 -1922
rect 6397 -1956 6420 -1922
rect 6340 -1989 6420 -1956
rect 6490 -1762 6570 -1739
rect 6490 -1796 6513 -1762
rect 6547 -1796 6570 -1762
rect 6490 -1842 6570 -1796
rect 6490 -1876 6513 -1842
rect 6547 -1876 6570 -1842
rect 6490 -1922 6570 -1876
rect 6490 -1956 6513 -1922
rect 6547 -1956 6570 -1922
rect 6490 -1989 6570 -1956
rect 6670 -1762 6750 -1739
rect 6670 -1796 6693 -1762
rect 6727 -1796 6750 -1762
rect 6670 -1842 6750 -1796
rect 6670 -1876 6693 -1842
rect 6727 -1876 6750 -1842
rect 6670 -1922 6750 -1876
rect 6670 -1956 6693 -1922
rect 6727 -1956 6750 -1922
rect 6670 -1989 6750 -1956
rect 6970 -1762 7050 -1739
rect 6970 -1796 6993 -1762
rect 7027 -1796 7050 -1762
rect 6970 -1842 7050 -1796
rect 6970 -1876 6993 -1842
rect 7027 -1876 7050 -1842
rect 6970 -1922 7050 -1876
rect 6970 -1956 6993 -1922
rect 7027 -1956 7050 -1922
rect 6970 -1989 7050 -1956
rect 4810 -2029 4850 -1989
rect 5430 -2029 5470 -1989
rect 5730 -2029 5770 -1989
rect 6061 -2029 6100 -1989
rect 3730 -2079 3810 -2059
rect 3850 -2069 4220 -2029
rect 2127 -2111 3505 -2079
rect 2070 -2119 3505 -2111
rect 3606 -2082 3810 -2079
rect 3606 -2116 3753 -2082
rect 3787 -2116 3810 -2082
rect 3606 -2119 3810 -2116
rect 2070 -2134 2150 -2119
rect 2170 -2199 2250 -2179
rect 1990 -2202 2250 -2199
rect 798 -2252 878 -2229
rect 1990 -2236 2193 -2202
rect 2227 -2236 2250 -2202
rect 1990 -2239 2250 -2236
rect 798 -2286 821 -2252
rect 855 -2269 878 -2252
rect 1090 -2269 1170 -2249
rect 1670 -2269 1750 -2249
rect 855 -2272 1750 -2269
rect 855 -2286 1113 -2272
rect 798 -2306 1113 -2286
rect 1147 -2306 1693 -2272
rect 1727 -2306 1750 -2272
rect 1990 -2289 2030 -2239
rect 2170 -2259 2250 -2239
rect 2290 -2289 2330 -2119
rect 2540 -2192 3380 -2169
rect 2540 -2226 2563 -2192
rect 2597 -2209 3323 -2192
rect 2597 -2226 2620 -2209
rect 2540 -2249 2620 -2226
rect 3300 -2226 3323 -2209
rect 3357 -2226 3380 -2192
rect 3300 -2249 3380 -2226
rect 2700 -2272 2780 -2249
rect 798 -2309 1750 -2306
rect 1090 -2329 1170 -2309
rect 1670 -2329 1750 -2309
rect 1820 -2322 1900 -2299
rect 684 -2352 764 -2329
rect 684 -2386 707 -2352
rect 741 -2369 764 -2352
rect 1540 -2369 1620 -2349
rect 741 -2372 1620 -2369
rect 741 -2386 1563 -2372
rect 684 -2406 1563 -2386
rect 1597 -2406 1620 -2372
rect 684 -2409 1620 -2406
rect 1540 -2429 1620 -2409
rect 1820 -2356 1843 -2322
rect 1877 -2356 1900 -2322
rect 1820 -2402 1900 -2356
rect 1820 -2436 1843 -2402
rect 1877 -2436 1900 -2402
rect 342 -2469 422 -2449
rect 1290 -2469 1370 -2449
rect 1670 -2469 1750 -2449
rect 342 -2472 1750 -2469
rect 342 -2506 365 -2472
rect 399 -2506 1313 -2472
rect 1347 -2506 1693 -2472
rect 1727 -2506 1750 -2472
rect 342 -2509 1750 -2506
rect 342 -2529 422 -2509
rect 1290 -2529 1370 -2509
rect 1670 -2529 1750 -2509
rect 1820 -2482 1900 -2436
rect 1820 -2516 1843 -2482
rect 1877 -2516 1900 -2482
rect 1820 -2549 1900 -2516
rect 1970 -2322 2050 -2289
rect 1970 -2356 1993 -2322
rect 2027 -2356 2050 -2322
rect 1970 -2402 2050 -2356
rect 1970 -2436 1993 -2402
rect 2027 -2436 2050 -2402
rect 1970 -2482 2050 -2436
rect 1970 -2516 1993 -2482
rect 2027 -2516 2050 -2482
rect 1970 -2549 2050 -2516
rect 2120 -2322 2200 -2299
rect 2120 -2356 2143 -2322
rect 2177 -2356 2200 -2322
rect 2120 -2402 2200 -2356
rect 2120 -2436 2143 -2402
rect 2177 -2436 2200 -2402
rect 2120 -2482 2200 -2436
rect 2120 -2516 2143 -2482
rect 2177 -2516 2200 -2482
rect 2120 -2549 2200 -2516
rect 2270 -2322 2350 -2289
rect 2270 -2356 2293 -2322
rect 2327 -2356 2350 -2322
rect 2270 -2402 2350 -2356
rect 2270 -2436 2293 -2402
rect 2327 -2436 2350 -2402
rect 2270 -2482 2350 -2436
rect 2270 -2516 2293 -2482
rect 2327 -2516 2350 -2482
rect 2270 -2549 2350 -2516
rect 2420 -2322 2500 -2299
rect 2420 -2356 2443 -2322
rect 2477 -2356 2500 -2322
rect 2700 -2306 2723 -2272
rect 2757 -2306 2780 -2272
rect 2700 -2329 2780 -2306
rect 2420 -2402 2500 -2356
rect 2420 -2436 2443 -2402
rect 2477 -2436 2500 -2402
rect 3150 -2372 3230 -2349
rect 3150 -2406 3173 -2372
rect 3207 -2406 3230 -2372
rect 3150 -2429 3230 -2406
rect 2420 -2482 2500 -2436
rect 2420 -2516 2443 -2482
rect 2477 -2516 2500 -2482
rect 2420 -2549 2500 -2516
rect 3000 -2472 3080 -2449
rect 3000 -2506 3023 -2472
rect 3057 -2506 3080 -2472
rect 3000 -2529 3080 -2506
rect 3465 -2501 3505 -2119
rect 3730 -2139 3810 -2119
rect 4180 -2199 4220 -2069
rect 4260 -2077 4340 -2054
rect 4260 -2111 4283 -2077
rect 4317 -2079 4340 -2077
rect 4480 -2069 5370 -2029
rect 5430 -2069 6100 -2029
rect 4480 -2079 4520 -2069
rect 4317 -2111 4520 -2079
rect 4260 -2119 4520 -2111
rect 4260 -2134 4340 -2119
rect 4360 -2199 4440 -2179
rect 4180 -2202 4440 -2199
rect 4180 -2236 4383 -2202
rect 4417 -2236 4440 -2202
rect 4180 -2239 4440 -2236
rect 4180 -2289 4220 -2239
rect 4360 -2259 4440 -2239
rect 4480 -2289 4520 -2119
rect 5330 -2149 5370 -2069
rect 5460 -2149 5540 -2129
rect 5330 -2152 5540 -2149
rect 4760 -2199 4840 -2179
rect 5330 -2186 5483 -2152
rect 5517 -2186 5540 -2152
rect 5330 -2189 5540 -2186
rect 4760 -2202 5235 -2199
rect 4760 -2236 4783 -2202
rect 4817 -2236 5235 -2202
rect 5460 -2209 5540 -2189
rect 6060 -2199 6100 -2069
rect 6140 -2077 6220 -2054
rect 6140 -2111 6163 -2077
rect 6197 -2079 6220 -2077
rect 6360 -2079 6400 -1989
rect 6690 -2079 6730 -1989
rect 7073 -2079 7153 -2059
rect 6197 -2082 7153 -2079
rect 6197 -2111 7096 -2082
rect 6140 -2116 7096 -2111
rect 7130 -2116 7153 -2082
rect 6140 -2119 7153 -2116
rect 6140 -2134 6220 -2119
rect 6240 -2199 6320 -2179
rect 6060 -2202 6320 -2199
rect 4760 -2239 5235 -2236
rect 4760 -2259 4840 -2239
rect 3860 -2319 3940 -2299
rect 3660 -2322 3940 -2319
rect 3660 -2356 3883 -2322
rect 3917 -2356 3940 -2322
rect 3660 -2359 3940 -2356
rect 3860 -2379 3940 -2359
rect 4010 -2322 4090 -2299
rect 4010 -2356 4033 -2322
rect 4067 -2356 4090 -2322
rect 4010 -2402 4090 -2356
rect 4010 -2436 4033 -2402
rect 4067 -2436 4090 -2402
rect 4010 -2482 4090 -2436
rect 3572 -2501 3652 -2483
rect 3465 -2506 3652 -2501
rect 3465 -2540 3595 -2506
rect 3629 -2540 3652 -2506
rect 3465 -2541 3652 -2540
rect 1410 -2569 1490 -2549
rect 1540 -2569 1620 -2549
rect 228 -2572 1620 -2569
rect 228 -2592 1433 -2572
rect 228 -2626 251 -2592
rect 285 -2606 1433 -2592
rect 1467 -2606 1563 -2572
rect 1597 -2606 1620 -2572
rect 285 -2609 1620 -2606
rect 285 -2626 308 -2609
rect 228 -2649 308 -2626
rect 1410 -2629 1490 -2609
rect 1540 -2629 1620 -2609
rect 2800 -2572 2880 -2549
rect 3572 -2563 3652 -2541
rect 4010 -2516 4033 -2482
rect 4067 -2516 4090 -2482
rect 4010 -2549 4090 -2516
rect 4160 -2322 4240 -2289
rect 4160 -2356 4183 -2322
rect 4217 -2356 4240 -2322
rect 4160 -2402 4240 -2356
rect 4160 -2436 4183 -2402
rect 4217 -2436 4240 -2402
rect 4160 -2482 4240 -2436
rect 4160 -2516 4183 -2482
rect 4217 -2516 4240 -2482
rect 4160 -2549 4240 -2516
rect 4310 -2322 4390 -2299
rect 4310 -2356 4333 -2322
rect 4367 -2356 4390 -2322
rect 4310 -2402 4390 -2356
rect 4310 -2436 4333 -2402
rect 4367 -2436 4390 -2402
rect 4310 -2482 4390 -2436
rect 4310 -2516 4333 -2482
rect 4367 -2516 4390 -2482
rect 4310 -2549 4390 -2516
rect 4460 -2322 4540 -2289
rect 4460 -2356 4483 -2322
rect 4517 -2356 4540 -2322
rect 4460 -2402 4540 -2356
rect 4460 -2436 4483 -2402
rect 4517 -2436 4540 -2402
rect 4460 -2482 4540 -2436
rect 4460 -2516 4483 -2482
rect 4517 -2516 4540 -2482
rect 4460 -2549 4540 -2516
rect 4610 -2322 4690 -2299
rect 4610 -2356 4633 -2322
rect 4667 -2356 4690 -2322
rect 4610 -2402 4690 -2356
rect 4760 -2319 4840 -2299
rect 4890 -2319 4970 -2299
rect 4760 -2322 4970 -2319
rect 4760 -2356 4783 -2322
rect 4817 -2356 4913 -2322
rect 4947 -2356 4970 -2322
rect 4760 -2359 4970 -2356
rect 4760 -2379 4840 -2359
rect 4890 -2379 4970 -2359
rect 5195 -2349 5235 -2239
rect 5310 -2249 5390 -2229
rect 5610 -2249 5690 -2229
rect 5310 -2252 5690 -2249
rect 5310 -2286 5333 -2252
rect 5367 -2286 5633 -2252
rect 5667 -2286 5690 -2252
rect 5310 -2289 5690 -2286
rect 6060 -2236 6263 -2202
rect 6297 -2236 6320 -2202
rect 6060 -2239 6320 -2236
rect 6060 -2289 6100 -2239
rect 6240 -2259 6320 -2239
rect 6360 -2289 6400 -2119
rect 7073 -2139 7153 -2119
rect 6640 -2199 6720 -2179
rect 6640 -2202 7144 -2199
rect 6640 -2236 6663 -2202
rect 6697 -2236 7144 -2202
rect 6640 -2239 7144 -2236
rect 6640 -2259 6720 -2239
rect 5310 -2309 5390 -2289
rect 5610 -2309 5690 -2289
rect 5890 -2322 5970 -2299
rect 5740 -2349 5820 -2329
rect 5195 -2352 5820 -2349
rect 5195 -2386 5763 -2352
rect 5797 -2386 5820 -2352
rect 5195 -2389 5820 -2386
rect 4610 -2436 4633 -2402
rect 4667 -2436 4690 -2402
rect 5740 -2409 5820 -2389
rect 5890 -2356 5913 -2322
rect 5947 -2356 5970 -2322
rect 5890 -2402 5970 -2356
rect 4610 -2482 4690 -2436
rect 5890 -2436 5913 -2402
rect 5947 -2436 5970 -2402
rect 4610 -2516 4633 -2482
rect 4667 -2516 4690 -2482
rect 4610 -2549 4690 -2516
rect 5310 -2469 5390 -2450
rect 5740 -2469 5820 -2449
rect 5310 -2472 5820 -2469
rect 5310 -2473 5763 -2472
rect 5310 -2507 5333 -2473
rect 5367 -2506 5763 -2473
rect 5797 -2506 5820 -2472
rect 5367 -2507 5820 -2506
rect 5310 -2509 5820 -2507
rect 5310 -2530 5390 -2509
rect 5740 -2529 5820 -2509
rect 5890 -2482 5970 -2436
rect 5890 -2516 5913 -2482
rect 5947 -2516 5970 -2482
rect 5890 -2549 5970 -2516
rect 6040 -2322 6120 -2289
rect 6040 -2356 6063 -2322
rect 6097 -2356 6120 -2322
rect 6040 -2402 6120 -2356
rect 6040 -2436 6063 -2402
rect 6097 -2436 6120 -2402
rect 6040 -2482 6120 -2436
rect 6040 -2516 6063 -2482
rect 6097 -2516 6120 -2482
rect 6040 -2549 6120 -2516
rect 6190 -2322 6270 -2299
rect 6190 -2356 6213 -2322
rect 6247 -2356 6270 -2322
rect 6190 -2402 6270 -2356
rect 6190 -2436 6213 -2402
rect 6247 -2436 6270 -2402
rect 6190 -2482 6270 -2436
rect 6190 -2516 6213 -2482
rect 6247 -2516 6270 -2482
rect 6190 -2549 6270 -2516
rect 6340 -2322 6420 -2289
rect 6340 -2356 6363 -2322
rect 6397 -2356 6420 -2322
rect 6340 -2402 6420 -2356
rect 6340 -2436 6363 -2402
rect 6397 -2436 6420 -2402
rect 6340 -2482 6420 -2436
rect 6340 -2516 6363 -2482
rect 6397 -2516 6420 -2482
rect 6340 -2549 6420 -2516
rect 6490 -2322 6570 -2299
rect 6490 -2356 6513 -2322
rect 6547 -2356 6570 -2322
rect 6490 -2402 6570 -2356
rect 6490 -2436 6513 -2402
rect 6547 -2436 6570 -2402
rect 6720 -2352 6800 -2329
rect 6720 -2386 6743 -2352
rect 6777 -2386 6800 -2352
rect 6720 -2409 6800 -2386
rect 6490 -2482 6570 -2436
rect 6490 -2516 6513 -2482
rect 6547 -2516 6570 -2482
rect 6490 -2549 6570 -2516
rect 6870 -2472 6950 -2449
rect 6870 -2506 6893 -2472
rect 6927 -2506 6950 -2472
rect 6870 -2529 6950 -2506
rect 2800 -2606 2823 -2572
rect 2857 -2606 2880 -2572
rect 2800 -2629 2880 -2606
rect 1020 -2702 3300 -2679
rect 1020 -2736 1103 -2702
rect 1137 -2736 1183 -2702
rect 1217 -2736 1263 -2702
rect 1297 -2736 1343 -2702
rect 1377 -2736 1423 -2702
rect 1457 -2736 1503 -2702
rect 1537 -2736 1583 -2702
rect 1617 -2736 1663 -2702
rect 1697 -2736 1743 -2702
rect 1777 -2736 1823 -2702
rect 1857 -2736 1903 -2702
rect 1937 -2736 1983 -2702
rect 2017 -2736 2063 -2702
rect 2097 -2736 2143 -2702
rect 2177 -2736 2223 -2702
rect 2257 -2736 2303 -2702
rect 2337 -2736 2383 -2702
rect 2417 -2736 2463 -2702
rect 2497 -2736 2543 -2702
rect 2577 -2736 2623 -2702
rect 2657 -2736 2703 -2702
rect 2737 -2736 2783 -2702
rect 2817 -2736 2863 -2702
rect 2897 -2736 2943 -2702
rect 2977 -2736 3023 -2702
rect 3057 -2736 3103 -2702
rect 3137 -2736 3183 -2702
rect 3217 -2736 3300 -2702
rect 1020 -2759 3300 -2736
rect 3660 -2702 5040 -2679
rect 3660 -2736 3693 -2702
rect 3727 -2736 3773 -2702
rect 3807 -2736 3853 -2702
rect 3887 -2736 3933 -2702
rect 3967 -2736 4013 -2702
rect 4047 -2736 4093 -2702
rect 4127 -2736 4173 -2702
rect 4207 -2736 4253 -2702
rect 4287 -2736 4333 -2702
rect 4367 -2736 4413 -2702
rect 4447 -2736 4493 -2702
rect 4527 -2736 4573 -2702
rect 4607 -2736 4653 -2702
rect 4687 -2736 4733 -2702
rect 4767 -2736 4813 -2702
rect 4847 -2736 4893 -2702
rect 4927 -2736 4973 -2702
rect 5007 -2736 5040 -2702
rect 3660 -2759 5040 -2736
rect 5390 -2702 7070 -2679
rect 5390 -2736 5413 -2702
rect 5447 -2736 5493 -2702
rect 5527 -2736 5573 -2702
rect 5607 -2736 5653 -2702
rect 5687 -2736 5733 -2702
rect 5767 -2736 5813 -2702
rect 5847 -2736 5893 -2702
rect 5927 -2736 5973 -2702
rect 6007 -2736 6053 -2702
rect 6087 -2736 6133 -2702
rect 6167 -2736 6213 -2702
rect 6247 -2736 6293 -2702
rect 6327 -2736 6373 -2702
rect 6407 -2736 6453 -2702
rect 6487 -2736 6533 -2702
rect 6567 -2736 6613 -2702
rect 6647 -2736 6693 -2702
rect 6727 -2736 6773 -2702
rect 6807 -2736 6853 -2702
rect 6887 -2736 6933 -2702
rect 6967 -2736 7013 -2702
rect 7047 -2736 7070 -2702
rect 5390 -2759 7070 -2736
rect 5398 -2933 5478 -2913
rect 5024 -2936 5478 -2933
rect 5024 -2970 5421 -2936
rect 5455 -2970 5478 -2936
rect 5024 -2973 5478 -2970
rect 1161 -3162 3161 -3139
rect 1161 -3196 1184 -3162
rect 1218 -3196 1264 -3162
rect 1298 -3196 1344 -3162
rect 1378 -3196 1424 -3162
rect 1458 -3196 1504 -3162
rect 1538 -3196 1584 -3162
rect 1618 -3196 1664 -3162
rect 1698 -3196 1744 -3162
rect 1778 -3196 1824 -3162
rect 1858 -3196 1904 -3162
rect 1938 -3196 1984 -3162
rect 2018 -3196 2064 -3162
rect 2098 -3196 2144 -3162
rect 2178 -3196 2224 -3162
rect 2258 -3196 2304 -3162
rect 2338 -3196 2384 -3162
rect 2418 -3196 2464 -3162
rect 2498 -3196 2544 -3162
rect 2578 -3196 2624 -3162
rect 2658 -3196 2704 -3162
rect 2738 -3196 2784 -3162
rect 2818 -3196 2864 -3162
rect 2898 -3196 2944 -3162
rect 2978 -3196 3024 -3162
rect 3058 -3196 3104 -3162
rect 3138 -3196 3161 -3162
rect 1161 -3219 3161 -3196
rect 3521 -3162 4901 -3139
rect 3521 -3196 3554 -3162
rect 3588 -3196 3634 -3162
rect 3668 -3196 3714 -3162
rect 3748 -3196 3794 -3162
rect 3828 -3196 3874 -3162
rect 3908 -3196 3954 -3162
rect 3988 -3196 4034 -3162
rect 4068 -3196 4114 -3162
rect 4148 -3196 4194 -3162
rect 4228 -3196 4274 -3162
rect 4308 -3196 4354 -3162
rect 4388 -3196 4434 -3162
rect 4468 -3196 4514 -3162
rect 4548 -3196 4594 -3162
rect 4628 -3196 4674 -3162
rect 4708 -3196 4754 -3162
rect 4788 -3196 4834 -3162
rect 4868 -3196 4901 -3162
rect 3521 -3219 4901 -3196
rect 798 -3262 878 -3239
rect 798 -3296 821 -3262
rect 855 -3279 878 -3262
rect 1581 -3279 1661 -3259
rect 855 -3282 1661 -3279
rect 855 -3296 1604 -3282
rect 798 -3316 1604 -3296
rect 1638 -3316 1661 -3282
rect 798 -3319 1661 -3316
rect 1581 -3339 1661 -3319
rect 2951 -3282 3031 -3259
rect 2951 -3316 2974 -3282
rect 3008 -3316 3031 -3282
rect 2951 -3339 3031 -3316
rect 5024 -3346 5064 -2973
rect 5398 -2993 5478 -2973
rect 7104 -3060 7144 -2239
rect 7187 -2967 7227 -879
rect 7343 -2967 7423 -2946
rect 7187 -2969 7423 -2967
rect 7187 -3003 7366 -2969
rect 7400 -3003 7423 -2969
rect 7187 -3007 7423 -3003
rect 7343 -3026 7423 -3007
rect 7104 -3100 7429 -3060
rect 5251 -3163 7251 -3140
rect 5251 -3197 5274 -3163
rect 5308 -3197 5354 -3163
rect 5388 -3197 5434 -3163
rect 5468 -3197 5514 -3163
rect 5548 -3197 5594 -3163
rect 5628 -3197 5674 -3163
rect 5708 -3197 5754 -3163
rect 5788 -3197 5834 -3163
rect 5868 -3197 5914 -3163
rect 5948 -3197 5994 -3163
rect 6028 -3197 6074 -3163
rect 6108 -3197 6154 -3163
rect 6188 -3197 6234 -3163
rect 6268 -3197 6314 -3163
rect 6348 -3197 6394 -3163
rect 6428 -3197 6474 -3163
rect 6508 -3197 6554 -3163
rect 6588 -3197 6634 -3163
rect 6668 -3197 6714 -3163
rect 6748 -3197 6794 -3163
rect 6828 -3197 6874 -3163
rect 6908 -3197 6954 -3163
rect 6988 -3197 7034 -3163
rect 7068 -3197 7114 -3163
rect 7148 -3197 7194 -3163
rect 7228 -3197 7251 -3163
rect 5251 -3220 7251 -3197
rect 5381 -3288 5461 -3265
rect 5381 -3322 5404 -3288
rect 5438 -3322 5461 -3288
rect 5381 -3345 5461 -3322
rect 6661 -3290 6741 -3270
rect 7229 -3290 7309 -3270
rect 6661 -3293 7309 -3290
rect 6661 -3327 6684 -3293
rect 6718 -3327 7252 -3293
rect 7286 -3327 7309 -3293
rect 6661 -3330 7309 -3327
rect 228 -3382 308 -3359
rect 228 -3416 251 -3382
rect 285 -3399 308 -3382
rect 1671 -3399 1751 -3379
rect 285 -3402 1751 -3399
rect 285 -3416 1694 -3402
rect 228 -3436 1694 -3416
rect 1728 -3436 1751 -3402
rect 228 -3439 1751 -3436
rect 1671 -3459 1751 -3439
rect 1821 -3382 1901 -3349
rect 1821 -3416 1844 -3382
rect 1878 -3416 1901 -3382
rect 1821 -3462 1901 -3416
rect 114 -3481 194 -3462
rect 114 -3485 838 -3481
rect 114 -3519 137 -3485
rect 171 -3509 838 -3485
rect 1821 -3496 1844 -3462
rect 1878 -3496 1901 -3462
rect 1641 -3509 1721 -3499
rect 171 -3519 1721 -3509
rect 114 -3521 1721 -3519
rect 114 -3542 194 -3521
rect 798 -3522 1721 -3521
rect 798 -3549 1664 -3522
rect 684 -3578 764 -3555
rect 684 -3612 707 -3578
rect 741 -3589 764 -3578
rect 1641 -3556 1664 -3549
rect 1698 -3556 1721 -3522
rect 1641 -3579 1721 -3556
rect 1821 -3542 1901 -3496
rect 1821 -3576 1844 -3542
rect 1878 -3576 1901 -3542
rect 741 -3612 1601 -3589
rect 1821 -3599 1901 -3576
rect 1971 -3382 2051 -3349
rect 1971 -3416 1994 -3382
rect 2028 -3416 2051 -3382
rect 1971 -3462 2051 -3416
rect 1971 -3496 1994 -3462
rect 2028 -3496 2051 -3462
rect 1971 -3542 2051 -3496
rect 1971 -3576 1994 -3542
rect 2028 -3576 2051 -3542
rect 1971 -3609 2051 -3576
rect 2121 -3382 2201 -3349
rect 2121 -3416 2144 -3382
rect 2178 -3416 2201 -3382
rect 2121 -3462 2201 -3416
rect 2121 -3496 2144 -3462
rect 2178 -3496 2201 -3462
rect 2121 -3542 2201 -3496
rect 2121 -3576 2144 -3542
rect 2178 -3576 2201 -3542
rect 2121 -3599 2201 -3576
rect 2271 -3382 2351 -3349
rect 2271 -3416 2294 -3382
rect 2328 -3416 2351 -3382
rect 2271 -3462 2351 -3416
rect 2271 -3496 2294 -3462
rect 2328 -3496 2351 -3462
rect 2271 -3542 2351 -3496
rect 2271 -3576 2294 -3542
rect 2328 -3576 2351 -3542
rect 2271 -3609 2351 -3576
rect 2421 -3382 2501 -3349
rect 2421 -3416 2444 -3382
rect 2478 -3416 2501 -3382
rect 2421 -3462 2501 -3416
rect 2801 -3402 2881 -3379
rect 2801 -3436 2824 -3402
rect 2858 -3436 2881 -3402
rect 2801 -3459 2881 -3436
rect 3871 -3382 3951 -3349
rect 3871 -3416 3894 -3382
rect 3928 -3416 3951 -3382
rect 2421 -3496 2444 -3462
rect 2478 -3496 2501 -3462
rect 2421 -3542 2501 -3496
rect 3871 -3462 3951 -3416
rect 3871 -3496 3894 -3462
rect 3928 -3496 3951 -3462
rect 2421 -3576 2444 -3542
rect 2478 -3576 2501 -3542
rect 2421 -3599 2501 -3576
rect 2671 -3522 2751 -3499
rect 2671 -3556 2694 -3522
rect 2728 -3556 2751 -3522
rect 2671 -3579 2751 -3556
rect 3433 -3539 3513 -3519
rect 3721 -3539 3801 -3519
rect 3433 -3542 3801 -3539
rect 3433 -3576 3456 -3542
rect 3490 -3576 3744 -3542
rect 3778 -3576 3801 -3542
rect 3433 -3579 3801 -3576
rect 3433 -3599 3513 -3579
rect 3721 -3599 3801 -3579
rect 3871 -3542 3951 -3496
rect 3871 -3576 3894 -3542
rect 3928 -3576 3951 -3542
rect 3871 -3599 3951 -3576
rect 4021 -3382 4101 -3349
rect 4021 -3416 4044 -3382
rect 4078 -3416 4101 -3382
rect 4021 -3462 4101 -3416
rect 4021 -3496 4044 -3462
rect 4078 -3496 4101 -3462
rect 4021 -3542 4101 -3496
rect 4021 -3576 4044 -3542
rect 4078 -3576 4101 -3542
rect 4021 -3609 4101 -3576
rect 4171 -3382 4251 -3349
rect 4171 -3416 4194 -3382
rect 4228 -3416 4251 -3382
rect 4171 -3462 4251 -3416
rect 4171 -3496 4194 -3462
rect 4228 -3496 4251 -3462
rect 4171 -3542 4251 -3496
rect 4171 -3576 4194 -3542
rect 4228 -3576 4251 -3542
rect 4171 -3599 4251 -3576
rect 4321 -3382 4401 -3349
rect 4321 -3416 4344 -3382
rect 4378 -3416 4401 -3382
rect 4321 -3462 4401 -3416
rect 4321 -3496 4344 -3462
rect 4378 -3496 4401 -3462
rect 4321 -3542 4401 -3496
rect 4321 -3576 4344 -3542
rect 4378 -3576 4401 -3542
rect 4321 -3609 4401 -3576
rect 4471 -3382 4551 -3349
rect 4471 -3416 4494 -3382
rect 4528 -3416 4551 -3382
rect 4471 -3462 4551 -3416
rect 5004 -3369 5084 -3346
rect 6661 -3350 6741 -3330
rect 7229 -3350 7309 -3330
rect 5004 -3403 5027 -3369
rect 5061 -3403 5084 -3369
rect 5911 -3383 5991 -3350
rect 5004 -3426 5084 -3403
rect 5481 -3413 5561 -3390
rect 4471 -3496 4494 -3462
rect 4528 -3496 4551 -3462
rect 5481 -3447 5504 -3413
rect 5538 -3447 5561 -3413
rect 5481 -3470 5561 -3447
rect 5911 -3417 5934 -3383
rect 5968 -3417 5991 -3383
rect 5911 -3463 5991 -3417
rect 4471 -3542 4551 -3496
rect 5681 -3503 5761 -3480
rect 4471 -3576 4494 -3542
rect 4528 -3576 4551 -3542
rect 4471 -3599 4551 -3576
rect 4621 -3539 4701 -3519
rect 4751 -3539 4831 -3519
rect 4621 -3542 4831 -3539
rect 5681 -3537 5704 -3503
rect 5738 -3537 5761 -3503
rect 4621 -3576 4644 -3542
rect 4678 -3576 4774 -3542
rect 4808 -3576 4831 -3542
rect 5180 -3562 5260 -3542
rect 5681 -3560 5761 -3537
rect 5911 -3497 5934 -3463
rect 5968 -3497 5991 -3463
rect 5911 -3543 5991 -3497
rect 4621 -3579 4831 -3576
rect 4621 -3599 4701 -3579
rect 4751 -3599 4831 -3579
rect 5066 -3565 5260 -3562
rect 5066 -3599 5203 -3565
rect 5237 -3599 5260 -3565
rect 5066 -3602 5260 -3599
rect 5911 -3577 5934 -3543
rect 5968 -3577 5991 -3543
rect 5911 -3600 5991 -3577
rect 6061 -3383 6141 -3350
rect 6061 -3417 6084 -3383
rect 6118 -3417 6141 -3383
rect 6061 -3463 6141 -3417
rect 6061 -3497 6084 -3463
rect 6118 -3497 6141 -3463
rect 6061 -3543 6141 -3497
rect 6061 -3577 6084 -3543
rect 6118 -3577 6141 -3543
rect 684 -3629 1601 -3612
rect 342 -3652 422 -3629
rect 684 -3635 764 -3629
rect 342 -3686 365 -3652
rect 399 -3669 422 -3652
rect 1541 -3649 1601 -3629
rect 399 -3686 1451 -3669
rect 342 -3692 1451 -3686
rect 342 -3709 1394 -3692
rect 1371 -3726 1394 -3709
rect 1428 -3726 1451 -3692
rect 0 -3752 80 -3729
rect 1371 -3749 1451 -3726
rect 1541 -3672 1621 -3649
rect 1541 -3706 1564 -3672
rect 1598 -3706 1621 -3672
rect 1541 -3729 1621 -3706
rect 1991 -3659 2031 -3609
rect 2171 -3659 2251 -3639
rect 1991 -3662 2251 -3659
rect 1991 -3696 2194 -3662
rect 2228 -3696 2251 -3662
rect 1991 -3699 2251 -3696
rect 0 -3786 23 -3752
rect 57 -3769 80 -3752
rect 1241 -3769 1321 -3749
rect 57 -3772 1321 -3769
rect 57 -3786 1264 -3772
rect 0 -3806 1264 -3786
rect 1298 -3806 1321 -3772
rect 0 -3809 1321 -3806
rect 1241 -3829 1321 -3809
rect 1991 -3829 2031 -3699
rect 2171 -3719 2251 -3699
rect 1361 -3869 2031 -3829
rect 2071 -3779 2151 -3764
rect 2291 -3779 2331 -3609
rect 2571 -3659 2651 -3639
rect 4041 -3659 4081 -3609
rect 4221 -3659 4301 -3639
rect 2571 -3662 3354 -3659
rect 2571 -3696 2594 -3662
rect 2628 -3696 3354 -3662
rect 2571 -3699 3354 -3696
rect 2571 -3719 2651 -3699
rect 3151 -3779 3231 -3758
rect 2071 -3781 3231 -3779
rect 2071 -3787 3174 -3781
rect 2071 -3821 2094 -3787
rect 2128 -3815 3174 -3787
rect 3208 -3815 3231 -3781
rect 2128 -3819 3231 -3815
rect 3314 -3779 3354 -3699
rect 4041 -3662 4301 -3659
rect 4041 -3696 4244 -3662
rect 4278 -3696 4301 -3662
rect 4041 -3699 4301 -3696
rect 3591 -3779 3671 -3759
rect 3314 -3782 3671 -3779
rect 3314 -3816 3614 -3782
rect 3648 -3816 3671 -3782
rect 3314 -3819 3671 -3816
rect 2128 -3821 2151 -3819
rect 2071 -3844 2151 -3821
rect 1361 -3909 1401 -3869
rect 1661 -3909 1701 -3869
rect 1991 -3909 2031 -3869
rect 2291 -3909 2331 -3819
rect 2621 -3909 2661 -3819
rect 3151 -3838 3231 -3819
rect 3591 -3839 3671 -3819
rect 4041 -3829 4081 -3699
rect 4221 -3719 4301 -3699
rect 3711 -3869 4081 -3829
rect 4121 -3779 4201 -3764
rect 4341 -3779 4381 -3609
rect 4621 -3659 4701 -3639
rect 5066 -3659 5106 -3602
rect 5180 -3622 5260 -3602
rect 6061 -3610 6141 -3577
rect 6211 -3383 6291 -3350
rect 6211 -3417 6234 -3383
rect 6268 -3417 6291 -3383
rect 6211 -3463 6291 -3417
rect 6211 -3497 6234 -3463
rect 6268 -3497 6291 -3463
rect 6211 -3543 6291 -3497
rect 6211 -3577 6234 -3543
rect 6268 -3577 6291 -3543
rect 6211 -3600 6291 -3577
rect 6361 -3383 6441 -3350
rect 6361 -3417 6384 -3383
rect 6418 -3417 6441 -3383
rect 6361 -3463 6441 -3417
rect 6361 -3497 6384 -3463
rect 6418 -3497 6441 -3463
rect 6361 -3543 6441 -3497
rect 6361 -3577 6384 -3543
rect 6418 -3577 6441 -3543
rect 6361 -3610 6441 -3577
rect 6511 -3383 6591 -3350
rect 6511 -3417 6534 -3383
rect 6568 -3417 6591 -3383
rect 6511 -3463 6591 -3417
rect 6781 -3400 6861 -3380
rect 7033 -3400 7113 -3380
rect 6781 -3403 7241 -3400
rect 6781 -3437 6804 -3403
rect 6838 -3437 7056 -3403
rect 7090 -3437 7241 -3403
rect 6781 -3440 7241 -3437
rect 6781 -3460 6861 -3440
rect 7033 -3460 7113 -3440
rect 6511 -3497 6534 -3463
rect 6568 -3497 6591 -3463
rect 6511 -3543 6591 -3497
rect 6511 -3577 6534 -3543
rect 6568 -3577 6591 -3543
rect 6661 -3500 6741 -3480
rect 6661 -3503 7241 -3500
rect 6661 -3537 6684 -3503
rect 6718 -3537 7241 -3503
rect 6661 -3540 7241 -3537
rect 6661 -3560 6741 -3540
rect 6511 -3600 6591 -3577
rect 7275 -3590 7355 -3568
rect 7081 -3591 7355 -3590
rect 4621 -3662 5106 -3659
rect 4621 -3696 4644 -3662
rect 4678 -3696 5106 -3662
rect 4621 -3699 5106 -3696
rect 5181 -3660 5261 -3656
rect 5761 -3660 5841 -3640
rect 5181 -3663 5841 -3660
rect 5181 -3679 5784 -3663
rect 4621 -3719 4701 -3699
rect 5181 -3713 5204 -3679
rect 5238 -3697 5784 -3679
rect 5818 -3697 5841 -3663
rect 5238 -3700 5841 -3697
rect 5238 -3713 5261 -3700
rect 5181 -3736 5261 -3713
rect 5761 -3720 5841 -3700
rect 4121 -3787 4381 -3779
rect 4121 -3821 4144 -3787
rect 4178 -3819 4381 -3787
rect 5181 -3780 5261 -3770
rect 6081 -3780 6121 -3610
rect 6161 -3660 6241 -3640
rect 6381 -3660 6421 -3610
rect 6161 -3663 6421 -3660
rect 6161 -3697 6184 -3663
rect 6218 -3697 6421 -3663
rect 7081 -3613 7298 -3591
rect 7081 -3647 7104 -3613
rect 7138 -3625 7298 -3613
rect 7332 -3625 7355 -3591
rect 7138 -3630 7355 -3625
rect 7138 -3647 7161 -3630
rect 7081 -3670 7161 -3647
rect 7275 -3648 7355 -3630
rect 6161 -3700 6421 -3697
rect 6161 -3720 6241 -3700
rect 6261 -3780 6341 -3765
rect 5181 -3788 6341 -3780
rect 5181 -3793 6284 -3788
rect 4178 -3821 4201 -3819
rect 4121 -3844 4201 -3821
rect 4341 -3829 4381 -3819
rect 4915 -3829 4995 -3809
rect 4341 -3832 4995 -3829
rect 4341 -3866 4938 -3832
rect 4972 -3866 4995 -3832
rect 5181 -3827 5204 -3793
rect 5238 -3820 6284 -3793
rect 5238 -3827 5261 -3820
rect 5181 -3850 5261 -3827
rect 4341 -3869 4995 -3866
rect 3711 -3909 3751 -3869
rect 4041 -3909 4081 -3869
rect 1191 -3942 1271 -3909
rect 1191 -3976 1214 -3942
rect 1248 -3976 1271 -3942
rect 1191 -4022 1271 -3976
rect 1191 -4056 1214 -4022
rect 1248 -4056 1271 -4022
rect 1191 -4102 1271 -4056
rect 1191 -4136 1214 -4102
rect 1248 -4136 1271 -4102
rect 1191 -4159 1271 -4136
rect 1341 -3942 1421 -3909
rect 1341 -3976 1364 -3942
rect 1398 -3976 1421 -3942
rect 1341 -4022 1421 -3976
rect 1341 -4056 1364 -4022
rect 1398 -4056 1421 -4022
rect 1341 -4102 1421 -4056
rect 1341 -4136 1364 -4102
rect 1398 -4136 1421 -4102
rect 1341 -4159 1421 -4136
rect 1491 -3942 1571 -3909
rect 1491 -3976 1514 -3942
rect 1548 -3976 1571 -3942
rect 1491 -4022 1571 -3976
rect 1491 -4056 1514 -4022
rect 1548 -4056 1571 -4022
rect 1491 -4102 1571 -4056
rect 1491 -4136 1514 -4102
rect 1548 -4136 1571 -4102
rect 1491 -4159 1571 -4136
rect 1641 -3942 1721 -3909
rect 1641 -3976 1664 -3942
rect 1698 -3976 1721 -3942
rect 1641 -4022 1721 -3976
rect 1641 -4056 1664 -4022
rect 1698 -4056 1721 -4022
rect 1641 -4102 1721 -4056
rect 1641 -4136 1664 -4102
rect 1698 -4136 1721 -4102
rect 1641 -4159 1721 -4136
rect 1821 -3942 1901 -3909
rect 1821 -3976 1844 -3942
rect 1878 -3976 1901 -3942
rect 1821 -4022 1901 -3976
rect 1821 -4056 1844 -4022
rect 1878 -4056 1901 -4022
rect 1821 -4102 1901 -4056
rect 1821 -4136 1844 -4102
rect 1878 -4136 1901 -4102
rect 1821 -4159 1901 -4136
rect 1971 -3942 2051 -3909
rect 1971 -3976 1994 -3942
rect 2028 -3976 2051 -3942
rect 1971 -4022 2051 -3976
rect 1971 -4056 1994 -4022
rect 2028 -4056 2051 -4022
rect 1971 -4102 2051 -4056
rect 1971 -4136 1994 -4102
rect 2028 -4136 2051 -4102
rect 1971 -4159 2051 -4136
rect 2121 -3942 2201 -3909
rect 2121 -3976 2144 -3942
rect 2178 -3976 2201 -3942
rect 2121 -4022 2201 -3976
rect 2121 -4056 2144 -4022
rect 2178 -4056 2201 -4022
rect 2121 -4102 2201 -4056
rect 2121 -4136 2144 -4102
rect 2178 -4136 2201 -4102
rect 2121 -4159 2201 -4136
rect 2271 -3942 2351 -3909
rect 2271 -3976 2294 -3942
rect 2328 -3976 2351 -3942
rect 2271 -4022 2351 -3976
rect 2271 -4056 2294 -4022
rect 2328 -4056 2351 -4022
rect 2271 -4102 2351 -4056
rect 2271 -4136 2294 -4102
rect 2328 -4136 2351 -4102
rect 2271 -4159 2351 -4136
rect 2421 -3942 2501 -3909
rect 2421 -3976 2444 -3942
rect 2478 -3976 2501 -3942
rect 2421 -4022 2501 -3976
rect 2421 -4056 2444 -4022
rect 2478 -4056 2501 -4022
rect 2421 -4102 2501 -4056
rect 2421 -4136 2444 -4102
rect 2478 -4136 2501 -4102
rect 2421 -4159 2501 -4136
rect 2601 -3942 2681 -3909
rect 2601 -3976 2624 -3942
rect 2658 -3976 2681 -3942
rect 2601 -4022 2681 -3976
rect 2601 -4056 2624 -4022
rect 2658 -4056 2681 -4022
rect 2601 -4102 2681 -4056
rect 2601 -4136 2624 -4102
rect 2658 -4136 2681 -4102
rect 2601 -4159 2681 -4136
rect 3051 -3942 3131 -3909
rect 3051 -3976 3074 -3942
rect 3108 -3976 3131 -3942
rect 3051 -4022 3131 -3976
rect 3051 -4056 3074 -4022
rect 3108 -4056 3131 -4022
rect 3051 -4102 3131 -4056
rect 3051 -4136 3074 -4102
rect 3108 -4136 3131 -4102
rect 3051 -4159 3131 -4136
rect 3541 -3942 3621 -3909
rect 3541 -3976 3564 -3942
rect 3598 -3976 3621 -3942
rect 3541 -4022 3621 -3976
rect 3541 -4056 3564 -4022
rect 3598 -4056 3621 -4022
rect 3541 -4102 3621 -4056
rect 3541 -4136 3564 -4102
rect 3598 -4136 3621 -4102
rect 3541 -4159 3621 -4136
rect 3691 -3942 3771 -3909
rect 3691 -3976 3714 -3942
rect 3748 -3976 3771 -3942
rect 3691 -4022 3771 -3976
rect 3691 -4056 3714 -4022
rect 3748 -4056 3771 -4022
rect 3691 -4102 3771 -4056
rect 3691 -4136 3714 -4102
rect 3748 -4136 3771 -4102
rect 3691 -4159 3771 -4136
rect 3871 -3942 3951 -3909
rect 3871 -3976 3894 -3942
rect 3928 -3976 3951 -3942
rect 3871 -4022 3951 -3976
rect 3871 -4056 3894 -4022
rect 3928 -4056 3951 -4022
rect 3871 -4102 3951 -4056
rect 3871 -4136 3894 -4102
rect 3928 -4136 3951 -4102
rect 3871 -4159 3951 -4136
rect 4021 -3942 4101 -3909
rect 4021 -3976 4044 -3942
rect 4078 -3976 4101 -3942
rect 4021 -4022 4101 -3976
rect 4021 -4056 4044 -4022
rect 4078 -4056 4101 -4022
rect 4021 -4102 4101 -4056
rect 4021 -4136 4044 -4102
rect 4078 -4136 4101 -4102
rect 4021 -4159 4101 -4136
rect 4171 -3942 4251 -3909
rect 4171 -3976 4194 -3942
rect 4228 -3976 4251 -3942
rect 4171 -4022 4251 -3976
rect 4171 -4056 4194 -4022
rect 4228 -4056 4251 -4022
rect 4171 -4102 4251 -4056
rect 4171 -4136 4194 -4102
rect 4228 -4136 4251 -4102
rect 4171 -4159 4251 -4136
rect 4321 -3942 4401 -3869
rect 4671 -3909 4711 -3869
rect 4915 -3889 4995 -3869
rect 4321 -3976 4344 -3942
rect 4378 -3976 4401 -3942
rect 4321 -4022 4401 -3976
rect 4321 -4056 4344 -4022
rect 4378 -4056 4401 -4022
rect 4321 -4102 4401 -4056
rect 4321 -4136 4344 -4102
rect 4378 -4136 4401 -4102
rect 4321 -4159 4401 -4136
rect 4471 -3942 4551 -3909
rect 4471 -3976 4494 -3942
rect 4528 -3976 4551 -3942
rect 4471 -4022 4551 -3976
rect 4471 -4056 4494 -4022
rect 4528 -4056 4551 -4022
rect 4471 -4102 4551 -4056
rect 4471 -4136 4494 -4102
rect 4528 -4136 4551 -4102
rect 4471 -4159 4551 -4136
rect 4651 -3942 4731 -3909
rect 4651 -3976 4674 -3942
rect 4708 -3976 4731 -3942
rect 4651 -4022 4731 -3976
rect 4651 -4056 4674 -4022
rect 4708 -4056 4731 -4022
rect 4651 -4102 4731 -4056
rect 4651 -4136 4674 -4102
rect 4708 -4136 4731 -4102
rect 4651 -4159 4731 -4136
rect 4801 -3942 4881 -3909
rect 5451 -3910 5491 -3820
rect 5751 -3910 5791 -3820
rect 6081 -3910 6121 -3820
rect 6261 -3822 6284 -3820
rect 6318 -3822 6341 -3788
rect 6261 -3845 6341 -3822
rect 6381 -3830 6421 -3700
rect 6941 -3710 7021 -3690
rect 7389 -3710 7429 -3100
rect 6941 -3713 7429 -3710
rect 6941 -3747 6964 -3713
rect 6998 -3747 7429 -3713
rect 6941 -3750 7429 -3747
rect 6941 -3770 7021 -3750
rect 6791 -3793 6871 -3770
rect 6791 -3827 6814 -3793
rect 6848 -3810 6871 -3793
rect 6848 -3827 7241 -3810
rect 6381 -3870 6731 -3830
rect 6791 -3850 7241 -3827
rect 6381 -3910 6421 -3870
rect 6691 -3910 6731 -3870
rect 4801 -3976 4824 -3942
rect 4858 -3976 4881 -3942
rect 4801 -4022 4881 -3976
rect 4998 -3946 5078 -3923
rect 4998 -3980 5021 -3946
rect 5055 -3980 5078 -3946
rect 4998 -4003 5078 -3980
rect 5281 -3943 5361 -3910
rect 5281 -3977 5304 -3943
rect 5338 -3977 5361 -3943
rect 4801 -4056 4824 -4022
rect 4858 -4056 4881 -4022
rect 4801 -4102 4881 -4056
rect 4801 -4136 4824 -4102
rect 4858 -4136 4881 -4102
rect 4801 -4159 4881 -4136
rect 1171 -4219 1251 -4199
rect 1921 -4219 2001 -4199
rect 2321 -4219 2401 -4199
rect 3971 -4219 4051 -4199
rect 4371 -4219 4451 -4199
rect 5018 -4219 5058 -4003
rect 5281 -4023 5361 -3977
rect 5281 -4057 5304 -4023
rect 5338 -4057 5361 -4023
rect 5281 -4103 5361 -4057
rect 5281 -4137 5304 -4103
rect 5338 -4137 5361 -4103
rect 5281 -4160 5361 -4137
rect 5431 -3943 5511 -3910
rect 5431 -3977 5454 -3943
rect 5488 -3977 5511 -3943
rect 5431 -4023 5511 -3977
rect 5431 -4057 5454 -4023
rect 5488 -4057 5511 -4023
rect 5431 -4103 5511 -4057
rect 5431 -4137 5454 -4103
rect 5488 -4137 5511 -4103
rect 5431 -4160 5511 -4137
rect 5581 -3943 5661 -3910
rect 5581 -3977 5604 -3943
rect 5638 -3977 5661 -3943
rect 5581 -4023 5661 -3977
rect 5581 -4057 5604 -4023
rect 5638 -4057 5661 -4023
rect 5581 -4103 5661 -4057
rect 5581 -4137 5604 -4103
rect 5638 -4137 5661 -4103
rect 5581 -4160 5661 -4137
rect 5731 -3943 5811 -3910
rect 5731 -3977 5754 -3943
rect 5788 -3977 5811 -3943
rect 5731 -4023 5811 -3977
rect 5731 -4057 5754 -4023
rect 5788 -4057 5811 -4023
rect 5731 -4103 5811 -4057
rect 5731 -4137 5754 -4103
rect 5788 -4137 5811 -4103
rect 5731 -4160 5811 -4137
rect 5911 -3943 5991 -3910
rect 5911 -3977 5934 -3943
rect 5968 -3977 5991 -3943
rect 5911 -4023 5991 -3977
rect 5911 -4057 5934 -4023
rect 5968 -4057 5991 -4023
rect 5911 -4103 5991 -4057
rect 5911 -4137 5934 -4103
rect 5968 -4137 5991 -4103
rect 5911 -4160 5991 -4137
rect 6061 -3943 6141 -3910
rect 6061 -3977 6084 -3943
rect 6118 -3977 6141 -3943
rect 6061 -4023 6141 -3977
rect 6061 -4057 6084 -4023
rect 6118 -4057 6141 -4023
rect 6061 -4103 6141 -4057
rect 6061 -4137 6084 -4103
rect 6118 -4137 6141 -4103
rect 6061 -4160 6141 -4137
rect 6211 -3943 6291 -3910
rect 6211 -3977 6234 -3943
rect 6268 -3977 6291 -3943
rect 6211 -4023 6291 -3977
rect 6211 -4057 6234 -4023
rect 6268 -4057 6291 -4023
rect 6211 -4103 6291 -4057
rect 6211 -4137 6234 -4103
rect 6268 -4137 6291 -4103
rect 6211 -4160 6291 -4137
rect 6361 -3943 6441 -3910
rect 6361 -3977 6384 -3943
rect 6418 -3977 6441 -3943
rect 6361 -4023 6441 -3977
rect 6361 -4057 6384 -4023
rect 6418 -4057 6441 -4023
rect 6361 -4103 6441 -4057
rect 6361 -4137 6384 -4103
rect 6418 -4137 6441 -4103
rect 6361 -4160 6441 -4137
rect 6511 -3943 6591 -3910
rect 6511 -3977 6534 -3943
rect 6568 -3977 6591 -3943
rect 6511 -4023 6591 -3977
rect 6511 -4057 6534 -4023
rect 6568 -4057 6591 -4023
rect 6511 -4103 6591 -4057
rect 6511 -4137 6534 -4103
rect 6568 -4137 6591 -4103
rect 6511 -4160 6591 -4137
rect 6691 -3943 6771 -3910
rect 6691 -3977 6714 -3943
rect 6748 -3977 6771 -3943
rect 6691 -4023 6771 -3977
rect 6691 -4057 6714 -4023
rect 6748 -4057 6771 -4023
rect 6691 -4103 6771 -4057
rect 6691 -4137 6714 -4103
rect 6748 -4137 6771 -4103
rect 6691 -4160 6771 -4137
rect 7141 -3943 7221 -3910
rect 7141 -3977 7164 -3943
rect 7198 -3977 7221 -3943
rect 7141 -4023 7221 -3977
rect 7141 -4057 7164 -4023
rect 7198 -4057 7221 -4023
rect 7141 -4103 7221 -4057
rect 7141 -4137 7164 -4103
rect 7198 -4137 7221 -4103
rect 7141 -4160 7221 -4137
rect 1171 -4222 2401 -4219
rect 1171 -4256 1194 -4222
rect 1228 -4256 1944 -4222
rect 1978 -4256 2344 -4222
rect 2378 -4256 2401 -4222
rect 1171 -4259 2401 -4256
rect 3521 -4222 5058 -4219
rect 3521 -4256 3994 -4222
rect 4028 -4256 4394 -4222
rect 4428 -4256 5058 -4222
rect 3521 -4259 5058 -4256
rect 5092 -4220 5172 -4201
rect 6011 -4220 6091 -4200
rect 6411 -4220 6491 -4200
rect 5092 -4223 7241 -4220
rect 5092 -4224 6034 -4223
rect 5092 -4258 5115 -4224
rect 5149 -4257 6034 -4224
rect 6068 -4257 6434 -4223
rect 6468 -4257 7241 -4223
rect 5149 -4258 7241 -4257
rect 1171 -4279 1251 -4259
rect 1921 -4279 2001 -4259
rect 2321 -4279 2401 -4259
rect 3971 -4279 4051 -4259
rect 4371 -4279 4451 -4259
rect 5092 -4260 7241 -4258
rect 5092 -4281 5172 -4260
rect 6011 -4280 6091 -4260
rect 6411 -4280 6491 -4260
rect 912 -4342 3360 -4319
rect 912 -4376 935 -4342
rect 969 -4376 1184 -4342
rect 1218 -4376 1264 -4342
rect 1298 -4376 1344 -4342
rect 1378 -4376 1424 -4342
rect 1458 -4376 1504 -4342
rect 1538 -4376 1584 -4342
rect 1618 -4376 1664 -4342
rect 1698 -4376 1744 -4342
rect 1778 -4376 1824 -4342
rect 1858 -4376 1904 -4342
rect 1938 -4376 1984 -4342
rect 2018 -4376 2064 -4342
rect 2098 -4376 2144 -4342
rect 2178 -4376 2224 -4342
rect 2258 -4376 2304 -4342
rect 2338 -4376 2384 -4342
rect 2418 -4376 2464 -4342
rect 2498 -4376 2544 -4342
rect 2578 -4376 2624 -4342
rect 2658 -4376 2704 -4342
rect 2738 -4376 2784 -4342
rect 2818 -4376 2864 -4342
rect 2898 -4376 2944 -4342
rect 2978 -4376 3024 -4342
rect 3058 -4376 3104 -4342
rect 3138 -4376 3184 -4342
rect 3218 -4376 3264 -4342
rect 3298 -4376 3360 -4342
rect 912 -4399 3360 -4376
rect 913 -4422 3360 -4399
rect 913 -4456 936 -4422
rect 970 -4456 1063 -4422
rect 1097 -4456 1143 -4422
rect 1177 -4456 1223 -4422
rect 1257 -4456 1303 -4422
rect 1337 -4456 1383 -4422
rect 1417 -4456 1463 -4422
rect 1497 -4456 1543 -4422
rect 1577 -4456 1623 -4422
rect 1657 -4456 1703 -4422
rect 1737 -4456 1783 -4422
rect 1817 -4456 1863 -4422
rect 1897 -4456 1943 -4422
rect 1977 -4456 2023 -4422
rect 2057 -4456 2103 -4422
rect 2137 -4456 2183 -4422
rect 2217 -4456 2263 -4422
rect 2297 -4456 2343 -4422
rect 2377 -4456 2423 -4422
rect 2457 -4456 2503 -4422
rect 2537 -4456 2583 -4422
rect 2617 -4456 2663 -4422
rect 2697 -4456 2743 -4422
rect 2777 -4456 2823 -4422
rect 2857 -4456 2903 -4422
rect 2937 -4456 2983 -4422
rect 3017 -4456 3063 -4422
rect 3097 -4456 3143 -4422
rect 3177 -4456 3223 -4422
rect 3257 -4456 3303 -4422
rect 3337 -4456 3360 -4422
rect 913 -4479 3360 -4456
rect 3521 -4342 5101 -4319
rect 7251 -4320 7470 -4319
rect 3521 -4376 3554 -4342
rect 3588 -4376 3634 -4342
rect 3668 -4376 3714 -4342
rect 3748 -4376 3794 -4342
rect 3828 -4376 3874 -4342
rect 3908 -4376 3954 -4342
rect 3988 -4376 4034 -4342
rect 4068 -4376 4114 -4342
rect 4148 -4376 4194 -4342
rect 4228 -4376 4274 -4342
rect 4308 -4376 4354 -4342
rect 4388 -4376 4434 -4342
rect 4468 -4376 4514 -4342
rect 4548 -4376 4594 -4342
rect 4628 -4376 4674 -4342
rect 4708 -4376 4754 -4342
rect 4788 -4376 4834 -4342
rect 4868 -4376 4914 -4342
rect 4948 -4376 4994 -4342
rect 5028 -4376 5101 -4342
rect 3521 -4423 5101 -4376
rect 3521 -4457 3594 -4423
rect 3628 -4457 3674 -4423
rect 3708 -4457 3754 -4423
rect 3788 -4457 3834 -4423
rect 3868 -4457 3914 -4423
rect 3948 -4457 3994 -4423
rect 4028 -4457 4074 -4423
rect 4108 -4457 4154 -4423
rect 4188 -4457 4234 -4423
rect 4268 -4457 4314 -4423
rect 4348 -4457 4394 -4423
rect 4428 -4457 4474 -4423
rect 4508 -4457 4554 -4423
rect 4588 -4457 4634 -4423
rect 4668 -4457 4714 -4423
rect 4748 -4457 4794 -4423
rect 4828 -4457 4874 -4423
rect 4908 -4457 4954 -4423
rect 4988 -4457 5034 -4423
rect 5068 -4457 5101 -4423
rect 3521 -4480 5101 -4457
rect 5251 -4342 7470 -4320
rect 5251 -4343 7274 -4342
rect 5251 -4377 5274 -4343
rect 5308 -4377 5354 -4343
rect 5388 -4377 5434 -4343
rect 5468 -4377 5514 -4343
rect 5548 -4377 5594 -4343
rect 5628 -4377 5674 -4343
rect 5708 -4377 5754 -4343
rect 5788 -4377 5834 -4343
rect 5868 -4377 5914 -4343
rect 5948 -4377 5994 -4343
rect 6028 -4377 6074 -4343
rect 6108 -4377 6154 -4343
rect 6188 -4377 6234 -4343
rect 6268 -4377 6314 -4343
rect 6348 -4377 6394 -4343
rect 6428 -4377 6474 -4343
rect 6508 -4377 6554 -4343
rect 6588 -4377 6634 -4343
rect 6668 -4377 6714 -4343
rect 6748 -4377 6794 -4343
rect 6828 -4377 6874 -4343
rect 6908 -4377 6954 -4343
rect 6988 -4377 7034 -4343
rect 7068 -4377 7114 -4343
rect 7148 -4377 7194 -4343
rect 7228 -4376 7274 -4343
rect 7308 -4376 7354 -4342
rect 7388 -4376 7470 -4342
rect 7228 -4377 7470 -4376
rect 5251 -4423 7470 -4377
rect 5251 -4457 5333 -4423
rect 5367 -4457 5413 -4423
rect 5447 -4457 5493 -4423
rect 5527 -4457 5573 -4423
rect 5607 -4457 5653 -4423
rect 5687 -4457 5733 -4423
rect 5767 -4457 5813 -4423
rect 5847 -4457 5893 -4423
rect 5927 -4457 5973 -4423
rect 6007 -4457 6053 -4423
rect 6087 -4457 6133 -4423
rect 6167 -4457 6213 -4423
rect 6247 -4457 6293 -4423
rect 6327 -4457 6373 -4423
rect 6407 -4457 6453 -4423
rect 6487 -4457 6533 -4423
rect 6567 -4457 6613 -4423
rect 6647 -4457 6693 -4423
rect 6727 -4457 6773 -4423
rect 6807 -4457 6853 -4423
rect 6887 -4457 6933 -4423
rect 6967 -4457 7013 -4423
rect 7047 -4457 7093 -4423
rect 7127 -4457 7173 -4423
rect 7207 -4457 7253 -4423
rect 7287 -4457 7333 -4423
rect 7367 -4457 7413 -4423
rect 7447 -4457 7470 -4423
rect 5251 -4480 7470 -4457
rect 1041 -4539 1121 -4522
rect 1960 -4539 2040 -4519
rect 2360 -4539 2440 -4519
rect 1041 -4542 2440 -4539
rect 4171 -4540 4251 -4520
rect 4571 -4540 4651 -4520
rect 5115 -4540 5195 -4520
rect 1041 -4545 1983 -4542
rect 1041 -4579 1064 -4545
rect 1098 -4576 1983 -4545
rect 2017 -4576 2383 -4542
rect 2417 -4576 2440 -4542
rect 1098 -4579 2440 -4576
rect 1041 -4602 1121 -4579
rect 1960 -4599 2040 -4579
rect 2360 -4599 2440 -4579
rect 3721 -4543 5195 -4540
rect 3721 -4577 4194 -4543
rect 4228 -4577 4594 -4543
rect 4628 -4577 5138 -4543
rect 5172 -4577 5195 -4543
rect 3721 -4580 5195 -4577
rect 4171 -4600 4251 -4580
rect 4571 -4600 4651 -4580
rect 5115 -4600 5195 -4580
rect 5312 -4540 5392 -4520
rect 6230 -4540 6310 -4520
rect 6630 -4540 6710 -4520
rect 5312 -4543 7460 -4540
rect 5312 -4577 5335 -4543
rect 5369 -4577 6253 -4543
rect 6287 -4577 6653 -4543
rect 6687 -4577 7460 -4543
rect 5312 -4580 7460 -4577
rect 5312 -4600 5392 -4580
rect 6230 -4600 6310 -4580
rect 6630 -4600 6710 -4580
rect 1080 -4662 1160 -4639
rect 1080 -4696 1103 -4662
rect 1137 -4696 1160 -4662
rect 1080 -4742 1160 -4696
rect 1080 -4776 1103 -4742
rect 1137 -4776 1160 -4742
rect 1080 -4822 1160 -4776
rect 1080 -4856 1103 -4822
rect 1137 -4856 1160 -4822
rect 1080 -4889 1160 -4856
rect 1230 -4662 1310 -4639
rect 1230 -4696 1253 -4662
rect 1287 -4696 1310 -4662
rect 1230 -4742 1310 -4696
rect 1230 -4776 1253 -4742
rect 1287 -4776 1310 -4742
rect 1230 -4822 1310 -4776
rect 1230 -4856 1253 -4822
rect 1287 -4856 1310 -4822
rect 1230 -4889 1310 -4856
rect 1380 -4662 1460 -4639
rect 1380 -4696 1403 -4662
rect 1437 -4696 1460 -4662
rect 1380 -4742 1460 -4696
rect 1380 -4776 1403 -4742
rect 1437 -4776 1460 -4742
rect 1380 -4822 1460 -4776
rect 1380 -4856 1403 -4822
rect 1437 -4856 1460 -4822
rect 1380 -4889 1460 -4856
rect 1530 -4662 1610 -4639
rect 1530 -4696 1553 -4662
rect 1587 -4696 1610 -4662
rect 1530 -4742 1610 -4696
rect 1530 -4776 1553 -4742
rect 1587 -4776 1610 -4742
rect 1530 -4822 1610 -4776
rect 1530 -4856 1553 -4822
rect 1587 -4856 1610 -4822
rect 1530 -4889 1610 -4856
rect 1680 -4662 1760 -4639
rect 1680 -4696 1703 -4662
rect 1737 -4696 1760 -4662
rect 1680 -4742 1760 -4696
rect 1680 -4776 1703 -4742
rect 1737 -4776 1760 -4742
rect 1680 -4822 1760 -4776
rect 1680 -4856 1703 -4822
rect 1737 -4856 1760 -4822
rect 1680 -4889 1760 -4856
rect 1860 -4662 1940 -4639
rect 1860 -4696 1883 -4662
rect 1917 -4696 1940 -4662
rect 1860 -4742 1940 -4696
rect 1860 -4776 1883 -4742
rect 1917 -4776 1940 -4742
rect 1860 -4822 1940 -4776
rect 1860 -4856 1883 -4822
rect 1917 -4856 1940 -4822
rect 1860 -4889 1940 -4856
rect 2010 -4662 2090 -4639
rect 2010 -4696 2033 -4662
rect 2067 -4696 2090 -4662
rect 2010 -4742 2090 -4696
rect 2010 -4776 2033 -4742
rect 2067 -4776 2090 -4742
rect 2010 -4822 2090 -4776
rect 2010 -4856 2033 -4822
rect 2067 -4856 2090 -4822
rect 2010 -4889 2090 -4856
rect 2160 -4662 2240 -4639
rect 2160 -4696 2183 -4662
rect 2217 -4696 2240 -4662
rect 2160 -4742 2240 -4696
rect 2160 -4776 2183 -4742
rect 2217 -4776 2240 -4742
rect 2160 -4822 2240 -4776
rect 2160 -4856 2183 -4822
rect 2217 -4856 2240 -4822
rect 2160 -4889 2240 -4856
rect 2310 -4662 2390 -4639
rect 2310 -4696 2333 -4662
rect 2367 -4696 2390 -4662
rect 2310 -4742 2390 -4696
rect 2310 -4776 2333 -4742
rect 2367 -4776 2390 -4742
rect 2310 -4822 2390 -4776
rect 2310 -4856 2333 -4822
rect 2367 -4856 2390 -4822
rect 2310 -4889 2390 -4856
rect 2460 -4662 2540 -4639
rect 2460 -4696 2483 -4662
rect 2517 -4696 2540 -4662
rect 2460 -4742 2540 -4696
rect 2460 -4776 2483 -4742
rect 2517 -4776 2540 -4742
rect 2460 -4822 2540 -4776
rect 2460 -4856 2483 -4822
rect 2517 -4856 2540 -4822
rect 2460 -4889 2540 -4856
rect 2640 -4662 2720 -4639
rect 2640 -4696 2663 -4662
rect 2697 -4696 2720 -4662
rect 2640 -4742 2720 -4696
rect 2640 -4776 2663 -4742
rect 2697 -4776 2720 -4742
rect 2640 -4822 2720 -4776
rect 2640 -4856 2663 -4822
rect 2697 -4856 2720 -4822
rect 2640 -4889 2720 -4856
rect 3240 -4662 3320 -4639
rect 3240 -4696 3263 -4662
rect 3297 -4696 3320 -4662
rect 3240 -4742 3320 -4696
rect 3240 -4776 3263 -4742
rect 3297 -4776 3320 -4742
rect 3240 -4822 3320 -4776
rect 3240 -4856 3263 -4822
rect 3297 -4856 3320 -4822
rect 3240 -4889 3320 -4856
rect 3741 -4663 3821 -4640
rect 3741 -4697 3764 -4663
rect 3798 -4697 3821 -4663
rect 3741 -4743 3821 -4697
rect 3741 -4777 3764 -4743
rect 3798 -4777 3821 -4743
rect 3741 -4823 3821 -4777
rect 3741 -4857 3764 -4823
rect 3798 -4857 3821 -4823
rect 1100 -4929 1140 -4889
rect 1400 -4929 1440 -4889
rect 1700 -4929 1740 -4889
rect 2030 -4929 2070 -4889
rect 1100 -4969 2070 -4929
rect 570 -5012 650 -4989
rect 570 -5046 593 -5012
rect 627 -5029 650 -5012
rect 1130 -5029 1210 -5009
rect 627 -5032 1210 -5029
rect 627 -5046 1153 -5032
rect 570 -5066 1153 -5046
rect 1187 -5066 1210 -5032
rect 570 -5069 1210 -5066
rect 1130 -5089 1210 -5069
rect 1280 -5129 1360 -5109
rect 114 -5132 1360 -5129
rect 114 -5152 1303 -5132
rect 114 -5186 137 -5152
rect 171 -5166 1303 -5152
rect 1337 -5166 1360 -5132
rect 171 -5169 1360 -5166
rect 171 -5186 194 -5169
rect 114 -5209 194 -5186
rect 1280 -5189 1360 -5169
rect 1430 -5229 1510 -5209
rect 342 -5232 1510 -5229
rect 342 -5252 1453 -5232
rect 342 -5286 365 -5252
rect 399 -5266 1453 -5252
rect 1487 -5266 1510 -5232
rect 399 -5269 1510 -5266
rect 399 -5286 422 -5269
rect 342 -5309 422 -5286
rect 1430 -5289 1510 -5269
rect 684 -5329 764 -5309
rect 1580 -5329 1660 -5309
rect 684 -5332 1660 -5329
rect 684 -5366 707 -5332
rect 741 -5366 1603 -5332
rect 1637 -5366 1660 -5332
rect 684 -5369 1660 -5366
rect 684 -5389 764 -5369
rect 1580 -5389 1660 -5369
rect 2030 -5329 2070 -4969
rect 2330 -4929 2370 -4889
rect 2640 -4929 2680 -4889
rect 3741 -4890 3821 -4857
rect 3891 -4663 3971 -4640
rect 3891 -4697 3914 -4663
rect 3948 -4697 3971 -4663
rect 3891 -4743 3971 -4697
rect 3891 -4777 3914 -4743
rect 3948 -4777 3971 -4743
rect 3891 -4823 3971 -4777
rect 3891 -4857 3914 -4823
rect 3948 -4857 3971 -4823
rect 3891 -4890 3971 -4857
rect 4071 -4663 4151 -4640
rect 4071 -4697 4094 -4663
rect 4128 -4697 4151 -4663
rect 4071 -4743 4151 -4697
rect 4071 -4777 4094 -4743
rect 4128 -4777 4151 -4743
rect 4071 -4823 4151 -4777
rect 4071 -4857 4094 -4823
rect 4128 -4857 4151 -4823
rect 4071 -4890 4151 -4857
rect 4221 -4663 4301 -4640
rect 4221 -4697 4244 -4663
rect 4278 -4697 4301 -4663
rect 4221 -4743 4301 -4697
rect 4221 -4777 4244 -4743
rect 4278 -4777 4301 -4743
rect 4221 -4823 4301 -4777
rect 4221 -4857 4244 -4823
rect 4278 -4857 4301 -4823
rect 4221 -4890 4301 -4857
rect 4371 -4663 4451 -4640
rect 4371 -4697 4394 -4663
rect 4428 -4697 4451 -4663
rect 4371 -4743 4451 -4697
rect 4371 -4777 4394 -4743
rect 4428 -4777 4451 -4743
rect 4371 -4823 4451 -4777
rect 4371 -4857 4394 -4823
rect 4428 -4857 4451 -4823
rect 4371 -4890 4451 -4857
rect 4521 -4663 4601 -4640
rect 4521 -4697 4544 -4663
rect 4578 -4697 4601 -4663
rect 4521 -4743 4601 -4697
rect 4521 -4777 4544 -4743
rect 4578 -4777 4601 -4743
rect 4521 -4823 4601 -4777
rect 4521 -4857 4544 -4823
rect 4578 -4857 4601 -4823
rect 2330 -4969 2680 -4929
rect 3911 -4930 3951 -4890
rect 4241 -4930 4281 -4890
rect 4521 -4930 4601 -4857
rect 4671 -4663 4751 -4640
rect 4671 -4697 4694 -4663
rect 4728 -4697 4751 -4663
rect 4671 -4743 4751 -4697
rect 4671 -4777 4694 -4743
rect 4728 -4777 4751 -4743
rect 4671 -4823 4751 -4777
rect 4671 -4857 4694 -4823
rect 4728 -4857 4751 -4823
rect 4671 -4890 4751 -4857
rect 4851 -4663 4931 -4640
rect 4851 -4697 4874 -4663
rect 4908 -4697 4931 -4663
rect 4851 -4743 4931 -4697
rect 4851 -4777 4874 -4743
rect 4908 -4777 4931 -4743
rect 4851 -4823 4931 -4777
rect 4851 -4857 4874 -4823
rect 4908 -4857 4931 -4823
rect 4851 -4890 4931 -4857
rect 5001 -4663 5081 -4640
rect 5001 -4697 5024 -4663
rect 5058 -4697 5081 -4663
rect 5001 -4743 5081 -4697
rect 5001 -4777 5024 -4743
rect 5058 -4777 5081 -4743
rect 5001 -4823 5081 -4777
rect 5001 -4857 5024 -4823
rect 5058 -4857 5081 -4823
rect 5001 -4890 5081 -4857
rect 5500 -4663 5580 -4640
rect 5500 -4697 5523 -4663
rect 5557 -4697 5580 -4663
rect 5500 -4743 5580 -4697
rect 5500 -4777 5523 -4743
rect 5557 -4777 5580 -4743
rect 5500 -4823 5580 -4777
rect 5500 -4857 5523 -4823
rect 5557 -4857 5580 -4823
rect 5500 -4890 5580 -4857
rect 5650 -4663 5730 -4640
rect 5650 -4697 5673 -4663
rect 5707 -4697 5730 -4663
rect 5650 -4743 5730 -4697
rect 5650 -4777 5673 -4743
rect 5707 -4777 5730 -4743
rect 5650 -4823 5730 -4777
rect 5650 -4857 5673 -4823
rect 5707 -4857 5730 -4823
rect 5650 -4890 5730 -4857
rect 5800 -4663 5880 -4640
rect 5800 -4697 5823 -4663
rect 5857 -4697 5880 -4663
rect 5800 -4743 5880 -4697
rect 5800 -4777 5823 -4743
rect 5857 -4777 5880 -4743
rect 5800 -4823 5880 -4777
rect 5800 -4857 5823 -4823
rect 5857 -4857 5880 -4823
rect 5800 -4890 5880 -4857
rect 5950 -4663 6030 -4640
rect 5950 -4697 5973 -4663
rect 6007 -4697 6030 -4663
rect 5950 -4743 6030 -4697
rect 5950 -4777 5973 -4743
rect 6007 -4777 6030 -4743
rect 5950 -4823 6030 -4777
rect 5950 -4857 5973 -4823
rect 6007 -4857 6030 -4823
rect 5950 -4890 6030 -4857
rect 6130 -4663 6210 -4640
rect 6130 -4697 6153 -4663
rect 6187 -4697 6210 -4663
rect 6130 -4743 6210 -4697
rect 6130 -4777 6153 -4743
rect 6187 -4777 6210 -4743
rect 6130 -4823 6210 -4777
rect 6130 -4857 6153 -4823
rect 6187 -4857 6210 -4823
rect 6130 -4890 6210 -4857
rect 6280 -4663 6360 -4640
rect 6280 -4697 6303 -4663
rect 6337 -4697 6360 -4663
rect 6280 -4743 6360 -4697
rect 6280 -4777 6303 -4743
rect 6337 -4777 6360 -4743
rect 6280 -4823 6360 -4777
rect 6280 -4857 6303 -4823
rect 6337 -4857 6360 -4823
rect 6280 -4890 6360 -4857
rect 6430 -4663 6510 -4640
rect 6430 -4697 6453 -4663
rect 6487 -4697 6510 -4663
rect 6430 -4743 6510 -4697
rect 6430 -4777 6453 -4743
rect 6487 -4777 6510 -4743
rect 6430 -4823 6510 -4777
rect 6430 -4857 6453 -4823
rect 6487 -4857 6510 -4823
rect 6430 -4890 6510 -4857
rect 6580 -4663 6660 -4640
rect 6580 -4697 6603 -4663
rect 6637 -4697 6660 -4663
rect 6580 -4743 6660 -4697
rect 6580 -4777 6603 -4743
rect 6637 -4777 6660 -4743
rect 6580 -4823 6660 -4777
rect 6580 -4857 6603 -4823
rect 6637 -4857 6660 -4823
rect 6580 -4890 6660 -4857
rect 6730 -4663 6810 -4640
rect 6730 -4697 6753 -4663
rect 6787 -4697 6810 -4663
rect 6730 -4743 6810 -4697
rect 6730 -4777 6753 -4743
rect 6787 -4777 6810 -4743
rect 6730 -4823 6810 -4777
rect 6730 -4857 6753 -4823
rect 6787 -4857 6810 -4823
rect 6730 -4890 6810 -4857
rect 6910 -4663 6990 -4640
rect 6910 -4697 6933 -4663
rect 6967 -4697 6990 -4663
rect 6910 -4743 6990 -4697
rect 6910 -4777 6933 -4743
rect 6967 -4777 6990 -4743
rect 6910 -4823 6990 -4777
rect 6910 -4857 6933 -4823
rect 6967 -4857 6990 -4823
rect 6910 -4890 6990 -4857
rect 7360 -4663 7440 -4640
rect 7360 -4697 7383 -4663
rect 7417 -4697 7440 -4663
rect 7360 -4743 7440 -4697
rect 7360 -4777 7383 -4743
rect 7417 -4777 7440 -4743
rect 7360 -4823 7440 -4777
rect 7360 -4857 7383 -4823
rect 7417 -4857 7440 -4823
rect 7360 -4890 7440 -4857
rect 4871 -4930 4911 -4890
rect 5115 -4930 5195 -4910
rect 2110 -5192 2190 -5169
rect 2110 -5226 2133 -5192
rect 2167 -5209 2190 -5192
rect 2330 -5209 2370 -4969
rect 3633 -4980 3713 -4960
rect 3791 -4980 3871 -4960
rect 3911 -4970 4281 -4930
rect 4541 -4933 5195 -4930
rect 3633 -4983 3871 -4980
rect 2690 -5032 2770 -5009
rect 2690 -5066 2713 -5032
rect 2747 -5066 2770 -5032
rect 2690 -5089 2770 -5066
rect 2840 -5032 2920 -5009
rect 2840 -5066 2863 -5032
rect 2897 -5066 2920 -5032
rect 2840 -5089 2920 -5066
rect 2990 -5032 3070 -5009
rect 2990 -5066 3013 -5032
rect 3047 -5066 3070 -5032
rect 2990 -5089 3070 -5066
rect 3140 -5032 3220 -5009
rect 3140 -5066 3163 -5032
rect 3197 -5066 3220 -5032
rect 3633 -5017 3656 -4983
rect 3690 -5017 3814 -4983
rect 3848 -5017 3871 -4983
rect 3633 -5020 3871 -5017
rect 3633 -5040 3713 -5020
rect 3791 -5040 3871 -5020
rect 3140 -5089 3220 -5066
rect 4241 -5100 4281 -4970
rect 4321 -4978 4401 -4955
rect 4321 -5012 4344 -4978
rect 4378 -4980 4401 -4978
rect 4541 -4967 5138 -4933
rect 5172 -4967 5195 -4933
rect 4541 -4970 5195 -4967
rect 4541 -4980 4581 -4970
rect 4378 -5012 4581 -4980
rect 5115 -4990 5195 -4970
rect 5400 -4963 5480 -4940
rect 4321 -5020 4581 -5012
rect 5400 -4997 5423 -4963
rect 5457 -4980 5480 -4963
rect 5670 -4980 5710 -4890
rect 5970 -4980 6010 -4890
rect 6300 -4980 6340 -4890
rect 6600 -4930 6640 -4890
rect 6910 -4930 6950 -4890
rect 6480 -4978 6560 -4955
rect 6480 -4980 6503 -4978
rect 5457 -4997 6503 -4980
rect 5400 -5012 6503 -4997
rect 6537 -5012 6560 -4978
rect 5400 -5020 6560 -5012
rect 4321 -5035 4401 -5020
rect 4421 -5100 4501 -5080
rect 4241 -5103 4501 -5100
rect 4241 -5137 4444 -5103
rect 4478 -5137 4501 -5103
rect 4241 -5140 4501 -5137
rect 4241 -5190 4281 -5140
rect 4421 -5160 4501 -5140
rect 4541 -5190 4581 -5020
rect 4821 -5100 4901 -5080
rect 5400 -5083 5480 -5060
rect 4821 -5103 5255 -5100
rect 4821 -5137 4844 -5103
rect 4878 -5137 5255 -5103
rect 4821 -5140 5255 -5137
rect 5400 -5117 5423 -5083
rect 5457 -5100 5480 -5083
rect 5980 -5100 6060 -5080
rect 5457 -5103 6060 -5100
rect 5457 -5117 6003 -5103
rect 5400 -5137 6003 -5117
rect 6037 -5137 6060 -5103
rect 5400 -5140 6060 -5137
rect 4821 -5160 4901 -5140
rect 2167 -5220 3553 -5209
rect 3921 -5220 4001 -5200
rect 2167 -5223 4001 -5220
rect 2167 -5226 3944 -5223
rect 2110 -5249 3944 -5226
rect 2210 -5329 2290 -5309
rect 2030 -5332 2290 -5329
rect 2030 -5366 2233 -5332
rect 2267 -5366 2290 -5332
rect 2030 -5369 2290 -5366
rect 456 -5412 536 -5389
rect 456 -5446 479 -5412
rect 513 -5429 536 -5412
rect 1130 -5429 1210 -5409
rect 513 -5432 1210 -5429
rect 513 -5446 1153 -5432
rect 456 -5466 1153 -5446
rect 1187 -5466 1210 -5432
rect 456 -5469 1210 -5466
rect 1130 -5489 1210 -5469
rect 2030 -5509 2070 -5369
rect 2210 -5389 2290 -5369
rect 2330 -5509 2370 -5249
rect 3513 -5257 3944 -5249
rect 3978 -5257 4001 -5223
rect 3513 -5260 4001 -5257
rect 3921 -5280 4001 -5260
rect 4071 -5223 4151 -5200
rect 4071 -5257 4094 -5223
rect 4128 -5257 4151 -5223
rect 4071 -5303 4151 -5257
rect 2410 -5329 2490 -5309
rect 3340 -5329 3420 -5310
rect 2410 -5332 3420 -5329
rect 2410 -5366 2433 -5332
rect 2467 -5333 3420 -5332
rect 2467 -5366 3363 -5333
rect 2410 -5367 3363 -5366
rect 3397 -5367 3420 -5333
rect 2410 -5369 3420 -5367
rect 2410 -5389 2490 -5369
rect 3340 -5390 3420 -5369
rect 4071 -5337 4094 -5303
rect 4128 -5337 4151 -5303
rect 4071 -5383 4151 -5337
rect 4071 -5417 4094 -5383
rect 4128 -5417 4151 -5383
rect 4071 -5450 4151 -5417
rect 4221 -5223 4301 -5190
rect 4221 -5257 4244 -5223
rect 4278 -5257 4301 -5223
rect 4221 -5303 4301 -5257
rect 4221 -5337 4244 -5303
rect 4278 -5337 4301 -5303
rect 4221 -5383 4301 -5337
rect 4221 -5417 4244 -5383
rect 4278 -5417 4301 -5383
rect 4221 -5450 4301 -5417
rect 4371 -5223 4451 -5200
rect 4371 -5257 4394 -5223
rect 4428 -5257 4451 -5223
rect 4371 -5303 4451 -5257
rect 4371 -5337 4394 -5303
rect 4428 -5337 4451 -5303
rect 4371 -5383 4451 -5337
rect 4371 -5417 4394 -5383
rect 4428 -5417 4451 -5383
rect 4371 -5450 4451 -5417
rect 4521 -5223 4601 -5190
rect 5215 -5192 5255 -5140
rect 5980 -5160 6060 -5140
rect 5400 -5192 5480 -5188
rect 6300 -5190 6340 -5020
rect 6480 -5035 6560 -5020
rect 6600 -4970 6950 -4930
rect 6380 -5100 6460 -5080
rect 6600 -5100 6640 -4970
rect 7010 -4973 7460 -4950
rect 7010 -5007 7033 -4973
rect 7067 -4990 7460 -4973
rect 7067 -5007 7090 -4990
rect 7010 -5030 7090 -5007
rect 6380 -5103 6640 -5100
rect 6380 -5137 6403 -5103
rect 6437 -5137 6640 -5103
rect 7160 -5050 7240 -5030
rect 7160 -5053 7648 -5050
rect 7160 -5087 7183 -5053
rect 7217 -5087 7648 -5053
rect 7160 -5090 7648 -5087
rect 7160 -5110 7240 -5090
rect 6380 -5140 6640 -5137
rect 6380 -5160 6460 -5140
rect 6600 -5190 6640 -5140
rect 7300 -5153 7380 -5130
rect 7300 -5187 7323 -5153
rect 7357 -5170 7380 -5153
rect 7494 -5170 7574 -5153
rect 7357 -5176 7574 -5170
rect 7357 -5187 7517 -5176
rect 4521 -5257 4544 -5223
rect 4578 -5257 4601 -5223
rect 4521 -5303 4601 -5257
rect 4521 -5337 4544 -5303
rect 4578 -5337 4601 -5303
rect 4521 -5383 4601 -5337
rect 4521 -5417 4544 -5383
rect 4578 -5417 4601 -5383
rect 4521 -5450 4601 -5417
rect 4671 -5223 4751 -5200
rect 4671 -5257 4694 -5223
rect 4728 -5257 4751 -5223
rect 4671 -5303 4751 -5257
rect 4821 -5220 4901 -5200
rect 4951 -5220 5031 -5200
rect 4821 -5223 5031 -5220
rect 4821 -5257 4844 -5223
rect 4878 -5257 4974 -5223
rect 5008 -5257 5031 -5223
rect 5215 -5211 5480 -5192
rect 5215 -5232 5423 -5211
rect 4821 -5260 5031 -5257
rect 4821 -5280 4901 -5260
rect 4951 -5280 5031 -5260
rect 5400 -5245 5423 -5232
rect 5457 -5245 5480 -5211
rect 6130 -5223 6210 -5200
rect 5400 -5268 5480 -5245
rect 5900 -5263 5980 -5240
rect 4671 -5337 4694 -5303
rect 4728 -5337 4751 -5303
rect 5900 -5297 5923 -5263
rect 5957 -5297 5980 -5263
rect 5900 -5320 5980 -5297
rect 6130 -5257 6153 -5223
rect 6187 -5257 6210 -5223
rect 6130 -5303 6210 -5257
rect 4671 -5383 4751 -5337
rect 5700 -5353 5780 -5330
rect 4671 -5417 4694 -5383
rect 4728 -5417 4751 -5383
rect 4671 -5450 4751 -5417
rect 5115 -5396 5195 -5373
rect 5115 -5430 5138 -5396
rect 5172 -5430 5195 -5396
rect 5700 -5387 5723 -5353
rect 5757 -5387 5780 -5353
rect 5700 -5410 5780 -5387
rect 6130 -5337 6153 -5303
rect 6187 -5337 6210 -5303
rect 6130 -5383 6210 -5337
rect 5115 -5453 5195 -5430
rect 6130 -5417 6153 -5383
rect 6187 -5417 6210 -5383
rect 6130 -5450 6210 -5417
rect 6280 -5223 6360 -5190
rect 6280 -5257 6303 -5223
rect 6337 -5257 6360 -5223
rect 6280 -5303 6360 -5257
rect 6280 -5337 6303 -5303
rect 6337 -5337 6360 -5303
rect 6280 -5383 6360 -5337
rect 6280 -5417 6303 -5383
rect 6337 -5417 6360 -5383
rect 6280 -5450 6360 -5417
rect 6430 -5223 6510 -5200
rect 6430 -5257 6453 -5223
rect 6487 -5257 6510 -5223
rect 6430 -5303 6510 -5257
rect 6430 -5337 6453 -5303
rect 6487 -5337 6510 -5303
rect 6430 -5383 6510 -5337
rect 6430 -5417 6453 -5383
rect 6487 -5417 6510 -5383
rect 6430 -5450 6510 -5417
rect 6580 -5223 6660 -5190
rect 6580 -5257 6603 -5223
rect 6637 -5257 6660 -5223
rect 6580 -5303 6660 -5257
rect 6580 -5337 6603 -5303
rect 6637 -5337 6660 -5303
rect 6580 -5383 6660 -5337
rect 6580 -5417 6603 -5383
rect 6637 -5417 6660 -5383
rect 6580 -5450 6660 -5417
rect 6730 -5223 6810 -5200
rect 7300 -5210 7517 -5187
rect 7551 -5210 7574 -5176
rect 6730 -5257 6753 -5223
rect 6787 -5257 6810 -5223
rect 7494 -5233 7574 -5210
rect 6730 -5303 6810 -5257
rect 6730 -5337 6753 -5303
rect 6787 -5337 6810 -5303
rect 6880 -5260 6960 -5240
rect 6880 -5263 7460 -5260
rect 6880 -5297 6903 -5263
rect 6937 -5297 7460 -5263
rect 7608 -5267 7648 -5090
rect 6880 -5300 7460 -5297
rect 6880 -5320 6960 -5300
rect 7514 -5307 7648 -5267
rect 6730 -5383 6810 -5337
rect 6730 -5417 6753 -5383
rect 6787 -5417 6810 -5383
rect 6730 -5450 6810 -5417
rect 7000 -5360 7080 -5340
rect 7132 -5360 7212 -5339
rect 7000 -5362 7460 -5360
rect 7000 -5363 7155 -5362
rect 7000 -5397 7023 -5363
rect 7057 -5396 7155 -5363
rect 7189 -5396 7460 -5362
rect 7057 -5397 7460 -5396
rect 7000 -5400 7460 -5397
rect 7000 -5420 7080 -5400
rect 7132 -5419 7212 -5400
rect 0 -5532 80 -5509
rect 0 -5566 23 -5532
rect 57 -5549 80 -5532
rect 1130 -5549 1210 -5529
rect 57 -5552 1210 -5549
rect 57 -5566 1153 -5552
rect 0 -5586 1153 -5566
rect 1187 -5586 1210 -5552
rect 0 -5589 1210 -5586
rect 1130 -5609 1210 -5589
rect 1860 -5542 1940 -5519
rect 1860 -5576 1883 -5542
rect 1917 -5576 1940 -5542
rect 1860 -5622 1940 -5576
rect 228 -5652 308 -5629
rect 228 -5686 251 -5652
rect 285 -5669 308 -5652
rect 1130 -5669 1210 -5649
rect 285 -5672 1210 -5669
rect 285 -5686 1153 -5672
rect 228 -5706 1153 -5686
rect 1187 -5706 1210 -5672
rect 228 -5709 1210 -5706
rect 1130 -5729 1210 -5709
rect 1860 -5656 1883 -5622
rect 1917 -5656 1940 -5622
rect 1860 -5702 1940 -5656
rect 1860 -5736 1883 -5702
rect 1917 -5736 1940 -5702
rect 1860 -5769 1940 -5736
rect 2010 -5542 2090 -5509
rect 2010 -5576 2033 -5542
rect 2067 -5576 2090 -5542
rect 2010 -5622 2090 -5576
rect 2010 -5656 2033 -5622
rect 2067 -5656 2090 -5622
rect 2010 -5702 2090 -5656
rect 2010 -5736 2033 -5702
rect 2067 -5736 2090 -5702
rect 2010 -5769 2090 -5736
rect 2160 -5542 2240 -5519
rect 2160 -5576 2183 -5542
rect 2217 -5576 2240 -5542
rect 2160 -5622 2240 -5576
rect 2160 -5656 2183 -5622
rect 2217 -5656 2240 -5622
rect 2160 -5702 2240 -5656
rect 2160 -5736 2183 -5702
rect 2217 -5736 2240 -5702
rect 2160 -5769 2240 -5736
rect 2310 -5542 2390 -5509
rect 2310 -5576 2333 -5542
rect 2367 -5576 2390 -5542
rect 2310 -5622 2390 -5576
rect 2310 -5656 2333 -5622
rect 2367 -5656 2390 -5622
rect 2310 -5702 2390 -5656
rect 2310 -5736 2333 -5702
rect 2367 -5736 2390 -5702
rect 2310 -5769 2390 -5736
rect 2460 -5542 2540 -5519
rect 2460 -5576 2483 -5542
rect 2517 -5576 2540 -5542
rect 2460 -5622 2540 -5576
rect 2460 -5656 2483 -5622
rect 2517 -5656 2540 -5622
rect 2460 -5702 2540 -5656
rect 3721 -5603 5101 -5580
rect 3721 -5637 3754 -5603
rect 3788 -5637 3834 -5603
rect 3868 -5637 3914 -5603
rect 3948 -5637 3994 -5603
rect 4028 -5637 4074 -5603
rect 4108 -5637 4154 -5603
rect 4188 -5637 4234 -5603
rect 4268 -5637 4314 -5603
rect 4348 -5637 4394 -5603
rect 4428 -5637 4474 -5603
rect 4508 -5637 4554 -5603
rect 4588 -5637 4634 -5603
rect 4668 -5637 4714 -5603
rect 4748 -5637 4794 -5603
rect 4828 -5637 4874 -5603
rect 4908 -5637 4954 -5603
rect 4988 -5637 5034 -5603
rect 5068 -5637 5101 -5603
rect 3721 -5660 5101 -5637
rect 2460 -5736 2483 -5702
rect 2517 -5736 2540 -5702
rect 2460 -5769 2540 -5736
rect 1130 -5789 1210 -5769
rect 798 -5792 1210 -5789
rect 798 -5812 1153 -5792
rect 798 -5846 821 -5812
rect 855 -5826 1153 -5812
rect 1187 -5826 1210 -5792
rect 855 -5829 1210 -5826
rect 855 -5846 878 -5829
rect 798 -5869 878 -5846
rect 1130 -5849 1210 -5829
rect 5135 -5826 5175 -5453
rect 5600 -5478 5680 -5455
rect 5600 -5512 5623 -5478
rect 5657 -5512 5680 -5478
rect 5600 -5535 5680 -5512
rect 6880 -5470 6960 -5450
rect 7270 -5470 7350 -5450
rect 6880 -5473 7460 -5470
rect 6880 -5507 6903 -5473
rect 6937 -5507 7293 -5473
rect 7327 -5507 7460 -5473
rect 6880 -5510 7460 -5507
rect 6880 -5530 6960 -5510
rect 7270 -5530 7350 -5510
rect 5470 -5603 7470 -5580
rect 5470 -5637 5493 -5603
rect 5527 -5637 5573 -5603
rect 5607 -5637 5653 -5603
rect 5687 -5637 5733 -5603
rect 5767 -5637 5813 -5603
rect 5847 -5637 5893 -5603
rect 5927 -5637 5973 -5603
rect 6007 -5637 6053 -5603
rect 6087 -5637 6133 -5603
rect 6167 -5637 6213 -5603
rect 6247 -5637 6293 -5603
rect 6327 -5637 6373 -5603
rect 6407 -5637 6453 -5603
rect 6487 -5637 6533 -5603
rect 6567 -5637 6613 -5603
rect 6647 -5637 6693 -5603
rect 6727 -5637 6773 -5603
rect 6807 -5637 6853 -5603
rect 6887 -5637 6933 -5603
rect 6967 -5637 7013 -5603
rect 7047 -5637 7093 -5603
rect 7127 -5637 7173 -5603
rect 7207 -5637 7253 -5603
rect 7287 -5637 7333 -5603
rect 7367 -5637 7413 -5603
rect 7447 -5637 7470 -5603
rect 5470 -5660 7470 -5637
rect 7514 -5699 7554 -5307
rect 7164 -5739 7554 -5699
rect 5458 -5826 5538 -5806
rect 5135 -5829 5538 -5826
rect 5135 -5863 5481 -5829
rect 5515 -5863 5538 -5829
rect 5135 -5866 5538 -5863
rect 5458 -5886 5538 -5866
rect 1040 -5922 3360 -5899
rect 1040 -5956 1063 -5922
rect 1097 -5956 1143 -5922
rect 1177 -5956 1223 -5922
rect 1257 -5956 1303 -5922
rect 1337 -5956 1383 -5922
rect 1417 -5956 1463 -5922
rect 1497 -5956 1543 -5922
rect 1577 -5956 1623 -5922
rect 1657 -5956 1703 -5922
rect 1737 -5956 1783 -5922
rect 1817 -5956 1863 -5922
rect 1897 -5956 1943 -5922
rect 1977 -5956 2023 -5922
rect 2057 -5956 2103 -5922
rect 2137 -5956 2183 -5922
rect 2217 -5956 2263 -5922
rect 2297 -5956 2343 -5922
rect 2377 -5956 2423 -5922
rect 2457 -5956 2503 -5922
rect 2537 -5956 2583 -5922
rect 2617 -5956 2663 -5922
rect 2697 -5956 2743 -5922
rect 2777 -5956 2823 -5922
rect 2857 -5956 2903 -5922
rect 2937 -5956 2983 -5922
rect 3017 -5956 3063 -5922
rect 3097 -5956 3143 -5922
rect 3177 -5956 3223 -5922
rect 3257 -5956 3303 -5922
rect 3337 -5956 3360 -5922
rect 1040 -6063 3360 -5956
rect 1040 -6097 1063 -6063
rect 1097 -6097 1143 -6063
rect 1177 -6097 1223 -6063
rect 1257 -6097 1303 -6063
rect 1337 -6097 1383 -6063
rect 1417 -6097 1463 -6063
rect 1497 -6097 1543 -6063
rect 1577 -6097 1623 -6063
rect 1657 -6097 1703 -6063
rect 1737 -6097 1783 -6063
rect 1817 -6097 1863 -6063
rect 1897 -6097 1943 -6063
rect 1977 -6097 2023 -6063
rect 2057 -6097 2103 -6063
rect 2137 -6097 2183 -6063
rect 2217 -6097 2263 -6063
rect 2297 -6097 2343 -6063
rect 2377 -6097 2423 -6063
rect 2457 -6097 2503 -6063
rect 2537 -6097 2583 -6063
rect 2617 -6097 2663 -6063
rect 2697 -6097 2743 -6063
rect 2777 -6097 2823 -6063
rect 2857 -6097 2903 -6063
rect 2937 -6097 2983 -6063
rect 3017 -6097 3063 -6063
rect 3097 -6097 3143 -6063
rect 3177 -6097 3223 -6063
rect 3257 -6097 3303 -6063
rect 3337 -6097 3360 -6063
rect 1040 -6120 3360 -6097
rect 3720 -6063 5100 -6040
rect 3720 -6097 3753 -6063
rect 3787 -6097 3833 -6063
rect 3867 -6097 3913 -6063
rect 3947 -6097 3993 -6063
rect 4027 -6097 4073 -6063
rect 4107 -6097 4153 -6063
rect 4187 -6097 4233 -6063
rect 4267 -6097 4313 -6063
rect 4347 -6097 4393 -6063
rect 4427 -6097 4473 -6063
rect 4507 -6097 4553 -6063
rect 4587 -6097 4633 -6063
rect 4667 -6097 4713 -6063
rect 4747 -6097 4793 -6063
rect 4827 -6097 4873 -6063
rect 4907 -6097 4953 -6063
rect 4987 -6097 5033 -6063
rect 5067 -6097 5100 -6063
rect 3720 -6120 5100 -6097
rect 5449 -6063 7129 -6040
rect 5449 -6097 5472 -6063
rect 5506 -6097 5552 -6063
rect 5586 -6097 5632 -6063
rect 5666 -6097 5712 -6063
rect 5746 -6097 5792 -6063
rect 5826 -6097 5872 -6063
rect 5906 -6097 5952 -6063
rect 5986 -6097 6032 -6063
rect 6066 -6097 6112 -6063
rect 6146 -6097 6192 -6063
rect 6226 -6097 6272 -6063
rect 6306 -6097 6352 -6063
rect 6386 -6097 6432 -6063
rect 6466 -6097 6512 -6063
rect 6546 -6097 6592 -6063
rect 6626 -6097 6672 -6063
rect 6706 -6097 6752 -6063
rect 6786 -6097 6832 -6063
rect 6866 -6097 6912 -6063
rect 6946 -6097 6992 -6063
rect 7026 -6097 7072 -6063
rect 7106 -6097 7129 -6063
rect 5449 -6120 7129 -6097
rect 228 -6173 308 -6150
rect 228 -6207 251 -6173
rect 285 -6190 308 -6173
rect 1450 -6190 1530 -6170
rect 1580 -6190 1660 -6170
rect 285 -6193 1660 -6190
rect 285 -6207 1473 -6193
rect 228 -6227 1473 -6207
rect 1507 -6227 1603 -6193
rect 1637 -6227 1660 -6193
rect 228 -6230 1660 -6227
rect 1450 -6250 1530 -6230
rect 1580 -6250 1660 -6230
rect 2840 -6193 2920 -6170
rect 2840 -6227 2863 -6193
rect 2897 -6227 2920 -6193
rect 2840 -6250 2920 -6227
rect 342 -6287 422 -6264
rect 342 -6321 365 -6287
rect 399 -6290 422 -6287
rect 1330 -6290 1410 -6270
rect 1710 -6290 1790 -6270
rect 399 -6293 1790 -6290
rect 399 -6321 1353 -6293
rect 342 -6327 1353 -6321
rect 1387 -6327 1733 -6293
rect 1767 -6327 1790 -6293
rect 342 -6330 1790 -6327
rect 342 -6344 422 -6330
rect 1330 -6350 1410 -6330
rect 1710 -6350 1790 -6330
rect 1860 -6283 1940 -6250
rect 1860 -6317 1883 -6283
rect 1917 -6317 1940 -6283
rect 1860 -6363 1940 -6317
rect 0 -6390 80 -6371
rect 1580 -6390 1660 -6370
rect 0 -6393 1660 -6390
rect 0 -6394 1603 -6393
rect 0 -6428 23 -6394
rect 57 -6427 1603 -6394
rect 1637 -6427 1660 -6393
rect 57 -6428 1660 -6427
rect 0 -6430 1660 -6428
rect 0 -6451 80 -6430
rect 1580 -6450 1660 -6430
rect 1860 -6397 1883 -6363
rect 1917 -6397 1940 -6363
rect 1860 -6443 1940 -6397
rect 1130 -6490 1210 -6470
rect 1710 -6490 1790 -6470
rect 114 -6493 1790 -6490
rect 114 -6513 1153 -6493
rect 114 -6547 137 -6513
rect 171 -6527 1153 -6513
rect 1187 -6527 1733 -6493
rect 1767 -6527 1790 -6493
rect 1860 -6477 1883 -6443
rect 1917 -6477 1940 -6443
rect 1860 -6500 1940 -6477
rect 2010 -6283 2090 -6250
rect 2010 -6317 2033 -6283
rect 2067 -6317 2090 -6283
rect 2010 -6363 2090 -6317
rect 2010 -6397 2033 -6363
rect 2067 -6397 2090 -6363
rect 2010 -6443 2090 -6397
rect 2010 -6477 2033 -6443
rect 2067 -6477 2090 -6443
rect 2010 -6510 2090 -6477
rect 2160 -6283 2240 -6250
rect 2160 -6317 2183 -6283
rect 2217 -6317 2240 -6283
rect 2160 -6363 2240 -6317
rect 2160 -6397 2183 -6363
rect 2217 -6397 2240 -6363
rect 2160 -6443 2240 -6397
rect 2160 -6477 2183 -6443
rect 2217 -6477 2240 -6443
rect 2160 -6500 2240 -6477
rect 2310 -6283 2390 -6250
rect 2310 -6317 2333 -6283
rect 2367 -6317 2390 -6283
rect 2310 -6363 2390 -6317
rect 2310 -6397 2333 -6363
rect 2367 -6397 2390 -6363
rect 2310 -6443 2390 -6397
rect 2310 -6477 2333 -6443
rect 2367 -6477 2390 -6443
rect 2310 -6510 2390 -6477
rect 2460 -6283 2540 -6250
rect 2460 -6317 2483 -6283
rect 2517 -6317 2540 -6283
rect 2460 -6363 2540 -6317
rect 3040 -6293 3120 -6270
rect 3632 -6290 3712 -6270
rect 3040 -6327 3063 -6293
rect 3097 -6327 3120 -6293
rect 3040 -6350 3120 -6327
rect 3479 -6293 3712 -6290
rect 3479 -6327 3655 -6293
rect 3689 -6327 3712 -6293
rect 3479 -6330 3712 -6327
rect 2460 -6397 2483 -6363
rect 2517 -6397 2540 -6363
rect 2460 -6443 2540 -6397
rect 2460 -6477 2483 -6443
rect 2517 -6477 2540 -6443
rect 3190 -6393 3270 -6370
rect 3190 -6427 3213 -6393
rect 3247 -6427 3270 -6393
rect 3190 -6450 3270 -6427
rect 2460 -6500 2540 -6477
rect 2740 -6493 2820 -6470
rect 171 -6530 1790 -6527
rect 171 -6547 194 -6530
rect 114 -6570 194 -6547
rect 1130 -6550 1210 -6530
rect 1710 -6550 1790 -6530
rect 2030 -6560 2070 -6510
rect 2210 -6560 2290 -6540
rect 2030 -6563 2290 -6560
rect 2030 -6597 2233 -6563
rect 2267 -6597 2290 -6563
rect 2030 -6600 2290 -6597
rect 2030 -6730 2070 -6600
rect 2210 -6620 2290 -6600
rect 1100 -6770 2070 -6730
rect 2110 -6680 2190 -6665
rect 2330 -6680 2370 -6510
rect 2740 -6527 2763 -6493
rect 2797 -6527 2820 -6493
rect 2740 -6550 2820 -6527
rect 2580 -6573 2660 -6550
rect 2580 -6607 2603 -6573
rect 2637 -6590 2660 -6573
rect 3340 -6573 3420 -6550
rect 3340 -6590 3363 -6573
rect 2637 -6607 3363 -6590
rect 3397 -6607 3420 -6573
rect 2580 -6630 3420 -6607
rect 3479 -6680 3519 -6330
rect 3632 -6350 3712 -6330
rect 4070 -6283 4150 -6250
rect 4070 -6317 4093 -6283
rect 4127 -6317 4150 -6283
rect 4070 -6363 4150 -6317
rect 4070 -6397 4093 -6363
rect 4127 -6397 4150 -6363
rect 3920 -6440 4000 -6420
rect 3720 -6443 4000 -6440
rect 3720 -6477 3943 -6443
rect 3977 -6477 4000 -6443
rect 3720 -6480 4000 -6477
rect 3920 -6500 4000 -6480
rect 4070 -6443 4150 -6397
rect 4070 -6477 4093 -6443
rect 4127 -6477 4150 -6443
rect 4070 -6500 4150 -6477
rect 4220 -6283 4300 -6250
rect 4220 -6317 4243 -6283
rect 4277 -6317 4300 -6283
rect 4220 -6363 4300 -6317
rect 4220 -6397 4243 -6363
rect 4277 -6397 4300 -6363
rect 4220 -6443 4300 -6397
rect 4220 -6477 4243 -6443
rect 4277 -6477 4300 -6443
rect 4220 -6510 4300 -6477
rect 4370 -6283 4450 -6250
rect 4370 -6317 4393 -6283
rect 4427 -6317 4450 -6283
rect 4370 -6363 4450 -6317
rect 4370 -6397 4393 -6363
rect 4427 -6397 4450 -6363
rect 4370 -6443 4450 -6397
rect 4370 -6477 4393 -6443
rect 4427 -6477 4450 -6443
rect 4370 -6500 4450 -6477
rect 4520 -6283 4600 -6250
rect 4520 -6317 4543 -6283
rect 4577 -6317 4600 -6283
rect 4520 -6363 4600 -6317
rect 4520 -6397 4543 -6363
rect 4577 -6397 4600 -6363
rect 4520 -6443 4600 -6397
rect 4520 -6477 4543 -6443
rect 4577 -6477 4600 -6443
rect 4520 -6510 4600 -6477
rect 4670 -6283 4750 -6250
rect 4670 -6317 4693 -6283
rect 4727 -6317 4750 -6283
rect 4670 -6363 4750 -6317
rect 4820 -6290 4900 -6270
rect 5799 -6290 5879 -6270
rect 4820 -6293 5879 -6290
rect 4820 -6327 4843 -6293
rect 4877 -6327 5822 -6293
rect 5856 -6327 5879 -6293
rect 4820 -6330 5879 -6327
rect 4820 -6350 4900 -6330
rect 5799 -6350 5879 -6330
rect 5949 -6283 6029 -6250
rect 5949 -6317 5972 -6283
rect 6006 -6317 6029 -6283
rect 4670 -6397 4693 -6363
rect 4727 -6397 4750 -6363
rect 5949 -6363 6029 -6317
rect 4670 -6443 4750 -6397
rect 5370 -6393 5450 -6370
rect 4670 -6477 4693 -6443
rect 4727 -6477 4750 -6443
rect 4670 -6500 4750 -6477
rect 4820 -6440 4900 -6420
rect 4950 -6440 5030 -6420
rect 4820 -6443 5030 -6440
rect 4820 -6477 4843 -6443
rect 4877 -6477 4973 -6443
rect 5007 -6477 5030 -6443
rect 5370 -6427 5393 -6393
rect 5427 -6410 5450 -6393
rect 5799 -6410 5879 -6390
rect 5427 -6413 5879 -6410
rect 5427 -6427 5822 -6413
rect 5370 -6447 5822 -6427
rect 5856 -6447 5879 -6413
rect 5370 -6450 5879 -6447
rect 5799 -6470 5879 -6450
rect 5949 -6397 5972 -6363
rect 6006 -6397 6029 -6363
rect 5949 -6443 6029 -6397
rect 4820 -6480 5030 -6477
rect 4820 -6500 4900 -6480
rect 4950 -6500 5030 -6480
rect 5949 -6477 5972 -6443
rect 6006 -6477 6029 -6443
rect 5370 -6510 5450 -6490
rect 5669 -6510 5749 -6490
rect 5949 -6500 6029 -6477
rect 6099 -6283 6179 -6250
rect 6099 -6317 6122 -6283
rect 6156 -6317 6179 -6283
rect 6099 -6363 6179 -6317
rect 6099 -6397 6122 -6363
rect 6156 -6397 6179 -6363
rect 6099 -6443 6179 -6397
rect 6099 -6477 6122 -6443
rect 6156 -6477 6179 -6443
rect 6099 -6510 6179 -6477
rect 6249 -6283 6329 -6250
rect 6249 -6317 6272 -6283
rect 6306 -6317 6329 -6283
rect 6249 -6363 6329 -6317
rect 6249 -6397 6272 -6363
rect 6306 -6397 6329 -6363
rect 6249 -6443 6329 -6397
rect 6249 -6477 6272 -6443
rect 6306 -6477 6329 -6443
rect 6249 -6500 6329 -6477
rect 6399 -6283 6479 -6250
rect 6399 -6317 6422 -6283
rect 6456 -6317 6479 -6283
rect 6399 -6363 6479 -6317
rect 6399 -6397 6422 -6363
rect 6456 -6397 6479 -6363
rect 6399 -6443 6479 -6397
rect 6399 -6477 6422 -6443
rect 6456 -6477 6479 -6443
rect 6399 -6510 6479 -6477
rect 6549 -6283 6629 -6250
rect 6549 -6317 6572 -6283
rect 6606 -6317 6629 -6283
rect 6549 -6363 6629 -6317
rect 6929 -6293 7009 -6270
rect 6929 -6327 6952 -6293
rect 6986 -6327 7009 -6293
rect 6929 -6350 7009 -6327
rect 6549 -6397 6572 -6363
rect 6606 -6397 6629 -6363
rect 6549 -6443 6629 -6397
rect 6549 -6477 6572 -6443
rect 6606 -6477 6629 -6443
rect 6779 -6413 6859 -6390
rect 6779 -6447 6802 -6413
rect 6836 -6447 6859 -6413
rect 6779 -6470 6859 -6447
rect 6549 -6500 6629 -6477
rect 4240 -6560 4280 -6510
rect 4420 -6560 4500 -6540
rect 4240 -6563 4500 -6560
rect 4240 -6597 4443 -6563
rect 4477 -6597 4500 -6563
rect 4240 -6600 4500 -6597
rect 3790 -6680 3870 -6660
rect 2110 -6688 3519 -6680
rect 2110 -6722 2133 -6688
rect 2167 -6720 3519 -6688
rect 3666 -6683 3870 -6680
rect 3666 -6717 3813 -6683
rect 3847 -6717 3870 -6683
rect 3666 -6720 3870 -6717
rect 2167 -6722 2190 -6720
rect 2110 -6745 2190 -6722
rect 1100 -6810 1140 -6770
rect 1700 -6810 1740 -6770
rect 2030 -6810 2070 -6770
rect 2330 -6810 2370 -6720
rect 2660 -6810 2700 -6720
rect 3260 -6810 3300 -6720
rect 1080 -6843 1160 -6810
rect 1080 -6877 1103 -6843
rect 1137 -6877 1160 -6843
rect 1080 -6923 1160 -6877
rect 1080 -6957 1103 -6923
rect 1137 -6957 1160 -6923
rect 1080 -7003 1160 -6957
rect 1080 -7037 1103 -7003
rect 1137 -7037 1160 -7003
rect 1080 -7060 1160 -7037
rect 1380 -6843 1460 -6810
rect 1380 -6877 1403 -6843
rect 1437 -6877 1460 -6843
rect 1380 -6923 1460 -6877
rect 1380 -6957 1403 -6923
rect 1437 -6957 1460 -6923
rect 1380 -7003 1460 -6957
rect 1380 -7037 1403 -7003
rect 1437 -7037 1460 -7003
rect 1380 -7060 1460 -7037
rect 1680 -6843 1760 -6810
rect 1680 -6877 1703 -6843
rect 1737 -6877 1760 -6843
rect 1680 -6923 1760 -6877
rect 1680 -6957 1703 -6923
rect 1737 -6957 1760 -6923
rect 1680 -7003 1760 -6957
rect 1680 -7037 1703 -7003
rect 1737 -7037 1760 -7003
rect 1680 -7060 1760 -7037
rect 1860 -6843 1940 -6810
rect 1860 -6877 1883 -6843
rect 1917 -6877 1940 -6843
rect 1860 -6923 1940 -6877
rect 1860 -6957 1883 -6923
rect 1917 -6957 1940 -6923
rect 1860 -7003 1940 -6957
rect 1860 -7037 1883 -7003
rect 1917 -7037 1940 -7003
rect 1860 -7060 1940 -7037
rect 2010 -6843 2090 -6810
rect 2010 -6877 2033 -6843
rect 2067 -6877 2090 -6843
rect 2010 -6923 2090 -6877
rect 2010 -6957 2033 -6923
rect 2067 -6957 2090 -6923
rect 2010 -7003 2090 -6957
rect 2010 -7037 2033 -7003
rect 2067 -7037 2090 -7003
rect 2010 -7060 2090 -7037
rect 2160 -6843 2240 -6810
rect 2160 -6877 2183 -6843
rect 2217 -6877 2240 -6843
rect 2160 -6923 2240 -6877
rect 2160 -6957 2183 -6923
rect 2217 -6957 2240 -6923
rect 2160 -7003 2240 -6957
rect 2160 -7037 2183 -7003
rect 2217 -7037 2240 -7003
rect 2160 -7060 2240 -7037
rect 2310 -6843 2390 -6810
rect 2310 -6877 2333 -6843
rect 2367 -6877 2390 -6843
rect 2310 -6923 2390 -6877
rect 2310 -6957 2333 -6923
rect 2367 -6957 2390 -6923
rect 2310 -7003 2390 -6957
rect 2310 -7037 2333 -7003
rect 2367 -7037 2390 -7003
rect 2310 -7060 2390 -7037
rect 2460 -6843 2540 -6810
rect 2460 -6877 2483 -6843
rect 2517 -6877 2540 -6843
rect 2460 -6923 2540 -6877
rect 2460 -6957 2483 -6923
rect 2517 -6957 2540 -6923
rect 2460 -7003 2540 -6957
rect 2460 -7037 2483 -7003
rect 2517 -7037 2540 -7003
rect 2460 -7060 2540 -7037
rect 2640 -6843 2720 -6810
rect 2640 -6877 2663 -6843
rect 2697 -6877 2720 -6843
rect 2640 -6923 2720 -6877
rect 2640 -6957 2663 -6923
rect 2697 -6957 2720 -6923
rect 2640 -7003 2720 -6957
rect 2640 -7037 2663 -7003
rect 2697 -7037 2720 -7003
rect 2640 -7060 2720 -7037
rect 2940 -6843 3020 -6810
rect 2940 -6877 2963 -6843
rect 2997 -6877 3020 -6843
rect 2940 -6923 3020 -6877
rect 2940 -6957 2963 -6923
rect 2997 -6957 3020 -6923
rect 2940 -7003 3020 -6957
rect 2940 -7037 2963 -7003
rect 2997 -7037 3020 -7003
rect 2940 -7060 3020 -7037
rect 3240 -6843 3320 -6810
rect 3240 -6877 3263 -6843
rect 3297 -6877 3320 -6843
rect 3240 -6923 3320 -6877
rect 3240 -6957 3263 -6923
rect 3297 -6957 3320 -6923
rect 3240 -7003 3320 -6957
rect 3354 -6920 3434 -6899
rect 3666 -6920 3706 -6720
rect 3790 -6740 3870 -6720
rect 4240 -6730 4280 -6600
rect 4420 -6620 4500 -6600
rect 3910 -6770 4280 -6730
rect 4320 -6680 4400 -6665
rect 4540 -6680 4580 -6510
rect 5370 -6513 5749 -6510
rect 4820 -6560 4900 -6540
rect 5370 -6547 5393 -6513
rect 5427 -6547 5692 -6513
rect 5726 -6547 5749 -6513
rect 5370 -6550 5749 -6547
rect 4820 -6563 5269 -6560
rect 4820 -6597 4843 -6563
rect 4877 -6597 5269 -6563
rect 5370 -6570 5450 -6550
rect 5669 -6570 5749 -6550
rect 6119 -6560 6159 -6510
rect 6299 -6560 6379 -6540
rect 6119 -6563 6379 -6560
rect 4820 -6600 5269 -6597
rect 4820 -6620 4900 -6600
rect 5229 -6610 5269 -6600
rect 5519 -6610 5599 -6590
rect 5229 -6613 5599 -6610
rect 5229 -6647 5542 -6613
rect 5576 -6647 5599 -6613
rect 5229 -6650 5599 -6647
rect 5519 -6670 5599 -6650
rect 6119 -6597 6322 -6563
rect 6356 -6597 6379 -6563
rect 6119 -6600 6379 -6597
rect 4320 -6688 4580 -6680
rect 4320 -6722 4343 -6688
rect 4377 -6720 4580 -6688
rect 4377 -6722 4400 -6720
rect 4320 -6745 4400 -6722
rect 4540 -6730 4580 -6720
rect 5108 -6730 5188 -6710
rect 6119 -6730 6159 -6600
rect 6299 -6620 6379 -6600
rect 4540 -6733 5188 -6730
rect 4540 -6767 5131 -6733
rect 5165 -6767 5188 -6733
rect 4540 -6770 5188 -6767
rect 3910 -6810 3950 -6770
rect 4240 -6810 4280 -6770
rect 3354 -6923 3706 -6920
rect 3354 -6957 3377 -6923
rect 3411 -6957 3706 -6923
rect 3354 -6960 3706 -6957
rect 3740 -6843 3820 -6810
rect 3740 -6877 3763 -6843
rect 3797 -6877 3820 -6843
rect 3740 -6923 3820 -6877
rect 3740 -6957 3763 -6923
rect 3797 -6957 3820 -6923
rect 3354 -6979 3434 -6960
rect 3240 -7037 3263 -7003
rect 3297 -7037 3320 -7003
rect 3240 -7060 3320 -7037
rect 3740 -7003 3820 -6957
rect 3740 -7037 3763 -7003
rect 3797 -7037 3820 -7003
rect 3740 -7060 3820 -7037
rect 3890 -6843 3970 -6810
rect 3890 -6877 3913 -6843
rect 3947 -6877 3970 -6843
rect 3890 -6923 3970 -6877
rect 3890 -6957 3913 -6923
rect 3947 -6957 3970 -6923
rect 3890 -7003 3970 -6957
rect 3890 -7037 3913 -7003
rect 3947 -7037 3970 -7003
rect 3890 -7060 3970 -7037
rect 4070 -6843 4150 -6810
rect 4070 -6877 4093 -6843
rect 4127 -6877 4150 -6843
rect 4070 -6923 4150 -6877
rect 4070 -6957 4093 -6923
rect 4127 -6957 4150 -6923
rect 4070 -7003 4150 -6957
rect 4070 -7037 4093 -7003
rect 4127 -7037 4150 -7003
rect 4070 -7060 4150 -7037
rect 4220 -6843 4300 -6810
rect 4220 -6877 4243 -6843
rect 4277 -6877 4300 -6843
rect 4220 -6923 4300 -6877
rect 4220 -6957 4243 -6923
rect 4277 -6957 4300 -6923
rect 4220 -7003 4300 -6957
rect 4220 -7037 4243 -7003
rect 4277 -7037 4300 -7003
rect 4220 -7060 4300 -7037
rect 4370 -6843 4450 -6810
rect 4370 -6877 4393 -6843
rect 4427 -6877 4450 -6843
rect 4370 -6923 4450 -6877
rect 4370 -6957 4393 -6923
rect 4427 -6957 4450 -6923
rect 4370 -7003 4450 -6957
rect 4370 -7037 4393 -7003
rect 4427 -7037 4450 -7003
rect 4370 -7060 4450 -7037
rect 4520 -6843 4600 -6770
rect 4870 -6810 4910 -6770
rect 5108 -6790 5188 -6770
rect 5489 -6770 6159 -6730
rect 6199 -6680 6279 -6665
rect 6419 -6680 6459 -6510
rect 6699 -6560 6779 -6540
rect 7164 -6560 7204 -5739
rect 7494 -5794 7574 -5774
rect 6699 -6563 7204 -6560
rect 6699 -6597 6722 -6563
rect 6756 -6597 7204 -6563
rect 6699 -6600 7204 -6597
rect 7282 -5797 7574 -5794
rect 7282 -5831 7517 -5797
rect 7551 -5831 7574 -5797
rect 7282 -5834 7574 -5831
rect 6699 -6620 6779 -6600
rect 7129 -6680 7209 -6660
rect 6199 -6683 7209 -6680
rect 6199 -6688 7152 -6683
rect 6199 -6722 6222 -6688
rect 6256 -6717 7152 -6688
rect 7186 -6717 7209 -6683
rect 6256 -6720 7209 -6717
rect 6256 -6722 6279 -6720
rect 6199 -6745 6279 -6722
rect 5489 -6810 5529 -6770
rect 5789 -6810 5829 -6770
rect 6120 -6810 6159 -6770
rect 6419 -6810 6459 -6720
rect 6749 -6810 6789 -6720
rect 7129 -6740 7209 -6720
rect 4520 -6877 4543 -6843
rect 4577 -6877 4600 -6843
rect 4520 -6923 4600 -6877
rect 4520 -6957 4543 -6923
rect 4577 -6957 4600 -6923
rect 4520 -7003 4600 -6957
rect 4520 -7037 4543 -7003
rect 4577 -7037 4600 -7003
rect 4520 -7060 4600 -7037
rect 4670 -6843 4750 -6810
rect 4670 -6877 4693 -6843
rect 4727 -6877 4750 -6843
rect 4670 -6923 4750 -6877
rect 4670 -6957 4693 -6923
rect 4727 -6957 4750 -6923
rect 4670 -7003 4750 -6957
rect 4670 -7037 4693 -7003
rect 4727 -7037 4750 -7003
rect 4670 -7060 4750 -7037
rect 4850 -6843 4930 -6810
rect 4850 -6877 4873 -6843
rect 4907 -6877 4930 -6843
rect 4850 -6923 4930 -6877
rect 4850 -6957 4873 -6923
rect 4907 -6957 4930 -6923
rect 4850 -7003 4930 -6957
rect 4850 -7037 4873 -7003
rect 4907 -7037 4930 -7003
rect 4850 -7060 4930 -7037
rect 5000 -6843 5080 -6810
rect 5000 -6877 5023 -6843
rect 5057 -6877 5080 -6843
rect 5000 -6923 5080 -6877
rect 5000 -6957 5023 -6923
rect 5057 -6957 5080 -6923
rect 5000 -7003 5080 -6957
rect 5000 -7037 5023 -7003
rect 5057 -7037 5080 -7003
rect 5000 -7060 5080 -7037
rect 5469 -6843 5549 -6810
rect 5469 -6877 5492 -6843
rect 5526 -6877 5549 -6843
rect 5469 -6923 5549 -6877
rect 5469 -6957 5492 -6923
rect 5526 -6957 5549 -6923
rect 5469 -7003 5549 -6957
rect 5469 -7037 5492 -7003
rect 5526 -7037 5549 -7003
rect 5469 -7060 5549 -7037
rect 5619 -6843 5699 -6810
rect 5619 -6877 5642 -6843
rect 5676 -6877 5699 -6843
rect 5619 -6923 5699 -6877
rect 5619 -6957 5642 -6923
rect 5676 -6957 5699 -6923
rect 5619 -7003 5699 -6957
rect 5619 -7037 5642 -7003
rect 5676 -7037 5699 -7003
rect 5619 -7060 5699 -7037
rect 5769 -6843 5849 -6810
rect 5769 -6877 5792 -6843
rect 5826 -6877 5849 -6843
rect 5769 -6923 5849 -6877
rect 5769 -6957 5792 -6923
rect 5826 -6957 5849 -6923
rect 5769 -7003 5849 -6957
rect 5769 -7037 5792 -7003
rect 5826 -7037 5849 -7003
rect 5769 -7060 5849 -7037
rect 5949 -6843 6029 -6810
rect 5949 -6877 5972 -6843
rect 6006 -6877 6029 -6843
rect 5949 -6923 6029 -6877
rect 5949 -6957 5972 -6923
rect 6006 -6957 6029 -6923
rect 5949 -7003 6029 -6957
rect 5949 -7037 5972 -7003
rect 6006 -7037 6029 -7003
rect 5949 -7060 6029 -7037
rect 6099 -6843 6179 -6810
rect 6099 -6877 6122 -6843
rect 6156 -6877 6179 -6843
rect 6099 -6923 6179 -6877
rect 6099 -6957 6122 -6923
rect 6156 -6957 6179 -6923
rect 6099 -7003 6179 -6957
rect 6099 -7037 6122 -7003
rect 6156 -7037 6179 -7003
rect 6099 -7060 6179 -7037
rect 6249 -6843 6329 -6810
rect 6249 -6877 6272 -6843
rect 6306 -6877 6329 -6843
rect 6249 -6923 6329 -6877
rect 6249 -6957 6272 -6923
rect 6306 -6957 6329 -6923
rect 6249 -7003 6329 -6957
rect 6249 -7037 6272 -7003
rect 6306 -7037 6329 -7003
rect 6249 -7060 6329 -7037
rect 6399 -6843 6479 -6810
rect 6399 -6877 6422 -6843
rect 6456 -6877 6479 -6843
rect 6399 -6923 6479 -6877
rect 6399 -6957 6422 -6923
rect 6456 -6957 6479 -6923
rect 6399 -7003 6479 -6957
rect 6399 -7037 6422 -7003
rect 6456 -7037 6479 -7003
rect 6399 -7060 6479 -7037
rect 6549 -6843 6629 -6810
rect 6549 -6877 6572 -6843
rect 6606 -6877 6629 -6843
rect 6549 -6923 6629 -6877
rect 6549 -6957 6572 -6923
rect 6606 -6957 6629 -6923
rect 6549 -7003 6629 -6957
rect 6549 -7037 6572 -7003
rect 6606 -7037 6629 -7003
rect 6549 -7060 6629 -7037
rect 6729 -6843 6809 -6810
rect 6729 -6877 6752 -6843
rect 6786 -6877 6809 -6843
rect 6729 -6923 6809 -6877
rect 6729 -6957 6752 -6923
rect 6786 -6957 6809 -6923
rect 6729 -7003 6809 -6957
rect 6729 -7037 6752 -7003
rect 6786 -7037 6809 -7003
rect 6729 -7060 6809 -7037
rect 7029 -6843 7109 -6810
rect 7029 -6877 7052 -6843
rect 7086 -6877 7109 -6843
rect 7029 -6923 7109 -6877
rect 7029 -6957 7052 -6923
rect 7086 -6957 7109 -6923
rect 7029 -7003 7109 -6957
rect 7029 -7037 7052 -7003
rect 7086 -7037 7109 -7003
rect 7029 -7060 7109 -7037
rect 1492 -7120 1572 -7100
rect 1960 -7120 2040 -7100
rect 2360 -7120 2440 -7100
rect 4170 -7120 4250 -7100
rect 4570 -7120 4650 -7100
rect 5456 -7120 5536 -7100
rect 6049 -7120 6129 -7100
rect 6449 -7120 6529 -7100
rect 1060 -7123 4650 -7120
rect 1060 -7157 1515 -7123
rect 1549 -7157 1983 -7123
rect 2017 -7157 2383 -7123
rect 2417 -7157 4193 -7123
rect 4227 -7157 4593 -7123
rect 4627 -7157 4650 -7123
rect 1060 -7160 4650 -7157
rect 5449 -7123 6529 -7120
rect 5449 -7157 5479 -7123
rect 5513 -7157 6072 -7123
rect 6106 -7157 6472 -7123
rect 6506 -7157 6529 -7123
rect 5449 -7160 6529 -7157
rect 1492 -7180 1572 -7160
rect 1960 -7180 2040 -7160
rect 2360 -7180 2440 -7160
rect 4170 -7180 4250 -7160
rect 4570 -7180 4650 -7160
rect 5456 -7180 5536 -7160
rect 6049 -7180 6129 -7160
rect 6449 -7180 6529 -7160
rect 912 -7243 3340 -7220
rect 912 -7277 935 -7243
rect 969 -7277 1143 -7243
rect 1177 -7277 1223 -7243
rect 1257 -7277 1303 -7243
rect 1337 -7277 1383 -7243
rect 1417 -7277 1463 -7243
rect 1497 -7277 1543 -7243
rect 1577 -7277 1623 -7243
rect 1657 -7277 1703 -7243
rect 1737 -7277 1783 -7243
rect 1817 -7277 1863 -7243
rect 1897 -7277 1943 -7243
rect 1977 -7277 2023 -7243
rect 2057 -7277 2103 -7243
rect 2137 -7277 2183 -7243
rect 2217 -7277 2263 -7243
rect 2297 -7277 2343 -7243
rect 2377 -7277 2423 -7243
rect 2457 -7277 2503 -7243
rect 2537 -7277 2583 -7243
rect 2617 -7277 2663 -7243
rect 2697 -7277 2743 -7243
rect 2777 -7277 2823 -7243
rect 2857 -7277 2903 -7243
rect 2937 -7277 2983 -7243
rect 3017 -7277 3063 -7243
rect 3097 -7277 3143 -7243
rect 3177 -7277 3223 -7243
rect 3257 -7277 3340 -7243
rect 912 -7300 3340 -7277
rect 3720 -7243 5100 -7220
rect 3720 -7277 3753 -7243
rect 3787 -7277 3833 -7243
rect 3867 -7277 3913 -7243
rect 3947 -7277 3993 -7243
rect 4027 -7277 4073 -7243
rect 4107 -7277 4153 -7243
rect 4187 -7277 4233 -7243
rect 4267 -7277 4313 -7243
rect 4347 -7277 4393 -7243
rect 4427 -7277 4473 -7243
rect 4507 -7277 4553 -7243
rect 4587 -7277 4633 -7243
rect 4667 -7277 4713 -7243
rect 4747 -7277 4793 -7243
rect 4827 -7277 4873 -7243
rect 4907 -7277 4953 -7243
rect 4987 -7277 5033 -7243
rect 5067 -7277 5100 -7243
rect 3720 -7300 5100 -7277
rect 5449 -7243 7129 -7220
rect 5449 -7277 5472 -7243
rect 5506 -7277 5552 -7243
rect 5586 -7277 5632 -7243
rect 5666 -7277 5712 -7243
rect 5746 -7277 5792 -7243
rect 5826 -7277 5872 -7243
rect 5906 -7277 5952 -7243
rect 5986 -7277 6032 -7243
rect 6066 -7277 6112 -7243
rect 6146 -7277 6192 -7243
rect 6226 -7277 6272 -7243
rect 6306 -7277 6352 -7243
rect 6386 -7277 6432 -7243
rect 6466 -7277 6512 -7243
rect 6546 -7277 6592 -7243
rect 6626 -7277 6672 -7243
rect 6706 -7277 6752 -7243
rect 6786 -7277 6832 -7243
rect 6866 -7277 6912 -7243
rect 6946 -7277 6992 -7243
rect 7026 -7277 7072 -7243
rect 7106 -7277 7129 -7243
rect 5449 -7300 7129 -7277
rect 1492 -7360 1572 -7340
rect 1960 -7360 2040 -7340
rect 2360 -7360 2440 -7340
rect 4170 -7360 4250 -7340
rect 4570 -7360 4650 -7340
rect 5458 -7360 5538 -7340
rect 6049 -7360 6129 -7340
rect 6449 -7360 6529 -7340
rect 1060 -7363 4650 -7360
rect 1060 -7397 1515 -7363
rect 1549 -7397 1983 -7363
rect 2017 -7397 2383 -7363
rect 2417 -7397 4193 -7363
rect 4227 -7397 4593 -7363
rect 4627 -7397 4650 -7363
rect 1060 -7400 4650 -7397
rect 5449 -7363 6529 -7360
rect 5449 -7397 5481 -7363
rect 5515 -7397 6072 -7363
rect 6106 -7397 6472 -7363
rect 6506 -7397 6529 -7363
rect 5449 -7400 6529 -7397
rect 1492 -7420 1572 -7400
rect 1960 -7420 2040 -7400
rect 2360 -7420 2440 -7400
rect 4170 -7420 4250 -7400
rect 4570 -7420 4650 -7400
rect 5458 -7420 5538 -7400
rect 6049 -7420 6129 -7400
rect 6449 -7420 6529 -7400
rect 1080 -7483 1160 -7460
rect 1080 -7517 1103 -7483
rect 1137 -7517 1160 -7483
rect 1080 -7563 1160 -7517
rect 1080 -7597 1103 -7563
rect 1137 -7597 1160 -7563
rect 1080 -7643 1160 -7597
rect 1080 -7677 1103 -7643
rect 1137 -7677 1160 -7643
rect 1080 -7710 1160 -7677
rect 1380 -7483 1460 -7460
rect 1380 -7517 1403 -7483
rect 1437 -7517 1460 -7483
rect 1380 -7563 1460 -7517
rect 1380 -7597 1403 -7563
rect 1437 -7597 1460 -7563
rect 1380 -7643 1460 -7597
rect 1380 -7677 1403 -7643
rect 1437 -7677 1460 -7643
rect 1380 -7710 1460 -7677
rect 1680 -7483 1760 -7460
rect 1680 -7517 1703 -7483
rect 1737 -7517 1760 -7483
rect 1680 -7563 1760 -7517
rect 1680 -7597 1703 -7563
rect 1737 -7597 1760 -7563
rect 1680 -7643 1760 -7597
rect 1680 -7677 1703 -7643
rect 1737 -7677 1760 -7643
rect 1680 -7710 1760 -7677
rect 1860 -7483 1940 -7460
rect 1860 -7517 1883 -7483
rect 1917 -7517 1940 -7483
rect 1860 -7563 1940 -7517
rect 1860 -7597 1883 -7563
rect 1917 -7597 1940 -7563
rect 1860 -7643 1940 -7597
rect 1860 -7677 1883 -7643
rect 1917 -7677 1940 -7643
rect 1860 -7710 1940 -7677
rect 2010 -7483 2090 -7460
rect 2010 -7517 2033 -7483
rect 2067 -7517 2090 -7483
rect 2010 -7563 2090 -7517
rect 2010 -7597 2033 -7563
rect 2067 -7597 2090 -7563
rect 2010 -7643 2090 -7597
rect 2010 -7677 2033 -7643
rect 2067 -7677 2090 -7643
rect 2010 -7710 2090 -7677
rect 2160 -7483 2240 -7460
rect 2160 -7517 2183 -7483
rect 2217 -7517 2240 -7483
rect 2160 -7563 2240 -7517
rect 2160 -7597 2183 -7563
rect 2217 -7597 2240 -7563
rect 2160 -7643 2240 -7597
rect 2160 -7677 2183 -7643
rect 2217 -7677 2240 -7643
rect 2160 -7710 2240 -7677
rect 2310 -7483 2390 -7460
rect 2310 -7517 2333 -7483
rect 2367 -7517 2390 -7483
rect 2310 -7563 2390 -7517
rect 2310 -7597 2333 -7563
rect 2367 -7597 2390 -7563
rect 2310 -7643 2390 -7597
rect 2310 -7677 2333 -7643
rect 2367 -7677 2390 -7643
rect 2310 -7710 2390 -7677
rect 2460 -7483 2540 -7460
rect 2460 -7517 2483 -7483
rect 2517 -7517 2540 -7483
rect 2460 -7563 2540 -7517
rect 2460 -7597 2483 -7563
rect 2517 -7597 2540 -7563
rect 2460 -7643 2540 -7597
rect 2460 -7677 2483 -7643
rect 2517 -7677 2540 -7643
rect 2460 -7710 2540 -7677
rect 2640 -7483 2720 -7460
rect 2640 -7517 2663 -7483
rect 2697 -7517 2720 -7483
rect 2640 -7563 2720 -7517
rect 2640 -7597 2663 -7563
rect 2697 -7597 2720 -7563
rect 2640 -7643 2720 -7597
rect 2640 -7677 2663 -7643
rect 2697 -7677 2720 -7643
rect 2640 -7710 2720 -7677
rect 2940 -7483 3020 -7460
rect 2940 -7517 2963 -7483
rect 2997 -7517 3020 -7483
rect 2940 -7563 3020 -7517
rect 2940 -7597 2963 -7563
rect 2997 -7597 3020 -7563
rect 2940 -7643 3020 -7597
rect 2940 -7677 2963 -7643
rect 2997 -7677 3020 -7643
rect 2940 -7710 3020 -7677
rect 3240 -7483 3320 -7460
rect 3240 -7517 3263 -7483
rect 3297 -7517 3320 -7483
rect 3240 -7563 3320 -7517
rect 3740 -7483 3820 -7460
rect 3740 -7517 3763 -7483
rect 3797 -7517 3820 -7483
rect 3240 -7597 3263 -7563
rect 3297 -7597 3320 -7563
rect 3240 -7643 3320 -7597
rect 3354 -7557 3434 -7537
rect 3354 -7561 3706 -7557
rect 3354 -7595 3377 -7561
rect 3411 -7595 3706 -7561
rect 3354 -7597 3706 -7595
rect 3354 -7617 3434 -7597
rect 3240 -7677 3263 -7643
rect 3297 -7677 3320 -7643
rect 3240 -7710 3320 -7677
rect 1100 -7750 1140 -7710
rect 1700 -7750 1740 -7710
rect 2030 -7750 2070 -7710
rect 1100 -7790 2070 -7750
rect 2030 -7920 2070 -7790
rect 2110 -7798 2190 -7775
rect 2110 -7832 2133 -7798
rect 2167 -7800 2190 -7798
rect 2330 -7800 2370 -7710
rect 2660 -7800 2700 -7710
rect 3260 -7800 3300 -7710
rect 3340 -7799 3420 -7776
rect 3340 -7800 3363 -7799
rect 2167 -7832 3363 -7800
rect 2110 -7833 3363 -7832
rect 3397 -7833 3420 -7799
rect 2110 -7840 3420 -7833
rect 3666 -7800 3706 -7597
rect 3740 -7563 3820 -7517
rect 3740 -7597 3763 -7563
rect 3797 -7597 3820 -7563
rect 3740 -7643 3820 -7597
rect 3740 -7677 3763 -7643
rect 3797 -7677 3820 -7643
rect 3740 -7710 3820 -7677
rect 3890 -7483 3970 -7460
rect 3890 -7517 3913 -7483
rect 3947 -7517 3970 -7483
rect 3890 -7563 3970 -7517
rect 3890 -7597 3913 -7563
rect 3947 -7597 3970 -7563
rect 3890 -7643 3970 -7597
rect 3890 -7677 3913 -7643
rect 3947 -7677 3970 -7643
rect 3890 -7710 3970 -7677
rect 4070 -7483 4150 -7460
rect 4070 -7517 4093 -7483
rect 4127 -7517 4150 -7483
rect 4070 -7563 4150 -7517
rect 4070 -7597 4093 -7563
rect 4127 -7597 4150 -7563
rect 4070 -7643 4150 -7597
rect 4070 -7677 4093 -7643
rect 4127 -7677 4150 -7643
rect 4070 -7710 4150 -7677
rect 4220 -7483 4300 -7460
rect 4220 -7517 4243 -7483
rect 4277 -7517 4300 -7483
rect 4220 -7563 4300 -7517
rect 4220 -7597 4243 -7563
rect 4277 -7597 4300 -7563
rect 4220 -7643 4300 -7597
rect 4220 -7677 4243 -7643
rect 4277 -7677 4300 -7643
rect 4220 -7710 4300 -7677
rect 4370 -7483 4450 -7460
rect 4370 -7517 4393 -7483
rect 4427 -7517 4450 -7483
rect 4370 -7563 4450 -7517
rect 4370 -7597 4393 -7563
rect 4427 -7597 4450 -7563
rect 4370 -7643 4450 -7597
rect 4370 -7677 4393 -7643
rect 4427 -7677 4450 -7643
rect 4370 -7710 4450 -7677
rect 4520 -7483 4600 -7460
rect 4520 -7517 4543 -7483
rect 4577 -7517 4600 -7483
rect 4520 -7563 4600 -7517
rect 4520 -7597 4543 -7563
rect 4577 -7597 4600 -7563
rect 4520 -7643 4600 -7597
rect 4520 -7677 4543 -7643
rect 4577 -7677 4600 -7643
rect 3910 -7750 3950 -7710
rect 4240 -7750 4280 -7710
rect 4520 -7750 4600 -7677
rect 4670 -7483 4750 -7460
rect 4670 -7517 4693 -7483
rect 4727 -7517 4750 -7483
rect 4670 -7563 4750 -7517
rect 4670 -7597 4693 -7563
rect 4727 -7597 4750 -7563
rect 4670 -7643 4750 -7597
rect 4670 -7677 4693 -7643
rect 4727 -7677 4750 -7643
rect 4670 -7710 4750 -7677
rect 4850 -7483 4930 -7460
rect 4850 -7517 4873 -7483
rect 4907 -7517 4930 -7483
rect 4850 -7563 4930 -7517
rect 4850 -7597 4873 -7563
rect 4907 -7597 4930 -7563
rect 4850 -7643 4930 -7597
rect 4850 -7677 4873 -7643
rect 4907 -7677 4930 -7643
rect 4850 -7710 4930 -7677
rect 5000 -7483 5080 -7460
rect 5000 -7517 5023 -7483
rect 5057 -7517 5080 -7483
rect 5000 -7563 5080 -7517
rect 5000 -7597 5023 -7563
rect 5057 -7597 5080 -7563
rect 5000 -7643 5080 -7597
rect 5000 -7677 5023 -7643
rect 5057 -7677 5080 -7643
rect 5000 -7710 5080 -7677
rect 5469 -7483 5549 -7460
rect 5469 -7517 5492 -7483
rect 5526 -7517 5549 -7483
rect 5469 -7563 5549 -7517
rect 5469 -7597 5492 -7563
rect 5526 -7597 5549 -7563
rect 5469 -7643 5549 -7597
rect 5469 -7677 5492 -7643
rect 5526 -7677 5549 -7643
rect 5469 -7710 5549 -7677
rect 5619 -7483 5699 -7460
rect 5619 -7517 5642 -7483
rect 5676 -7517 5699 -7483
rect 5619 -7563 5699 -7517
rect 5619 -7597 5642 -7563
rect 5676 -7597 5699 -7563
rect 5619 -7643 5699 -7597
rect 5619 -7677 5642 -7643
rect 5676 -7677 5699 -7643
rect 5619 -7710 5699 -7677
rect 5769 -7483 5849 -7460
rect 5769 -7517 5792 -7483
rect 5826 -7517 5849 -7483
rect 5769 -7563 5849 -7517
rect 5769 -7597 5792 -7563
rect 5826 -7597 5849 -7563
rect 5769 -7643 5849 -7597
rect 5769 -7677 5792 -7643
rect 5826 -7677 5849 -7643
rect 5769 -7710 5849 -7677
rect 5949 -7483 6029 -7460
rect 5949 -7517 5972 -7483
rect 6006 -7517 6029 -7483
rect 5949 -7563 6029 -7517
rect 5949 -7597 5972 -7563
rect 6006 -7597 6029 -7563
rect 5949 -7643 6029 -7597
rect 5949 -7677 5972 -7643
rect 6006 -7677 6029 -7643
rect 5949 -7710 6029 -7677
rect 6099 -7483 6179 -7460
rect 6099 -7517 6122 -7483
rect 6156 -7517 6179 -7483
rect 6099 -7563 6179 -7517
rect 6099 -7597 6122 -7563
rect 6156 -7597 6179 -7563
rect 6099 -7643 6179 -7597
rect 6099 -7677 6122 -7643
rect 6156 -7677 6179 -7643
rect 6099 -7710 6179 -7677
rect 6249 -7483 6329 -7460
rect 6249 -7517 6272 -7483
rect 6306 -7517 6329 -7483
rect 6249 -7563 6329 -7517
rect 6249 -7597 6272 -7563
rect 6306 -7597 6329 -7563
rect 6249 -7643 6329 -7597
rect 6249 -7677 6272 -7643
rect 6306 -7677 6329 -7643
rect 6249 -7710 6329 -7677
rect 6399 -7483 6479 -7460
rect 6399 -7517 6422 -7483
rect 6456 -7517 6479 -7483
rect 6399 -7563 6479 -7517
rect 6399 -7597 6422 -7563
rect 6456 -7597 6479 -7563
rect 6399 -7643 6479 -7597
rect 6399 -7677 6422 -7643
rect 6456 -7677 6479 -7643
rect 6399 -7710 6479 -7677
rect 6549 -7483 6629 -7460
rect 6549 -7517 6572 -7483
rect 6606 -7517 6629 -7483
rect 6549 -7563 6629 -7517
rect 6549 -7597 6572 -7563
rect 6606 -7597 6629 -7563
rect 6549 -7643 6629 -7597
rect 6549 -7677 6572 -7643
rect 6606 -7677 6629 -7643
rect 6549 -7710 6629 -7677
rect 6729 -7483 6809 -7460
rect 6729 -7517 6752 -7483
rect 6786 -7517 6809 -7483
rect 6729 -7563 6809 -7517
rect 6729 -7597 6752 -7563
rect 6786 -7597 6809 -7563
rect 6729 -7643 6809 -7597
rect 6729 -7677 6752 -7643
rect 6786 -7677 6809 -7643
rect 6729 -7710 6809 -7677
rect 7029 -7483 7109 -7460
rect 7029 -7517 7052 -7483
rect 7086 -7517 7109 -7483
rect 7029 -7563 7109 -7517
rect 7029 -7597 7052 -7563
rect 7086 -7597 7109 -7563
rect 7029 -7643 7109 -7597
rect 7029 -7677 7052 -7643
rect 7086 -7677 7109 -7643
rect 7029 -7710 7109 -7677
rect 4870 -7750 4910 -7710
rect 5489 -7750 5529 -7710
rect 5789 -7750 5829 -7710
rect 6120 -7750 6159 -7710
rect 3790 -7800 3870 -7780
rect 3910 -7790 4280 -7750
rect 4540 -7773 5188 -7750
rect 3666 -7803 3870 -7800
rect 3666 -7837 3813 -7803
rect 3847 -7837 3870 -7803
rect 3666 -7840 3870 -7837
rect 2110 -7855 2190 -7840
rect 2210 -7920 2290 -7900
rect 2030 -7923 2290 -7920
rect 570 -7973 650 -7950
rect 2030 -7957 2233 -7923
rect 2267 -7957 2290 -7923
rect 2030 -7960 2290 -7957
rect 570 -8007 593 -7973
rect 627 -7990 650 -7973
rect 1130 -7990 1210 -7970
rect 1710 -7990 1790 -7970
rect 627 -7993 1790 -7990
rect 627 -8007 1153 -7993
rect 570 -8027 1153 -8007
rect 1187 -8027 1733 -7993
rect 1767 -8027 1790 -7993
rect 2030 -8010 2070 -7960
rect 2210 -7980 2290 -7960
rect 2330 -8010 2370 -7840
rect 3340 -7856 3420 -7840
rect 3790 -7860 3870 -7840
rect 2580 -7913 3344 -7890
rect 2580 -7947 2603 -7913
rect 2637 -7930 3344 -7913
rect 2637 -7947 2660 -7930
rect 2580 -7970 2660 -7947
rect 2740 -7993 2820 -7970
rect 570 -8030 1790 -8027
rect 1130 -8050 1210 -8030
rect 1710 -8050 1790 -8030
rect 1860 -8043 1940 -8020
rect 456 -8073 536 -8050
rect 456 -8107 479 -8073
rect 513 -8090 536 -8073
rect 1580 -8090 1660 -8070
rect 513 -8093 1660 -8090
rect 513 -8107 1603 -8093
rect 456 -8127 1603 -8107
rect 1637 -8127 1660 -8093
rect 456 -8130 1660 -8127
rect 1580 -8150 1660 -8130
rect 1860 -8077 1883 -8043
rect 1917 -8077 1940 -8043
rect 1860 -8123 1940 -8077
rect 1860 -8157 1883 -8123
rect 1917 -8157 1940 -8123
rect 798 -8190 878 -8168
rect 1330 -8190 1410 -8170
rect 1710 -8190 1790 -8170
rect 798 -8191 1790 -8190
rect 798 -8225 821 -8191
rect 855 -8193 1790 -8191
rect 855 -8225 1353 -8193
rect 798 -8227 1353 -8225
rect 1387 -8227 1733 -8193
rect 1767 -8227 1790 -8193
rect 798 -8230 1790 -8227
rect 798 -8248 878 -8230
rect 1330 -8250 1410 -8230
rect 1710 -8250 1790 -8230
rect 1860 -8203 1940 -8157
rect 1860 -8237 1883 -8203
rect 1917 -8237 1940 -8203
rect 684 -8273 764 -8250
rect 1860 -8270 1940 -8237
rect 2010 -8043 2090 -8010
rect 2010 -8077 2033 -8043
rect 2067 -8077 2090 -8043
rect 2010 -8123 2090 -8077
rect 2010 -8157 2033 -8123
rect 2067 -8157 2090 -8123
rect 2010 -8203 2090 -8157
rect 2010 -8237 2033 -8203
rect 2067 -8237 2090 -8203
rect 2010 -8270 2090 -8237
rect 2160 -8043 2240 -8020
rect 2160 -8077 2183 -8043
rect 2217 -8077 2240 -8043
rect 2160 -8123 2240 -8077
rect 2160 -8157 2183 -8123
rect 2217 -8157 2240 -8123
rect 2160 -8203 2240 -8157
rect 2160 -8237 2183 -8203
rect 2217 -8237 2240 -8203
rect 2160 -8270 2240 -8237
rect 2310 -8043 2390 -8010
rect 2310 -8077 2333 -8043
rect 2367 -8077 2390 -8043
rect 2310 -8123 2390 -8077
rect 2310 -8157 2333 -8123
rect 2367 -8157 2390 -8123
rect 2310 -8203 2390 -8157
rect 2310 -8237 2333 -8203
rect 2367 -8237 2390 -8203
rect 2310 -8270 2390 -8237
rect 2460 -8043 2540 -8020
rect 2460 -8077 2483 -8043
rect 2517 -8077 2540 -8043
rect 2740 -8027 2763 -7993
rect 2797 -8027 2820 -7993
rect 2740 -8050 2820 -8027
rect 2460 -8123 2540 -8077
rect 2460 -8157 2483 -8123
rect 2517 -8157 2540 -8123
rect 3190 -8093 3270 -8070
rect 3190 -8127 3213 -8093
rect 3247 -8127 3270 -8093
rect 3190 -8150 3270 -8127
rect 2460 -8203 2540 -8157
rect 2460 -8237 2483 -8203
rect 2517 -8237 2540 -8203
rect 2460 -8270 2540 -8237
rect 3040 -8193 3120 -8170
rect 3040 -8227 3063 -8193
rect 3097 -8227 3120 -8193
rect 3040 -8250 3120 -8227
rect 3304 -8224 3344 -7930
rect 4240 -7920 4280 -7790
rect 4320 -7798 4400 -7775
rect 4320 -7832 4343 -7798
rect 4377 -7800 4400 -7798
rect 4540 -7790 5131 -7773
rect 4540 -7800 4580 -7790
rect 4377 -7832 4580 -7800
rect 5108 -7807 5131 -7790
rect 5165 -7807 5188 -7773
rect 5489 -7790 6159 -7750
rect 5108 -7830 5188 -7807
rect 4320 -7840 4580 -7832
rect 4320 -7855 4400 -7840
rect 4420 -7920 4500 -7900
rect 4240 -7923 4500 -7920
rect 4240 -7957 4443 -7923
rect 4477 -7957 4500 -7923
rect 4240 -7960 4500 -7957
rect 4240 -8010 4280 -7960
rect 4420 -7980 4500 -7960
rect 4540 -8010 4580 -7840
rect 5519 -7870 5599 -7850
rect 5242 -7873 5599 -7870
rect 4820 -7920 4900 -7900
rect 5242 -7907 5542 -7873
rect 5576 -7907 5599 -7873
rect 5242 -7910 5599 -7907
rect 5242 -7920 5282 -7910
rect 4820 -7923 5282 -7920
rect 4820 -7957 4843 -7923
rect 4877 -7957 5282 -7923
rect 5519 -7930 5599 -7910
rect 6119 -7920 6159 -7790
rect 6199 -7798 6279 -7775
rect 6199 -7832 6222 -7798
rect 6256 -7800 6279 -7798
rect 6419 -7800 6459 -7710
rect 6749 -7800 6789 -7710
rect 7133 -7800 7213 -7781
rect 6256 -7804 7213 -7800
rect 6256 -7832 7156 -7804
rect 6199 -7838 7156 -7832
rect 7190 -7838 7213 -7804
rect 6199 -7840 7213 -7838
rect 6199 -7855 6279 -7840
rect 6299 -7920 6379 -7900
rect 6119 -7923 6379 -7920
rect 4820 -7960 5282 -7957
rect 4820 -7980 4900 -7960
rect 5669 -7970 5749 -7950
rect 5316 -7973 5749 -7970
rect 5316 -7994 5692 -7973
rect 5129 -8007 5692 -7994
rect 5726 -8007 5749 -7973
rect 5129 -8010 5749 -8007
rect 6119 -7957 6322 -7923
rect 6356 -7957 6379 -7923
rect 6119 -7960 6379 -7957
rect 6119 -8010 6159 -7960
rect 6299 -7980 6379 -7960
rect 6419 -8010 6459 -7840
rect 7133 -7861 7213 -7840
rect 6699 -7920 6779 -7900
rect 7282 -7920 7322 -5834
rect 7494 -5854 7574 -5834
rect 6699 -7923 7322 -7920
rect 6699 -7957 6722 -7923
rect 6756 -7957 7322 -7923
rect 6699 -7960 7322 -7957
rect 6699 -7980 6779 -7960
rect 3920 -8040 4000 -8020
rect 3720 -8043 4000 -8040
rect 3720 -8077 3943 -8043
rect 3977 -8077 4000 -8043
rect 3720 -8080 4000 -8077
rect 3920 -8100 4000 -8080
rect 4070 -8043 4150 -8020
rect 4070 -8077 4093 -8043
rect 4127 -8077 4150 -8043
rect 4070 -8123 4150 -8077
rect 4070 -8157 4093 -8123
rect 4127 -8157 4150 -8123
rect 4070 -8203 4150 -8157
rect 3632 -8224 3712 -8204
rect 3304 -8227 3712 -8224
rect 3304 -8261 3655 -8227
rect 3689 -8261 3712 -8227
rect 3304 -8264 3712 -8261
rect 684 -8307 707 -8273
rect 741 -8290 764 -8273
rect 1450 -8290 1530 -8270
rect 1580 -8290 1660 -8270
rect 741 -8293 1660 -8290
rect 741 -8307 1473 -8293
rect 684 -8327 1473 -8307
rect 1507 -8327 1603 -8293
rect 1637 -8327 1660 -8293
rect 684 -8330 1660 -8327
rect 1450 -8350 1530 -8330
rect 1580 -8350 1660 -8330
rect 2840 -8293 2920 -8270
rect 3632 -8284 3712 -8264
rect 4070 -8237 4093 -8203
rect 4127 -8237 4150 -8203
rect 4070 -8270 4150 -8237
rect 4220 -8043 4300 -8010
rect 4220 -8077 4243 -8043
rect 4277 -8077 4300 -8043
rect 4220 -8123 4300 -8077
rect 4220 -8157 4243 -8123
rect 4277 -8157 4300 -8123
rect 4220 -8203 4300 -8157
rect 4220 -8237 4243 -8203
rect 4277 -8237 4300 -8203
rect 4220 -8270 4300 -8237
rect 4370 -8043 4450 -8020
rect 4370 -8077 4393 -8043
rect 4427 -8077 4450 -8043
rect 4370 -8123 4450 -8077
rect 4370 -8157 4393 -8123
rect 4427 -8157 4450 -8123
rect 4370 -8203 4450 -8157
rect 4370 -8237 4393 -8203
rect 4427 -8237 4450 -8203
rect 4370 -8270 4450 -8237
rect 4520 -8043 4600 -8010
rect 4520 -8077 4543 -8043
rect 4577 -8077 4600 -8043
rect 4520 -8123 4600 -8077
rect 4520 -8157 4543 -8123
rect 4577 -8157 4600 -8123
rect 4520 -8203 4600 -8157
rect 4520 -8237 4543 -8203
rect 4577 -8237 4600 -8203
rect 4520 -8270 4600 -8237
rect 4670 -8043 4750 -8020
rect 4670 -8077 4693 -8043
rect 4727 -8077 4750 -8043
rect 4670 -8123 4750 -8077
rect 4820 -8040 4900 -8020
rect 4950 -8040 5030 -8020
rect 4820 -8043 5030 -8040
rect 4820 -8077 4843 -8043
rect 4877 -8077 4973 -8043
rect 5007 -8077 5030 -8043
rect 4820 -8080 5030 -8077
rect 4820 -8100 4900 -8080
rect 4950 -8100 5030 -8080
rect 5129 -8034 5356 -8010
rect 5669 -8030 5749 -8010
rect 5129 -8089 5169 -8034
rect 5949 -8043 6029 -8020
rect 5799 -8070 5879 -8050
rect 5370 -8073 5879 -8070
rect 4670 -8157 4693 -8123
rect 4727 -8157 4750 -8123
rect 4670 -8203 4750 -8157
rect 5108 -8112 5188 -8089
rect 5108 -8146 5131 -8112
rect 5165 -8146 5188 -8112
rect 5108 -8169 5188 -8146
rect 5370 -8093 5822 -8073
rect 5370 -8127 5393 -8093
rect 5427 -8107 5822 -8093
rect 5856 -8107 5879 -8073
rect 5427 -8110 5879 -8107
rect 5427 -8127 5450 -8110
rect 5370 -8150 5450 -8127
rect 5799 -8130 5879 -8110
rect 5949 -8077 5972 -8043
rect 6006 -8077 6029 -8043
rect 5949 -8123 6029 -8077
rect 5949 -8157 5972 -8123
rect 6006 -8157 6029 -8123
rect 5799 -8190 5879 -8170
rect 4670 -8237 4693 -8203
rect 4727 -8237 4750 -8203
rect 5430 -8193 5879 -8190
rect 5430 -8204 5822 -8193
rect 4670 -8270 4750 -8237
rect 5108 -8227 5822 -8204
rect 5856 -8227 5879 -8193
rect 5108 -8261 5131 -8227
rect 5165 -8230 5879 -8227
rect 5165 -8244 5470 -8230
rect 5165 -8261 5188 -8244
rect 5799 -8250 5879 -8230
rect 5949 -8203 6029 -8157
rect 5949 -8237 5972 -8203
rect 6006 -8237 6029 -8203
rect 5108 -8284 5188 -8261
rect 5949 -8270 6029 -8237
rect 6099 -8043 6179 -8010
rect 6099 -8077 6122 -8043
rect 6156 -8077 6179 -8043
rect 6099 -8123 6179 -8077
rect 6099 -8157 6122 -8123
rect 6156 -8157 6179 -8123
rect 6099 -8203 6179 -8157
rect 6099 -8237 6122 -8203
rect 6156 -8237 6179 -8203
rect 6099 -8270 6179 -8237
rect 6249 -8043 6329 -8020
rect 6249 -8077 6272 -8043
rect 6306 -8077 6329 -8043
rect 6249 -8123 6329 -8077
rect 6249 -8157 6272 -8123
rect 6306 -8157 6329 -8123
rect 6249 -8203 6329 -8157
rect 6249 -8237 6272 -8203
rect 6306 -8237 6329 -8203
rect 6249 -8270 6329 -8237
rect 6399 -8043 6479 -8010
rect 6399 -8077 6422 -8043
rect 6456 -8077 6479 -8043
rect 6399 -8123 6479 -8077
rect 6399 -8157 6422 -8123
rect 6456 -8157 6479 -8123
rect 6399 -8203 6479 -8157
rect 6399 -8237 6422 -8203
rect 6456 -8237 6479 -8203
rect 6399 -8270 6479 -8237
rect 6549 -8043 6629 -8020
rect 6549 -8077 6572 -8043
rect 6606 -8077 6629 -8043
rect 6549 -8123 6629 -8077
rect 6549 -8157 6572 -8123
rect 6606 -8157 6629 -8123
rect 6779 -8073 6859 -8050
rect 6779 -8107 6802 -8073
rect 6836 -8107 6859 -8073
rect 6779 -8130 6859 -8107
rect 6549 -8203 6629 -8157
rect 6549 -8237 6572 -8203
rect 6606 -8237 6629 -8203
rect 6549 -8270 6629 -8237
rect 6929 -8193 7009 -8170
rect 6929 -8227 6952 -8193
rect 6986 -8227 7009 -8193
rect 6929 -8250 7009 -8227
rect 2840 -8327 2863 -8293
rect 2897 -8327 2920 -8293
rect 2840 -8350 2920 -8327
rect 1060 -8423 3340 -8400
rect 1060 -8457 1143 -8423
rect 1177 -8457 1223 -8423
rect 1257 -8457 1303 -8423
rect 1337 -8457 1383 -8423
rect 1417 -8457 1463 -8423
rect 1497 -8457 1543 -8423
rect 1577 -8457 1623 -8423
rect 1657 -8457 1703 -8423
rect 1737 -8457 1783 -8423
rect 1817 -8457 1863 -8423
rect 1897 -8457 1943 -8423
rect 1977 -8457 2023 -8423
rect 2057 -8457 2103 -8423
rect 2137 -8457 2183 -8423
rect 2217 -8457 2263 -8423
rect 2297 -8457 2343 -8423
rect 2377 -8457 2423 -8423
rect 2457 -8457 2503 -8423
rect 2537 -8457 2583 -8423
rect 2617 -8457 2663 -8423
rect 2697 -8457 2743 -8423
rect 2777 -8457 2823 -8423
rect 2857 -8457 2903 -8423
rect 2937 -8457 2983 -8423
rect 3017 -8457 3063 -8423
rect 3097 -8457 3143 -8423
rect 3177 -8457 3223 -8423
rect 3257 -8457 3340 -8423
rect 1060 -8480 3340 -8457
rect 3720 -8423 5100 -8400
rect 3720 -8457 3753 -8423
rect 3787 -8457 3833 -8423
rect 3867 -8457 3913 -8423
rect 3947 -8457 3993 -8423
rect 4027 -8457 4073 -8423
rect 4107 -8457 4153 -8423
rect 4187 -8457 4233 -8423
rect 4267 -8457 4313 -8423
rect 4347 -8457 4393 -8423
rect 4427 -8457 4473 -8423
rect 4507 -8457 4553 -8423
rect 4587 -8457 4633 -8423
rect 4667 -8457 4713 -8423
rect 4747 -8457 4793 -8423
rect 4827 -8457 4873 -8423
rect 4907 -8457 4953 -8423
rect 4987 -8457 5033 -8423
rect 5067 -8457 5100 -8423
rect 3720 -8480 5100 -8457
rect 5449 -8423 7129 -8400
rect 5449 -8457 5472 -8423
rect 5506 -8457 5552 -8423
rect 5586 -8457 5632 -8423
rect 5666 -8457 5712 -8423
rect 5746 -8457 5792 -8423
rect 5826 -8457 5872 -8423
rect 5906 -8457 5952 -8423
rect 5986 -8457 6032 -8423
rect 6066 -8457 6112 -8423
rect 6146 -8457 6192 -8423
rect 6226 -8457 6272 -8423
rect 6306 -8457 6352 -8423
rect 6386 -8457 6432 -8423
rect 6466 -8457 6512 -8423
rect 6546 -8457 6592 -8423
rect 6626 -8457 6672 -8423
rect 6706 -8457 6752 -8423
rect 6786 -8457 6832 -8423
rect 6866 -8457 6912 -8423
rect 6946 -8457 6992 -8423
rect 7026 -8457 7072 -8423
rect 7106 -8457 7129 -8423
rect 5449 -8480 7129 -8457
rect 1020 -8883 3300 -8860
rect 1020 -8917 1103 -8883
rect 1137 -8917 1183 -8883
rect 1217 -8917 1263 -8883
rect 1297 -8917 1343 -8883
rect 1377 -8917 1423 -8883
rect 1457 -8917 1503 -8883
rect 1537 -8917 1583 -8883
rect 1617 -8917 1663 -8883
rect 1697 -8917 1743 -8883
rect 1777 -8917 1823 -8883
rect 1857 -8917 1903 -8883
rect 1937 -8917 1983 -8883
rect 2017 -8917 2063 -8883
rect 2097 -8917 2143 -8883
rect 2177 -8917 2223 -8883
rect 2257 -8917 2303 -8883
rect 2337 -8917 2383 -8883
rect 2417 -8917 2463 -8883
rect 2497 -8917 2543 -8883
rect 2577 -8917 2623 -8883
rect 2657 -8917 2703 -8883
rect 2737 -8917 2783 -8883
rect 2817 -8917 2863 -8883
rect 2897 -8917 2943 -8883
rect 2977 -8917 3023 -8883
rect 3057 -8917 3103 -8883
rect 3137 -8917 3183 -8883
rect 3217 -8917 3300 -8883
rect 1020 -8940 3300 -8917
rect 3660 -8883 5040 -8860
rect 3660 -8917 3693 -8883
rect 3727 -8917 3773 -8883
rect 3807 -8917 3853 -8883
rect 3887 -8917 3933 -8883
rect 3967 -8917 4013 -8883
rect 4047 -8917 4093 -8883
rect 4127 -8917 4173 -8883
rect 4207 -8917 4253 -8883
rect 4287 -8917 4333 -8883
rect 4367 -8917 4413 -8883
rect 4447 -8917 4493 -8883
rect 4527 -8917 4573 -8883
rect 4607 -8917 4653 -8883
rect 4687 -8917 4733 -8883
rect 4767 -8917 4813 -8883
rect 4847 -8917 4893 -8883
rect 4927 -8917 4973 -8883
rect 5007 -8917 5040 -8883
rect 3660 -8940 5040 -8917
rect 5390 -8883 7070 -8860
rect 5390 -8917 5413 -8883
rect 5447 -8917 5493 -8883
rect 5527 -8917 5573 -8883
rect 5607 -8917 5653 -8883
rect 5687 -8917 5733 -8883
rect 5767 -8917 5813 -8883
rect 5847 -8917 5893 -8883
rect 5927 -8917 5973 -8883
rect 6007 -8917 6053 -8883
rect 6087 -8917 6133 -8883
rect 6167 -8917 6213 -8883
rect 6247 -8917 6293 -8883
rect 6327 -8917 6373 -8883
rect 6407 -8917 6453 -8883
rect 6487 -8917 6533 -8883
rect 6567 -8917 6613 -8883
rect 6647 -8917 6693 -8883
rect 6727 -8917 6773 -8883
rect 6807 -8917 6853 -8883
rect 6887 -8917 6933 -8883
rect 6967 -8917 7013 -8883
rect 7047 -8917 7070 -8883
rect 5390 -8940 7070 -8917
rect 228 -9010 308 -8990
rect 1410 -9010 1490 -8990
rect 1540 -9010 1620 -8990
rect 228 -9013 1620 -9010
rect 228 -9047 251 -9013
rect 285 -9047 1433 -9013
rect 1467 -9047 1563 -9013
rect 1597 -9047 1620 -9013
rect 228 -9050 1620 -9047
rect 228 -9070 308 -9050
rect 1410 -9070 1490 -9050
rect 1540 -9070 1620 -9050
rect 2800 -9013 2880 -8990
rect 2800 -9047 2823 -9013
rect 2857 -9047 2880 -9013
rect 2800 -9070 2880 -9047
rect 342 -9110 422 -9090
rect 1290 -9110 1370 -9090
rect 1670 -9110 1750 -9090
rect 342 -9113 1750 -9110
rect 342 -9147 365 -9113
rect 399 -9147 1313 -9113
rect 1347 -9147 1693 -9113
rect 1727 -9147 1750 -9113
rect 342 -9150 1750 -9147
rect 342 -9170 422 -9150
rect 1290 -9170 1370 -9150
rect 1670 -9170 1750 -9150
rect 1820 -9103 1900 -9070
rect 1820 -9137 1843 -9103
rect 1877 -9137 1900 -9103
rect 1820 -9183 1900 -9137
rect 0 -9210 80 -9190
rect 1540 -9210 1620 -9190
rect 0 -9213 1620 -9210
rect 0 -9247 23 -9213
rect 57 -9247 1563 -9213
rect 1597 -9247 1620 -9213
rect 0 -9250 1620 -9247
rect 0 -9270 80 -9250
rect 1540 -9270 1620 -9250
rect 1820 -9217 1843 -9183
rect 1877 -9217 1900 -9183
rect 1820 -9263 1900 -9217
rect 114 -9310 194 -9290
rect 1090 -9310 1170 -9290
rect 1670 -9310 1750 -9290
rect 114 -9313 1750 -9310
rect 114 -9347 137 -9313
rect 171 -9347 1113 -9313
rect 1147 -9347 1693 -9313
rect 1727 -9347 1750 -9313
rect 1820 -9297 1843 -9263
rect 1877 -9297 1900 -9263
rect 1820 -9320 1900 -9297
rect 1970 -9103 2050 -9070
rect 1970 -9137 1993 -9103
rect 2027 -9137 2050 -9103
rect 1970 -9183 2050 -9137
rect 1970 -9217 1993 -9183
rect 2027 -9217 2050 -9183
rect 1970 -9263 2050 -9217
rect 1970 -9297 1993 -9263
rect 2027 -9297 2050 -9263
rect 1970 -9330 2050 -9297
rect 2120 -9103 2200 -9070
rect 2120 -9137 2143 -9103
rect 2177 -9137 2200 -9103
rect 2120 -9183 2200 -9137
rect 2120 -9217 2143 -9183
rect 2177 -9217 2200 -9183
rect 2120 -9263 2200 -9217
rect 2120 -9297 2143 -9263
rect 2177 -9297 2200 -9263
rect 2120 -9320 2200 -9297
rect 2270 -9103 2350 -9070
rect 2270 -9137 2293 -9103
rect 2327 -9137 2350 -9103
rect 2270 -9183 2350 -9137
rect 2270 -9217 2293 -9183
rect 2327 -9217 2350 -9183
rect 2270 -9263 2350 -9217
rect 2270 -9297 2293 -9263
rect 2327 -9297 2350 -9263
rect 2270 -9330 2350 -9297
rect 2420 -9103 2500 -9070
rect 3572 -9078 3652 -9056
rect 3299 -9079 3652 -9078
rect 2420 -9137 2443 -9103
rect 2477 -9137 2500 -9103
rect 2420 -9183 2500 -9137
rect 3000 -9113 3080 -9090
rect 3000 -9147 3023 -9113
rect 3057 -9147 3080 -9113
rect 3000 -9170 3080 -9147
rect 3299 -9113 3595 -9079
rect 3629 -9113 3652 -9079
rect 3299 -9118 3652 -9113
rect 2420 -9217 2443 -9183
rect 2477 -9217 2500 -9183
rect 2420 -9263 2500 -9217
rect 2420 -9297 2443 -9263
rect 2477 -9297 2500 -9263
rect 3150 -9213 3230 -9190
rect 3150 -9247 3173 -9213
rect 3207 -9247 3230 -9213
rect 3150 -9270 3230 -9247
rect 2420 -9320 2500 -9297
rect 2700 -9313 2780 -9290
rect 114 -9350 1750 -9347
rect 114 -9370 194 -9350
rect 1090 -9370 1170 -9350
rect 1670 -9370 1750 -9350
rect 1990 -9380 2030 -9330
rect 2170 -9380 2250 -9360
rect 1990 -9383 2250 -9380
rect 1990 -9417 2193 -9383
rect 2227 -9417 2250 -9383
rect 1990 -9420 2250 -9417
rect 1990 -9550 2030 -9420
rect 2170 -9440 2250 -9420
rect 1060 -9590 2030 -9550
rect 2070 -9500 2150 -9485
rect 2290 -9500 2330 -9330
rect 2700 -9347 2723 -9313
rect 2757 -9347 2780 -9313
rect 2700 -9370 2780 -9347
rect 2540 -9393 2620 -9370
rect 2540 -9427 2563 -9393
rect 2597 -9410 2620 -9393
rect 3299 -9410 3339 -9118
rect 3572 -9136 3652 -9118
rect 4010 -9103 4090 -9070
rect 4010 -9137 4033 -9103
rect 4067 -9137 4090 -9103
rect 4010 -9183 4090 -9137
rect 4010 -9217 4033 -9183
rect 4067 -9217 4090 -9183
rect 3860 -9260 3940 -9240
rect 3660 -9263 3940 -9260
rect 3660 -9297 3883 -9263
rect 3917 -9297 3940 -9263
rect 3660 -9300 3940 -9297
rect 3860 -9320 3940 -9300
rect 4010 -9263 4090 -9217
rect 4010 -9297 4033 -9263
rect 4067 -9297 4090 -9263
rect 4010 -9320 4090 -9297
rect 4160 -9103 4240 -9070
rect 4160 -9137 4183 -9103
rect 4217 -9137 4240 -9103
rect 4160 -9183 4240 -9137
rect 4160 -9217 4183 -9183
rect 4217 -9217 4240 -9183
rect 4160 -9263 4240 -9217
rect 4160 -9297 4183 -9263
rect 4217 -9297 4240 -9263
rect 4160 -9330 4240 -9297
rect 4310 -9103 4390 -9070
rect 4310 -9137 4333 -9103
rect 4367 -9137 4390 -9103
rect 4310 -9183 4390 -9137
rect 4310 -9217 4333 -9183
rect 4367 -9217 4390 -9183
rect 4310 -9263 4390 -9217
rect 4310 -9297 4333 -9263
rect 4367 -9297 4390 -9263
rect 4310 -9320 4390 -9297
rect 4460 -9103 4540 -9070
rect 4460 -9137 4483 -9103
rect 4517 -9137 4540 -9103
rect 4460 -9183 4540 -9137
rect 4460 -9217 4483 -9183
rect 4517 -9217 4540 -9183
rect 4460 -9263 4540 -9217
rect 4460 -9297 4483 -9263
rect 4517 -9297 4540 -9263
rect 4460 -9330 4540 -9297
rect 4610 -9103 4690 -9070
rect 4610 -9137 4633 -9103
rect 4667 -9137 4690 -9103
rect 4610 -9183 4690 -9137
rect 5310 -9110 5390 -9090
rect 5740 -9110 5820 -9090
rect 5310 -9113 5820 -9110
rect 5310 -9147 5333 -9113
rect 5367 -9147 5763 -9113
rect 5797 -9147 5820 -9113
rect 5310 -9150 5820 -9147
rect 5310 -9170 5390 -9150
rect 5740 -9170 5820 -9150
rect 5890 -9103 5970 -9070
rect 5890 -9137 5913 -9103
rect 5947 -9137 5970 -9103
rect 4610 -9217 4633 -9183
rect 4667 -9217 4690 -9183
rect 5890 -9183 5970 -9137
rect 4610 -9263 4690 -9217
rect 5162 -9230 5551 -9225
rect 5740 -9230 5820 -9210
rect 5162 -9233 5820 -9230
rect 4610 -9297 4633 -9263
rect 4667 -9297 4690 -9263
rect 4610 -9320 4690 -9297
rect 4760 -9260 4840 -9240
rect 4890 -9260 4970 -9240
rect 4760 -9263 4970 -9260
rect 4760 -9297 4783 -9263
rect 4817 -9297 4913 -9263
rect 4947 -9297 4970 -9263
rect 4760 -9300 4970 -9297
rect 4760 -9320 4840 -9300
rect 4890 -9320 4970 -9300
rect 5162 -9265 5763 -9233
rect 2597 -9427 3339 -9410
rect 2540 -9450 3339 -9427
rect 4180 -9380 4220 -9330
rect 4360 -9380 4440 -9360
rect 4180 -9383 4440 -9380
rect 4180 -9417 4383 -9383
rect 4417 -9417 4440 -9383
rect 4180 -9420 4440 -9417
rect 3300 -9500 3380 -9484
rect 3730 -9500 3810 -9480
rect 2070 -9507 3380 -9500
rect 2070 -9508 3323 -9507
rect 2070 -9542 2093 -9508
rect 2127 -9540 3323 -9508
rect 2127 -9542 2150 -9540
rect 2070 -9565 2150 -9542
rect 1060 -9630 1100 -9590
rect 1660 -9630 1700 -9590
rect 1990 -9630 2030 -9590
rect 2290 -9630 2330 -9540
rect 2620 -9630 2660 -9540
rect 3220 -9630 3260 -9540
rect 3300 -9541 3323 -9540
rect 3357 -9541 3380 -9507
rect 3300 -9564 3380 -9541
rect 3606 -9503 3810 -9500
rect 3606 -9537 3753 -9503
rect 3787 -9537 3810 -9503
rect 3606 -9540 3810 -9537
rect 1040 -9663 1120 -9630
rect 1040 -9697 1063 -9663
rect 1097 -9697 1120 -9663
rect 1040 -9743 1120 -9697
rect 1040 -9777 1063 -9743
rect 1097 -9777 1120 -9743
rect 1040 -9823 1120 -9777
rect 1040 -9857 1063 -9823
rect 1097 -9857 1120 -9823
rect 1040 -9880 1120 -9857
rect 1340 -9663 1420 -9630
rect 1340 -9697 1363 -9663
rect 1397 -9697 1420 -9663
rect 1340 -9743 1420 -9697
rect 1340 -9777 1363 -9743
rect 1397 -9777 1420 -9743
rect 1340 -9823 1420 -9777
rect 1340 -9857 1363 -9823
rect 1397 -9857 1420 -9823
rect 1340 -9880 1420 -9857
rect 1640 -9663 1720 -9630
rect 1640 -9697 1663 -9663
rect 1697 -9697 1720 -9663
rect 1640 -9743 1720 -9697
rect 1640 -9777 1663 -9743
rect 1697 -9777 1720 -9743
rect 1640 -9823 1720 -9777
rect 1640 -9857 1663 -9823
rect 1697 -9857 1720 -9823
rect 1640 -9880 1720 -9857
rect 1820 -9663 1900 -9630
rect 1820 -9697 1843 -9663
rect 1877 -9697 1900 -9663
rect 1820 -9743 1900 -9697
rect 1820 -9777 1843 -9743
rect 1877 -9777 1900 -9743
rect 1820 -9823 1900 -9777
rect 1820 -9857 1843 -9823
rect 1877 -9857 1900 -9823
rect 1820 -9880 1900 -9857
rect 1970 -9663 2050 -9630
rect 1970 -9697 1993 -9663
rect 2027 -9697 2050 -9663
rect 1970 -9743 2050 -9697
rect 1970 -9777 1993 -9743
rect 2027 -9777 2050 -9743
rect 1970 -9823 2050 -9777
rect 1970 -9857 1993 -9823
rect 2027 -9857 2050 -9823
rect 1970 -9880 2050 -9857
rect 2120 -9663 2200 -9630
rect 2120 -9697 2143 -9663
rect 2177 -9697 2200 -9663
rect 2120 -9743 2200 -9697
rect 2120 -9777 2143 -9743
rect 2177 -9777 2200 -9743
rect 2120 -9823 2200 -9777
rect 2120 -9857 2143 -9823
rect 2177 -9857 2200 -9823
rect 2120 -9880 2200 -9857
rect 2270 -9663 2350 -9630
rect 2270 -9697 2293 -9663
rect 2327 -9697 2350 -9663
rect 2270 -9743 2350 -9697
rect 2270 -9777 2293 -9743
rect 2327 -9777 2350 -9743
rect 2270 -9823 2350 -9777
rect 2270 -9857 2293 -9823
rect 2327 -9857 2350 -9823
rect 2270 -9880 2350 -9857
rect 2420 -9663 2500 -9630
rect 2420 -9697 2443 -9663
rect 2477 -9697 2500 -9663
rect 2420 -9743 2500 -9697
rect 2420 -9777 2443 -9743
rect 2477 -9777 2500 -9743
rect 2420 -9823 2500 -9777
rect 2420 -9857 2443 -9823
rect 2477 -9857 2500 -9823
rect 2420 -9880 2500 -9857
rect 2600 -9663 2680 -9630
rect 2600 -9697 2623 -9663
rect 2657 -9697 2680 -9663
rect 2600 -9743 2680 -9697
rect 2600 -9777 2623 -9743
rect 2657 -9777 2680 -9743
rect 2600 -9823 2680 -9777
rect 2600 -9857 2623 -9823
rect 2657 -9857 2680 -9823
rect 2600 -9880 2680 -9857
rect 2900 -9663 2980 -9630
rect 2900 -9697 2923 -9663
rect 2957 -9697 2980 -9663
rect 2900 -9743 2980 -9697
rect 2900 -9777 2923 -9743
rect 2957 -9777 2980 -9743
rect 2900 -9823 2980 -9777
rect 2900 -9857 2923 -9823
rect 2957 -9857 2980 -9823
rect 2900 -9880 2980 -9857
rect 3200 -9663 3280 -9630
rect 3200 -9697 3223 -9663
rect 3257 -9697 3280 -9663
rect 3200 -9743 3280 -9697
rect 3200 -9777 3223 -9743
rect 3257 -9777 3280 -9743
rect 3314 -9708 3394 -9689
rect 3606 -9708 3646 -9540
rect 3730 -9560 3810 -9540
rect 4180 -9550 4220 -9420
rect 4360 -9440 4440 -9420
rect 3850 -9590 4220 -9550
rect 4260 -9500 4340 -9485
rect 4480 -9500 4520 -9330
rect 4760 -9380 4840 -9360
rect 5048 -9380 5128 -9366
rect 4760 -9383 5128 -9380
rect 4760 -9417 4783 -9383
rect 4817 -9389 5128 -9383
rect 4817 -9417 5071 -9389
rect 4760 -9420 5071 -9417
rect 4760 -9440 4840 -9420
rect 5048 -9423 5071 -9420
rect 5105 -9423 5128 -9389
rect 5048 -9446 5128 -9423
rect 4260 -9508 4520 -9500
rect 4260 -9542 4283 -9508
rect 4317 -9540 4520 -9508
rect 4317 -9542 4340 -9540
rect 4260 -9565 4340 -9542
rect 4480 -9550 4520 -9540
rect 5162 -9550 5202 -9265
rect 5390 -9267 5763 -9265
rect 5797 -9267 5820 -9233
rect 5390 -9270 5820 -9267
rect 5740 -9290 5820 -9270
rect 5890 -9217 5913 -9183
rect 5947 -9217 5970 -9183
rect 5890 -9263 5970 -9217
rect 5890 -9297 5913 -9263
rect 5947 -9297 5970 -9263
rect 5310 -9330 5390 -9310
rect 5610 -9330 5690 -9310
rect 5890 -9320 5970 -9297
rect 6040 -9103 6120 -9070
rect 6040 -9137 6063 -9103
rect 6097 -9137 6120 -9103
rect 6040 -9183 6120 -9137
rect 6040 -9217 6063 -9183
rect 6097 -9217 6120 -9183
rect 6040 -9263 6120 -9217
rect 6040 -9297 6063 -9263
rect 6097 -9297 6120 -9263
rect 6040 -9330 6120 -9297
rect 6190 -9103 6270 -9070
rect 6190 -9137 6213 -9103
rect 6247 -9137 6270 -9103
rect 6190 -9183 6270 -9137
rect 6190 -9217 6213 -9183
rect 6247 -9217 6270 -9183
rect 6190 -9263 6270 -9217
rect 6190 -9297 6213 -9263
rect 6247 -9297 6270 -9263
rect 6190 -9320 6270 -9297
rect 6340 -9103 6420 -9070
rect 6340 -9137 6363 -9103
rect 6397 -9137 6420 -9103
rect 6340 -9183 6420 -9137
rect 6340 -9217 6363 -9183
rect 6397 -9217 6420 -9183
rect 6340 -9263 6420 -9217
rect 6340 -9297 6363 -9263
rect 6397 -9297 6420 -9263
rect 6340 -9330 6420 -9297
rect 6490 -9103 6570 -9070
rect 6490 -9137 6513 -9103
rect 6547 -9137 6570 -9103
rect 6490 -9183 6570 -9137
rect 6870 -9113 6950 -9090
rect 6870 -9147 6893 -9113
rect 6927 -9147 6950 -9113
rect 6870 -9170 6950 -9147
rect 6490 -9217 6513 -9183
rect 6547 -9217 6570 -9183
rect 6490 -9263 6570 -9217
rect 6490 -9297 6513 -9263
rect 6547 -9297 6570 -9263
rect 6720 -9233 6800 -9210
rect 6720 -9267 6743 -9233
rect 6777 -9267 6800 -9233
rect 6720 -9290 6800 -9267
rect 6490 -9320 6570 -9297
rect 5310 -9333 5690 -9330
rect 5310 -9367 5333 -9333
rect 5367 -9367 5633 -9333
rect 5667 -9367 5690 -9333
rect 5310 -9370 5690 -9367
rect 5310 -9390 5390 -9370
rect 5610 -9390 5690 -9370
rect 6060 -9380 6100 -9330
rect 6240 -9380 6320 -9360
rect 6060 -9383 6320 -9380
rect 5460 -9430 5540 -9410
rect 5310 -9433 5540 -9430
rect 5310 -9453 5483 -9433
rect 5310 -9487 5333 -9453
rect 5367 -9467 5483 -9453
rect 5517 -9467 5540 -9433
rect 5367 -9470 5540 -9467
rect 5367 -9487 5390 -9470
rect 5310 -9510 5390 -9487
rect 5460 -9490 5540 -9470
rect 6060 -9417 6263 -9383
rect 6297 -9417 6320 -9383
rect 6060 -9420 6320 -9417
rect 6060 -9550 6100 -9420
rect 6240 -9440 6320 -9420
rect 4480 -9590 5202 -9550
rect 5430 -9590 6100 -9550
rect 6140 -9500 6220 -9485
rect 6360 -9500 6400 -9330
rect 6640 -9380 6720 -9360
rect 6640 -9383 7227 -9380
rect 6640 -9417 6663 -9383
rect 6697 -9417 7227 -9383
rect 6640 -9420 7227 -9417
rect 6640 -9440 6720 -9420
rect 7073 -9500 7153 -9480
rect 6140 -9503 7153 -9500
rect 6140 -9508 7096 -9503
rect 6140 -9542 6163 -9508
rect 6197 -9537 7096 -9508
rect 7130 -9537 7153 -9503
rect 6197 -9540 7153 -9537
rect 6197 -9542 6220 -9540
rect 6140 -9565 6220 -9542
rect 3850 -9630 3890 -9590
rect 4180 -9630 4220 -9590
rect 3314 -9711 3646 -9708
rect 3314 -9745 3337 -9711
rect 3371 -9745 3646 -9711
rect 3314 -9748 3646 -9745
rect 3680 -9663 3760 -9630
rect 3680 -9697 3703 -9663
rect 3737 -9697 3760 -9663
rect 3680 -9743 3760 -9697
rect 3314 -9769 3394 -9748
rect 3200 -9823 3280 -9777
rect 3200 -9857 3223 -9823
rect 3257 -9857 3280 -9823
rect 3200 -9880 3280 -9857
rect 3680 -9777 3703 -9743
rect 3737 -9777 3760 -9743
rect 3680 -9823 3760 -9777
rect 3680 -9857 3703 -9823
rect 3737 -9857 3760 -9823
rect 3680 -9880 3760 -9857
rect 3830 -9663 3910 -9630
rect 3830 -9697 3853 -9663
rect 3887 -9697 3910 -9663
rect 3830 -9743 3910 -9697
rect 3830 -9777 3853 -9743
rect 3887 -9777 3910 -9743
rect 3830 -9823 3910 -9777
rect 3830 -9857 3853 -9823
rect 3887 -9857 3910 -9823
rect 3830 -9880 3910 -9857
rect 4010 -9663 4090 -9630
rect 4010 -9697 4033 -9663
rect 4067 -9697 4090 -9663
rect 4010 -9743 4090 -9697
rect 4010 -9777 4033 -9743
rect 4067 -9777 4090 -9743
rect 4010 -9823 4090 -9777
rect 4010 -9857 4033 -9823
rect 4067 -9857 4090 -9823
rect 4010 -9880 4090 -9857
rect 4160 -9663 4240 -9630
rect 4160 -9697 4183 -9663
rect 4217 -9697 4240 -9663
rect 4160 -9743 4240 -9697
rect 4160 -9777 4183 -9743
rect 4217 -9777 4240 -9743
rect 4160 -9823 4240 -9777
rect 4160 -9857 4183 -9823
rect 4217 -9857 4240 -9823
rect 4160 -9880 4240 -9857
rect 4310 -9663 4390 -9630
rect 4310 -9697 4333 -9663
rect 4367 -9697 4390 -9663
rect 4310 -9743 4390 -9697
rect 4310 -9777 4333 -9743
rect 4367 -9777 4390 -9743
rect 4310 -9823 4390 -9777
rect 4310 -9857 4333 -9823
rect 4367 -9857 4390 -9823
rect 4310 -9880 4390 -9857
rect 4460 -9663 4540 -9590
rect 4810 -9630 4850 -9590
rect 5430 -9630 5470 -9590
rect 5730 -9630 5770 -9590
rect 6061 -9630 6100 -9590
rect 6360 -9630 6400 -9540
rect 6690 -9630 6730 -9540
rect 7073 -9560 7153 -9540
rect 4460 -9697 4483 -9663
rect 4517 -9697 4540 -9663
rect 4460 -9743 4540 -9697
rect 4460 -9777 4483 -9743
rect 4517 -9777 4540 -9743
rect 4460 -9823 4540 -9777
rect 4460 -9857 4483 -9823
rect 4517 -9857 4540 -9823
rect 4460 -9880 4540 -9857
rect 4610 -9663 4690 -9630
rect 4610 -9697 4633 -9663
rect 4667 -9697 4690 -9663
rect 4610 -9743 4690 -9697
rect 4610 -9777 4633 -9743
rect 4667 -9777 4690 -9743
rect 4610 -9823 4690 -9777
rect 4610 -9857 4633 -9823
rect 4667 -9857 4690 -9823
rect 4610 -9880 4690 -9857
rect 4790 -9663 4870 -9630
rect 4790 -9697 4813 -9663
rect 4847 -9697 4870 -9663
rect 4790 -9743 4870 -9697
rect 4790 -9777 4813 -9743
rect 4847 -9777 4870 -9743
rect 4790 -9823 4870 -9777
rect 4790 -9857 4813 -9823
rect 4847 -9857 4870 -9823
rect 4790 -9880 4870 -9857
rect 4940 -9663 5020 -9630
rect 4940 -9697 4963 -9663
rect 4997 -9697 5020 -9663
rect 4940 -9743 5020 -9697
rect 4940 -9777 4963 -9743
rect 4997 -9777 5020 -9743
rect 4940 -9823 5020 -9777
rect 4940 -9857 4963 -9823
rect 4997 -9857 5020 -9823
rect 4940 -9880 5020 -9857
rect 5410 -9663 5490 -9630
rect 5410 -9697 5433 -9663
rect 5467 -9697 5490 -9663
rect 5410 -9743 5490 -9697
rect 5410 -9777 5433 -9743
rect 5467 -9777 5490 -9743
rect 5410 -9823 5490 -9777
rect 5410 -9857 5433 -9823
rect 5467 -9857 5490 -9823
rect 5410 -9880 5490 -9857
rect 5560 -9663 5640 -9630
rect 5560 -9697 5583 -9663
rect 5617 -9697 5640 -9663
rect 5560 -9743 5640 -9697
rect 5560 -9777 5583 -9743
rect 5617 -9777 5640 -9743
rect 5560 -9823 5640 -9777
rect 5560 -9857 5583 -9823
rect 5617 -9857 5640 -9823
rect 5560 -9880 5640 -9857
rect 5710 -9663 5790 -9630
rect 5710 -9697 5733 -9663
rect 5767 -9697 5790 -9663
rect 5710 -9743 5790 -9697
rect 5710 -9777 5733 -9743
rect 5767 -9777 5790 -9743
rect 5710 -9823 5790 -9777
rect 5710 -9857 5733 -9823
rect 5767 -9857 5790 -9823
rect 5710 -9880 5790 -9857
rect 5890 -9663 5970 -9630
rect 5890 -9697 5913 -9663
rect 5947 -9697 5970 -9663
rect 5890 -9743 5970 -9697
rect 5890 -9777 5913 -9743
rect 5947 -9777 5970 -9743
rect 5890 -9823 5970 -9777
rect 5890 -9857 5913 -9823
rect 5947 -9857 5970 -9823
rect 5890 -9880 5970 -9857
rect 6040 -9663 6120 -9630
rect 6040 -9697 6063 -9663
rect 6097 -9697 6120 -9663
rect 6040 -9743 6120 -9697
rect 6040 -9777 6063 -9743
rect 6097 -9777 6120 -9743
rect 6040 -9823 6120 -9777
rect 6040 -9857 6063 -9823
rect 6097 -9857 6120 -9823
rect 6040 -9880 6120 -9857
rect 6190 -9663 6270 -9630
rect 6190 -9697 6213 -9663
rect 6247 -9697 6270 -9663
rect 6190 -9743 6270 -9697
rect 6190 -9777 6213 -9743
rect 6247 -9777 6270 -9743
rect 6190 -9823 6270 -9777
rect 6190 -9857 6213 -9823
rect 6247 -9857 6270 -9823
rect 6190 -9880 6270 -9857
rect 6340 -9663 6420 -9630
rect 6340 -9697 6363 -9663
rect 6397 -9697 6420 -9663
rect 6340 -9743 6420 -9697
rect 6340 -9777 6363 -9743
rect 6397 -9777 6420 -9743
rect 6340 -9823 6420 -9777
rect 6340 -9857 6363 -9823
rect 6397 -9857 6420 -9823
rect 6340 -9880 6420 -9857
rect 6490 -9663 6570 -9630
rect 6490 -9697 6513 -9663
rect 6547 -9697 6570 -9663
rect 6490 -9743 6570 -9697
rect 6490 -9777 6513 -9743
rect 6547 -9777 6570 -9743
rect 6490 -9823 6570 -9777
rect 6490 -9857 6513 -9823
rect 6547 -9857 6570 -9823
rect 6490 -9880 6570 -9857
rect 6670 -9663 6750 -9630
rect 6670 -9697 6693 -9663
rect 6727 -9697 6750 -9663
rect 6670 -9743 6750 -9697
rect 6670 -9777 6693 -9743
rect 6727 -9777 6750 -9743
rect 6670 -9823 6750 -9777
rect 6670 -9857 6693 -9823
rect 6727 -9857 6750 -9823
rect 6670 -9880 6750 -9857
rect 6970 -9663 7050 -9630
rect 6970 -9697 6993 -9663
rect 7027 -9697 7050 -9663
rect 6970 -9743 7050 -9697
rect 6970 -9777 6993 -9743
rect 7027 -9777 7050 -9743
rect 6970 -9823 7050 -9777
rect 6970 -9857 6993 -9823
rect 7027 -9857 7050 -9823
rect 6970 -9880 7050 -9857
rect 1171 -9940 1251 -9920
rect 1920 -9940 2000 -9920
rect 2320 -9940 2400 -9920
rect 4110 -9940 4190 -9920
rect 4510 -9940 4590 -9920
rect 5398 -9940 5478 -9920
rect 5990 -9940 6070 -9920
rect 6390 -9940 6470 -9920
rect 1020 -9943 4590 -9940
rect 1020 -9977 1194 -9943
rect 1228 -9977 1943 -9943
rect 1977 -9977 2343 -9943
rect 2377 -9977 4133 -9943
rect 4167 -9977 4533 -9943
rect 4567 -9977 4590 -9943
rect 1020 -9980 4590 -9977
rect 5390 -9943 6470 -9940
rect 5390 -9977 5421 -9943
rect 5455 -9977 6013 -9943
rect 6047 -9977 6413 -9943
rect 6447 -9977 6470 -9943
rect 5390 -9980 6470 -9977
rect 1171 -10000 1251 -9980
rect 1920 -10000 2000 -9980
rect 2320 -10000 2400 -9980
rect 4110 -10000 4190 -9980
rect 4510 -10000 4590 -9980
rect 5398 -10000 5478 -9980
rect 5990 -10000 6070 -9980
rect 6390 -10000 6470 -9980
rect 912 -10063 3300 -10040
rect 912 -10097 935 -10063
rect 969 -10097 1103 -10063
rect 1137 -10097 1183 -10063
rect 1217 -10097 1263 -10063
rect 1297 -10097 1343 -10063
rect 1377 -10097 1423 -10063
rect 1457 -10097 1503 -10063
rect 1537 -10097 1583 -10063
rect 1617 -10097 1663 -10063
rect 1697 -10097 1743 -10063
rect 1777 -10097 1823 -10063
rect 1857 -10097 1903 -10063
rect 1937 -10097 1983 -10063
rect 2017 -10097 2063 -10063
rect 2097 -10097 2143 -10063
rect 2177 -10097 2223 -10063
rect 2257 -10097 2303 -10063
rect 2337 -10097 2383 -10063
rect 2417 -10097 2463 -10063
rect 2497 -10097 2543 -10063
rect 2577 -10097 2623 -10063
rect 2657 -10097 2703 -10063
rect 2737 -10097 2783 -10063
rect 2817 -10097 2863 -10063
rect 2897 -10097 2943 -10063
rect 2977 -10097 3023 -10063
rect 3057 -10097 3103 -10063
rect 3137 -10097 3183 -10063
rect 3217 -10097 3300 -10063
rect 912 -10120 3300 -10097
rect 3660 -10063 5040 -10040
rect 3660 -10097 3693 -10063
rect 3727 -10097 3773 -10063
rect 3807 -10097 3853 -10063
rect 3887 -10097 3933 -10063
rect 3967 -10097 4013 -10063
rect 4047 -10097 4093 -10063
rect 4127 -10097 4173 -10063
rect 4207 -10097 4253 -10063
rect 4287 -10097 4333 -10063
rect 4367 -10097 4413 -10063
rect 4447 -10097 4493 -10063
rect 4527 -10097 4573 -10063
rect 4607 -10097 4653 -10063
rect 4687 -10097 4733 -10063
rect 4767 -10097 4813 -10063
rect 4847 -10097 4893 -10063
rect 4927 -10097 4973 -10063
rect 5007 -10097 5040 -10063
rect 3660 -10120 5040 -10097
rect 5390 -10063 7070 -10040
rect 5390 -10097 5413 -10063
rect 5447 -10097 5493 -10063
rect 5527 -10097 5573 -10063
rect 5607 -10097 5653 -10063
rect 5687 -10097 5733 -10063
rect 5767 -10097 5813 -10063
rect 5847 -10097 5893 -10063
rect 5927 -10097 5973 -10063
rect 6007 -10097 6053 -10063
rect 6087 -10097 6133 -10063
rect 6167 -10097 6213 -10063
rect 6247 -10097 6293 -10063
rect 6327 -10097 6373 -10063
rect 6407 -10097 6453 -10063
rect 6487 -10097 6533 -10063
rect 6567 -10097 6613 -10063
rect 6647 -10097 6693 -10063
rect 6727 -10097 6773 -10063
rect 6807 -10097 6853 -10063
rect 6887 -10097 6933 -10063
rect 6967 -10097 7013 -10063
rect 7047 -10097 7070 -10063
rect 5390 -10120 7070 -10097
rect 1171 -10180 1251 -10160
rect 1920 -10180 2000 -10160
rect 2320 -10180 2400 -10160
rect 4110 -10180 4190 -10160
rect 4510 -10180 4590 -10160
rect 5398 -10180 5478 -10159
rect 5990 -10180 6070 -10160
rect 6390 -10180 6470 -10160
rect 1020 -10183 4590 -10180
rect 1020 -10217 1194 -10183
rect 1228 -10217 1943 -10183
rect 1977 -10217 2343 -10183
rect 2377 -10217 4133 -10183
rect 4167 -10217 4533 -10183
rect 4567 -10217 4590 -10183
rect 1020 -10220 4590 -10217
rect 5390 -10182 6470 -10180
rect 5390 -10216 5421 -10182
rect 5455 -10183 6470 -10182
rect 5455 -10216 6013 -10183
rect 5390 -10217 6013 -10216
rect 6047 -10217 6413 -10183
rect 6447 -10217 6470 -10183
rect 5390 -10220 6470 -10217
rect 1171 -10240 1251 -10220
rect 1920 -10240 2000 -10220
rect 2320 -10240 2400 -10220
rect 4110 -10240 4190 -10220
rect 4510 -10240 4590 -10220
rect 5398 -10239 5478 -10220
rect 5990 -10240 6070 -10220
rect 6390 -10240 6470 -10220
rect 1040 -10303 1120 -10280
rect 1040 -10337 1063 -10303
rect 1097 -10337 1120 -10303
rect 1040 -10383 1120 -10337
rect 1040 -10417 1063 -10383
rect 1097 -10417 1120 -10383
rect 1040 -10463 1120 -10417
rect 1040 -10497 1063 -10463
rect 1097 -10497 1120 -10463
rect 1040 -10530 1120 -10497
rect 1340 -10303 1420 -10280
rect 1340 -10337 1363 -10303
rect 1397 -10337 1420 -10303
rect 1340 -10383 1420 -10337
rect 1340 -10417 1363 -10383
rect 1397 -10417 1420 -10383
rect 1340 -10463 1420 -10417
rect 1340 -10497 1363 -10463
rect 1397 -10497 1420 -10463
rect 1340 -10530 1420 -10497
rect 1640 -10303 1720 -10280
rect 1640 -10337 1663 -10303
rect 1697 -10337 1720 -10303
rect 1640 -10383 1720 -10337
rect 1640 -10417 1663 -10383
rect 1697 -10417 1720 -10383
rect 1640 -10463 1720 -10417
rect 1640 -10497 1663 -10463
rect 1697 -10497 1720 -10463
rect 1640 -10530 1720 -10497
rect 1820 -10303 1900 -10280
rect 1820 -10337 1843 -10303
rect 1877 -10337 1900 -10303
rect 1820 -10383 1900 -10337
rect 1820 -10417 1843 -10383
rect 1877 -10417 1900 -10383
rect 1820 -10463 1900 -10417
rect 1820 -10497 1843 -10463
rect 1877 -10497 1900 -10463
rect 1820 -10530 1900 -10497
rect 1970 -10303 2050 -10280
rect 1970 -10337 1993 -10303
rect 2027 -10337 2050 -10303
rect 1970 -10383 2050 -10337
rect 1970 -10417 1993 -10383
rect 2027 -10417 2050 -10383
rect 1970 -10463 2050 -10417
rect 1970 -10497 1993 -10463
rect 2027 -10497 2050 -10463
rect 1970 -10530 2050 -10497
rect 2120 -10303 2200 -10280
rect 2120 -10337 2143 -10303
rect 2177 -10337 2200 -10303
rect 2120 -10383 2200 -10337
rect 2120 -10417 2143 -10383
rect 2177 -10417 2200 -10383
rect 2120 -10463 2200 -10417
rect 2120 -10497 2143 -10463
rect 2177 -10497 2200 -10463
rect 2120 -10530 2200 -10497
rect 2270 -10303 2350 -10280
rect 2270 -10337 2293 -10303
rect 2327 -10337 2350 -10303
rect 2270 -10383 2350 -10337
rect 2270 -10417 2293 -10383
rect 2327 -10417 2350 -10383
rect 2270 -10463 2350 -10417
rect 2270 -10497 2293 -10463
rect 2327 -10497 2350 -10463
rect 2270 -10530 2350 -10497
rect 2420 -10303 2500 -10280
rect 2420 -10337 2443 -10303
rect 2477 -10337 2500 -10303
rect 2420 -10383 2500 -10337
rect 2420 -10417 2443 -10383
rect 2477 -10417 2500 -10383
rect 2420 -10463 2500 -10417
rect 2420 -10497 2443 -10463
rect 2477 -10497 2500 -10463
rect 2420 -10530 2500 -10497
rect 2600 -10303 2680 -10280
rect 2600 -10337 2623 -10303
rect 2657 -10337 2680 -10303
rect 2600 -10383 2680 -10337
rect 2600 -10417 2623 -10383
rect 2657 -10417 2680 -10383
rect 2600 -10463 2680 -10417
rect 2600 -10497 2623 -10463
rect 2657 -10497 2680 -10463
rect 2600 -10530 2680 -10497
rect 2900 -10303 2980 -10280
rect 2900 -10337 2923 -10303
rect 2957 -10337 2980 -10303
rect 2900 -10383 2980 -10337
rect 2900 -10417 2923 -10383
rect 2957 -10417 2980 -10383
rect 2900 -10463 2980 -10417
rect 2900 -10497 2923 -10463
rect 2957 -10497 2980 -10463
rect 2900 -10530 2980 -10497
rect 3200 -10303 3280 -10280
rect 3200 -10337 3223 -10303
rect 3257 -10337 3280 -10303
rect 3200 -10383 3280 -10337
rect 3200 -10417 3223 -10383
rect 3257 -10417 3280 -10383
rect 3680 -10303 3760 -10280
rect 3680 -10337 3703 -10303
rect 3737 -10337 3760 -10303
rect 3680 -10383 3760 -10337
rect 3200 -10463 3280 -10417
rect 3200 -10497 3223 -10463
rect 3257 -10497 3280 -10463
rect 3314 -10403 3394 -10384
rect 3314 -10406 3646 -10403
rect 3314 -10440 3337 -10406
rect 3371 -10440 3646 -10406
rect 3314 -10443 3646 -10440
rect 3314 -10464 3394 -10443
rect 3200 -10530 3280 -10497
rect 1060 -10570 1100 -10530
rect 1660 -10570 1700 -10530
rect 1990 -10570 2030 -10530
rect 1060 -10610 2030 -10570
rect 1990 -10740 2030 -10610
rect 2070 -10618 2150 -10595
rect 2070 -10652 2093 -10618
rect 2127 -10620 2150 -10618
rect 2290 -10620 2330 -10530
rect 2620 -10620 2660 -10530
rect 3220 -10620 3260 -10530
rect 3606 -10620 3646 -10443
rect 3680 -10417 3703 -10383
rect 3737 -10417 3760 -10383
rect 3680 -10463 3760 -10417
rect 3680 -10497 3703 -10463
rect 3737 -10497 3760 -10463
rect 3680 -10530 3760 -10497
rect 3830 -10303 3910 -10280
rect 3830 -10337 3853 -10303
rect 3887 -10337 3910 -10303
rect 3830 -10383 3910 -10337
rect 3830 -10417 3853 -10383
rect 3887 -10417 3910 -10383
rect 3830 -10463 3910 -10417
rect 3830 -10497 3853 -10463
rect 3887 -10497 3910 -10463
rect 3830 -10530 3910 -10497
rect 4010 -10303 4090 -10280
rect 4010 -10337 4033 -10303
rect 4067 -10337 4090 -10303
rect 4010 -10383 4090 -10337
rect 4010 -10417 4033 -10383
rect 4067 -10417 4090 -10383
rect 4010 -10463 4090 -10417
rect 4010 -10497 4033 -10463
rect 4067 -10497 4090 -10463
rect 4010 -10530 4090 -10497
rect 4160 -10303 4240 -10280
rect 4160 -10337 4183 -10303
rect 4217 -10337 4240 -10303
rect 4160 -10383 4240 -10337
rect 4160 -10417 4183 -10383
rect 4217 -10417 4240 -10383
rect 4160 -10463 4240 -10417
rect 4160 -10497 4183 -10463
rect 4217 -10497 4240 -10463
rect 4160 -10530 4240 -10497
rect 4310 -10303 4390 -10280
rect 4310 -10337 4333 -10303
rect 4367 -10337 4390 -10303
rect 4310 -10383 4390 -10337
rect 4310 -10417 4333 -10383
rect 4367 -10417 4390 -10383
rect 4310 -10463 4390 -10417
rect 4310 -10497 4333 -10463
rect 4367 -10497 4390 -10463
rect 4310 -10530 4390 -10497
rect 4460 -10303 4540 -10280
rect 4460 -10337 4483 -10303
rect 4517 -10337 4540 -10303
rect 4460 -10383 4540 -10337
rect 4460 -10417 4483 -10383
rect 4517 -10417 4540 -10383
rect 4460 -10463 4540 -10417
rect 4460 -10497 4483 -10463
rect 4517 -10497 4540 -10463
rect 3850 -10570 3890 -10530
rect 4180 -10570 4220 -10530
rect 4460 -10570 4540 -10497
rect 4610 -10303 4690 -10280
rect 4610 -10337 4633 -10303
rect 4667 -10337 4690 -10303
rect 4610 -10383 4690 -10337
rect 4610 -10417 4633 -10383
rect 4667 -10417 4690 -10383
rect 4610 -10463 4690 -10417
rect 4610 -10497 4633 -10463
rect 4667 -10497 4690 -10463
rect 4610 -10530 4690 -10497
rect 4790 -10303 4870 -10280
rect 4790 -10337 4813 -10303
rect 4847 -10337 4870 -10303
rect 4790 -10383 4870 -10337
rect 4790 -10417 4813 -10383
rect 4847 -10417 4870 -10383
rect 4790 -10463 4870 -10417
rect 4790 -10497 4813 -10463
rect 4847 -10497 4870 -10463
rect 4790 -10530 4870 -10497
rect 4940 -10303 5020 -10280
rect 4940 -10337 4963 -10303
rect 4997 -10337 5020 -10303
rect 4940 -10383 5020 -10337
rect 4940 -10417 4963 -10383
rect 4997 -10417 5020 -10383
rect 4940 -10463 5020 -10417
rect 4940 -10497 4963 -10463
rect 4997 -10497 5020 -10463
rect 4940 -10530 5020 -10497
rect 5410 -10303 5490 -10280
rect 5410 -10337 5433 -10303
rect 5467 -10337 5490 -10303
rect 5410 -10383 5490 -10337
rect 5410 -10417 5433 -10383
rect 5467 -10417 5490 -10383
rect 5410 -10463 5490 -10417
rect 5410 -10497 5433 -10463
rect 5467 -10497 5490 -10463
rect 5410 -10530 5490 -10497
rect 5560 -10303 5640 -10280
rect 5560 -10337 5583 -10303
rect 5617 -10337 5640 -10303
rect 5560 -10383 5640 -10337
rect 5560 -10417 5583 -10383
rect 5617 -10417 5640 -10383
rect 5560 -10463 5640 -10417
rect 5560 -10497 5583 -10463
rect 5617 -10497 5640 -10463
rect 5560 -10530 5640 -10497
rect 5710 -10303 5790 -10280
rect 5710 -10337 5733 -10303
rect 5767 -10337 5790 -10303
rect 5710 -10383 5790 -10337
rect 5710 -10417 5733 -10383
rect 5767 -10417 5790 -10383
rect 5710 -10463 5790 -10417
rect 5710 -10497 5733 -10463
rect 5767 -10497 5790 -10463
rect 5710 -10530 5790 -10497
rect 5890 -10303 5970 -10280
rect 5890 -10337 5913 -10303
rect 5947 -10337 5970 -10303
rect 5890 -10383 5970 -10337
rect 5890 -10417 5913 -10383
rect 5947 -10417 5970 -10383
rect 5890 -10463 5970 -10417
rect 5890 -10497 5913 -10463
rect 5947 -10497 5970 -10463
rect 5890 -10530 5970 -10497
rect 6040 -10303 6120 -10280
rect 6040 -10337 6063 -10303
rect 6097 -10337 6120 -10303
rect 6040 -10383 6120 -10337
rect 6040 -10417 6063 -10383
rect 6097 -10417 6120 -10383
rect 6040 -10463 6120 -10417
rect 6040 -10497 6063 -10463
rect 6097 -10497 6120 -10463
rect 6040 -10530 6120 -10497
rect 6190 -10303 6270 -10280
rect 6190 -10337 6213 -10303
rect 6247 -10337 6270 -10303
rect 6190 -10383 6270 -10337
rect 6190 -10417 6213 -10383
rect 6247 -10417 6270 -10383
rect 6190 -10463 6270 -10417
rect 6190 -10497 6213 -10463
rect 6247 -10497 6270 -10463
rect 6190 -10530 6270 -10497
rect 6340 -10303 6420 -10280
rect 6340 -10337 6363 -10303
rect 6397 -10337 6420 -10303
rect 6340 -10383 6420 -10337
rect 6340 -10417 6363 -10383
rect 6397 -10417 6420 -10383
rect 6340 -10463 6420 -10417
rect 6340 -10497 6363 -10463
rect 6397 -10497 6420 -10463
rect 6340 -10530 6420 -10497
rect 6490 -10303 6570 -10280
rect 6490 -10337 6513 -10303
rect 6547 -10337 6570 -10303
rect 6490 -10383 6570 -10337
rect 6490 -10417 6513 -10383
rect 6547 -10417 6570 -10383
rect 6490 -10463 6570 -10417
rect 6490 -10497 6513 -10463
rect 6547 -10497 6570 -10463
rect 6490 -10530 6570 -10497
rect 6670 -10303 6750 -10280
rect 6670 -10337 6693 -10303
rect 6727 -10337 6750 -10303
rect 6670 -10383 6750 -10337
rect 6670 -10417 6693 -10383
rect 6727 -10417 6750 -10383
rect 6670 -10463 6750 -10417
rect 6670 -10497 6693 -10463
rect 6727 -10497 6750 -10463
rect 6670 -10530 6750 -10497
rect 6970 -10303 7050 -10280
rect 6970 -10337 6993 -10303
rect 7027 -10337 7050 -10303
rect 6970 -10383 7050 -10337
rect 6970 -10417 6993 -10383
rect 7027 -10417 7050 -10383
rect 6970 -10463 7050 -10417
rect 6970 -10497 6993 -10463
rect 7027 -10497 7050 -10463
rect 6970 -10530 7050 -10497
rect 4810 -10570 4850 -10530
rect 5048 -10570 5128 -10550
rect 3730 -10620 3810 -10600
rect 3850 -10610 4220 -10570
rect 4480 -10573 5128 -10570
rect 2127 -10652 3505 -10620
rect 2070 -10660 3505 -10652
rect 3606 -10623 3810 -10620
rect 3606 -10657 3753 -10623
rect 3787 -10657 3810 -10623
rect 3606 -10660 3810 -10657
rect 2070 -10675 2150 -10660
rect 2170 -10740 2250 -10720
rect 1990 -10743 2250 -10740
rect 1990 -10777 2193 -10743
rect 2227 -10777 2250 -10743
rect 1990 -10780 2250 -10777
rect 798 -10810 878 -10790
rect 1090 -10810 1170 -10790
rect 1670 -10810 1750 -10790
rect 798 -10813 1750 -10810
rect 798 -10847 821 -10813
rect 855 -10847 1113 -10813
rect 1147 -10847 1693 -10813
rect 1727 -10847 1750 -10813
rect 1990 -10830 2030 -10780
rect 2170 -10800 2250 -10780
rect 2290 -10830 2330 -10660
rect 2540 -10733 3380 -10710
rect 2540 -10767 2563 -10733
rect 2597 -10750 3323 -10733
rect 2597 -10767 2620 -10750
rect 2540 -10790 2620 -10767
rect 3300 -10767 3323 -10750
rect 3357 -10767 3380 -10733
rect 3300 -10790 3380 -10767
rect 2700 -10813 2780 -10790
rect 798 -10850 1750 -10847
rect 798 -10870 878 -10850
rect 1090 -10870 1170 -10850
rect 1670 -10870 1750 -10850
rect 1820 -10863 1900 -10840
rect 684 -10910 764 -10890
rect 1540 -10910 1620 -10890
rect 684 -10913 1620 -10910
rect 684 -10947 707 -10913
rect 741 -10947 1563 -10913
rect 1597 -10947 1620 -10913
rect 684 -10950 1620 -10947
rect 684 -10970 764 -10950
rect 1540 -10970 1620 -10950
rect 1820 -10897 1843 -10863
rect 1877 -10897 1900 -10863
rect 1820 -10943 1900 -10897
rect 1820 -10977 1843 -10943
rect 1877 -10977 1900 -10943
rect 570 -11010 650 -10990
rect 1290 -11010 1370 -10990
rect 1670 -11010 1750 -10990
rect 570 -11013 1750 -11010
rect 570 -11047 593 -11013
rect 627 -11047 1313 -11013
rect 1347 -11047 1693 -11013
rect 1727 -11047 1750 -11013
rect 570 -11050 1750 -11047
rect 570 -11070 650 -11050
rect 1290 -11070 1370 -11050
rect 1670 -11070 1750 -11050
rect 1820 -11023 1900 -10977
rect 1820 -11057 1843 -11023
rect 1877 -11057 1900 -11023
rect 1820 -11090 1900 -11057
rect 1970 -10863 2050 -10830
rect 1970 -10897 1993 -10863
rect 2027 -10897 2050 -10863
rect 1970 -10943 2050 -10897
rect 1970 -10977 1993 -10943
rect 2027 -10977 2050 -10943
rect 1970 -11023 2050 -10977
rect 1970 -11057 1993 -11023
rect 2027 -11057 2050 -11023
rect 1970 -11090 2050 -11057
rect 2120 -10863 2200 -10840
rect 2120 -10897 2143 -10863
rect 2177 -10897 2200 -10863
rect 2120 -10943 2200 -10897
rect 2120 -10977 2143 -10943
rect 2177 -10977 2200 -10943
rect 2120 -11023 2200 -10977
rect 2120 -11057 2143 -11023
rect 2177 -11057 2200 -11023
rect 2120 -11090 2200 -11057
rect 2270 -10863 2350 -10830
rect 2270 -10897 2293 -10863
rect 2327 -10897 2350 -10863
rect 2270 -10943 2350 -10897
rect 2270 -10977 2293 -10943
rect 2327 -10977 2350 -10943
rect 2270 -11023 2350 -10977
rect 2270 -11057 2293 -11023
rect 2327 -11057 2350 -11023
rect 2270 -11090 2350 -11057
rect 2420 -10863 2500 -10840
rect 2420 -10897 2443 -10863
rect 2477 -10897 2500 -10863
rect 2700 -10847 2723 -10813
rect 2757 -10847 2780 -10813
rect 2700 -10870 2780 -10847
rect 2420 -10943 2500 -10897
rect 2420 -10977 2443 -10943
rect 2477 -10977 2500 -10943
rect 3150 -10913 3230 -10890
rect 3150 -10947 3173 -10913
rect 3207 -10947 3230 -10913
rect 3150 -10970 3230 -10947
rect 2420 -11023 2500 -10977
rect 2420 -11057 2443 -11023
rect 2477 -11057 2500 -11023
rect 2420 -11090 2500 -11057
rect 3000 -11013 3080 -10990
rect 3000 -11047 3023 -11013
rect 3057 -11047 3080 -11013
rect 3000 -11070 3080 -11047
rect 3465 -11042 3505 -10660
rect 3730 -10680 3810 -10660
rect 4180 -10740 4220 -10610
rect 4260 -10618 4340 -10595
rect 4260 -10652 4283 -10618
rect 4317 -10620 4340 -10618
rect 4480 -10607 5071 -10573
rect 5105 -10607 5128 -10573
rect 4480 -10610 5128 -10607
rect 5430 -10570 5470 -10530
rect 5730 -10570 5770 -10530
rect 6061 -10570 6100 -10530
rect 5430 -10610 6100 -10570
rect 4480 -10620 4520 -10610
rect 4317 -10652 4520 -10620
rect 5048 -10630 5128 -10610
rect 4260 -10660 4520 -10652
rect 4260 -10675 4340 -10660
rect 4360 -10740 4440 -10720
rect 4180 -10743 4440 -10740
rect 4180 -10777 4383 -10743
rect 4417 -10777 4440 -10743
rect 4180 -10780 4440 -10777
rect 4180 -10830 4220 -10780
rect 4360 -10800 4440 -10780
rect 4480 -10830 4520 -10660
rect 5460 -10690 5540 -10670
rect 5020 -10693 5540 -10690
rect 4760 -10740 4840 -10720
rect 5020 -10727 5483 -10693
rect 5517 -10727 5540 -10693
rect 5020 -10730 5540 -10727
rect 5020 -10740 5060 -10730
rect 4760 -10743 5060 -10740
rect 4760 -10777 4783 -10743
rect 4817 -10777 5060 -10743
rect 5460 -10750 5540 -10730
rect 6060 -10740 6100 -10610
rect 6140 -10618 6220 -10595
rect 6140 -10652 6163 -10618
rect 6197 -10620 6220 -10618
rect 6360 -10620 6400 -10530
rect 6690 -10620 6730 -10530
rect 7073 -10620 7153 -10600
rect 6197 -10623 7153 -10620
rect 6197 -10652 7096 -10623
rect 6140 -10657 7096 -10652
rect 7130 -10657 7153 -10623
rect 6140 -10660 7153 -10657
rect 6140 -10675 6220 -10660
rect 6240 -10740 6320 -10720
rect 6060 -10743 6320 -10740
rect 4760 -10780 5060 -10777
rect 4760 -10800 4840 -10780
rect 5610 -10790 5690 -10770
rect 5162 -10793 5690 -10790
rect 5162 -10827 5633 -10793
rect 5667 -10827 5690 -10793
rect 5162 -10830 5690 -10827
rect 6060 -10777 6263 -10743
rect 6297 -10777 6320 -10743
rect 6060 -10780 6320 -10777
rect 6060 -10830 6100 -10780
rect 6240 -10800 6320 -10780
rect 6360 -10830 6400 -10660
rect 7073 -10680 7153 -10660
rect 6640 -10740 6720 -10720
rect 6640 -10743 7144 -10740
rect 6640 -10777 6663 -10743
rect 6697 -10777 7144 -10743
rect 6640 -10780 7144 -10777
rect 6640 -10800 6720 -10780
rect 3860 -10860 3940 -10840
rect 3660 -10863 3940 -10860
rect 3660 -10897 3883 -10863
rect 3917 -10897 3940 -10863
rect 3660 -10900 3940 -10897
rect 3860 -10920 3940 -10900
rect 4010 -10863 4090 -10840
rect 4010 -10897 4033 -10863
rect 4067 -10897 4090 -10863
rect 4010 -10943 4090 -10897
rect 4010 -10977 4033 -10943
rect 4067 -10977 4090 -10943
rect 4010 -11023 4090 -10977
rect 3572 -11042 3652 -11024
rect 3465 -11047 3652 -11042
rect 3465 -11081 3595 -11047
rect 3629 -11081 3652 -11047
rect 3465 -11082 3652 -11081
rect 456 -11110 536 -11090
rect 1410 -11110 1490 -11090
rect 1540 -11110 1620 -11090
rect 456 -11113 1620 -11110
rect 456 -11147 479 -11113
rect 513 -11147 1433 -11113
rect 1467 -11147 1563 -11113
rect 1597 -11147 1620 -11113
rect 456 -11150 1620 -11147
rect 456 -11170 536 -11150
rect 1410 -11170 1490 -11150
rect 1540 -11170 1620 -11150
rect 2800 -11113 2880 -11090
rect 3572 -11104 3652 -11082
rect 4010 -11057 4033 -11023
rect 4067 -11057 4090 -11023
rect 4010 -11090 4090 -11057
rect 4160 -10863 4240 -10830
rect 4160 -10897 4183 -10863
rect 4217 -10897 4240 -10863
rect 4160 -10943 4240 -10897
rect 4160 -10977 4183 -10943
rect 4217 -10977 4240 -10943
rect 4160 -11023 4240 -10977
rect 4160 -11057 4183 -11023
rect 4217 -11057 4240 -11023
rect 4160 -11090 4240 -11057
rect 4310 -10863 4390 -10840
rect 4310 -10897 4333 -10863
rect 4367 -10897 4390 -10863
rect 4310 -10943 4390 -10897
rect 4310 -10977 4333 -10943
rect 4367 -10977 4390 -10943
rect 4310 -11023 4390 -10977
rect 4310 -11057 4333 -11023
rect 4367 -11057 4390 -11023
rect 4310 -11090 4390 -11057
rect 4460 -10863 4540 -10830
rect 4460 -10897 4483 -10863
rect 4517 -10897 4540 -10863
rect 4460 -10943 4540 -10897
rect 4460 -10977 4483 -10943
rect 4517 -10977 4540 -10943
rect 4460 -11023 4540 -10977
rect 4460 -11057 4483 -11023
rect 4517 -11057 4540 -11023
rect 4460 -11090 4540 -11057
rect 4610 -10863 4690 -10840
rect 4610 -10897 4633 -10863
rect 4667 -10897 4690 -10863
rect 4610 -10943 4690 -10897
rect 4760 -10860 4840 -10840
rect 4890 -10860 4970 -10840
rect 4760 -10863 4970 -10860
rect 4760 -10897 4783 -10863
rect 4817 -10897 4913 -10863
rect 4947 -10897 4970 -10863
rect 4760 -10900 4970 -10897
rect 4760 -10920 4840 -10900
rect 4890 -10920 4970 -10900
rect 5048 -10898 5128 -10878
rect 5162 -10898 5202 -10830
rect 5610 -10850 5690 -10830
rect 5890 -10863 5970 -10840
rect 5048 -10901 5202 -10898
rect 4610 -10977 4633 -10943
rect 4667 -10977 4690 -10943
rect 5048 -10935 5071 -10901
rect 5105 -10935 5202 -10901
rect 5048 -10938 5202 -10935
rect 5310 -10890 5390 -10870
rect 5740 -10890 5820 -10870
rect 5310 -10893 5820 -10890
rect 5310 -10927 5333 -10893
rect 5367 -10927 5763 -10893
rect 5797 -10927 5820 -10893
rect 5310 -10930 5820 -10927
rect 5048 -10958 5128 -10938
rect 5310 -10950 5390 -10930
rect 5740 -10950 5820 -10930
rect 5890 -10897 5913 -10863
rect 5947 -10897 5970 -10863
rect 5890 -10943 5970 -10897
rect 4610 -11023 4690 -10977
rect 5890 -10977 5913 -10943
rect 5947 -10977 5970 -10943
rect 4610 -11057 4633 -11023
rect 4667 -11057 4690 -11023
rect 4610 -11090 4690 -11057
rect 5310 -11010 5390 -10991
rect 5740 -11010 5820 -10990
rect 5310 -11013 5820 -11010
rect 5310 -11014 5763 -11013
rect 5310 -11048 5333 -11014
rect 5367 -11047 5763 -11014
rect 5797 -11047 5820 -11013
rect 5367 -11048 5820 -11047
rect 5310 -11050 5820 -11048
rect 5310 -11071 5390 -11050
rect 5740 -11070 5820 -11050
rect 5890 -11023 5970 -10977
rect 5890 -11057 5913 -11023
rect 5947 -11057 5970 -11023
rect 5890 -11090 5970 -11057
rect 6040 -10863 6120 -10830
rect 6040 -10897 6063 -10863
rect 6097 -10897 6120 -10863
rect 6040 -10943 6120 -10897
rect 6040 -10977 6063 -10943
rect 6097 -10977 6120 -10943
rect 6040 -11023 6120 -10977
rect 6040 -11057 6063 -11023
rect 6097 -11057 6120 -11023
rect 6040 -11090 6120 -11057
rect 6190 -10863 6270 -10840
rect 6190 -10897 6213 -10863
rect 6247 -10897 6270 -10863
rect 6190 -10943 6270 -10897
rect 6190 -10977 6213 -10943
rect 6247 -10977 6270 -10943
rect 6190 -11023 6270 -10977
rect 6190 -11057 6213 -11023
rect 6247 -11057 6270 -11023
rect 6190 -11090 6270 -11057
rect 6340 -10863 6420 -10830
rect 6340 -10897 6363 -10863
rect 6397 -10897 6420 -10863
rect 6340 -10943 6420 -10897
rect 6340 -10977 6363 -10943
rect 6397 -10977 6420 -10943
rect 6340 -11023 6420 -10977
rect 6340 -11057 6363 -11023
rect 6397 -11057 6420 -11023
rect 6340 -11090 6420 -11057
rect 6490 -10863 6570 -10840
rect 6490 -10897 6513 -10863
rect 6547 -10897 6570 -10863
rect 6490 -10943 6570 -10897
rect 6490 -10977 6513 -10943
rect 6547 -10977 6570 -10943
rect 6720 -10893 6800 -10870
rect 6720 -10927 6743 -10893
rect 6777 -10927 6800 -10893
rect 6720 -10950 6800 -10927
rect 6490 -11023 6570 -10977
rect 6490 -11057 6513 -11023
rect 6547 -11057 6570 -11023
rect 6490 -11090 6570 -11057
rect 6870 -11013 6950 -10990
rect 6870 -11047 6893 -11013
rect 6927 -11047 6950 -11013
rect 6870 -11070 6950 -11047
rect 2800 -11147 2823 -11113
rect 2857 -11147 2880 -11113
rect 2800 -11170 2880 -11147
rect 1020 -11243 3300 -11220
rect 1020 -11277 1103 -11243
rect 1137 -11277 1183 -11243
rect 1217 -11277 1263 -11243
rect 1297 -11277 1343 -11243
rect 1377 -11277 1423 -11243
rect 1457 -11277 1503 -11243
rect 1537 -11277 1583 -11243
rect 1617 -11277 1663 -11243
rect 1697 -11277 1743 -11243
rect 1777 -11277 1823 -11243
rect 1857 -11277 1903 -11243
rect 1937 -11277 1983 -11243
rect 2017 -11277 2063 -11243
rect 2097 -11277 2143 -11243
rect 2177 -11277 2223 -11243
rect 2257 -11277 2303 -11243
rect 2337 -11277 2383 -11243
rect 2417 -11277 2463 -11243
rect 2497 -11277 2543 -11243
rect 2577 -11277 2623 -11243
rect 2657 -11277 2703 -11243
rect 2737 -11277 2783 -11243
rect 2817 -11277 2863 -11243
rect 2897 -11277 2943 -11243
rect 2977 -11277 3023 -11243
rect 3057 -11277 3103 -11243
rect 3137 -11277 3183 -11243
rect 3217 -11277 3300 -11243
rect 1020 -11300 3300 -11277
rect 3660 -11243 5040 -11220
rect 3660 -11277 3693 -11243
rect 3727 -11277 3773 -11243
rect 3807 -11277 3853 -11243
rect 3887 -11277 3933 -11243
rect 3967 -11277 4013 -11243
rect 4047 -11277 4093 -11243
rect 4127 -11277 4173 -11243
rect 4207 -11277 4253 -11243
rect 4287 -11277 4333 -11243
rect 4367 -11277 4413 -11243
rect 4447 -11277 4493 -11243
rect 4527 -11277 4573 -11243
rect 4607 -11277 4653 -11243
rect 4687 -11277 4733 -11243
rect 4767 -11277 4813 -11243
rect 4847 -11277 4893 -11243
rect 4927 -11277 4973 -11243
rect 5007 -11277 5040 -11243
rect 3660 -11300 5040 -11277
rect 5390 -11243 7070 -11220
rect 5390 -11277 5413 -11243
rect 5447 -11277 5493 -11243
rect 5527 -11277 5573 -11243
rect 5607 -11277 5653 -11243
rect 5687 -11277 5733 -11243
rect 5767 -11277 5813 -11243
rect 5847 -11277 5893 -11243
rect 5927 -11277 5973 -11243
rect 6007 -11277 6053 -11243
rect 6087 -11277 6133 -11243
rect 6167 -11277 6213 -11243
rect 6247 -11277 6293 -11243
rect 6327 -11277 6373 -11243
rect 6407 -11277 6453 -11243
rect 6487 -11277 6533 -11243
rect 6567 -11277 6613 -11243
rect 6647 -11277 6693 -11243
rect 6727 -11277 6773 -11243
rect 6807 -11277 6853 -11243
rect 6887 -11277 6933 -11243
rect 6967 -11277 7013 -11243
rect 7047 -11277 7070 -11243
rect 5390 -11300 7070 -11277
rect 5398 -11474 5478 -11454
rect 5024 -11477 5478 -11474
rect 5024 -11511 5421 -11477
rect 5455 -11511 5478 -11477
rect 5024 -11514 5478 -11511
rect 1161 -11703 3161 -11680
rect 1161 -11737 1184 -11703
rect 1218 -11737 1264 -11703
rect 1298 -11737 1344 -11703
rect 1378 -11737 1424 -11703
rect 1458 -11737 1504 -11703
rect 1538 -11737 1584 -11703
rect 1618 -11737 1664 -11703
rect 1698 -11737 1744 -11703
rect 1778 -11737 1824 -11703
rect 1858 -11737 1904 -11703
rect 1938 -11737 1984 -11703
rect 2018 -11737 2064 -11703
rect 2098 -11737 2144 -11703
rect 2178 -11737 2224 -11703
rect 2258 -11737 2304 -11703
rect 2338 -11737 2384 -11703
rect 2418 -11737 2464 -11703
rect 2498 -11737 2544 -11703
rect 2578 -11737 2624 -11703
rect 2658 -11737 2704 -11703
rect 2738 -11737 2784 -11703
rect 2818 -11737 2864 -11703
rect 2898 -11737 2944 -11703
rect 2978 -11737 3024 -11703
rect 3058 -11737 3104 -11703
rect 3138 -11737 3161 -11703
rect 1161 -11760 3161 -11737
rect 3521 -11703 4901 -11680
rect 3521 -11737 3554 -11703
rect 3588 -11737 3634 -11703
rect 3668 -11737 3714 -11703
rect 3748 -11737 3794 -11703
rect 3828 -11737 3874 -11703
rect 3908 -11737 3954 -11703
rect 3988 -11737 4034 -11703
rect 4068 -11737 4114 -11703
rect 4148 -11737 4194 -11703
rect 4228 -11737 4274 -11703
rect 4308 -11737 4354 -11703
rect 4388 -11737 4434 -11703
rect 4468 -11737 4514 -11703
rect 4548 -11737 4594 -11703
rect 4628 -11737 4674 -11703
rect 4708 -11737 4754 -11703
rect 4788 -11737 4834 -11703
rect 4868 -11737 4901 -11703
rect 3521 -11760 4901 -11737
rect 570 -11820 650 -11800
rect 1581 -11820 1661 -11800
rect 570 -11823 1661 -11820
rect 570 -11857 593 -11823
rect 627 -11857 1604 -11823
rect 1638 -11857 1661 -11823
rect 570 -11860 1661 -11857
rect 570 -11880 650 -11860
rect 1581 -11880 1661 -11860
rect 2951 -11823 3031 -11800
rect 2951 -11857 2974 -11823
rect 3008 -11857 3031 -11823
rect 2951 -11880 3031 -11857
rect 5024 -11887 5064 -11514
rect 5398 -11534 5478 -11514
rect 7104 -11601 7144 -10780
rect 7187 -11508 7227 -9420
rect 7343 -11508 7423 -11487
rect 7187 -11510 7423 -11508
rect 7187 -11544 7366 -11510
rect 7400 -11544 7423 -11510
rect 7187 -11548 7423 -11544
rect 7343 -11567 7423 -11548
rect 7104 -11641 7429 -11601
rect 5251 -11704 7251 -11681
rect 5251 -11738 5274 -11704
rect 5308 -11738 5354 -11704
rect 5388 -11738 5434 -11704
rect 5468 -11738 5514 -11704
rect 5548 -11738 5594 -11704
rect 5628 -11738 5674 -11704
rect 5708 -11738 5754 -11704
rect 5788 -11738 5834 -11704
rect 5868 -11738 5914 -11704
rect 5948 -11738 5994 -11704
rect 6028 -11738 6074 -11704
rect 6108 -11738 6154 -11704
rect 6188 -11738 6234 -11704
rect 6268 -11738 6314 -11704
rect 6348 -11738 6394 -11704
rect 6428 -11738 6474 -11704
rect 6508 -11738 6554 -11704
rect 6588 -11738 6634 -11704
rect 6668 -11738 6714 -11704
rect 6748 -11738 6794 -11704
rect 6828 -11738 6874 -11704
rect 6908 -11738 6954 -11704
rect 6988 -11738 7034 -11704
rect 7068 -11738 7114 -11704
rect 7148 -11738 7194 -11704
rect 7228 -11738 7251 -11704
rect 5251 -11761 7251 -11738
rect 5381 -11829 5461 -11806
rect 5381 -11863 5404 -11829
rect 5438 -11863 5461 -11829
rect 5381 -11886 5461 -11863
rect 6661 -11831 6741 -11811
rect 7229 -11831 7309 -11811
rect 6661 -11834 7309 -11831
rect 6661 -11868 6684 -11834
rect 6718 -11868 7252 -11834
rect 7286 -11868 7309 -11834
rect 6661 -11871 7309 -11868
rect 0 -11940 80 -11920
rect 1671 -11940 1751 -11920
rect 0 -11943 1751 -11940
rect 0 -11977 23 -11943
rect 57 -11977 1694 -11943
rect 1728 -11977 1751 -11943
rect 0 -11980 1751 -11977
rect 0 -12000 80 -11980
rect 1671 -12000 1751 -11980
rect 1821 -11923 1901 -11890
rect 1821 -11957 1844 -11923
rect 1878 -11957 1901 -11923
rect 1821 -12003 1901 -11957
rect 684 -12039 764 -12016
rect 684 -12073 707 -12039
rect 741 -12050 764 -12039
rect 1821 -12037 1844 -12003
rect 1878 -12037 1901 -12003
rect 1641 -12050 1721 -12040
rect 741 -12063 1721 -12050
rect 741 -12073 1664 -12063
rect 684 -12090 1664 -12073
rect 684 -12096 764 -12090
rect 456 -12119 536 -12096
rect 456 -12153 479 -12119
rect 513 -12130 536 -12119
rect 1641 -12097 1664 -12090
rect 1698 -12097 1721 -12063
rect 1641 -12120 1721 -12097
rect 1821 -12083 1901 -12037
rect 1821 -12117 1844 -12083
rect 1878 -12117 1901 -12083
rect 513 -12153 1601 -12130
rect 1821 -12140 1901 -12117
rect 1971 -11923 2051 -11890
rect 1971 -11957 1994 -11923
rect 2028 -11957 2051 -11923
rect 1971 -12003 2051 -11957
rect 1971 -12037 1994 -12003
rect 2028 -12037 2051 -12003
rect 1971 -12083 2051 -12037
rect 1971 -12117 1994 -12083
rect 2028 -12117 2051 -12083
rect 1971 -12150 2051 -12117
rect 2121 -11923 2201 -11890
rect 2121 -11957 2144 -11923
rect 2178 -11957 2201 -11923
rect 2121 -12003 2201 -11957
rect 2121 -12037 2144 -12003
rect 2178 -12037 2201 -12003
rect 2121 -12083 2201 -12037
rect 2121 -12117 2144 -12083
rect 2178 -12117 2201 -12083
rect 2121 -12140 2201 -12117
rect 2271 -11923 2351 -11890
rect 2271 -11957 2294 -11923
rect 2328 -11957 2351 -11923
rect 2271 -12003 2351 -11957
rect 2271 -12037 2294 -12003
rect 2328 -12037 2351 -12003
rect 2271 -12083 2351 -12037
rect 2271 -12117 2294 -12083
rect 2328 -12117 2351 -12083
rect 2271 -12150 2351 -12117
rect 2421 -11923 2501 -11890
rect 2421 -11957 2444 -11923
rect 2478 -11957 2501 -11923
rect 2421 -12003 2501 -11957
rect 2801 -11943 2881 -11920
rect 2801 -11977 2824 -11943
rect 2858 -11977 2881 -11943
rect 2801 -12000 2881 -11977
rect 3871 -11923 3951 -11890
rect 3871 -11957 3894 -11923
rect 3928 -11957 3951 -11923
rect 2421 -12037 2444 -12003
rect 2478 -12037 2501 -12003
rect 2421 -12083 2501 -12037
rect 3871 -12003 3951 -11957
rect 3871 -12037 3894 -12003
rect 3928 -12037 3951 -12003
rect 2421 -12117 2444 -12083
rect 2478 -12117 2501 -12083
rect 2421 -12140 2501 -12117
rect 2671 -12063 2751 -12040
rect 2671 -12097 2694 -12063
rect 2728 -12097 2751 -12063
rect 2671 -12120 2751 -12097
rect 3433 -12080 3513 -12060
rect 3721 -12080 3801 -12060
rect 3433 -12083 3801 -12080
rect 3433 -12117 3456 -12083
rect 3490 -12117 3744 -12083
rect 3778 -12117 3801 -12083
rect 3433 -12120 3801 -12117
rect 3433 -12140 3513 -12120
rect 3721 -12140 3801 -12120
rect 3871 -12083 3951 -12037
rect 3871 -12117 3894 -12083
rect 3928 -12117 3951 -12083
rect 3871 -12140 3951 -12117
rect 4021 -11923 4101 -11890
rect 4021 -11957 4044 -11923
rect 4078 -11957 4101 -11923
rect 4021 -12003 4101 -11957
rect 4021 -12037 4044 -12003
rect 4078 -12037 4101 -12003
rect 4021 -12083 4101 -12037
rect 4021 -12117 4044 -12083
rect 4078 -12117 4101 -12083
rect 4021 -12150 4101 -12117
rect 4171 -11923 4251 -11890
rect 4171 -11957 4194 -11923
rect 4228 -11957 4251 -11923
rect 4171 -12003 4251 -11957
rect 4171 -12037 4194 -12003
rect 4228 -12037 4251 -12003
rect 4171 -12083 4251 -12037
rect 4171 -12117 4194 -12083
rect 4228 -12117 4251 -12083
rect 4171 -12140 4251 -12117
rect 4321 -11923 4401 -11890
rect 4321 -11957 4344 -11923
rect 4378 -11957 4401 -11923
rect 4321 -12003 4401 -11957
rect 4321 -12037 4344 -12003
rect 4378 -12037 4401 -12003
rect 4321 -12083 4401 -12037
rect 4321 -12117 4344 -12083
rect 4378 -12117 4401 -12083
rect 4321 -12150 4401 -12117
rect 4471 -11923 4551 -11890
rect 4471 -11957 4494 -11923
rect 4528 -11957 4551 -11923
rect 4471 -12003 4551 -11957
rect 5004 -11910 5084 -11887
rect 6661 -11891 6741 -11871
rect 7229 -11891 7309 -11871
rect 5004 -11944 5027 -11910
rect 5061 -11944 5084 -11910
rect 5911 -11924 5991 -11891
rect 5004 -11967 5084 -11944
rect 5481 -11954 5561 -11931
rect 4471 -12037 4494 -12003
rect 4528 -12037 4551 -12003
rect 5481 -11988 5504 -11954
rect 5538 -11988 5561 -11954
rect 5481 -12011 5561 -11988
rect 5911 -11958 5934 -11924
rect 5968 -11958 5991 -11924
rect 5911 -12004 5991 -11958
rect 4471 -12083 4551 -12037
rect 5681 -12044 5761 -12021
rect 4471 -12117 4494 -12083
rect 4528 -12117 4551 -12083
rect 4471 -12140 4551 -12117
rect 4621 -12080 4701 -12060
rect 4751 -12080 4831 -12060
rect 4621 -12083 4831 -12080
rect 5681 -12078 5704 -12044
rect 5738 -12078 5761 -12044
rect 4621 -12117 4644 -12083
rect 4678 -12117 4774 -12083
rect 4808 -12117 4831 -12083
rect 5180 -12103 5260 -12083
rect 5681 -12101 5761 -12078
rect 5911 -12038 5934 -12004
rect 5968 -12038 5991 -12004
rect 5911 -12084 5991 -12038
rect 4621 -12120 4831 -12117
rect 4621 -12140 4701 -12120
rect 4751 -12140 4831 -12120
rect 5066 -12106 5260 -12103
rect 5066 -12140 5203 -12106
rect 5237 -12140 5260 -12106
rect 5066 -12143 5260 -12140
rect 5911 -12118 5934 -12084
rect 5968 -12118 5991 -12084
rect 5911 -12141 5991 -12118
rect 6061 -11924 6141 -11891
rect 6061 -11958 6084 -11924
rect 6118 -11958 6141 -11924
rect 6061 -12004 6141 -11958
rect 6061 -12038 6084 -12004
rect 6118 -12038 6141 -12004
rect 6061 -12084 6141 -12038
rect 6061 -12118 6084 -12084
rect 6118 -12118 6141 -12084
rect 456 -12170 1601 -12153
rect 456 -12176 536 -12170
rect 1541 -12190 1601 -12170
rect 114 -12210 194 -12190
rect 114 -12213 1451 -12210
rect 114 -12247 137 -12213
rect 171 -12233 1451 -12213
rect 171 -12247 1394 -12233
rect 114 -12250 1394 -12247
rect 114 -12270 194 -12250
rect 1371 -12267 1394 -12250
rect 1428 -12267 1451 -12233
rect 1371 -12290 1451 -12267
rect 1541 -12213 1621 -12190
rect 1541 -12247 1564 -12213
rect 1598 -12247 1621 -12213
rect 1541 -12270 1621 -12247
rect 1991 -12200 2031 -12150
rect 2171 -12200 2251 -12180
rect 1991 -12203 2251 -12200
rect 1991 -12237 2194 -12203
rect 2228 -12237 2251 -12203
rect 1991 -12240 2251 -12237
rect 798 -12310 878 -12290
rect 1241 -12310 1321 -12290
rect 798 -12313 1321 -12310
rect 798 -12347 821 -12313
rect 855 -12347 1264 -12313
rect 1298 -12347 1321 -12313
rect 798 -12350 1321 -12347
rect 798 -12370 878 -12350
rect 1241 -12370 1321 -12350
rect 1991 -12370 2031 -12240
rect 2171 -12260 2251 -12240
rect 1361 -12410 2031 -12370
rect 2071 -12320 2151 -12305
rect 2291 -12320 2331 -12150
rect 2571 -12200 2651 -12180
rect 4041 -12200 4081 -12150
rect 4221 -12200 4301 -12180
rect 2571 -12203 3354 -12200
rect 2571 -12237 2594 -12203
rect 2628 -12237 3354 -12203
rect 2571 -12240 3354 -12237
rect 2571 -12260 2651 -12240
rect 3151 -12320 3231 -12299
rect 2071 -12322 3231 -12320
rect 2071 -12328 3174 -12322
rect 2071 -12362 2094 -12328
rect 2128 -12356 3174 -12328
rect 3208 -12356 3231 -12322
rect 2128 -12360 3231 -12356
rect 3314 -12320 3354 -12240
rect 4041 -12203 4301 -12200
rect 4041 -12237 4244 -12203
rect 4278 -12237 4301 -12203
rect 4041 -12240 4301 -12237
rect 3591 -12320 3671 -12300
rect 3314 -12323 3671 -12320
rect 3314 -12357 3614 -12323
rect 3648 -12357 3671 -12323
rect 3314 -12360 3671 -12357
rect 2128 -12362 2151 -12360
rect 2071 -12385 2151 -12362
rect 1361 -12450 1401 -12410
rect 1661 -12450 1701 -12410
rect 1991 -12450 2031 -12410
rect 2291 -12450 2331 -12360
rect 2621 -12450 2661 -12360
rect 3151 -12379 3231 -12360
rect 3591 -12380 3671 -12360
rect 4041 -12370 4081 -12240
rect 4221 -12260 4301 -12240
rect 3711 -12410 4081 -12370
rect 4121 -12320 4201 -12305
rect 4341 -12320 4381 -12150
rect 4621 -12200 4701 -12180
rect 5066 -12200 5106 -12143
rect 5180 -12163 5260 -12143
rect 6061 -12151 6141 -12118
rect 6211 -11924 6291 -11891
rect 6211 -11958 6234 -11924
rect 6268 -11958 6291 -11924
rect 6211 -12004 6291 -11958
rect 6211 -12038 6234 -12004
rect 6268 -12038 6291 -12004
rect 6211 -12084 6291 -12038
rect 6211 -12118 6234 -12084
rect 6268 -12118 6291 -12084
rect 6211 -12141 6291 -12118
rect 6361 -11924 6441 -11891
rect 6361 -11958 6384 -11924
rect 6418 -11958 6441 -11924
rect 6361 -12004 6441 -11958
rect 6361 -12038 6384 -12004
rect 6418 -12038 6441 -12004
rect 6361 -12084 6441 -12038
rect 6361 -12118 6384 -12084
rect 6418 -12118 6441 -12084
rect 6361 -12151 6441 -12118
rect 6511 -11924 6591 -11891
rect 6511 -11958 6534 -11924
rect 6568 -11958 6591 -11924
rect 6511 -12004 6591 -11958
rect 6781 -11941 6861 -11921
rect 7033 -11941 7113 -11921
rect 6781 -11944 7241 -11941
rect 6781 -11978 6804 -11944
rect 6838 -11978 7056 -11944
rect 7090 -11978 7241 -11944
rect 6781 -11981 7241 -11978
rect 6781 -12001 6861 -11981
rect 7033 -12001 7113 -11981
rect 6511 -12038 6534 -12004
rect 6568 -12038 6591 -12004
rect 6511 -12084 6591 -12038
rect 6511 -12118 6534 -12084
rect 6568 -12118 6591 -12084
rect 6661 -12041 6741 -12021
rect 6661 -12044 7241 -12041
rect 6661 -12078 6684 -12044
rect 6718 -12078 7241 -12044
rect 6661 -12081 7241 -12078
rect 6661 -12101 6741 -12081
rect 6511 -12141 6591 -12118
rect 7275 -12131 7355 -12109
rect 7081 -12132 7355 -12131
rect 4621 -12203 5106 -12200
rect 4621 -12237 4644 -12203
rect 4678 -12237 5106 -12203
rect 4621 -12240 5106 -12237
rect 5181 -12201 5261 -12197
rect 5761 -12201 5841 -12181
rect 5181 -12204 5841 -12201
rect 5181 -12220 5784 -12204
rect 4621 -12260 4701 -12240
rect 5181 -12254 5204 -12220
rect 5238 -12238 5784 -12220
rect 5818 -12238 5841 -12204
rect 5238 -12241 5841 -12238
rect 5238 -12254 5261 -12241
rect 5181 -12277 5261 -12254
rect 5761 -12261 5841 -12241
rect 4121 -12328 4381 -12320
rect 4121 -12362 4144 -12328
rect 4178 -12360 4381 -12328
rect 5181 -12321 5261 -12311
rect 6081 -12321 6121 -12151
rect 6161 -12201 6241 -12181
rect 6381 -12201 6421 -12151
rect 6161 -12204 6421 -12201
rect 6161 -12238 6184 -12204
rect 6218 -12238 6421 -12204
rect 7081 -12154 7298 -12132
rect 7081 -12188 7104 -12154
rect 7138 -12166 7298 -12154
rect 7332 -12166 7355 -12132
rect 7138 -12171 7355 -12166
rect 7138 -12188 7161 -12171
rect 7081 -12211 7161 -12188
rect 7275 -12189 7355 -12171
rect 6161 -12241 6421 -12238
rect 6161 -12261 6241 -12241
rect 6261 -12321 6341 -12306
rect 5181 -12329 6341 -12321
rect 5181 -12334 6284 -12329
rect 4178 -12362 4201 -12360
rect 4121 -12385 4201 -12362
rect 4341 -12370 4381 -12360
rect 4915 -12370 4995 -12350
rect 4341 -12373 4995 -12370
rect 4341 -12407 4938 -12373
rect 4972 -12407 4995 -12373
rect 5181 -12368 5204 -12334
rect 5238 -12361 6284 -12334
rect 5238 -12368 5261 -12361
rect 5181 -12391 5261 -12368
rect 4341 -12410 4995 -12407
rect 3711 -12450 3751 -12410
rect 4041 -12450 4081 -12410
rect 1191 -12483 1271 -12450
rect 1191 -12517 1214 -12483
rect 1248 -12517 1271 -12483
rect 1191 -12563 1271 -12517
rect 1191 -12597 1214 -12563
rect 1248 -12597 1271 -12563
rect 1191 -12643 1271 -12597
rect 1191 -12677 1214 -12643
rect 1248 -12677 1271 -12643
rect 1191 -12700 1271 -12677
rect 1341 -12483 1421 -12450
rect 1341 -12517 1364 -12483
rect 1398 -12517 1421 -12483
rect 1341 -12563 1421 -12517
rect 1341 -12597 1364 -12563
rect 1398 -12597 1421 -12563
rect 1341 -12643 1421 -12597
rect 1341 -12677 1364 -12643
rect 1398 -12677 1421 -12643
rect 1341 -12700 1421 -12677
rect 1491 -12483 1571 -12450
rect 1491 -12517 1514 -12483
rect 1548 -12517 1571 -12483
rect 1491 -12563 1571 -12517
rect 1491 -12597 1514 -12563
rect 1548 -12597 1571 -12563
rect 1491 -12643 1571 -12597
rect 1491 -12677 1514 -12643
rect 1548 -12677 1571 -12643
rect 1491 -12700 1571 -12677
rect 1641 -12483 1721 -12450
rect 1641 -12517 1664 -12483
rect 1698 -12517 1721 -12483
rect 1641 -12563 1721 -12517
rect 1641 -12597 1664 -12563
rect 1698 -12597 1721 -12563
rect 1641 -12643 1721 -12597
rect 1641 -12677 1664 -12643
rect 1698 -12677 1721 -12643
rect 1641 -12700 1721 -12677
rect 1821 -12483 1901 -12450
rect 1821 -12517 1844 -12483
rect 1878 -12517 1901 -12483
rect 1821 -12563 1901 -12517
rect 1821 -12597 1844 -12563
rect 1878 -12597 1901 -12563
rect 1821 -12643 1901 -12597
rect 1821 -12677 1844 -12643
rect 1878 -12677 1901 -12643
rect 1821 -12700 1901 -12677
rect 1971 -12483 2051 -12450
rect 1971 -12517 1994 -12483
rect 2028 -12517 2051 -12483
rect 1971 -12563 2051 -12517
rect 1971 -12597 1994 -12563
rect 2028 -12597 2051 -12563
rect 1971 -12643 2051 -12597
rect 1971 -12677 1994 -12643
rect 2028 -12677 2051 -12643
rect 1971 -12700 2051 -12677
rect 2121 -12483 2201 -12450
rect 2121 -12517 2144 -12483
rect 2178 -12517 2201 -12483
rect 2121 -12563 2201 -12517
rect 2121 -12597 2144 -12563
rect 2178 -12597 2201 -12563
rect 2121 -12643 2201 -12597
rect 2121 -12677 2144 -12643
rect 2178 -12677 2201 -12643
rect 2121 -12700 2201 -12677
rect 2271 -12483 2351 -12450
rect 2271 -12517 2294 -12483
rect 2328 -12517 2351 -12483
rect 2271 -12563 2351 -12517
rect 2271 -12597 2294 -12563
rect 2328 -12597 2351 -12563
rect 2271 -12643 2351 -12597
rect 2271 -12677 2294 -12643
rect 2328 -12677 2351 -12643
rect 2271 -12700 2351 -12677
rect 2421 -12483 2501 -12450
rect 2421 -12517 2444 -12483
rect 2478 -12517 2501 -12483
rect 2421 -12563 2501 -12517
rect 2421 -12597 2444 -12563
rect 2478 -12597 2501 -12563
rect 2421 -12643 2501 -12597
rect 2421 -12677 2444 -12643
rect 2478 -12677 2501 -12643
rect 2421 -12700 2501 -12677
rect 2601 -12483 2681 -12450
rect 2601 -12517 2624 -12483
rect 2658 -12517 2681 -12483
rect 2601 -12563 2681 -12517
rect 2601 -12597 2624 -12563
rect 2658 -12597 2681 -12563
rect 2601 -12643 2681 -12597
rect 2601 -12677 2624 -12643
rect 2658 -12677 2681 -12643
rect 2601 -12700 2681 -12677
rect 3051 -12483 3131 -12450
rect 3051 -12517 3074 -12483
rect 3108 -12517 3131 -12483
rect 3051 -12563 3131 -12517
rect 3051 -12597 3074 -12563
rect 3108 -12597 3131 -12563
rect 3051 -12643 3131 -12597
rect 3051 -12677 3074 -12643
rect 3108 -12677 3131 -12643
rect 3051 -12700 3131 -12677
rect 3541 -12483 3621 -12450
rect 3541 -12517 3564 -12483
rect 3598 -12517 3621 -12483
rect 3541 -12563 3621 -12517
rect 3541 -12597 3564 -12563
rect 3598 -12597 3621 -12563
rect 3541 -12643 3621 -12597
rect 3541 -12677 3564 -12643
rect 3598 -12677 3621 -12643
rect 3541 -12700 3621 -12677
rect 3691 -12483 3771 -12450
rect 3691 -12517 3714 -12483
rect 3748 -12517 3771 -12483
rect 3691 -12563 3771 -12517
rect 3691 -12597 3714 -12563
rect 3748 -12597 3771 -12563
rect 3691 -12643 3771 -12597
rect 3691 -12677 3714 -12643
rect 3748 -12677 3771 -12643
rect 3691 -12700 3771 -12677
rect 3871 -12483 3951 -12450
rect 3871 -12517 3894 -12483
rect 3928 -12517 3951 -12483
rect 3871 -12563 3951 -12517
rect 3871 -12597 3894 -12563
rect 3928 -12597 3951 -12563
rect 3871 -12643 3951 -12597
rect 3871 -12677 3894 -12643
rect 3928 -12677 3951 -12643
rect 3871 -12700 3951 -12677
rect 4021 -12483 4101 -12450
rect 4021 -12517 4044 -12483
rect 4078 -12517 4101 -12483
rect 4021 -12563 4101 -12517
rect 4021 -12597 4044 -12563
rect 4078 -12597 4101 -12563
rect 4021 -12643 4101 -12597
rect 4021 -12677 4044 -12643
rect 4078 -12677 4101 -12643
rect 4021 -12700 4101 -12677
rect 4171 -12483 4251 -12450
rect 4171 -12517 4194 -12483
rect 4228 -12517 4251 -12483
rect 4171 -12563 4251 -12517
rect 4171 -12597 4194 -12563
rect 4228 -12597 4251 -12563
rect 4171 -12643 4251 -12597
rect 4171 -12677 4194 -12643
rect 4228 -12677 4251 -12643
rect 4171 -12700 4251 -12677
rect 4321 -12483 4401 -12410
rect 4671 -12450 4711 -12410
rect 4915 -12430 4995 -12410
rect 4321 -12517 4344 -12483
rect 4378 -12517 4401 -12483
rect 4321 -12563 4401 -12517
rect 4321 -12597 4344 -12563
rect 4378 -12597 4401 -12563
rect 4321 -12643 4401 -12597
rect 4321 -12677 4344 -12643
rect 4378 -12677 4401 -12643
rect 4321 -12700 4401 -12677
rect 4471 -12483 4551 -12450
rect 4471 -12517 4494 -12483
rect 4528 -12517 4551 -12483
rect 4471 -12563 4551 -12517
rect 4471 -12597 4494 -12563
rect 4528 -12597 4551 -12563
rect 4471 -12643 4551 -12597
rect 4471 -12677 4494 -12643
rect 4528 -12677 4551 -12643
rect 4471 -12700 4551 -12677
rect 4651 -12483 4731 -12450
rect 4651 -12517 4674 -12483
rect 4708 -12517 4731 -12483
rect 4651 -12563 4731 -12517
rect 4651 -12597 4674 -12563
rect 4708 -12597 4731 -12563
rect 4651 -12643 4731 -12597
rect 4651 -12677 4674 -12643
rect 4708 -12677 4731 -12643
rect 4651 -12700 4731 -12677
rect 4801 -12483 4881 -12450
rect 5451 -12451 5491 -12361
rect 5751 -12451 5791 -12361
rect 6081 -12451 6121 -12361
rect 6261 -12363 6284 -12361
rect 6318 -12363 6341 -12329
rect 6261 -12386 6341 -12363
rect 6381 -12371 6421 -12241
rect 6941 -12251 7021 -12231
rect 7389 -12251 7429 -11641
rect 6941 -12254 7429 -12251
rect 6941 -12288 6964 -12254
rect 6998 -12288 7429 -12254
rect 6941 -12291 7429 -12288
rect 6941 -12311 7021 -12291
rect 6791 -12334 6871 -12311
rect 6791 -12368 6814 -12334
rect 6848 -12351 6871 -12334
rect 6848 -12368 7241 -12351
rect 6381 -12411 6731 -12371
rect 6791 -12391 7241 -12368
rect 6381 -12451 6421 -12411
rect 6691 -12451 6731 -12411
rect 4801 -12517 4824 -12483
rect 4858 -12517 4881 -12483
rect 4801 -12563 4881 -12517
rect 4998 -12487 5078 -12464
rect 4998 -12521 5021 -12487
rect 5055 -12521 5078 -12487
rect 4998 -12544 5078 -12521
rect 5281 -12484 5361 -12451
rect 5281 -12518 5304 -12484
rect 5338 -12518 5361 -12484
rect 4801 -12597 4824 -12563
rect 4858 -12597 4881 -12563
rect 4801 -12643 4881 -12597
rect 4801 -12677 4824 -12643
rect 4858 -12677 4881 -12643
rect 4801 -12700 4881 -12677
rect 1171 -12760 1251 -12740
rect 1921 -12760 2001 -12740
rect 2321 -12760 2401 -12740
rect 3971 -12760 4051 -12740
rect 4371 -12760 4451 -12740
rect 5018 -12760 5058 -12544
rect 5281 -12564 5361 -12518
rect 5281 -12598 5304 -12564
rect 5338 -12598 5361 -12564
rect 5281 -12644 5361 -12598
rect 5281 -12678 5304 -12644
rect 5338 -12678 5361 -12644
rect 5281 -12701 5361 -12678
rect 5431 -12484 5511 -12451
rect 5431 -12518 5454 -12484
rect 5488 -12518 5511 -12484
rect 5431 -12564 5511 -12518
rect 5431 -12598 5454 -12564
rect 5488 -12598 5511 -12564
rect 5431 -12644 5511 -12598
rect 5431 -12678 5454 -12644
rect 5488 -12678 5511 -12644
rect 5431 -12701 5511 -12678
rect 5581 -12484 5661 -12451
rect 5581 -12518 5604 -12484
rect 5638 -12518 5661 -12484
rect 5581 -12564 5661 -12518
rect 5581 -12598 5604 -12564
rect 5638 -12598 5661 -12564
rect 5581 -12644 5661 -12598
rect 5581 -12678 5604 -12644
rect 5638 -12678 5661 -12644
rect 5581 -12701 5661 -12678
rect 5731 -12484 5811 -12451
rect 5731 -12518 5754 -12484
rect 5788 -12518 5811 -12484
rect 5731 -12564 5811 -12518
rect 5731 -12598 5754 -12564
rect 5788 -12598 5811 -12564
rect 5731 -12644 5811 -12598
rect 5731 -12678 5754 -12644
rect 5788 -12678 5811 -12644
rect 5731 -12701 5811 -12678
rect 5911 -12484 5991 -12451
rect 5911 -12518 5934 -12484
rect 5968 -12518 5991 -12484
rect 5911 -12564 5991 -12518
rect 5911 -12598 5934 -12564
rect 5968 -12598 5991 -12564
rect 5911 -12644 5991 -12598
rect 5911 -12678 5934 -12644
rect 5968 -12678 5991 -12644
rect 5911 -12701 5991 -12678
rect 6061 -12484 6141 -12451
rect 6061 -12518 6084 -12484
rect 6118 -12518 6141 -12484
rect 6061 -12564 6141 -12518
rect 6061 -12598 6084 -12564
rect 6118 -12598 6141 -12564
rect 6061 -12644 6141 -12598
rect 6061 -12678 6084 -12644
rect 6118 -12678 6141 -12644
rect 6061 -12701 6141 -12678
rect 6211 -12484 6291 -12451
rect 6211 -12518 6234 -12484
rect 6268 -12518 6291 -12484
rect 6211 -12564 6291 -12518
rect 6211 -12598 6234 -12564
rect 6268 -12598 6291 -12564
rect 6211 -12644 6291 -12598
rect 6211 -12678 6234 -12644
rect 6268 -12678 6291 -12644
rect 6211 -12701 6291 -12678
rect 6361 -12484 6441 -12451
rect 6361 -12518 6384 -12484
rect 6418 -12518 6441 -12484
rect 6361 -12564 6441 -12518
rect 6361 -12598 6384 -12564
rect 6418 -12598 6441 -12564
rect 6361 -12644 6441 -12598
rect 6361 -12678 6384 -12644
rect 6418 -12678 6441 -12644
rect 6361 -12701 6441 -12678
rect 6511 -12484 6591 -12451
rect 6511 -12518 6534 -12484
rect 6568 -12518 6591 -12484
rect 6511 -12564 6591 -12518
rect 6511 -12598 6534 -12564
rect 6568 -12598 6591 -12564
rect 6511 -12644 6591 -12598
rect 6511 -12678 6534 -12644
rect 6568 -12678 6591 -12644
rect 6511 -12701 6591 -12678
rect 6691 -12484 6771 -12451
rect 6691 -12518 6714 -12484
rect 6748 -12518 6771 -12484
rect 6691 -12564 6771 -12518
rect 6691 -12598 6714 -12564
rect 6748 -12598 6771 -12564
rect 6691 -12644 6771 -12598
rect 6691 -12678 6714 -12644
rect 6748 -12678 6771 -12644
rect 6691 -12701 6771 -12678
rect 7141 -12484 7221 -12451
rect 7141 -12518 7164 -12484
rect 7198 -12518 7221 -12484
rect 7141 -12564 7221 -12518
rect 7141 -12598 7164 -12564
rect 7198 -12598 7221 -12564
rect 7141 -12644 7221 -12598
rect 7141 -12678 7164 -12644
rect 7198 -12678 7221 -12644
rect 7141 -12701 7221 -12678
rect 1171 -12763 2401 -12760
rect 1171 -12797 1194 -12763
rect 1228 -12797 1944 -12763
rect 1978 -12797 2344 -12763
rect 2378 -12797 2401 -12763
rect 1171 -12800 2401 -12797
rect 3521 -12763 5058 -12760
rect 3521 -12797 3994 -12763
rect 4028 -12797 4394 -12763
rect 4428 -12797 5058 -12763
rect 3521 -12800 5058 -12797
rect 5092 -12761 5172 -12742
rect 6011 -12761 6091 -12741
rect 6411 -12761 6491 -12741
rect 5092 -12764 7241 -12761
rect 5092 -12765 6034 -12764
rect 5092 -12799 5115 -12765
rect 5149 -12798 6034 -12765
rect 6068 -12798 6434 -12764
rect 6468 -12798 7241 -12764
rect 5149 -12799 7241 -12798
rect 1171 -12820 1251 -12800
rect 1921 -12820 2001 -12800
rect 2321 -12820 2401 -12800
rect 3971 -12820 4051 -12800
rect 4371 -12820 4451 -12800
rect 5092 -12801 7241 -12799
rect 5092 -12822 5172 -12801
rect 6011 -12821 6091 -12801
rect 6411 -12821 6491 -12801
rect 912 -12883 3161 -12860
rect 912 -12917 935 -12883
rect 969 -12917 1184 -12883
rect 1218 -12917 1264 -12883
rect 1298 -12917 1344 -12883
rect 1378 -12917 1424 -12883
rect 1458 -12917 1504 -12883
rect 1538 -12917 1584 -12883
rect 1618 -12917 1664 -12883
rect 1698 -12917 1744 -12883
rect 1778 -12917 1824 -12883
rect 1858 -12917 1904 -12883
rect 1938 -12917 1984 -12883
rect 2018 -12917 2064 -12883
rect 2098 -12917 2144 -12883
rect 2178 -12917 2224 -12883
rect 2258 -12917 2304 -12883
rect 2338 -12917 2384 -12883
rect 2418 -12917 2464 -12883
rect 2498 -12917 2544 -12883
rect 2578 -12917 2624 -12883
rect 2658 -12917 2704 -12883
rect 2738 -12917 2784 -12883
rect 2818 -12917 2864 -12883
rect 2898 -12917 2944 -12883
rect 2978 -12917 3024 -12883
rect 3058 -12917 3104 -12883
rect 3138 -12917 3161 -12883
rect 912 -12940 3161 -12917
rect 3521 -12883 4901 -12860
rect 3521 -12917 3554 -12883
rect 3588 -12917 3634 -12883
rect 3668 -12917 3714 -12883
rect 3748 -12917 3794 -12883
rect 3828 -12917 3874 -12883
rect 3908 -12917 3954 -12883
rect 3988 -12917 4034 -12883
rect 4068 -12917 4114 -12883
rect 4148 -12917 4194 -12883
rect 4228 -12917 4274 -12883
rect 4308 -12917 4354 -12883
rect 4388 -12917 4434 -12883
rect 4468 -12917 4514 -12883
rect 4548 -12917 4594 -12883
rect 4628 -12917 4674 -12883
rect 4708 -12917 4754 -12883
rect 4788 -12917 4834 -12883
rect 4868 -12917 4901 -12883
rect 3521 -12940 4901 -12917
rect 5251 -12884 7251 -12861
rect 5251 -12918 5274 -12884
rect 5308 -12918 5354 -12884
rect 5388 -12918 5434 -12884
rect 5468 -12918 5514 -12884
rect 5548 -12918 5594 -12884
rect 5628 -12918 5674 -12884
rect 5708 -12918 5754 -12884
rect 5788 -12918 5834 -12884
rect 5868 -12918 5914 -12884
rect 5948 -12918 5994 -12884
rect 6028 -12918 6074 -12884
rect 6108 -12918 6154 -12884
rect 6188 -12918 6234 -12884
rect 6268 -12918 6314 -12884
rect 6348 -12918 6394 -12884
rect 6428 -12918 6474 -12884
rect 6508 -12918 6554 -12884
rect 6588 -12918 6634 -12884
rect 6668 -12918 6714 -12884
rect 6748 -12918 6794 -12884
rect 6828 -12918 6874 -12884
rect 6908 -12918 6954 -12884
rect 6988 -12918 7034 -12884
rect 7068 -12918 7114 -12884
rect 7148 -12918 7194 -12884
rect 7228 -12918 7251 -12884
rect 5251 -12941 7251 -12918
<< viali >>
rect 1103 2444 1137 2478
rect 1183 2444 1217 2478
rect 1263 2444 1297 2478
rect 1343 2444 1377 2478
rect 1423 2444 1457 2478
rect 1503 2444 1537 2478
rect 1583 2444 1617 2478
rect 1663 2444 1697 2478
rect 1743 2444 1777 2478
rect 1823 2444 1857 2478
rect 1903 2444 1937 2478
rect 1983 2444 2017 2478
rect 2063 2444 2097 2478
rect 2143 2444 2177 2478
rect 2223 2444 2257 2478
rect 2303 2444 2337 2478
rect 2383 2444 2417 2478
rect 2463 2444 2497 2478
rect 2543 2444 2577 2478
rect 2623 2444 2657 2478
rect 2703 2444 2737 2478
rect 2783 2444 2817 2478
rect 2863 2444 2897 2478
rect 2943 2444 2977 2478
rect 3023 2444 3057 2478
rect 3103 2444 3137 2478
rect 3183 2444 3217 2478
rect 3663 2444 3697 2478
rect 3743 2444 3777 2478
rect 3823 2444 3857 2478
rect 3903 2444 3937 2478
rect 3983 2444 4017 2478
rect 4063 2444 4097 2478
rect 4143 2444 4177 2478
rect 4223 2444 4257 2478
rect 4303 2444 4337 2478
rect 4383 2444 4417 2478
rect 4463 2444 4497 2478
rect 4543 2444 4577 2478
rect 4623 2444 4657 2478
rect 4703 2444 4737 2478
rect 4783 2444 4817 2478
rect 4863 2444 4897 2478
rect 4943 2444 4977 2478
rect 5023 2444 5057 2478
rect 5103 2444 5137 2478
rect 5183 2444 5217 2478
rect 5263 2444 5297 2478
rect 5683 2444 5717 2478
rect 5763 2444 5797 2478
rect 5843 2444 5877 2478
rect 5923 2444 5957 2478
rect 6003 2444 6037 2478
rect 6083 2444 6117 2478
rect 6163 2444 6197 2478
rect 6243 2444 6277 2478
rect 6323 2444 6357 2478
rect 6403 2444 6437 2478
rect 6483 2444 6517 2478
rect 6563 2444 6597 2478
rect 6643 2444 6677 2478
rect 6723 2444 6757 2478
rect 6803 2444 6837 2478
rect 6883 2444 6917 2478
rect 6963 2444 6997 2478
rect 7043 2444 7077 2478
rect 7123 2444 7157 2478
rect 7203 2444 7237 2478
rect 7283 2444 7317 2478
rect 23 2294 57 2328
rect 1563 2314 1597 2348
rect 2823 2314 2857 2348
rect 137 2194 171 2228
rect 1693 2214 1727 2248
rect 1843 2224 1877 2258
rect 707 2094 741 2128
rect 1563 2114 1597 2148
rect 1843 2144 1877 2178
rect 821 1994 855 2028
rect 1693 2014 1727 2048
rect 1843 2064 1877 2098
rect 2143 2224 2177 2258
rect 2143 2144 2177 2178
rect 2143 2064 2177 2098
rect 2443 2224 2477 2258
rect 3023 2214 3057 2248
rect 3583 2204 3617 2238
rect 4013 2184 4047 2218
rect 2443 2144 2477 2178
rect 2443 2064 2477 2098
rect 4163 2224 4197 2258
rect 3173 2114 3207 2148
rect 4163 2144 4197 2178
rect 3583 2084 3617 2118
rect 2193 1944 2227 1978
rect 2723 2014 2757 2048
rect 4013 2064 4047 2098
rect 3323 2022 3357 2056
rect 4163 2064 4197 2098
rect 4463 2224 4497 2258
rect 4463 2144 4497 2178
rect 4463 2064 4497 2098
rect 4763 2224 4797 2258
rect 4763 2144 4797 2178
rect 5193 2184 5227 2218
rect 5603 2214 5637 2248
rect 6033 2214 6067 2248
rect 6183 2224 6217 2258
rect 4763 2064 4797 2098
rect 4993 2064 5027 2098
rect 5273 2070 5307 2104
rect 6033 2094 6067 2128
rect 6183 2144 6217 2178
rect 6183 2064 6217 2098
rect 6483 2224 6517 2258
rect 6483 2144 6517 2178
rect 6483 2064 6517 2098
rect 6783 2224 6817 2258
rect 7163 2214 7197 2248
rect 6783 2144 6817 2178
rect 6783 2064 6817 2098
rect 7013 2094 7047 2128
rect 2563 1934 2597 1968
rect 3077 1934 3111 1968
rect 3583 1964 3617 1998
rect 4513 1944 4547 1978
rect 3323 1820 3357 1854
rect 3583 1844 3617 1878
rect 5603 1993 5637 2027
rect 4913 1944 4947 1978
rect 5273 1844 5307 1878
rect 6533 1944 6567 1978
rect 6933 1944 6967 1978
rect 7363 1944 7397 1978
rect 1363 1664 1397 1698
rect 1363 1584 1397 1618
rect 1363 1504 1397 1538
rect 1843 1664 1877 1698
rect 1843 1584 1877 1618
rect 1843 1504 1877 1538
rect 2143 1664 2177 1698
rect 2143 1584 2177 1618
rect 2143 1504 2177 1538
rect 2443 1664 2477 1698
rect 2443 1584 2477 1618
rect 2443 1504 2477 1538
rect 2923 1664 2957 1698
rect 2923 1584 2957 1618
rect 2923 1504 2957 1538
rect 3683 1664 3717 1698
rect 3683 1584 3717 1618
rect 3683 1504 3717 1538
rect 4163 1664 4197 1698
rect 4163 1584 4197 1618
rect 4163 1504 4197 1538
rect 4463 1664 4497 1698
rect 4463 1584 4497 1618
rect 4463 1504 4497 1538
rect 4763 1664 4797 1698
rect 4763 1584 4797 1618
rect 4763 1504 4797 1538
rect 5093 1664 5127 1698
rect 5093 1584 5127 1618
rect 5093 1504 5127 1538
rect 5853 1664 5887 1698
rect 5853 1584 5887 1618
rect 5853 1504 5887 1538
rect 6183 1664 6217 1698
rect 6183 1584 6217 1618
rect 6183 1504 6217 1538
rect 6483 1664 6517 1698
rect 6483 1584 6517 1618
rect 6483 1504 6517 1538
rect 6783 1664 6817 1698
rect 6783 1584 6817 1618
rect 6783 1504 6817 1538
rect 7263 1664 7297 1698
rect 7263 1584 7297 1618
rect 7263 1504 7297 1538
rect 1152 1384 1186 1418
rect 5765 1384 5799 1418
rect 935 1264 969 1298
rect 1103 1264 1137 1298
rect 1183 1264 1217 1298
rect 1263 1264 1297 1298
rect 1343 1264 1377 1298
rect 1423 1264 1457 1298
rect 1503 1264 1537 1298
rect 1583 1264 1617 1298
rect 1663 1264 1697 1298
rect 1743 1264 1777 1298
rect 1823 1264 1857 1298
rect 1903 1264 1937 1298
rect 1983 1264 2017 1298
rect 2063 1264 2097 1298
rect 2143 1264 2177 1298
rect 2223 1264 2257 1298
rect 2303 1264 2337 1298
rect 2383 1264 2417 1298
rect 2463 1264 2497 1298
rect 2543 1264 2577 1298
rect 2623 1264 2657 1298
rect 2703 1264 2737 1298
rect 2783 1264 2817 1298
rect 2863 1264 2897 1298
rect 2943 1264 2977 1298
rect 3023 1264 3057 1298
rect 3103 1264 3137 1298
rect 3183 1264 3217 1298
rect 3663 1264 3697 1298
rect 3743 1264 3777 1298
rect 3823 1264 3857 1298
rect 3903 1264 3937 1298
rect 3983 1264 4017 1298
rect 4063 1264 4097 1298
rect 4143 1264 4177 1298
rect 4223 1264 4257 1298
rect 4303 1264 4337 1298
rect 4383 1264 4417 1298
rect 4463 1264 4497 1298
rect 4543 1264 4577 1298
rect 4623 1264 4657 1298
rect 4703 1264 4737 1298
rect 4783 1264 4817 1298
rect 4863 1264 4897 1298
rect 4943 1264 4977 1298
rect 5023 1264 5057 1298
rect 5103 1264 5137 1298
rect 5183 1264 5217 1298
rect 5263 1264 5297 1298
rect 5683 1264 5717 1298
rect 5763 1264 5797 1298
rect 5843 1264 5877 1298
rect 5923 1264 5957 1298
rect 6003 1264 6037 1298
rect 6083 1264 6117 1298
rect 6163 1264 6197 1298
rect 6243 1264 6277 1298
rect 6323 1264 6357 1298
rect 6403 1264 6437 1298
rect 6483 1264 6517 1298
rect 6563 1264 6597 1298
rect 6643 1264 6677 1298
rect 6723 1264 6757 1298
rect 6803 1264 6837 1298
rect 6883 1264 6917 1298
rect 6963 1264 6997 1298
rect 7043 1264 7077 1298
rect 7123 1264 7157 1298
rect 7203 1264 7237 1298
rect 7283 1264 7317 1298
rect 1151 1144 1185 1178
rect 5096 1145 5130 1179
rect 5945 1144 5979 1178
rect 1513 1024 1547 1058
rect 1513 944 1547 978
rect 1513 864 1547 898
rect 1843 1024 1877 1058
rect 1843 944 1877 978
rect 1843 864 1877 898
rect 2143 1024 2177 1058
rect 2143 944 2177 978
rect 2143 864 2177 898
rect 2443 1024 2477 1058
rect 2443 944 2477 978
rect 2443 864 2477 898
rect 2923 1024 2957 1058
rect 2923 944 2957 978
rect 2923 864 2957 898
rect 3833 1024 3867 1058
rect 3833 944 3867 978
rect 3833 864 3867 898
rect 4163 1024 4197 1058
rect 4163 944 4197 978
rect 4163 864 4197 898
rect 4463 1024 4497 1058
rect 4463 944 4497 978
rect 4463 864 4497 898
rect 4763 1024 4797 1058
rect 4763 944 4797 978
rect 4763 864 4797 898
rect 5243 1024 5277 1058
rect 5243 944 5277 978
rect 5243 864 5277 898
rect 5853 1024 5887 1058
rect 5853 944 5887 978
rect 5853 864 5887 898
rect 6183 1024 6217 1058
rect 6183 944 6217 978
rect 6183 864 6217 898
rect 6483 1024 6517 1058
rect 6483 944 6517 978
rect 6483 864 6517 898
rect 6783 1024 6817 1058
rect 6783 944 6817 978
rect 6783 864 6817 898
rect 7263 1024 7297 1058
rect 7263 944 7297 978
rect 7113 854 7147 888
rect 7263 864 7297 898
rect 251 654 285 688
rect 3023 704 3057 738
rect 593 540 627 574
rect 2193 584 2227 618
rect 2593 584 2627 618
rect 3583 534 3617 568
rect 4513 584 4547 618
rect 4913 584 4947 618
rect 5494 584 5528 618
rect 365 434 399 468
rect 1693 434 1727 468
rect 1843 464 1877 498
rect 1843 384 1877 418
rect 479 314 513 348
rect 1693 314 1727 348
rect 1843 304 1877 338
rect 2143 464 2177 498
rect 2143 384 2177 418
rect 2143 304 2177 338
rect 2443 464 2477 498
rect 2443 384 2477 418
rect 2673 434 2707 468
rect 3023 454 3057 488
rect 4013 434 4047 468
rect 4163 464 4197 498
rect 4163 384 4197 418
rect 2443 304 2477 338
rect 2823 314 2857 348
rect 3077 314 3111 348
rect 4013 314 4047 348
rect 4163 304 4197 338
rect 4463 464 4497 498
rect 4463 384 4497 418
rect 4463 304 4497 338
rect 4763 464 4797 498
rect 5683 704 5717 738
rect 5683 584 5717 618
rect 6033 584 6067 618
rect 7357 665 7391 699
rect 6433 584 6467 618
rect 4763 384 4797 418
rect 4993 434 5027 468
rect 5953 464 5987 498
rect 6183 464 6217 498
rect 4763 304 4797 338
rect 5143 314 5177 348
rect 5753 344 5787 378
rect 6183 384 6217 418
rect 6183 304 6217 338
rect 6483 464 6517 498
rect 6483 384 6517 418
rect 6483 304 6517 338
rect 6783 464 6817 498
rect 6933 464 6967 498
rect 6783 384 6817 418
rect 6783 304 6817 338
rect 6933 344 6967 378
rect 1343 84 1377 118
rect 1423 84 1457 118
rect 1503 84 1537 118
rect 1583 84 1617 118
rect 1663 84 1697 118
rect 1743 84 1777 118
rect 1823 84 1857 118
rect 1903 84 1937 118
rect 1983 84 2017 118
rect 2063 84 2097 118
rect 2143 84 2177 118
rect 2223 84 2257 118
rect 2303 84 2337 118
rect 2383 84 2417 118
rect 2463 84 2497 118
rect 2543 84 2577 118
rect 2623 84 2657 118
rect 2703 84 2737 118
rect 2783 84 2817 118
rect 2863 84 2897 118
rect 2943 84 2977 118
rect 3663 84 3697 118
rect 3743 84 3777 118
rect 3823 84 3857 118
rect 3903 84 3937 118
rect 3983 84 4017 118
rect 4063 84 4097 118
rect 4143 84 4177 118
rect 4223 84 4257 118
rect 4303 84 4337 118
rect 4383 84 4417 118
rect 4463 84 4497 118
rect 4543 84 4577 118
rect 4623 84 4657 118
rect 4703 84 4737 118
rect 4783 84 4817 118
rect 4863 84 4897 118
rect 4943 84 4977 118
rect 5023 84 5057 118
rect 5103 84 5137 118
rect 5183 84 5217 118
rect 5263 84 5297 118
rect 5683 84 5717 118
rect 5763 84 5797 118
rect 5843 84 5877 118
rect 5923 84 5957 118
rect 6003 84 6037 118
rect 6083 84 6117 118
rect 6163 84 6197 118
rect 6243 84 6277 118
rect 6323 84 6357 118
rect 6403 84 6437 118
rect 6483 84 6517 118
rect 6563 84 6597 118
rect 6643 84 6677 118
rect 6723 84 6757 118
rect 6803 84 6837 118
rect 6883 84 6917 118
rect 6963 84 6997 118
rect 7043 84 7077 118
rect 7123 84 7157 118
rect 7203 84 7237 118
rect 7283 84 7317 118
rect 1103 -376 1137 -342
rect 1183 -376 1217 -342
rect 1263 -376 1297 -342
rect 1343 -376 1377 -342
rect 1423 -376 1457 -342
rect 1503 -376 1537 -342
rect 1583 -376 1617 -342
rect 1663 -376 1697 -342
rect 1743 -376 1777 -342
rect 1823 -376 1857 -342
rect 1903 -376 1937 -342
rect 1983 -376 2017 -342
rect 2063 -376 2097 -342
rect 2143 -376 2177 -342
rect 2223 -376 2257 -342
rect 2303 -376 2337 -342
rect 2383 -376 2417 -342
rect 2463 -376 2497 -342
rect 2543 -376 2577 -342
rect 2623 -376 2657 -342
rect 2703 -376 2737 -342
rect 2783 -376 2817 -342
rect 2863 -376 2897 -342
rect 2943 -376 2977 -342
rect 3023 -376 3057 -342
rect 3103 -376 3137 -342
rect 3183 -376 3217 -342
rect 3693 -376 3727 -342
rect 3773 -376 3807 -342
rect 3853 -376 3887 -342
rect 3933 -376 3967 -342
rect 4013 -376 4047 -342
rect 4093 -376 4127 -342
rect 4173 -376 4207 -342
rect 4253 -376 4287 -342
rect 4333 -376 4367 -342
rect 4413 -376 4447 -342
rect 4493 -376 4527 -342
rect 4573 -376 4607 -342
rect 4653 -376 4687 -342
rect 4733 -376 4767 -342
rect 4813 -376 4847 -342
rect 4893 -376 4927 -342
rect 4973 -376 5007 -342
rect 5413 -376 5447 -342
rect 5493 -376 5527 -342
rect 5573 -376 5607 -342
rect 5653 -376 5687 -342
rect 5733 -376 5767 -342
rect 5813 -376 5847 -342
rect 5893 -376 5927 -342
rect 5973 -376 6007 -342
rect 6053 -376 6087 -342
rect 6133 -376 6167 -342
rect 6213 -376 6247 -342
rect 6293 -376 6327 -342
rect 6373 -376 6407 -342
rect 6453 -376 6487 -342
rect 6533 -376 6567 -342
rect 6613 -376 6647 -342
rect 6693 -376 6727 -342
rect 6773 -376 6807 -342
rect 6853 -376 6887 -342
rect 6933 -376 6967 -342
rect 7013 -376 7047 -342
rect 479 -526 513 -492
rect 1563 -506 1597 -472
rect 2823 -506 2857 -472
rect 5274 -492 5308 -458
rect 5495 -494 5529 -460
rect 593 -606 627 -572
rect 1693 -606 1727 -572
rect 1843 -596 1877 -562
rect 23 -706 57 -672
rect 1563 -706 1597 -672
rect 1843 -676 1877 -642
rect 137 -827 171 -793
rect 1693 -806 1727 -772
rect 1843 -756 1877 -722
rect 2143 -596 2177 -562
rect 2143 -676 2177 -642
rect 2143 -756 2177 -722
rect 2443 -596 2477 -562
rect 3023 -606 3057 -572
rect 3595 -572 3629 -538
rect 2443 -676 2477 -642
rect 2443 -756 2477 -722
rect 3173 -706 3207 -672
rect 2193 -876 2227 -842
rect 2723 -806 2757 -772
rect 2563 -886 2597 -852
rect 4033 -596 4067 -562
rect 4033 -676 4067 -642
rect 3883 -756 3917 -722
rect 4033 -756 4067 -722
rect 4333 -596 4367 -562
rect 4333 -676 4367 -642
rect 4333 -756 4367 -722
rect 4633 -596 4667 -562
rect 5333 -606 5367 -572
rect 5763 -606 5797 -572
rect 5913 -596 5947 -562
rect 4633 -676 4667 -642
rect 4633 -756 4667 -722
rect 4783 -756 4817 -722
rect 4383 -876 4417 -842
rect 3323 -1000 3357 -966
rect 1363 -1156 1397 -1122
rect 1363 -1236 1397 -1202
rect 1363 -1316 1397 -1282
rect 1843 -1156 1877 -1122
rect 1843 -1236 1877 -1202
rect 1843 -1316 1877 -1282
rect 2143 -1156 2177 -1122
rect 2143 -1236 2177 -1202
rect 2143 -1316 2177 -1282
rect 2443 -1156 2477 -1122
rect 2443 -1236 2477 -1202
rect 2443 -1316 2477 -1282
rect 2923 -1156 2957 -1122
rect 2923 -1236 2957 -1202
rect 2923 -1316 2957 -1282
rect 4783 -876 4817 -842
rect 5071 -882 5105 -848
rect 5763 -726 5797 -692
rect 5913 -676 5947 -642
rect 5913 -756 5947 -722
rect 6213 -596 6247 -562
rect 6213 -676 6247 -642
rect 6213 -756 6247 -722
rect 6513 -596 6547 -562
rect 6893 -606 6927 -572
rect 6513 -676 6547 -642
rect 6513 -756 6547 -722
rect 6743 -726 6777 -692
rect 5333 -826 5367 -792
rect 5333 -946 5367 -912
rect 6263 -876 6297 -842
rect 6663 -876 6697 -842
rect 7096 -996 7130 -962
rect 3337 -1204 3371 -1170
rect 3703 -1156 3737 -1122
rect 3703 -1236 3737 -1202
rect 3703 -1316 3737 -1282
rect 4033 -1156 4067 -1122
rect 4033 -1236 4067 -1202
rect 4033 -1316 4067 -1282
rect 4333 -1156 4367 -1122
rect 4333 -1236 4367 -1202
rect 4333 -1316 4367 -1282
rect 4633 -1156 4667 -1122
rect 4633 -1236 4667 -1202
rect 4633 -1316 4667 -1282
rect 4963 -1156 4997 -1122
rect 4963 -1236 4997 -1202
rect 4963 -1316 4997 -1282
rect 5583 -1156 5617 -1122
rect 5583 -1236 5617 -1202
rect 5583 -1316 5617 -1282
rect 5913 -1156 5947 -1122
rect 5913 -1236 5947 -1202
rect 5913 -1316 5947 -1282
rect 6213 -1156 6247 -1122
rect 6213 -1236 6247 -1202
rect 6213 -1316 6247 -1282
rect 6513 -1156 6547 -1122
rect 6513 -1236 6547 -1202
rect 6513 -1316 6547 -1282
rect 6993 -1156 7027 -1122
rect 6993 -1236 7027 -1202
rect 6993 -1316 7027 -1282
rect 1194 -1436 1228 -1402
rect 5421 -1436 5455 -1402
rect 935 -1556 969 -1522
rect 1103 -1556 1137 -1522
rect 1183 -1556 1217 -1522
rect 1263 -1556 1297 -1522
rect 1343 -1556 1377 -1522
rect 1423 -1556 1457 -1522
rect 1503 -1556 1537 -1522
rect 1583 -1556 1617 -1522
rect 1663 -1556 1697 -1522
rect 1743 -1556 1777 -1522
rect 1823 -1556 1857 -1522
rect 1903 -1556 1937 -1522
rect 1983 -1556 2017 -1522
rect 2063 -1556 2097 -1522
rect 2143 -1556 2177 -1522
rect 2223 -1556 2257 -1522
rect 2303 -1556 2337 -1522
rect 2383 -1556 2417 -1522
rect 2463 -1556 2497 -1522
rect 2543 -1556 2577 -1522
rect 2623 -1556 2657 -1522
rect 2703 -1556 2737 -1522
rect 2783 -1556 2817 -1522
rect 2863 -1556 2897 -1522
rect 2943 -1556 2977 -1522
rect 3023 -1556 3057 -1522
rect 3103 -1556 3137 -1522
rect 3183 -1556 3217 -1522
rect 3693 -1556 3727 -1522
rect 3773 -1556 3807 -1522
rect 3853 -1556 3887 -1522
rect 3933 -1556 3967 -1522
rect 4013 -1556 4047 -1522
rect 4093 -1556 4127 -1522
rect 4173 -1556 4207 -1522
rect 4253 -1556 4287 -1522
rect 4333 -1556 4367 -1522
rect 4413 -1556 4447 -1522
rect 4493 -1556 4527 -1522
rect 4573 -1556 4607 -1522
rect 4653 -1556 4687 -1522
rect 4733 -1556 4767 -1522
rect 4813 -1556 4847 -1522
rect 4893 -1556 4927 -1522
rect 4973 -1556 5007 -1522
rect 5413 -1556 5447 -1522
rect 5493 -1556 5527 -1522
rect 5573 -1556 5607 -1522
rect 5653 -1556 5687 -1522
rect 5733 -1556 5767 -1522
rect 5813 -1556 5847 -1522
rect 5893 -1556 5927 -1522
rect 5973 -1556 6007 -1522
rect 6053 -1556 6087 -1522
rect 6133 -1556 6167 -1522
rect 6213 -1556 6247 -1522
rect 6293 -1556 6327 -1522
rect 6373 -1556 6407 -1522
rect 6453 -1556 6487 -1522
rect 6533 -1556 6567 -1522
rect 6613 -1556 6647 -1522
rect 6693 -1556 6727 -1522
rect 6773 -1556 6807 -1522
rect 6853 -1556 6887 -1522
rect 6933 -1556 6967 -1522
rect 7013 -1556 7047 -1522
rect 1194 -1676 1228 -1642
rect 5421 -1675 5455 -1641
rect 1363 -1796 1397 -1762
rect 1363 -1876 1397 -1842
rect 1363 -1956 1397 -1922
rect 1843 -1796 1877 -1762
rect 1843 -1876 1877 -1842
rect 1843 -1956 1877 -1922
rect 2143 -1796 2177 -1762
rect 2143 -1876 2177 -1842
rect 2143 -1956 2177 -1922
rect 2443 -1796 2477 -1762
rect 2443 -1876 2477 -1842
rect 2443 -1956 2477 -1922
rect 2923 -1796 2957 -1762
rect 2923 -1876 2957 -1842
rect 2923 -1956 2957 -1922
rect 3703 -1796 3737 -1762
rect 3337 -1899 3371 -1865
rect 3703 -1876 3737 -1842
rect 3703 -1956 3737 -1922
rect 4033 -1796 4067 -1762
rect 4033 -1876 4067 -1842
rect 4033 -1956 4067 -1922
rect 4333 -1796 4367 -1762
rect 4333 -1876 4367 -1842
rect 4333 -1956 4367 -1922
rect 4633 -1796 4667 -1762
rect 4633 -1876 4667 -1842
rect 4633 -1956 4667 -1922
rect 4963 -1796 4997 -1762
rect 4963 -1876 4997 -1842
rect 4963 -1956 4997 -1922
rect 5583 -1796 5617 -1762
rect 5583 -1876 5617 -1842
rect 5583 -1956 5617 -1922
rect 5913 -1796 5947 -1762
rect 5913 -1876 5947 -1842
rect 5913 -1956 5947 -1922
rect 6213 -1796 6247 -1762
rect 6213 -1876 6247 -1842
rect 6213 -1956 6247 -1922
rect 6513 -1796 6547 -1762
rect 6513 -1876 6547 -1842
rect 6513 -1956 6547 -1922
rect 6993 -1796 7027 -1762
rect 6993 -1876 7027 -1842
rect 6993 -1956 7027 -1922
rect 2193 -2236 2227 -2202
rect 821 -2286 855 -2252
rect 1693 -2306 1727 -2272
rect 2563 -2226 2597 -2192
rect 3323 -2226 3357 -2192
rect 707 -2386 741 -2352
rect 1563 -2406 1597 -2372
rect 1843 -2356 1877 -2322
rect 1843 -2436 1877 -2402
rect 365 -2506 399 -2472
rect 1693 -2506 1727 -2472
rect 1843 -2516 1877 -2482
rect 2143 -2356 2177 -2322
rect 2143 -2436 2177 -2402
rect 2143 -2516 2177 -2482
rect 2443 -2356 2477 -2322
rect 2723 -2306 2757 -2272
rect 2443 -2436 2477 -2402
rect 3173 -2406 3207 -2372
rect 2443 -2516 2477 -2482
rect 3023 -2506 3057 -2472
rect 4383 -2236 4417 -2202
rect 4783 -2236 4817 -2202
rect 7096 -2116 7130 -2082
rect 3883 -2356 3917 -2322
rect 4033 -2356 4067 -2322
rect 4033 -2436 4067 -2402
rect 3595 -2540 3629 -2506
rect 251 -2626 285 -2592
rect 1563 -2606 1597 -2572
rect 4033 -2516 4067 -2482
rect 4333 -2356 4367 -2322
rect 4333 -2436 4367 -2402
rect 4333 -2516 4367 -2482
rect 4633 -2356 4667 -2322
rect 4783 -2356 4817 -2322
rect 5333 -2286 5367 -2252
rect 6263 -2236 6297 -2202
rect 6663 -2236 6697 -2202
rect 5763 -2386 5797 -2352
rect 4633 -2436 4667 -2402
rect 5913 -2356 5947 -2322
rect 5913 -2436 5947 -2402
rect 4633 -2516 4667 -2482
rect 5333 -2507 5367 -2473
rect 5763 -2506 5797 -2472
rect 5913 -2516 5947 -2482
rect 6213 -2356 6247 -2322
rect 6213 -2436 6247 -2402
rect 6213 -2516 6247 -2482
rect 6513 -2356 6547 -2322
rect 6513 -2436 6547 -2402
rect 6743 -2386 6777 -2352
rect 6513 -2516 6547 -2482
rect 6893 -2506 6927 -2472
rect 2823 -2606 2857 -2572
rect 1103 -2736 1137 -2702
rect 1183 -2736 1217 -2702
rect 1263 -2736 1297 -2702
rect 1343 -2736 1377 -2702
rect 1423 -2736 1457 -2702
rect 1503 -2736 1537 -2702
rect 1583 -2736 1617 -2702
rect 1663 -2736 1697 -2702
rect 1743 -2736 1777 -2702
rect 1823 -2736 1857 -2702
rect 1903 -2736 1937 -2702
rect 1983 -2736 2017 -2702
rect 2063 -2736 2097 -2702
rect 2143 -2736 2177 -2702
rect 2223 -2736 2257 -2702
rect 2303 -2736 2337 -2702
rect 2383 -2736 2417 -2702
rect 2463 -2736 2497 -2702
rect 2543 -2736 2577 -2702
rect 2623 -2736 2657 -2702
rect 2703 -2736 2737 -2702
rect 2783 -2736 2817 -2702
rect 2863 -2736 2897 -2702
rect 2943 -2736 2977 -2702
rect 3023 -2736 3057 -2702
rect 3103 -2736 3137 -2702
rect 3183 -2736 3217 -2702
rect 3693 -2736 3727 -2702
rect 3773 -2736 3807 -2702
rect 3853 -2736 3887 -2702
rect 3933 -2736 3967 -2702
rect 4013 -2736 4047 -2702
rect 4093 -2736 4127 -2702
rect 4173 -2736 4207 -2702
rect 4253 -2736 4287 -2702
rect 4333 -2736 4367 -2702
rect 4413 -2736 4447 -2702
rect 4493 -2736 4527 -2702
rect 4573 -2736 4607 -2702
rect 4653 -2736 4687 -2702
rect 4733 -2736 4767 -2702
rect 4813 -2736 4847 -2702
rect 4893 -2736 4927 -2702
rect 4973 -2736 5007 -2702
rect 5413 -2736 5447 -2702
rect 5493 -2736 5527 -2702
rect 5573 -2736 5607 -2702
rect 5653 -2736 5687 -2702
rect 5733 -2736 5767 -2702
rect 5813 -2736 5847 -2702
rect 5893 -2736 5927 -2702
rect 5973 -2736 6007 -2702
rect 6053 -2736 6087 -2702
rect 6133 -2736 6167 -2702
rect 6213 -2736 6247 -2702
rect 6293 -2736 6327 -2702
rect 6373 -2736 6407 -2702
rect 6453 -2736 6487 -2702
rect 6533 -2736 6567 -2702
rect 6613 -2736 6647 -2702
rect 6693 -2736 6727 -2702
rect 6773 -2736 6807 -2702
rect 6853 -2736 6887 -2702
rect 6933 -2736 6967 -2702
rect 7013 -2736 7047 -2702
rect 5421 -2970 5455 -2936
rect 1184 -3196 1218 -3162
rect 1264 -3196 1298 -3162
rect 1344 -3196 1378 -3162
rect 1424 -3196 1458 -3162
rect 1504 -3196 1538 -3162
rect 1584 -3196 1618 -3162
rect 1664 -3196 1698 -3162
rect 1744 -3196 1778 -3162
rect 1824 -3196 1858 -3162
rect 1904 -3196 1938 -3162
rect 1984 -3196 2018 -3162
rect 2064 -3196 2098 -3162
rect 2144 -3196 2178 -3162
rect 2224 -3196 2258 -3162
rect 2304 -3196 2338 -3162
rect 2384 -3196 2418 -3162
rect 2464 -3196 2498 -3162
rect 2544 -3196 2578 -3162
rect 2624 -3196 2658 -3162
rect 2704 -3196 2738 -3162
rect 2784 -3196 2818 -3162
rect 2864 -3196 2898 -3162
rect 2944 -3196 2978 -3162
rect 3024 -3196 3058 -3162
rect 3104 -3196 3138 -3162
rect 3554 -3196 3588 -3162
rect 3634 -3196 3668 -3162
rect 3714 -3196 3748 -3162
rect 3794 -3196 3828 -3162
rect 3874 -3196 3908 -3162
rect 3954 -3196 3988 -3162
rect 4034 -3196 4068 -3162
rect 4114 -3196 4148 -3162
rect 4194 -3196 4228 -3162
rect 4274 -3196 4308 -3162
rect 4354 -3196 4388 -3162
rect 4434 -3196 4468 -3162
rect 4514 -3196 4548 -3162
rect 4594 -3196 4628 -3162
rect 4674 -3196 4708 -3162
rect 4754 -3196 4788 -3162
rect 4834 -3196 4868 -3162
rect 821 -3296 855 -3262
rect 1604 -3316 1638 -3282
rect 2974 -3316 3008 -3282
rect 7366 -3003 7400 -2969
rect 5274 -3197 5308 -3163
rect 5354 -3197 5388 -3163
rect 5434 -3197 5468 -3163
rect 5514 -3197 5548 -3163
rect 5594 -3197 5628 -3163
rect 5674 -3197 5708 -3163
rect 5754 -3197 5788 -3163
rect 5834 -3197 5868 -3163
rect 5914 -3197 5948 -3163
rect 5994 -3197 6028 -3163
rect 6074 -3197 6108 -3163
rect 6154 -3197 6188 -3163
rect 6234 -3197 6268 -3163
rect 6314 -3197 6348 -3163
rect 6394 -3197 6428 -3163
rect 6474 -3197 6508 -3163
rect 6554 -3197 6588 -3163
rect 6634 -3197 6668 -3163
rect 6714 -3197 6748 -3163
rect 6794 -3197 6828 -3163
rect 6874 -3197 6908 -3163
rect 6954 -3197 6988 -3163
rect 7034 -3197 7068 -3163
rect 7114 -3197 7148 -3163
rect 7194 -3197 7228 -3163
rect 5404 -3322 5438 -3288
rect 6684 -3327 6718 -3293
rect 7252 -3327 7286 -3293
rect 251 -3416 285 -3382
rect 1694 -3436 1728 -3402
rect 1844 -3416 1878 -3382
rect 137 -3519 171 -3485
rect 1844 -3496 1878 -3462
rect 707 -3612 741 -3578
rect 1664 -3556 1698 -3522
rect 1844 -3576 1878 -3542
rect 2144 -3416 2178 -3382
rect 2144 -3496 2178 -3462
rect 2144 -3576 2178 -3542
rect 2444 -3416 2478 -3382
rect 2824 -3436 2858 -3402
rect 3894 -3416 3928 -3382
rect 2444 -3496 2478 -3462
rect 3894 -3496 3928 -3462
rect 2444 -3576 2478 -3542
rect 2694 -3556 2728 -3522
rect 3456 -3576 3490 -3542
rect 3744 -3576 3778 -3542
rect 3894 -3576 3928 -3542
rect 4194 -3416 4228 -3382
rect 4194 -3496 4228 -3462
rect 4194 -3576 4228 -3542
rect 4494 -3416 4528 -3382
rect 5027 -3403 5061 -3369
rect 4494 -3496 4528 -3462
rect 5504 -3447 5538 -3413
rect 5934 -3417 5968 -3383
rect 4494 -3576 4528 -3542
rect 5704 -3537 5738 -3503
rect 4644 -3576 4678 -3542
rect 5934 -3497 5968 -3463
rect 5203 -3599 5237 -3565
rect 5934 -3577 5968 -3543
rect 365 -3686 399 -3652
rect 2194 -3696 2228 -3662
rect 23 -3786 57 -3752
rect 2594 -3696 2628 -3662
rect 3174 -3815 3208 -3781
rect 4244 -3696 4278 -3662
rect 6234 -3417 6268 -3383
rect 6234 -3497 6268 -3463
rect 6234 -3577 6268 -3543
rect 6534 -3417 6568 -3383
rect 6804 -3437 6838 -3403
rect 7056 -3437 7090 -3403
rect 6534 -3497 6568 -3463
rect 6534 -3577 6568 -3543
rect 6684 -3537 6718 -3503
rect 4644 -3696 4678 -3662
rect 5204 -3713 5238 -3679
rect 5784 -3697 5818 -3663
rect 6184 -3697 6218 -3663
rect 7298 -3625 7332 -3591
rect 4938 -3866 4972 -3832
rect 5204 -3827 5238 -3793
rect 1214 -3976 1248 -3942
rect 1214 -4056 1248 -4022
rect 1214 -4136 1248 -4102
rect 1514 -3976 1548 -3942
rect 1514 -4056 1548 -4022
rect 1514 -4136 1548 -4102
rect 1844 -3976 1878 -3942
rect 1844 -4056 1878 -4022
rect 1844 -4136 1878 -4102
rect 2144 -3976 2178 -3942
rect 2144 -4056 2178 -4022
rect 2144 -4136 2178 -4102
rect 2444 -3976 2478 -3942
rect 2444 -4056 2478 -4022
rect 2444 -4136 2478 -4102
rect 3074 -3976 3108 -3942
rect 3074 -4056 3108 -4022
rect 3074 -4136 3108 -4102
rect 3564 -3976 3598 -3942
rect 3564 -4056 3598 -4022
rect 3564 -4136 3598 -4102
rect 3894 -3976 3928 -3942
rect 3894 -4056 3928 -4022
rect 3894 -4136 3928 -4102
rect 4194 -3976 4228 -3942
rect 4194 -4056 4228 -4022
rect 4194 -4136 4228 -4102
rect 4494 -3976 4528 -3942
rect 4494 -4056 4528 -4022
rect 4494 -4136 4528 -4102
rect 6814 -3827 6848 -3793
rect 4824 -3976 4858 -3942
rect 5021 -3980 5055 -3946
rect 5304 -3977 5338 -3943
rect 4824 -4056 4858 -4022
rect 4824 -4136 4858 -4102
rect 5304 -4057 5338 -4023
rect 5304 -4137 5338 -4103
rect 5604 -3977 5638 -3943
rect 5604 -4057 5638 -4023
rect 5604 -4137 5638 -4103
rect 5934 -3977 5968 -3943
rect 5934 -4057 5968 -4023
rect 5934 -4137 5968 -4103
rect 6234 -3977 6268 -3943
rect 6234 -4057 6268 -4023
rect 6234 -4137 6268 -4103
rect 6534 -3977 6568 -3943
rect 6534 -4057 6568 -4023
rect 6534 -4137 6568 -4103
rect 7164 -3977 7198 -3943
rect 7164 -4057 7198 -4023
rect 7164 -4137 7198 -4103
rect 1194 -4256 1228 -4222
rect 5115 -4258 5149 -4224
rect 935 -4376 969 -4342
rect 1184 -4376 1218 -4342
rect 1264 -4376 1298 -4342
rect 1344 -4376 1378 -4342
rect 1424 -4376 1458 -4342
rect 1504 -4376 1538 -4342
rect 1584 -4376 1618 -4342
rect 1664 -4376 1698 -4342
rect 1744 -4376 1778 -4342
rect 1824 -4376 1858 -4342
rect 1904 -4376 1938 -4342
rect 1984 -4376 2018 -4342
rect 2064 -4376 2098 -4342
rect 2144 -4376 2178 -4342
rect 2224 -4376 2258 -4342
rect 2304 -4376 2338 -4342
rect 2384 -4376 2418 -4342
rect 2464 -4376 2498 -4342
rect 2544 -4376 2578 -4342
rect 2624 -4376 2658 -4342
rect 2704 -4376 2738 -4342
rect 2784 -4376 2818 -4342
rect 2864 -4376 2898 -4342
rect 2944 -4376 2978 -4342
rect 3024 -4376 3058 -4342
rect 3104 -4376 3138 -4342
rect 3184 -4376 3218 -4342
rect 3264 -4376 3298 -4342
rect 936 -4456 970 -4422
rect 1063 -4456 1097 -4422
rect 1143 -4456 1177 -4422
rect 1223 -4456 1257 -4422
rect 1303 -4456 1337 -4422
rect 1383 -4456 1417 -4422
rect 1463 -4456 1497 -4422
rect 1543 -4456 1577 -4422
rect 1623 -4456 1657 -4422
rect 1703 -4456 1737 -4422
rect 1783 -4456 1817 -4422
rect 1863 -4456 1897 -4422
rect 1943 -4456 1977 -4422
rect 2023 -4456 2057 -4422
rect 2103 -4456 2137 -4422
rect 2183 -4456 2217 -4422
rect 2263 -4456 2297 -4422
rect 2343 -4456 2377 -4422
rect 2423 -4456 2457 -4422
rect 2503 -4456 2537 -4422
rect 2583 -4456 2617 -4422
rect 2663 -4456 2697 -4422
rect 2743 -4456 2777 -4422
rect 2823 -4456 2857 -4422
rect 2903 -4456 2937 -4422
rect 2983 -4456 3017 -4422
rect 3063 -4456 3097 -4422
rect 3143 -4456 3177 -4422
rect 3223 -4456 3257 -4422
rect 3303 -4456 3337 -4422
rect 3554 -4376 3588 -4342
rect 3634 -4376 3668 -4342
rect 3714 -4376 3748 -4342
rect 3794 -4376 3828 -4342
rect 3874 -4376 3908 -4342
rect 3954 -4376 3988 -4342
rect 4034 -4376 4068 -4342
rect 4114 -4376 4148 -4342
rect 4194 -4376 4228 -4342
rect 4274 -4376 4308 -4342
rect 4354 -4376 4388 -4342
rect 4434 -4376 4468 -4342
rect 4514 -4376 4548 -4342
rect 4594 -4376 4628 -4342
rect 4674 -4376 4708 -4342
rect 4754 -4376 4788 -4342
rect 4834 -4376 4868 -4342
rect 4914 -4376 4948 -4342
rect 4994 -4376 5028 -4342
rect 3594 -4457 3628 -4423
rect 3674 -4457 3708 -4423
rect 3754 -4457 3788 -4423
rect 3834 -4457 3868 -4423
rect 3914 -4457 3948 -4423
rect 3994 -4457 4028 -4423
rect 4074 -4457 4108 -4423
rect 4154 -4457 4188 -4423
rect 4234 -4457 4268 -4423
rect 4314 -4457 4348 -4423
rect 4394 -4457 4428 -4423
rect 4474 -4457 4508 -4423
rect 4554 -4457 4588 -4423
rect 4634 -4457 4668 -4423
rect 4714 -4457 4748 -4423
rect 4794 -4457 4828 -4423
rect 4874 -4457 4908 -4423
rect 4954 -4457 4988 -4423
rect 5034 -4457 5068 -4423
rect 5274 -4377 5308 -4343
rect 5354 -4377 5388 -4343
rect 5434 -4377 5468 -4343
rect 5514 -4377 5548 -4343
rect 5594 -4377 5628 -4343
rect 5674 -4377 5708 -4343
rect 5754 -4377 5788 -4343
rect 5834 -4377 5868 -4343
rect 5914 -4377 5948 -4343
rect 5994 -4377 6028 -4343
rect 6074 -4377 6108 -4343
rect 6154 -4377 6188 -4343
rect 6234 -4377 6268 -4343
rect 6314 -4377 6348 -4343
rect 6394 -4377 6428 -4343
rect 6474 -4377 6508 -4343
rect 6554 -4377 6588 -4343
rect 6634 -4377 6668 -4343
rect 6714 -4377 6748 -4343
rect 6794 -4377 6828 -4343
rect 6874 -4377 6908 -4343
rect 6954 -4377 6988 -4343
rect 7034 -4377 7068 -4343
rect 7114 -4377 7148 -4343
rect 7194 -4377 7228 -4343
rect 7274 -4376 7308 -4342
rect 7354 -4376 7388 -4342
rect 5333 -4457 5367 -4423
rect 5413 -4457 5447 -4423
rect 5493 -4457 5527 -4423
rect 5573 -4457 5607 -4423
rect 5653 -4457 5687 -4423
rect 5733 -4457 5767 -4423
rect 5813 -4457 5847 -4423
rect 5893 -4457 5927 -4423
rect 5973 -4457 6007 -4423
rect 6053 -4457 6087 -4423
rect 6133 -4457 6167 -4423
rect 6213 -4457 6247 -4423
rect 6293 -4457 6327 -4423
rect 6373 -4457 6407 -4423
rect 6453 -4457 6487 -4423
rect 6533 -4457 6567 -4423
rect 6613 -4457 6647 -4423
rect 6693 -4457 6727 -4423
rect 6773 -4457 6807 -4423
rect 6853 -4457 6887 -4423
rect 6933 -4457 6967 -4423
rect 7013 -4457 7047 -4423
rect 7093 -4457 7127 -4423
rect 7173 -4457 7207 -4423
rect 7253 -4457 7287 -4423
rect 7333 -4457 7367 -4423
rect 7413 -4457 7447 -4423
rect 1064 -4579 1098 -4545
rect 5138 -4577 5172 -4543
rect 5335 -4577 5369 -4543
rect 1253 -4696 1287 -4662
rect 1253 -4776 1287 -4742
rect 1253 -4856 1287 -4822
rect 1553 -4696 1587 -4662
rect 1553 -4776 1587 -4742
rect 1553 -4856 1587 -4822
rect 1883 -4696 1917 -4662
rect 1883 -4776 1917 -4742
rect 1883 -4856 1917 -4822
rect 2183 -4696 2217 -4662
rect 2183 -4776 2217 -4742
rect 2183 -4856 2217 -4822
rect 2483 -4696 2517 -4662
rect 2483 -4776 2517 -4742
rect 2483 -4856 2517 -4822
rect 3263 -4696 3297 -4662
rect 3263 -4776 3297 -4742
rect 3263 -4856 3297 -4822
rect 3764 -4697 3798 -4663
rect 3764 -4777 3798 -4743
rect 3764 -4857 3798 -4823
rect 593 -5046 627 -5012
rect 137 -5186 171 -5152
rect 365 -5286 399 -5252
rect 707 -5366 741 -5332
rect 4094 -4697 4128 -4663
rect 4094 -4777 4128 -4743
rect 4094 -4857 4128 -4823
rect 4394 -4697 4428 -4663
rect 4394 -4777 4428 -4743
rect 4394 -4857 4428 -4823
rect 4694 -4697 4728 -4663
rect 4694 -4777 4728 -4743
rect 4694 -4857 4728 -4823
rect 5024 -4697 5058 -4663
rect 5024 -4777 5058 -4743
rect 5024 -4857 5058 -4823
rect 5523 -4697 5557 -4663
rect 5523 -4777 5557 -4743
rect 5523 -4857 5557 -4823
rect 5823 -4697 5857 -4663
rect 5823 -4777 5857 -4743
rect 5823 -4857 5857 -4823
rect 6153 -4697 6187 -4663
rect 6153 -4777 6187 -4743
rect 6153 -4857 6187 -4823
rect 6453 -4697 6487 -4663
rect 6453 -4777 6487 -4743
rect 6453 -4857 6487 -4823
rect 6753 -4697 6787 -4663
rect 6753 -4777 6787 -4743
rect 6753 -4857 6787 -4823
rect 7383 -4697 7417 -4663
rect 7383 -4777 7417 -4743
rect 7383 -4857 7417 -4823
rect 2713 -5066 2747 -5032
rect 2863 -5066 2897 -5032
rect 3013 -5066 3047 -5032
rect 3163 -5066 3197 -5032
rect 3656 -5017 3690 -4983
rect 5138 -4967 5172 -4933
rect 5423 -4997 5457 -4963
rect 4444 -5137 4478 -5103
rect 4844 -5137 4878 -5103
rect 5423 -5117 5457 -5083
rect 6003 -5137 6037 -5103
rect 2233 -5366 2267 -5332
rect 479 -5446 513 -5412
rect 1153 -5466 1187 -5432
rect 3944 -5257 3978 -5223
rect 4094 -5257 4128 -5223
rect 2433 -5366 2467 -5332
rect 3363 -5367 3397 -5333
rect 4094 -5337 4128 -5303
rect 4094 -5417 4128 -5383
rect 4394 -5257 4428 -5223
rect 4394 -5337 4428 -5303
rect 4394 -5417 4428 -5383
rect 7033 -5007 7067 -4973
rect 6403 -5137 6437 -5103
rect 4694 -5257 4728 -5223
rect 4844 -5257 4878 -5223
rect 5423 -5245 5457 -5211
rect 4694 -5337 4728 -5303
rect 5923 -5297 5957 -5263
rect 6153 -5257 6187 -5223
rect 4694 -5417 4728 -5383
rect 5138 -5430 5172 -5396
rect 5723 -5387 5757 -5353
rect 6153 -5337 6187 -5303
rect 6153 -5417 6187 -5383
rect 6453 -5257 6487 -5223
rect 6453 -5337 6487 -5303
rect 6453 -5417 6487 -5383
rect 7517 -5210 7551 -5176
rect 6753 -5257 6787 -5223
rect 6753 -5337 6787 -5303
rect 6903 -5297 6937 -5263
rect 6753 -5417 6787 -5383
rect 7023 -5397 7057 -5363
rect 7155 -5396 7189 -5362
rect 23 -5566 57 -5532
rect 1153 -5586 1187 -5552
rect 1883 -5576 1917 -5542
rect 251 -5686 285 -5652
rect 1153 -5706 1187 -5672
rect 1883 -5656 1917 -5622
rect 1883 -5736 1917 -5702
rect 2183 -5576 2217 -5542
rect 2183 -5656 2217 -5622
rect 2183 -5736 2217 -5702
rect 2483 -5576 2517 -5542
rect 2483 -5656 2517 -5622
rect 3754 -5637 3788 -5603
rect 3834 -5637 3868 -5603
rect 3914 -5637 3948 -5603
rect 3994 -5637 4028 -5603
rect 4074 -5637 4108 -5603
rect 4154 -5637 4188 -5603
rect 4234 -5637 4268 -5603
rect 4314 -5637 4348 -5603
rect 4394 -5637 4428 -5603
rect 4474 -5637 4508 -5603
rect 4554 -5637 4588 -5603
rect 4634 -5637 4668 -5603
rect 4714 -5637 4748 -5603
rect 4794 -5637 4828 -5603
rect 4874 -5637 4908 -5603
rect 4954 -5637 4988 -5603
rect 5034 -5637 5068 -5603
rect 2483 -5736 2517 -5702
rect 821 -5846 855 -5812
rect 1153 -5826 1187 -5792
rect 5623 -5512 5657 -5478
rect 6903 -5507 6937 -5473
rect 7293 -5507 7327 -5473
rect 5493 -5637 5527 -5603
rect 5573 -5637 5607 -5603
rect 5653 -5637 5687 -5603
rect 5733 -5637 5767 -5603
rect 5813 -5637 5847 -5603
rect 5893 -5637 5927 -5603
rect 5973 -5637 6007 -5603
rect 6053 -5637 6087 -5603
rect 6133 -5637 6167 -5603
rect 6213 -5637 6247 -5603
rect 6293 -5637 6327 -5603
rect 6373 -5637 6407 -5603
rect 6453 -5637 6487 -5603
rect 6533 -5637 6567 -5603
rect 6613 -5637 6647 -5603
rect 6693 -5637 6727 -5603
rect 6773 -5637 6807 -5603
rect 6853 -5637 6887 -5603
rect 6933 -5637 6967 -5603
rect 7013 -5637 7047 -5603
rect 7093 -5637 7127 -5603
rect 7173 -5637 7207 -5603
rect 7253 -5637 7287 -5603
rect 7333 -5637 7367 -5603
rect 7413 -5637 7447 -5603
rect 5481 -5863 5515 -5829
rect 1063 -5956 1097 -5922
rect 1143 -5956 1177 -5922
rect 1223 -5956 1257 -5922
rect 1303 -5956 1337 -5922
rect 1383 -5956 1417 -5922
rect 1463 -5956 1497 -5922
rect 1543 -5956 1577 -5922
rect 1623 -5956 1657 -5922
rect 1703 -5956 1737 -5922
rect 1783 -5956 1817 -5922
rect 1863 -5956 1897 -5922
rect 1943 -5956 1977 -5922
rect 2023 -5956 2057 -5922
rect 2103 -5956 2137 -5922
rect 2183 -5956 2217 -5922
rect 2263 -5956 2297 -5922
rect 2343 -5956 2377 -5922
rect 2423 -5956 2457 -5922
rect 2503 -5956 2537 -5922
rect 2583 -5956 2617 -5922
rect 2663 -5956 2697 -5922
rect 2743 -5956 2777 -5922
rect 2823 -5956 2857 -5922
rect 2903 -5956 2937 -5922
rect 2983 -5956 3017 -5922
rect 3063 -5956 3097 -5922
rect 3143 -5956 3177 -5922
rect 3223 -5956 3257 -5922
rect 3303 -5956 3337 -5922
rect 1063 -6097 1097 -6063
rect 1143 -6097 1177 -6063
rect 1223 -6097 1257 -6063
rect 1303 -6097 1337 -6063
rect 1383 -6097 1417 -6063
rect 1463 -6097 1497 -6063
rect 1543 -6097 1577 -6063
rect 1623 -6097 1657 -6063
rect 1703 -6097 1737 -6063
rect 1783 -6097 1817 -6063
rect 1863 -6097 1897 -6063
rect 1943 -6097 1977 -6063
rect 2023 -6097 2057 -6063
rect 2103 -6097 2137 -6063
rect 2183 -6097 2217 -6063
rect 2263 -6097 2297 -6063
rect 2343 -6097 2377 -6063
rect 2423 -6097 2457 -6063
rect 2503 -6097 2537 -6063
rect 2583 -6097 2617 -6063
rect 2663 -6097 2697 -6063
rect 2743 -6097 2777 -6063
rect 2823 -6097 2857 -6063
rect 2903 -6097 2937 -6063
rect 2983 -6097 3017 -6063
rect 3063 -6097 3097 -6063
rect 3143 -6097 3177 -6063
rect 3223 -6097 3257 -6063
rect 3303 -6097 3337 -6063
rect 3753 -6097 3787 -6063
rect 3833 -6097 3867 -6063
rect 3913 -6097 3947 -6063
rect 3993 -6097 4027 -6063
rect 4073 -6097 4107 -6063
rect 4153 -6097 4187 -6063
rect 4233 -6097 4267 -6063
rect 4313 -6097 4347 -6063
rect 4393 -6097 4427 -6063
rect 4473 -6097 4507 -6063
rect 4553 -6097 4587 -6063
rect 4633 -6097 4667 -6063
rect 4713 -6097 4747 -6063
rect 4793 -6097 4827 -6063
rect 4873 -6097 4907 -6063
rect 4953 -6097 4987 -6063
rect 5033 -6097 5067 -6063
rect 5472 -6097 5506 -6063
rect 5552 -6097 5586 -6063
rect 5632 -6097 5666 -6063
rect 5712 -6097 5746 -6063
rect 5792 -6097 5826 -6063
rect 5872 -6097 5906 -6063
rect 5952 -6097 5986 -6063
rect 6032 -6097 6066 -6063
rect 6112 -6097 6146 -6063
rect 6192 -6097 6226 -6063
rect 6272 -6097 6306 -6063
rect 6352 -6097 6386 -6063
rect 6432 -6097 6466 -6063
rect 6512 -6097 6546 -6063
rect 6592 -6097 6626 -6063
rect 6672 -6097 6706 -6063
rect 6752 -6097 6786 -6063
rect 6832 -6097 6866 -6063
rect 6912 -6097 6946 -6063
rect 6992 -6097 7026 -6063
rect 7072 -6097 7106 -6063
rect 251 -6207 285 -6173
rect 1603 -6227 1637 -6193
rect 2863 -6227 2897 -6193
rect 365 -6321 399 -6287
rect 1733 -6327 1767 -6293
rect 1883 -6317 1917 -6283
rect 23 -6428 57 -6394
rect 1603 -6427 1637 -6393
rect 1883 -6397 1917 -6363
rect 137 -6547 171 -6513
rect 1733 -6527 1767 -6493
rect 1883 -6477 1917 -6443
rect 2183 -6317 2217 -6283
rect 2183 -6397 2217 -6363
rect 2183 -6477 2217 -6443
rect 2483 -6317 2517 -6283
rect 3063 -6327 3097 -6293
rect 3655 -6327 3689 -6293
rect 2483 -6397 2517 -6363
rect 2483 -6477 2517 -6443
rect 3213 -6427 3247 -6393
rect 2233 -6597 2267 -6563
rect 2763 -6527 2797 -6493
rect 2603 -6607 2637 -6573
rect 3363 -6607 3397 -6573
rect 4093 -6317 4127 -6283
rect 4093 -6397 4127 -6363
rect 3943 -6477 3977 -6443
rect 4093 -6477 4127 -6443
rect 4393 -6317 4427 -6283
rect 4393 -6397 4427 -6363
rect 4393 -6477 4427 -6443
rect 4693 -6317 4727 -6283
rect 4843 -6327 4877 -6293
rect 5822 -6327 5856 -6293
rect 5972 -6317 6006 -6283
rect 4693 -6397 4727 -6363
rect 4693 -6477 4727 -6443
rect 4843 -6477 4877 -6443
rect 5393 -6427 5427 -6393
rect 5822 -6447 5856 -6413
rect 5972 -6397 6006 -6363
rect 5972 -6477 6006 -6443
rect 6272 -6317 6306 -6283
rect 6272 -6397 6306 -6363
rect 6272 -6477 6306 -6443
rect 6572 -6317 6606 -6283
rect 6952 -6327 6986 -6293
rect 6572 -6397 6606 -6363
rect 6572 -6477 6606 -6443
rect 6802 -6447 6836 -6413
rect 4443 -6597 4477 -6563
rect 1403 -6877 1437 -6843
rect 1403 -6957 1437 -6923
rect 1403 -7037 1437 -7003
rect 1883 -6877 1917 -6843
rect 1883 -6957 1917 -6923
rect 1883 -7037 1917 -7003
rect 2183 -6877 2217 -6843
rect 2183 -6957 2217 -6923
rect 2183 -7037 2217 -7003
rect 2483 -6877 2517 -6843
rect 2483 -6957 2517 -6923
rect 2483 -7037 2517 -7003
rect 2963 -6877 2997 -6843
rect 2963 -6957 2997 -6923
rect 2963 -7037 2997 -7003
rect 5393 -6547 5427 -6513
rect 4843 -6597 4877 -6563
rect 6322 -6597 6356 -6563
rect 5131 -6767 5165 -6733
rect 3377 -6957 3411 -6923
rect 3763 -6877 3797 -6843
rect 3763 -6957 3797 -6923
rect 3763 -7037 3797 -7003
rect 4093 -6877 4127 -6843
rect 4093 -6957 4127 -6923
rect 4093 -7037 4127 -7003
rect 4393 -6877 4427 -6843
rect 4393 -6957 4427 -6923
rect 4393 -7037 4427 -7003
rect 6722 -6597 6756 -6563
rect 7517 -5831 7551 -5797
rect 7152 -6717 7186 -6683
rect 4693 -6877 4727 -6843
rect 4693 -6957 4727 -6923
rect 4693 -7037 4727 -7003
rect 5023 -6877 5057 -6843
rect 5023 -6957 5057 -6923
rect 5023 -7037 5057 -7003
rect 5642 -6877 5676 -6843
rect 5642 -6957 5676 -6923
rect 5642 -7037 5676 -7003
rect 5972 -6877 6006 -6843
rect 5972 -6957 6006 -6923
rect 5972 -7037 6006 -7003
rect 6272 -6877 6306 -6843
rect 6272 -6957 6306 -6923
rect 6272 -7037 6306 -7003
rect 6572 -6877 6606 -6843
rect 6572 -6957 6606 -6923
rect 6572 -7037 6606 -7003
rect 7052 -6877 7086 -6843
rect 7052 -6957 7086 -6923
rect 7052 -7037 7086 -7003
rect 1515 -7157 1549 -7123
rect 5479 -7157 5513 -7123
rect 935 -7277 969 -7243
rect 1143 -7277 1177 -7243
rect 1223 -7277 1257 -7243
rect 1303 -7277 1337 -7243
rect 1383 -7277 1417 -7243
rect 1463 -7277 1497 -7243
rect 1543 -7277 1577 -7243
rect 1623 -7277 1657 -7243
rect 1703 -7277 1737 -7243
rect 1783 -7277 1817 -7243
rect 1863 -7277 1897 -7243
rect 1943 -7277 1977 -7243
rect 2023 -7277 2057 -7243
rect 2103 -7277 2137 -7243
rect 2183 -7277 2217 -7243
rect 2263 -7277 2297 -7243
rect 2343 -7277 2377 -7243
rect 2423 -7277 2457 -7243
rect 2503 -7277 2537 -7243
rect 2583 -7277 2617 -7243
rect 2663 -7277 2697 -7243
rect 2743 -7277 2777 -7243
rect 2823 -7277 2857 -7243
rect 2903 -7277 2937 -7243
rect 2983 -7277 3017 -7243
rect 3063 -7277 3097 -7243
rect 3143 -7277 3177 -7243
rect 3223 -7277 3257 -7243
rect 3753 -7277 3787 -7243
rect 3833 -7277 3867 -7243
rect 3913 -7277 3947 -7243
rect 3993 -7277 4027 -7243
rect 4073 -7277 4107 -7243
rect 4153 -7277 4187 -7243
rect 4233 -7277 4267 -7243
rect 4313 -7277 4347 -7243
rect 4393 -7277 4427 -7243
rect 4473 -7277 4507 -7243
rect 4553 -7277 4587 -7243
rect 4633 -7277 4667 -7243
rect 4713 -7277 4747 -7243
rect 4793 -7277 4827 -7243
rect 4873 -7277 4907 -7243
rect 4953 -7277 4987 -7243
rect 5033 -7277 5067 -7243
rect 5472 -7277 5506 -7243
rect 5552 -7277 5586 -7243
rect 5632 -7277 5666 -7243
rect 5712 -7277 5746 -7243
rect 5792 -7277 5826 -7243
rect 5872 -7277 5906 -7243
rect 5952 -7277 5986 -7243
rect 6032 -7277 6066 -7243
rect 6112 -7277 6146 -7243
rect 6192 -7277 6226 -7243
rect 6272 -7277 6306 -7243
rect 6352 -7277 6386 -7243
rect 6432 -7277 6466 -7243
rect 6512 -7277 6546 -7243
rect 6592 -7277 6626 -7243
rect 6672 -7277 6706 -7243
rect 6752 -7277 6786 -7243
rect 6832 -7277 6866 -7243
rect 6912 -7277 6946 -7243
rect 6992 -7277 7026 -7243
rect 7072 -7277 7106 -7243
rect 1515 -7397 1549 -7363
rect 5481 -7397 5515 -7363
rect 1403 -7517 1437 -7483
rect 1403 -7597 1437 -7563
rect 1403 -7677 1437 -7643
rect 1883 -7517 1917 -7483
rect 1883 -7597 1917 -7563
rect 1883 -7677 1917 -7643
rect 2183 -7517 2217 -7483
rect 2183 -7597 2217 -7563
rect 2183 -7677 2217 -7643
rect 2483 -7517 2517 -7483
rect 2483 -7597 2517 -7563
rect 2483 -7677 2517 -7643
rect 2963 -7517 2997 -7483
rect 2963 -7597 2997 -7563
rect 2963 -7677 2997 -7643
rect 3763 -7517 3797 -7483
rect 3377 -7595 3411 -7561
rect 3363 -7833 3397 -7799
rect 3763 -7597 3797 -7563
rect 3763 -7677 3797 -7643
rect 4093 -7517 4127 -7483
rect 4093 -7597 4127 -7563
rect 4093 -7677 4127 -7643
rect 4393 -7517 4427 -7483
rect 4393 -7597 4427 -7563
rect 4393 -7677 4427 -7643
rect 4693 -7517 4727 -7483
rect 4693 -7597 4727 -7563
rect 4693 -7677 4727 -7643
rect 5023 -7517 5057 -7483
rect 5023 -7597 5057 -7563
rect 5023 -7677 5057 -7643
rect 5642 -7517 5676 -7483
rect 5642 -7597 5676 -7563
rect 5642 -7677 5676 -7643
rect 5972 -7517 6006 -7483
rect 5972 -7597 6006 -7563
rect 5972 -7677 6006 -7643
rect 6272 -7517 6306 -7483
rect 6272 -7597 6306 -7563
rect 6272 -7677 6306 -7643
rect 6572 -7517 6606 -7483
rect 6572 -7597 6606 -7563
rect 6572 -7677 6606 -7643
rect 7052 -7517 7086 -7483
rect 7052 -7597 7086 -7563
rect 7052 -7677 7086 -7643
rect 2233 -7957 2267 -7923
rect 593 -8007 627 -7973
rect 1733 -8027 1767 -7993
rect 2603 -7947 2637 -7913
rect 479 -8107 513 -8073
rect 1603 -8127 1637 -8093
rect 1883 -8077 1917 -8043
rect 1883 -8157 1917 -8123
rect 821 -8225 855 -8191
rect 1733 -8227 1767 -8193
rect 1883 -8237 1917 -8203
rect 2183 -8077 2217 -8043
rect 2183 -8157 2217 -8123
rect 2183 -8237 2217 -8203
rect 2483 -8077 2517 -8043
rect 2763 -8027 2797 -7993
rect 2483 -8157 2517 -8123
rect 3213 -8127 3247 -8093
rect 2483 -8237 2517 -8203
rect 3063 -8227 3097 -8193
rect 5131 -7807 5165 -7773
rect 4443 -7957 4477 -7923
rect 4843 -7957 4877 -7923
rect 7156 -7838 7190 -7804
rect 6322 -7957 6356 -7923
rect 6722 -7957 6756 -7923
rect 3943 -8077 3977 -8043
rect 4093 -8077 4127 -8043
rect 4093 -8157 4127 -8123
rect 3655 -8261 3689 -8227
rect 707 -8307 741 -8273
rect 1603 -8327 1637 -8293
rect 4093 -8237 4127 -8203
rect 4393 -8077 4427 -8043
rect 4393 -8157 4427 -8123
rect 4393 -8237 4427 -8203
rect 4693 -8077 4727 -8043
rect 4843 -8077 4877 -8043
rect 4693 -8157 4727 -8123
rect 5131 -8146 5165 -8112
rect 5393 -8127 5427 -8093
rect 5822 -8107 5856 -8073
rect 5972 -8077 6006 -8043
rect 5972 -8157 6006 -8123
rect 4693 -8237 4727 -8203
rect 5822 -8227 5856 -8193
rect 5131 -8261 5165 -8227
rect 5972 -8237 6006 -8203
rect 6272 -8077 6306 -8043
rect 6272 -8157 6306 -8123
rect 6272 -8237 6306 -8203
rect 6572 -8077 6606 -8043
rect 6572 -8157 6606 -8123
rect 6802 -8107 6836 -8073
rect 6572 -8237 6606 -8203
rect 6952 -8227 6986 -8193
rect 2863 -8327 2897 -8293
rect 1143 -8457 1177 -8423
rect 1223 -8457 1257 -8423
rect 1303 -8457 1337 -8423
rect 1383 -8457 1417 -8423
rect 1463 -8457 1497 -8423
rect 1543 -8457 1577 -8423
rect 1623 -8457 1657 -8423
rect 1703 -8457 1737 -8423
rect 1783 -8457 1817 -8423
rect 1863 -8457 1897 -8423
rect 1943 -8457 1977 -8423
rect 2023 -8457 2057 -8423
rect 2103 -8457 2137 -8423
rect 2183 -8457 2217 -8423
rect 2263 -8457 2297 -8423
rect 2343 -8457 2377 -8423
rect 2423 -8457 2457 -8423
rect 2503 -8457 2537 -8423
rect 2583 -8457 2617 -8423
rect 2663 -8457 2697 -8423
rect 2743 -8457 2777 -8423
rect 2823 -8457 2857 -8423
rect 2903 -8457 2937 -8423
rect 2983 -8457 3017 -8423
rect 3063 -8457 3097 -8423
rect 3143 -8457 3177 -8423
rect 3223 -8457 3257 -8423
rect 3753 -8457 3787 -8423
rect 3833 -8457 3867 -8423
rect 3913 -8457 3947 -8423
rect 3993 -8457 4027 -8423
rect 4073 -8457 4107 -8423
rect 4153 -8457 4187 -8423
rect 4233 -8457 4267 -8423
rect 4313 -8457 4347 -8423
rect 4393 -8457 4427 -8423
rect 4473 -8457 4507 -8423
rect 4553 -8457 4587 -8423
rect 4633 -8457 4667 -8423
rect 4713 -8457 4747 -8423
rect 4793 -8457 4827 -8423
rect 4873 -8457 4907 -8423
rect 4953 -8457 4987 -8423
rect 5033 -8457 5067 -8423
rect 5472 -8457 5506 -8423
rect 5552 -8457 5586 -8423
rect 5632 -8457 5666 -8423
rect 5712 -8457 5746 -8423
rect 5792 -8457 5826 -8423
rect 5872 -8457 5906 -8423
rect 5952 -8457 5986 -8423
rect 6032 -8457 6066 -8423
rect 6112 -8457 6146 -8423
rect 6192 -8457 6226 -8423
rect 6272 -8457 6306 -8423
rect 6352 -8457 6386 -8423
rect 6432 -8457 6466 -8423
rect 6512 -8457 6546 -8423
rect 6592 -8457 6626 -8423
rect 6672 -8457 6706 -8423
rect 6752 -8457 6786 -8423
rect 6832 -8457 6866 -8423
rect 6912 -8457 6946 -8423
rect 6992 -8457 7026 -8423
rect 7072 -8457 7106 -8423
rect 1103 -8917 1137 -8883
rect 1183 -8917 1217 -8883
rect 1263 -8917 1297 -8883
rect 1343 -8917 1377 -8883
rect 1423 -8917 1457 -8883
rect 1503 -8917 1537 -8883
rect 1583 -8917 1617 -8883
rect 1663 -8917 1697 -8883
rect 1743 -8917 1777 -8883
rect 1823 -8917 1857 -8883
rect 1903 -8917 1937 -8883
rect 1983 -8917 2017 -8883
rect 2063 -8917 2097 -8883
rect 2143 -8917 2177 -8883
rect 2223 -8917 2257 -8883
rect 2303 -8917 2337 -8883
rect 2383 -8917 2417 -8883
rect 2463 -8917 2497 -8883
rect 2543 -8917 2577 -8883
rect 2623 -8917 2657 -8883
rect 2703 -8917 2737 -8883
rect 2783 -8917 2817 -8883
rect 2863 -8917 2897 -8883
rect 2943 -8917 2977 -8883
rect 3023 -8917 3057 -8883
rect 3103 -8917 3137 -8883
rect 3183 -8917 3217 -8883
rect 3693 -8917 3727 -8883
rect 3773 -8917 3807 -8883
rect 3853 -8917 3887 -8883
rect 3933 -8917 3967 -8883
rect 4013 -8917 4047 -8883
rect 4093 -8917 4127 -8883
rect 4173 -8917 4207 -8883
rect 4253 -8917 4287 -8883
rect 4333 -8917 4367 -8883
rect 4413 -8917 4447 -8883
rect 4493 -8917 4527 -8883
rect 4573 -8917 4607 -8883
rect 4653 -8917 4687 -8883
rect 4733 -8917 4767 -8883
rect 4813 -8917 4847 -8883
rect 4893 -8917 4927 -8883
rect 4973 -8917 5007 -8883
rect 5413 -8917 5447 -8883
rect 5493 -8917 5527 -8883
rect 5573 -8917 5607 -8883
rect 5653 -8917 5687 -8883
rect 5733 -8917 5767 -8883
rect 5813 -8917 5847 -8883
rect 5893 -8917 5927 -8883
rect 5973 -8917 6007 -8883
rect 6053 -8917 6087 -8883
rect 6133 -8917 6167 -8883
rect 6213 -8917 6247 -8883
rect 6293 -8917 6327 -8883
rect 6373 -8917 6407 -8883
rect 6453 -8917 6487 -8883
rect 6533 -8917 6567 -8883
rect 6613 -8917 6647 -8883
rect 6693 -8917 6727 -8883
rect 6773 -8917 6807 -8883
rect 6853 -8917 6887 -8883
rect 6933 -8917 6967 -8883
rect 7013 -8917 7047 -8883
rect 251 -9047 285 -9013
rect 1563 -9047 1597 -9013
rect 2823 -9047 2857 -9013
rect 365 -9147 399 -9113
rect 1693 -9147 1727 -9113
rect 1843 -9137 1877 -9103
rect 23 -9247 57 -9213
rect 1563 -9247 1597 -9213
rect 1843 -9217 1877 -9183
rect 137 -9347 171 -9313
rect 1693 -9347 1727 -9313
rect 1843 -9297 1877 -9263
rect 2143 -9137 2177 -9103
rect 2143 -9217 2177 -9183
rect 2143 -9297 2177 -9263
rect 2443 -9137 2477 -9103
rect 3023 -9147 3057 -9113
rect 3595 -9113 3629 -9079
rect 2443 -9217 2477 -9183
rect 2443 -9297 2477 -9263
rect 3173 -9247 3207 -9213
rect 2193 -9417 2227 -9383
rect 2723 -9347 2757 -9313
rect 2563 -9427 2597 -9393
rect 4033 -9137 4067 -9103
rect 4033 -9217 4067 -9183
rect 3883 -9297 3917 -9263
rect 4033 -9297 4067 -9263
rect 4333 -9137 4367 -9103
rect 4333 -9217 4367 -9183
rect 4333 -9297 4367 -9263
rect 4633 -9137 4667 -9103
rect 5333 -9147 5367 -9113
rect 5763 -9147 5797 -9113
rect 5913 -9137 5947 -9103
rect 4633 -9217 4667 -9183
rect 4633 -9297 4667 -9263
rect 4783 -9297 4817 -9263
rect 4383 -9417 4417 -9383
rect 3323 -9541 3357 -9507
rect 1363 -9697 1397 -9663
rect 1363 -9777 1397 -9743
rect 1363 -9857 1397 -9823
rect 1843 -9697 1877 -9663
rect 1843 -9777 1877 -9743
rect 1843 -9857 1877 -9823
rect 2143 -9697 2177 -9663
rect 2143 -9777 2177 -9743
rect 2143 -9857 2177 -9823
rect 2443 -9697 2477 -9663
rect 2443 -9777 2477 -9743
rect 2443 -9857 2477 -9823
rect 2923 -9697 2957 -9663
rect 2923 -9777 2957 -9743
rect 2923 -9857 2957 -9823
rect 4783 -9417 4817 -9383
rect 5071 -9423 5105 -9389
rect 5763 -9267 5797 -9233
rect 5913 -9217 5947 -9183
rect 5913 -9297 5947 -9263
rect 6213 -9137 6247 -9103
rect 6213 -9217 6247 -9183
rect 6213 -9297 6247 -9263
rect 6513 -9137 6547 -9103
rect 6893 -9147 6927 -9113
rect 6513 -9217 6547 -9183
rect 6513 -9297 6547 -9263
rect 6743 -9267 6777 -9233
rect 5333 -9367 5367 -9333
rect 5333 -9487 5367 -9453
rect 6263 -9417 6297 -9383
rect 6663 -9417 6697 -9383
rect 7096 -9537 7130 -9503
rect 3337 -9745 3371 -9711
rect 3703 -9697 3737 -9663
rect 3703 -9777 3737 -9743
rect 3703 -9857 3737 -9823
rect 4033 -9697 4067 -9663
rect 4033 -9777 4067 -9743
rect 4033 -9857 4067 -9823
rect 4333 -9697 4367 -9663
rect 4333 -9777 4367 -9743
rect 4333 -9857 4367 -9823
rect 4633 -9697 4667 -9663
rect 4633 -9777 4667 -9743
rect 4633 -9857 4667 -9823
rect 4963 -9697 4997 -9663
rect 4963 -9777 4997 -9743
rect 4963 -9857 4997 -9823
rect 5583 -9697 5617 -9663
rect 5583 -9777 5617 -9743
rect 5583 -9857 5617 -9823
rect 5913 -9697 5947 -9663
rect 5913 -9777 5947 -9743
rect 5913 -9857 5947 -9823
rect 6213 -9697 6247 -9663
rect 6213 -9777 6247 -9743
rect 6213 -9857 6247 -9823
rect 6513 -9697 6547 -9663
rect 6513 -9777 6547 -9743
rect 6513 -9857 6547 -9823
rect 6993 -9697 7027 -9663
rect 6993 -9777 7027 -9743
rect 6993 -9857 7027 -9823
rect 1194 -9977 1228 -9943
rect 5421 -9977 5455 -9943
rect 935 -10097 969 -10063
rect 1103 -10097 1137 -10063
rect 1183 -10097 1217 -10063
rect 1263 -10097 1297 -10063
rect 1343 -10097 1377 -10063
rect 1423 -10097 1457 -10063
rect 1503 -10097 1537 -10063
rect 1583 -10097 1617 -10063
rect 1663 -10097 1697 -10063
rect 1743 -10097 1777 -10063
rect 1823 -10097 1857 -10063
rect 1903 -10097 1937 -10063
rect 1983 -10097 2017 -10063
rect 2063 -10097 2097 -10063
rect 2143 -10097 2177 -10063
rect 2223 -10097 2257 -10063
rect 2303 -10097 2337 -10063
rect 2383 -10097 2417 -10063
rect 2463 -10097 2497 -10063
rect 2543 -10097 2577 -10063
rect 2623 -10097 2657 -10063
rect 2703 -10097 2737 -10063
rect 2783 -10097 2817 -10063
rect 2863 -10097 2897 -10063
rect 2943 -10097 2977 -10063
rect 3023 -10097 3057 -10063
rect 3103 -10097 3137 -10063
rect 3183 -10097 3217 -10063
rect 3693 -10097 3727 -10063
rect 3773 -10097 3807 -10063
rect 3853 -10097 3887 -10063
rect 3933 -10097 3967 -10063
rect 4013 -10097 4047 -10063
rect 4093 -10097 4127 -10063
rect 4173 -10097 4207 -10063
rect 4253 -10097 4287 -10063
rect 4333 -10097 4367 -10063
rect 4413 -10097 4447 -10063
rect 4493 -10097 4527 -10063
rect 4573 -10097 4607 -10063
rect 4653 -10097 4687 -10063
rect 4733 -10097 4767 -10063
rect 4813 -10097 4847 -10063
rect 4893 -10097 4927 -10063
rect 4973 -10097 5007 -10063
rect 5413 -10097 5447 -10063
rect 5493 -10097 5527 -10063
rect 5573 -10097 5607 -10063
rect 5653 -10097 5687 -10063
rect 5733 -10097 5767 -10063
rect 5813 -10097 5847 -10063
rect 5893 -10097 5927 -10063
rect 5973 -10097 6007 -10063
rect 6053 -10097 6087 -10063
rect 6133 -10097 6167 -10063
rect 6213 -10097 6247 -10063
rect 6293 -10097 6327 -10063
rect 6373 -10097 6407 -10063
rect 6453 -10097 6487 -10063
rect 6533 -10097 6567 -10063
rect 6613 -10097 6647 -10063
rect 6693 -10097 6727 -10063
rect 6773 -10097 6807 -10063
rect 6853 -10097 6887 -10063
rect 6933 -10097 6967 -10063
rect 7013 -10097 7047 -10063
rect 1194 -10217 1228 -10183
rect 5421 -10216 5455 -10182
rect 1363 -10337 1397 -10303
rect 1363 -10417 1397 -10383
rect 1363 -10497 1397 -10463
rect 1843 -10337 1877 -10303
rect 1843 -10417 1877 -10383
rect 1843 -10497 1877 -10463
rect 2143 -10337 2177 -10303
rect 2143 -10417 2177 -10383
rect 2143 -10497 2177 -10463
rect 2443 -10337 2477 -10303
rect 2443 -10417 2477 -10383
rect 2443 -10497 2477 -10463
rect 2923 -10337 2957 -10303
rect 2923 -10417 2957 -10383
rect 2923 -10497 2957 -10463
rect 3703 -10337 3737 -10303
rect 3337 -10440 3371 -10406
rect 3703 -10417 3737 -10383
rect 3703 -10497 3737 -10463
rect 4033 -10337 4067 -10303
rect 4033 -10417 4067 -10383
rect 4033 -10497 4067 -10463
rect 4333 -10337 4367 -10303
rect 4333 -10417 4367 -10383
rect 4333 -10497 4367 -10463
rect 4633 -10337 4667 -10303
rect 4633 -10417 4667 -10383
rect 4633 -10497 4667 -10463
rect 4963 -10337 4997 -10303
rect 4963 -10417 4997 -10383
rect 4963 -10497 4997 -10463
rect 5583 -10337 5617 -10303
rect 5583 -10417 5617 -10383
rect 5583 -10497 5617 -10463
rect 5913 -10337 5947 -10303
rect 5913 -10417 5947 -10383
rect 5913 -10497 5947 -10463
rect 6213 -10337 6247 -10303
rect 6213 -10417 6247 -10383
rect 6213 -10497 6247 -10463
rect 6513 -10337 6547 -10303
rect 6513 -10417 6547 -10383
rect 6513 -10497 6547 -10463
rect 6993 -10337 7027 -10303
rect 6993 -10417 7027 -10383
rect 6993 -10497 7027 -10463
rect 2193 -10777 2227 -10743
rect 821 -10847 855 -10813
rect 1693 -10847 1727 -10813
rect 2563 -10767 2597 -10733
rect 3323 -10767 3357 -10733
rect 707 -10947 741 -10913
rect 1563 -10947 1597 -10913
rect 1843 -10897 1877 -10863
rect 1843 -10977 1877 -10943
rect 593 -11047 627 -11013
rect 1693 -11047 1727 -11013
rect 1843 -11057 1877 -11023
rect 2143 -10897 2177 -10863
rect 2143 -10977 2177 -10943
rect 2143 -11057 2177 -11023
rect 2443 -10897 2477 -10863
rect 2723 -10847 2757 -10813
rect 2443 -10977 2477 -10943
rect 3173 -10947 3207 -10913
rect 2443 -11057 2477 -11023
rect 3023 -11047 3057 -11013
rect 5071 -10607 5105 -10573
rect 4383 -10777 4417 -10743
rect 4783 -10777 4817 -10743
rect 7096 -10657 7130 -10623
rect 6263 -10777 6297 -10743
rect 6663 -10777 6697 -10743
rect 3883 -10897 3917 -10863
rect 4033 -10897 4067 -10863
rect 4033 -10977 4067 -10943
rect 3595 -11081 3629 -11047
rect 479 -11147 513 -11113
rect 1563 -11147 1597 -11113
rect 4033 -11057 4067 -11023
rect 4333 -10897 4367 -10863
rect 4333 -10977 4367 -10943
rect 4333 -11057 4367 -11023
rect 4633 -10897 4667 -10863
rect 4783 -10897 4817 -10863
rect 4633 -10977 4667 -10943
rect 5071 -10935 5105 -10901
rect 5333 -10927 5367 -10893
rect 5763 -10927 5797 -10893
rect 5913 -10897 5947 -10863
rect 5913 -10977 5947 -10943
rect 4633 -11057 4667 -11023
rect 5333 -11048 5367 -11014
rect 5763 -11047 5797 -11013
rect 5913 -11057 5947 -11023
rect 6213 -10897 6247 -10863
rect 6213 -10977 6247 -10943
rect 6213 -11057 6247 -11023
rect 6513 -10897 6547 -10863
rect 6513 -10977 6547 -10943
rect 6743 -10927 6777 -10893
rect 6513 -11057 6547 -11023
rect 6893 -11047 6927 -11013
rect 2823 -11147 2857 -11113
rect 1103 -11277 1137 -11243
rect 1183 -11277 1217 -11243
rect 1263 -11277 1297 -11243
rect 1343 -11277 1377 -11243
rect 1423 -11277 1457 -11243
rect 1503 -11277 1537 -11243
rect 1583 -11277 1617 -11243
rect 1663 -11277 1697 -11243
rect 1743 -11277 1777 -11243
rect 1823 -11277 1857 -11243
rect 1903 -11277 1937 -11243
rect 1983 -11277 2017 -11243
rect 2063 -11277 2097 -11243
rect 2143 -11277 2177 -11243
rect 2223 -11277 2257 -11243
rect 2303 -11277 2337 -11243
rect 2383 -11277 2417 -11243
rect 2463 -11277 2497 -11243
rect 2543 -11277 2577 -11243
rect 2623 -11277 2657 -11243
rect 2703 -11277 2737 -11243
rect 2783 -11277 2817 -11243
rect 2863 -11277 2897 -11243
rect 2943 -11277 2977 -11243
rect 3023 -11277 3057 -11243
rect 3103 -11277 3137 -11243
rect 3183 -11277 3217 -11243
rect 3693 -11277 3727 -11243
rect 3773 -11277 3807 -11243
rect 3853 -11277 3887 -11243
rect 3933 -11277 3967 -11243
rect 4013 -11277 4047 -11243
rect 4093 -11277 4127 -11243
rect 4173 -11277 4207 -11243
rect 4253 -11277 4287 -11243
rect 4333 -11277 4367 -11243
rect 4413 -11277 4447 -11243
rect 4493 -11277 4527 -11243
rect 4573 -11277 4607 -11243
rect 4653 -11277 4687 -11243
rect 4733 -11277 4767 -11243
rect 4813 -11277 4847 -11243
rect 4893 -11277 4927 -11243
rect 4973 -11277 5007 -11243
rect 5413 -11277 5447 -11243
rect 5493 -11277 5527 -11243
rect 5573 -11277 5607 -11243
rect 5653 -11277 5687 -11243
rect 5733 -11277 5767 -11243
rect 5813 -11277 5847 -11243
rect 5893 -11277 5927 -11243
rect 5973 -11277 6007 -11243
rect 6053 -11277 6087 -11243
rect 6133 -11277 6167 -11243
rect 6213 -11277 6247 -11243
rect 6293 -11277 6327 -11243
rect 6373 -11277 6407 -11243
rect 6453 -11277 6487 -11243
rect 6533 -11277 6567 -11243
rect 6613 -11277 6647 -11243
rect 6693 -11277 6727 -11243
rect 6773 -11277 6807 -11243
rect 6853 -11277 6887 -11243
rect 6933 -11277 6967 -11243
rect 7013 -11277 7047 -11243
rect 5421 -11511 5455 -11477
rect 1184 -11737 1218 -11703
rect 1264 -11737 1298 -11703
rect 1344 -11737 1378 -11703
rect 1424 -11737 1458 -11703
rect 1504 -11737 1538 -11703
rect 1584 -11737 1618 -11703
rect 1664 -11737 1698 -11703
rect 1744 -11737 1778 -11703
rect 1824 -11737 1858 -11703
rect 1904 -11737 1938 -11703
rect 1984 -11737 2018 -11703
rect 2064 -11737 2098 -11703
rect 2144 -11737 2178 -11703
rect 2224 -11737 2258 -11703
rect 2304 -11737 2338 -11703
rect 2384 -11737 2418 -11703
rect 2464 -11737 2498 -11703
rect 2544 -11737 2578 -11703
rect 2624 -11737 2658 -11703
rect 2704 -11737 2738 -11703
rect 2784 -11737 2818 -11703
rect 2864 -11737 2898 -11703
rect 2944 -11737 2978 -11703
rect 3024 -11737 3058 -11703
rect 3104 -11737 3138 -11703
rect 3554 -11737 3588 -11703
rect 3634 -11737 3668 -11703
rect 3714 -11737 3748 -11703
rect 3794 -11737 3828 -11703
rect 3874 -11737 3908 -11703
rect 3954 -11737 3988 -11703
rect 4034 -11737 4068 -11703
rect 4114 -11737 4148 -11703
rect 4194 -11737 4228 -11703
rect 4274 -11737 4308 -11703
rect 4354 -11737 4388 -11703
rect 4434 -11737 4468 -11703
rect 4514 -11737 4548 -11703
rect 4594 -11737 4628 -11703
rect 4674 -11737 4708 -11703
rect 4754 -11737 4788 -11703
rect 4834 -11737 4868 -11703
rect 593 -11857 627 -11823
rect 1604 -11857 1638 -11823
rect 2974 -11857 3008 -11823
rect 7366 -11544 7400 -11510
rect 5274 -11738 5308 -11704
rect 5354 -11738 5388 -11704
rect 5434 -11738 5468 -11704
rect 5514 -11738 5548 -11704
rect 5594 -11738 5628 -11704
rect 5674 -11738 5708 -11704
rect 5754 -11738 5788 -11704
rect 5834 -11738 5868 -11704
rect 5914 -11738 5948 -11704
rect 5994 -11738 6028 -11704
rect 6074 -11738 6108 -11704
rect 6154 -11738 6188 -11704
rect 6234 -11738 6268 -11704
rect 6314 -11738 6348 -11704
rect 6394 -11738 6428 -11704
rect 6474 -11738 6508 -11704
rect 6554 -11738 6588 -11704
rect 6634 -11738 6668 -11704
rect 6714 -11738 6748 -11704
rect 6794 -11738 6828 -11704
rect 6874 -11738 6908 -11704
rect 6954 -11738 6988 -11704
rect 7034 -11738 7068 -11704
rect 7114 -11738 7148 -11704
rect 7194 -11738 7228 -11704
rect 5404 -11863 5438 -11829
rect 6684 -11868 6718 -11834
rect 7252 -11868 7286 -11834
rect 23 -11977 57 -11943
rect 1694 -11977 1728 -11943
rect 1844 -11957 1878 -11923
rect 707 -12073 741 -12039
rect 1844 -12037 1878 -12003
rect 479 -12153 513 -12119
rect 1664 -12097 1698 -12063
rect 1844 -12117 1878 -12083
rect 2144 -11957 2178 -11923
rect 2144 -12037 2178 -12003
rect 2144 -12117 2178 -12083
rect 2444 -11957 2478 -11923
rect 2824 -11977 2858 -11943
rect 3894 -11957 3928 -11923
rect 2444 -12037 2478 -12003
rect 3894 -12037 3928 -12003
rect 2444 -12117 2478 -12083
rect 2694 -12097 2728 -12063
rect 3456 -12117 3490 -12083
rect 3744 -12117 3778 -12083
rect 3894 -12117 3928 -12083
rect 4194 -11957 4228 -11923
rect 4194 -12037 4228 -12003
rect 4194 -12117 4228 -12083
rect 4494 -11957 4528 -11923
rect 5027 -11944 5061 -11910
rect 4494 -12037 4528 -12003
rect 5504 -11988 5538 -11954
rect 5934 -11958 5968 -11924
rect 4494 -12117 4528 -12083
rect 5704 -12078 5738 -12044
rect 4644 -12117 4678 -12083
rect 5934 -12038 5968 -12004
rect 5203 -12140 5237 -12106
rect 5934 -12118 5968 -12084
rect 137 -12247 171 -12213
rect 2194 -12237 2228 -12203
rect 821 -12347 855 -12313
rect 2594 -12237 2628 -12203
rect 3174 -12356 3208 -12322
rect 4244 -12237 4278 -12203
rect 6234 -11958 6268 -11924
rect 6234 -12038 6268 -12004
rect 6234 -12118 6268 -12084
rect 6534 -11958 6568 -11924
rect 6804 -11978 6838 -11944
rect 7056 -11978 7090 -11944
rect 6534 -12038 6568 -12004
rect 6534 -12118 6568 -12084
rect 6684 -12078 6718 -12044
rect 4644 -12237 4678 -12203
rect 5204 -12254 5238 -12220
rect 5784 -12238 5818 -12204
rect 6184 -12238 6218 -12204
rect 7298 -12166 7332 -12132
rect 4938 -12407 4972 -12373
rect 5204 -12368 5238 -12334
rect 1214 -12517 1248 -12483
rect 1214 -12597 1248 -12563
rect 1214 -12677 1248 -12643
rect 1514 -12517 1548 -12483
rect 1514 -12597 1548 -12563
rect 1514 -12677 1548 -12643
rect 1844 -12517 1878 -12483
rect 1844 -12597 1878 -12563
rect 1844 -12677 1878 -12643
rect 2144 -12517 2178 -12483
rect 2144 -12597 2178 -12563
rect 2144 -12677 2178 -12643
rect 2444 -12517 2478 -12483
rect 2444 -12597 2478 -12563
rect 2444 -12677 2478 -12643
rect 3074 -12517 3108 -12483
rect 3074 -12597 3108 -12563
rect 3074 -12677 3108 -12643
rect 3564 -12517 3598 -12483
rect 3564 -12597 3598 -12563
rect 3564 -12677 3598 -12643
rect 3894 -12517 3928 -12483
rect 3894 -12597 3928 -12563
rect 3894 -12677 3928 -12643
rect 4194 -12517 4228 -12483
rect 4194 -12597 4228 -12563
rect 4194 -12677 4228 -12643
rect 4494 -12517 4528 -12483
rect 4494 -12597 4528 -12563
rect 4494 -12677 4528 -12643
rect 6814 -12368 6848 -12334
rect 4824 -12517 4858 -12483
rect 5021 -12521 5055 -12487
rect 5304 -12518 5338 -12484
rect 4824 -12597 4858 -12563
rect 4824 -12677 4858 -12643
rect 5304 -12598 5338 -12564
rect 5304 -12678 5338 -12644
rect 5604 -12518 5638 -12484
rect 5604 -12598 5638 -12564
rect 5604 -12678 5638 -12644
rect 5934 -12518 5968 -12484
rect 5934 -12598 5968 -12564
rect 5934 -12678 5968 -12644
rect 6234 -12518 6268 -12484
rect 6234 -12598 6268 -12564
rect 6234 -12678 6268 -12644
rect 6534 -12518 6568 -12484
rect 6534 -12598 6568 -12564
rect 6534 -12678 6568 -12644
rect 7164 -12518 7198 -12484
rect 7164 -12598 7198 -12564
rect 7164 -12678 7198 -12644
rect 1194 -12797 1228 -12763
rect 5115 -12799 5149 -12765
rect 935 -12917 969 -12883
rect 1184 -12917 1218 -12883
rect 1264 -12917 1298 -12883
rect 1344 -12917 1378 -12883
rect 1424 -12917 1458 -12883
rect 1504 -12917 1538 -12883
rect 1584 -12917 1618 -12883
rect 1664 -12917 1698 -12883
rect 1744 -12917 1778 -12883
rect 1824 -12917 1858 -12883
rect 1904 -12917 1938 -12883
rect 1984 -12917 2018 -12883
rect 2064 -12917 2098 -12883
rect 2144 -12917 2178 -12883
rect 2224 -12917 2258 -12883
rect 2304 -12917 2338 -12883
rect 2384 -12917 2418 -12883
rect 2464 -12917 2498 -12883
rect 2544 -12917 2578 -12883
rect 2624 -12917 2658 -12883
rect 2704 -12917 2738 -12883
rect 2784 -12917 2818 -12883
rect 2864 -12917 2898 -12883
rect 2944 -12917 2978 -12883
rect 3024 -12917 3058 -12883
rect 3104 -12917 3138 -12883
rect 3554 -12917 3588 -12883
rect 3634 -12917 3668 -12883
rect 3714 -12917 3748 -12883
rect 3794 -12917 3828 -12883
rect 3874 -12917 3908 -12883
rect 3954 -12917 3988 -12883
rect 4034 -12917 4068 -12883
rect 4114 -12917 4148 -12883
rect 4194 -12917 4228 -12883
rect 4274 -12917 4308 -12883
rect 4354 -12917 4388 -12883
rect 4434 -12917 4468 -12883
rect 4514 -12917 4548 -12883
rect 4594 -12917 4628 -12883
rect 4674 -12917 4708 -12883
rect 4754 -12917 4788 -12883
rect 4834 -12917 4868 -12883
rect 5274 -12918 5308 -12884
rect 5354 -12918 5388 -12884
rect 5434 -12918 5468 -12884
rect 5514 -12918 5548 -12884
rect 5594 -12918 5628 -12884
rect 5674 -12918 5708 -12884
rect 5754 -12918 5788 -12884
rect 5834 -12918 5868 -12884
rect 5914 -12918 5948 -12884
rect 5994 -12918 6028 -12884
rect 6074 -12918 6108 -12884
rect 6154 -12918 6188 -12884
rect 6234 -12918 6268 -12884
rect 6314 -12918 6348 -12884
rect 6394 -12918 6428 -12884
rect 6474 -12918 6508 -12884
rect 6554 -12918 6588 -12884
rect 6634 -12918 6668 -12884
rect 6714 -12918 6748 -12884
rect 6794 -12918 6828 -12884
rect 6874 -12918 6908 -12884
rect 6954 -12918 6988 -12884
rect 7034 -12918 7068 -12884
rect 7114 -12918 7148 -12884
rect 7194 -12918 7228 -12884
<< metal1 >>
rect 1020 2487 5320 2511
rect 1020 2435 1034 2487
rect 1086 2478 5320 2487
rect 1086 2444 1103 2478
rect 1137 2444 1183 2478
rect 1217 2444 1263 2478
rect 1297 2444 1343 2478
rect 1377 2444 1423 2478
rect 1457 2444 1503 2478
rect 1537 2444 1583 2478
rect 1617 2444 1663 2478
rect 1697 2444 1743 2478
rect 1777 2444 1823 2478
rect 1857 2444 1903 2478
rect 1937 2444 1983 2478
rect 2017 2444 2063 2478
rect 2097 2444 2143 2478
rect 2177 2444 2223 2478
rect 2257 2444 2303 2478
rect 2337 2444 2383 2478
rect 2417 2444 2463 2478
rect 2497 2444 2543 2478
rect 2577 2444 2623 2478
rect 2657 2444 2703 2478
rect 2737 2444 2783 2478
rect 2817 2444 2863 2478
rect 2897 2444 2943 2478
rect 2977 2444 3023 2478
rect 3057 2444 3103 2478
rect 3137 2444 3183 2478
rect 3217 2444 3663 2478
rect 3697 2444 3743 2478
rect 3777 2444 3823 2478
rect 3857 2444 3903 2478
rect 3937 2444 3983 2478
rect 4017 2444 4063 2478
rect 4097 2444 4143 2478
rect 4177 2444 4223 2478
rect 4257 2444 4303 2478
rect 4337 2444 4383 2478
rect 4417 2444 4463 2478
rect 4497 2444 4543 2478
rect 4577 2444 4623 2478
rect 4657 2444 4703 2478
rect 4737 2444 4783 2478
rect 4817 2444 4863 2478
rect 4897 2444 4943 2478
rect 4977 2444 5023 2478
rect 5057 2444 5103 2478
rect 5137 2444 5183 2478
rect 5217 2444 5263 2478
rect 5297 2444 5320 2478
rect 1086 2435 5320 2444
rect 1020 2411 5320 2435
rect 5660 2487 7340 2511
rect 5660 2478 5844 2487
rect 5896 2478 7340 2487
rect 5660 2444 5683 2478
rect 5717 2444 5763 2478
rect 5797 2444 5843 2478
rect 5896 2444 5923 2478
rect 5957 2444 6003 2478
rect 6037 2444 6083 2478
rect 6117 2444 6163 2478
rect 6197 2444 6243 2478
rect 6277 2444 6323 2478
rect 6357 2444 6403 2478
rect 6437 2444 6483 2478
rect 6517 2444 6563 2478
rect 6597 2444 6643 2478
rect 6677 2444 6723 2478
rect 6757 2444 6803 2478
rect 6837 2444 6883 2478
rect 6917 2444 6963 2478
rect 6997 2444 7043 2478
rect 7077 2444 7123 2478
rect 7157 2444 7203 2478
rect 7237 2444 7283 2478
rect 7317 2444 7340 2478
rect 5660 2435 5844 2444
rect 5896 2435 7340 2444
rect 5660 2411 7340 2435
rect 228 2370 308 2383
rect 0 2328 80 2351
rect 0 2294 23 2328
rect 57 2294 80 2328
rect 0 -672 80 2294
rect 0 -706 23 -672
rect 57 -706 80 -672
rect 0 -3752 80 -706
rect 0 -3786 23 -3752
rect 57 -3786 80 -3752
rect 0 -5532 80 -3786
rect 0 -5566 23 -5532
rect 57 -5566 80 -5532
rect 0 -6394 80 -5566
rect 0 -6428 23 -6394
rect 57 -6428 80 -6394
rect 0 -9213 80 -6428
rect 0 -9247 23 -9213
rect 57 -9247 80 -9213
rect 0 -11943 80 -9247
rect 0 -11977 23 -11943
rect 57 -11977 80 -11943
rect 0 -12957 80 -11977
rect 114 2228 194 2351
rect 114 2194 137 2228
rect 171 2194 194 2228
rect 114 -793 194 2194
rect 114 -827 137 -793
rect 171 -827 194 -793
rect 114 -3485 194 -827
rect 114 -3519 137 -3485
rect 171 -3519 194 -3485
rect 114 -5152 194 -3519
rect 114 -5186 137 -5152
rect 171 -5186 194 -5152
rect 114 -6513 194 -5186
rect 114 -6547 137 -6513
rect 171 -6547 194 -6513
rect 114 -9313 194 -6547
rect 114 -9347 137 -9313
rect 171 -9347 194 -9313
rect 114 -12213 194 -9347
rect 114 -12247 137 -12213
rect 171 -12247 194 -12213
rect 114 -12957 194 -12247
rect 228 2318 242 2370
rect 294 2318 308 2370
rect 228 688 308 2318
rect 228 654 251 688
rect 285 654 308 688
rect 228 -2592 308 654
rect 228 -2626 251 -2592
rect 285 -2626 308 -2592
rect 228 -3382 308 -2626
rect 228 -3416 251 -3382
rect 285 -3416 308 -3382
rect 228 -5652 308 -3416
rect 228 -5686 251 -5652
rect 285 -5686 308 -5652
rect 228 -6173 308 -5686
rect 228 -6207 251 -6173
rect 285 -6207 308 -6173
rect 228 -7552 308 -6207
rect 228 -7604 242 -7552
rect 294 -7604 308 -7552
rect 228 -9013 308 -7604
rect 228 -9047 251 -9013
rect 285 -9047 308 -9013
rect 228 -11105 308 -9047
rect 228 -11157 242 -11105
rect 294 -11157 308 -11105
rect 228 -12957 308 -11157
rect 342 1536 422 2351
rect 342 1484 356 1536
rect 408 1484 422 1536
rect 342 468 422 1484
rect 342 434 365 468
rect 399 434 422 468
rect 342 -2472 422 434
rect 342 -2506 365 -2472
rect 399 -2506 422 -2472
rect 342 -3652 422 -2506
rect 342 -3686 365 -3652
rect 399 -3686 422 -3652
rect 342 -5252 422 -3686
rect 342 -5286 365 -5252
rect 399 -5286 422 -5252
rect 342 -6287 422 -5286
rect 342 -6321 365 -6287
rect 399 -6321 422 -6287
rect 342 -8287 422 -6321
rect 342 -8339 356 -8287
rect 408 -8339 422 -8287
rect 342 -9113 422 -8339
rect 342 -9147 365 -9113
rect 399 -9147 422 -9113
rect 342 -10398 422 -9147
rect 342 -10450 356 -10398
rect 408 -10450 422 -10398
rect 342 -12957 422 -10450
rect 456 1696 536 2351
rect 456 1644 470 1696
rect 522 1644 536 1696
rect 456 348 536 1644
rect 456 314 479 348
rect 513 314 536 348
rect 456 -492 536 314
rect 456 -526 479 -492
rect 513 -526 536 -492
rect 456 -2564 536 -526
rect 570 2227 650 2351
rect 570 2175 584 2227
rect 636 2175 650 2227
rect 570 574 650 2175
rect 570 540 593 574
rect 627 540 650 574
rect 570 -572 650 540
rect 570 -606 593 -572
rect 627 -606 650 -572
rect 570 -1844 650 -606
rect 568 -1857 650 -1844
rect 568 -1909 582 -1857
rect 634 -1909 650 -1857
rect 568 -1924 650 -1909
rect 456 -2616 470 -2564
rect 522 -2616 536 -2564
rect 456 -5412 536 -2616
rect 456 -5446 479 -5412
rect 513 -5446 536 -5412
rect 456 -6914 536 -5446
rect 456 -6966 470 -6914
rect 522 -6966 536 -6914
rect 456 -8073 536 -6966
rect 456 -8107 479 -8073
rect 513 -8107 536 -8073
rect 456 -11113 536 -8107
rect 456 -11147 479 -11113
rect 513 -11147 536 -11113
rect 456 -12119 536 -11147
rect 456 -12153 479 -12119
rect 513 -12153 536 -12119
rect 456 -12957 536 -12153
rect 570 -5012 650 -1924
rect 570 -5046 593 -5012
rect 627 -5046 650 -5012
rect 570 -6183 650 -5046
rect 570 -6235 584 -6183
rect 636 -6235 650 -6183
rect 570 -7973 650 -6235
rect 570 -8007 593 -7973
rect 627 -8007 650 -7973
rect 570 -11013 650 -8007
rect 570 -11047 593 -11013
rect 627 -11047 650 -11013
rect 570 -11823 650 -11047
rect 570 -11857 593 -11823
rect 627 -11857 650 -11823
rect 570 -12957 650 -11857
rect 684 2128 764 2351
rect 684 2094 707 2128
rect 741 2094 764 2128
rect 684 -460 764 2094
rect 684 -512 698 -460
rect 750 -512 764 -460
rect 684 -2352 764 -512
rect 684 -2386 707 -2352
rect 741 -2386 764 -2352
rect 684 -3578 764 -2386
rect 684 -3612 707 -3578
rect 741 -3612 764 -3578
rect 684 -5332 764 -3612
rect 684 -5366 707 -5332
rect 741 -5366 764 -5332
rect 684 -8273 764 -5366
rect 684 -8307 707 -8273
rect 741 -8307 764 -8273
rect 684 -9702 764 -8307
rect 684 -9754 698 -9702
rect 750 -9754 764 -9702
rect 684 -10913 764 -9754
rect 684 -10947 707 -10913
rect 741 -10947 764 -10913
rect 684 -12039 764 -10947
rect 684 -12073 707 -12039
rect 741 -12073 764 -12039
rect 684 -12957 764 -12073
rect 798 2028 878 2351
rect 798 1994 821 2028
rect 855 1994 878 2028
rect 798 -1161 878 1994
rect 798 -1213 812 -1161
rect 864 -1213 878 -1161
rect 798 -2252 878 -1213
rect 798 -2286 821 -2252
rect 855 -2286 878 -2252
rect 798 -3262 878 -2286
rect 798 -3296 821 -3262
rect 855 -3296 878 -3262
rect 798 -5812 878 -3296
rect 798 -5846 821 -5812
rect 855 -5846 878 -5812
rect 798 -8191 878 -5846
rect 798 -8225 821 -8191
rect 855 -8225 878 -8191
rect 798 -9002 878 -8225
rect 798 -9054 812 -9002
rect 864 -9054 878 -9002
rect 798 -10813 878 -9054
rect 798 -10847 821 -10813
rect 855 -10847 878 -10813
rect 798 -12313 878 -10847
rect 798 -12347 821 -12313
rect 855 -12347 878 -12313
rect 798 -12956 878 -12347
rect 912 1298 992 2351
rect 1360 1731 1400 2411
rect 1540 2357 1620 2371
rect 1540 2305 1554 2357
rect 1606 2305 1620 2357
rect 1540 2291 1620 2305
rect 1670 2257 1750 2271
rect 1670 2205 1684 2257
rect 1736 2205 1750 2257
rect 1670 2191 1750 2205
rect 1820 2258 1900 2411
rect 1820 2224 1843 2258
rect 1877 2224 1900 2258
rect 1820 2178 1900 2224
rect 1540 2157 1620 2171
rect 1540 2105 1554 2157
rect 1606 2105 1620 2157
rect 1540 2091 1620 2105
rect 1820 2144 1843 2178
rect 1877 2144 1900 2178
rect 1820 2098 1900 2144
rect 1670 2057 1750 2071
rect 1670 2005 1684 2057
rect 1736 2005 1750 2057
rect 1820 2064 1843 2098
rect 1877 2064 1900 2098
rect 1820 2041 1900 2064
rect 2120 2258 2200 2411
rect 2120 2224 2143 2258
rect 2177 2224 2200 2258
rect 2120 2178 2200 2224
rect 2120 2144 2143 2178
rect 2177 2144 2200 2178
rect 2120 2098 2200 2144
rect 2120 2064 2143 2098
rect 2177 2064 2200 2098
rect 2120 2041 2200 2064
rect 2420 2258 2500 2411
rect 2800 2357 2880 2371
rect 2800 2305 2814 2357
rect 2866 2305 2880 2357
rect 2800 2291 2880 2305
rect 2420 2224 2443 2258
rect 2477 2224 2500 2258
rect 2420 2178 2500 2224
rect 2420 2144 2443 2178
rect 2477 2144 2500 2178
rect 2420 2098 2500 2144
rect 2420 2064 2443 2098
rect 2477 2064 2500 2098
rect 2420 2041 2500 2064
rect 2700 2057 2780 2071
rect 1670 1991 1750 2005
rect 2700 2005 2714 2057
rect 2766 2005 2780 2057
rect 2170 1978 2250 2001
rect 2700 1991 2780 2005
rect 2170 1944 2193 1978
rect 2227 1961 2250 1978
rect 2540 1968 2620 1991
rect 2540 1961 2563 1968
rect 2227 1944 2563 1961
rect 2170 1934 2563 1944
rect 2597 1934 2620 1968
rect 2170 1921 2620 1934
rect 2540 1911 2620 1921
rect 2920 1731 2960 2411
rect 2988 2370 3068 2383
rect 2988 2318 3002 2370
rect 3054 2363 3068 2370
rect 3054 2323 3620 2363
rect 3054 2318 3068 2323
rect 2988 2303 3068 2318
rect 3000 2257 3080 2271
rect 3580 2261 3620 2323
rect 3000 2205 3014 2257
rect 3066 2205 3080 2257
rect 3000 2191 3080 2205
rect 3268 2230 3348 2243
rect 3268 2178 3282 2230
rect 3334 2223 3348 2230
rect 3560 2238 3640 2261
rect 3334 2183 3532 2223
rect 3334 2178 3348 2183
rect 3150 2157 3230 2171
rect 3268 2163 3348 2178
rect 3150 2105 3164 2157
rect 3216 2105 3230 2157
rect 3150 2091 3230 2105
rect 3492 2121 3532 2183
rect 3560 2204 3583 2238
rect 3617 2204 3640 2238
rect 3560 2181 3640 2204
rect 3560 2121 3640 2141
rect 3492 2118 3640 2121
rect 3492 2084 3583 2118
rect 3617 2084 3640 2118
rect 3492 2081 3640 2084
rect 3300 2065 3380 2079
rect 3300 2013 3314 2065
rect 3366 2013 3380 2065
rect 3560 2061 3640 2081
rect 3300 1999 3380 2013
rect 3560 2001 3640 2021
rect 3492 1998 3640 2001
rect 3054 1977 3134 1991
rect 3054 1925 3068 1977
rect 3120 1925 3134 1977
rect 3054 1911 3134 1925
rect 3492 1964 3583 1998
rect 3617 1964 3640 1998
rect 3492 1961 3640 1964
rect 3300 1863 3380 1877
rect 3300 1811 3314 1863
rect 3366 1811 3380 1863
rect 3300 1797 3380 1811
rect 1340 1698 1420 1731
rect 1340 1664 1363 1698
rect 1397 1664 1420 1698
rect 1340 1618 1420 1664
rect 1340 1584 1363 1618
rect 1397 1584 1420 1618
rect 1340 1538 1420 1584
rect 1340 1504 1363 1538
rect 1397 1504 1420 1538
rect 1340 1481 1420 1504
rect 1820 1698 1900 1731
rect 1820 1664 1843 1698
rect 1877 1664 1900 1698
rect 1820 1618 1900 1664
rect 1820 1584 1843 1618
rect 1877 1584 1900 1618
rect 1820 1538 1900 1584
rect 1820 1504 1843 1538
rect 1877 1504 1900 1538
rect 1820 1481 1900 1504
rect 2120 1698 2200 1731
rect 2120 1664 2143 1698
rect 2177 1664 2200 1698
rect 2120 1618 2200 1664
rect 2120 1584 2143 1618
rect 2177 1584 2200 1618
rect 2120 1538 2200 1584
rect 2120 1504 2143 1538
rect 2177 1504 2200 1538
rect 2120 1481 2200 1504
rect 2420 1698 2500 1731
rect 2420 1664 2443 1698
rect 2477 1664 2500 1698
rect 2420 1618 2500 1664
rect 2420 1584 2443 1618
rect 2477 1584 2500 1618
rect 2420 1538 2500 1584
rect 2420 1504 2443 1538
rect 2477 1504 2500 1538
rect 2420 1481 2500 1504
rect 2900 1698 2980 1731
rect 2900 1664 2923 1698
rect 2957 1664 2980 1698
rect 2900 1618 2980 1664
rect 3335 1696 3415 1709
rect 3335 1644 3349 1696
rect 3401 1689 3415 1696
rect 3492 1689 3532 1961
rect 3560 1941 3640 1961
rect 3560 1878 3640 1901
rect 3560 1844 3583 1878
rect 3617 1844 3640 1878
rect 3560 1821 3640 1844
rect 3401 1649 3532 1689
rect 3401 1644 3415 1649
rect 3335 1629 3415 1644
rect 2900 1584 2923 1618
rect 2957 1584 2980 1618
rect 2900 1538 2980 1584
rect 2900 1504 2923 1538
rect 2957 1504 2980 1538
rect 2900 1481 2980 1504
rect 3335 1536 3415 1549
rect 3335 1484 3349 1536
rect 3401 1529 3415 1536
rect 3580 1529 3620 1821
rect 3680 1731 3720 2411
rect 4140 2258 4220 2411
rect 3990 2227 4070 2241
rect 3990 2175 4004 2227
rect 4056 2175 4070 2227
rect 3990 2161 4070 2175
rect 4140 2224 4163 2258
rect 4197 2224 4220 2258
rect 4140 2178 4220 2224
rect 4140 2144 4163 2178
rect 4197 2144 4220 2178
rect 3990 2107 4070 2121
rect 3990 2055 4004 2107
rect 4056 2055 4070 2107
rect 3990 2041 4070 2055
rect 4140 2098 4220 2144
rect 4140 2064 4163 2098
rect 4197 2064 4220 2098
rect 4140 2041 4220 2064
rect 4440 2258 4520 2411
rect 4440 2224 4463 2258
rect 4497 2224 4520 2258
rect 4440 2178 4520 2224
rect 4440 2144 4463 2178
rect 4497 2144 4520 2178
rect 4440 2098 4520 2144
rect 4440 2064 4463 2098
rect 4497 2064 4520 2098
rect 4440 2041 4520 2064
rect 4740 2258 4820 2411
rect 4740 2224 4763 2258
rect 4797 2224 4820 2258
rect 4740 2178 4820 2224
rect 4740 2144 4763 2178
rect 4797 2144 4820 2178
rect 4740 2098 4820 2144
rect 4740 2064 4763 2098
rect 4797 2064 4820 2098
rect 4740 2041 4820 2064
rect 4970 2107 5050 2121
rect 4970 2055 4984 2107
rect 5036 2055 5050 2107
rect 4970 2041 5050 2055
rect 4490 1981 4570 2001
rect 4890 1981 4970 2001
rect 4490 1978 4970 1981
rect 4490 1944 4513 1978
rect 4547 1944 4913 1978
rect 4947 1944 4970 1978
rect 4490 1941 4970 1944
rect 4490 1921 4570 1941
rect 4890 1921 4970 1941
rect 5090 1731 5130 2411
rect 5284 2335 5364 2349
rect 5284 2283 5298 2335
rect 5350 2283 5364 2335
rect 5284 2251 5364 2283
rect 5580 2251 5660 2271
rect 5284 2248 5660 2251
rect 5170 2227 5250 2241
rect 5170 2175 5184 2227
rect 5236 2175 5250 2227
rect 5284 2214 5603 2248
rect 5637 2214 5660 2248
rect 5284 2211 5660 2214
rect 5580 2191 5660 2211
rect 5170 2161 5250 2175
rect 5250 2104 5330 2127
rect 5250 2070 5273 2104
rect 5307 2070 5330 2104
rect 5250 2047 5330 2070
rect 5269 1901 5309 2047
rect 5580 2027 5660 2050
rect 5580 2010 5603 2027
rect 5370 1996 5603 2010
rect 5370 1944 5384 1996
rect 5436 1993 5603 1996
rect 5637 1993 5660 2027
rect 5436 1970 5660 1993
rect 5436 1944 5450 1970
rect 5370 1930 5450 1944
rect 5250 1878 5330 1901
rect 5250 1844 5273 1878
rect 5307 1844 5330 1878
rect 5250 1821 5330 1844
rect 5850 1731 5890 2411
rect 6010 2257 6090 2271
rect 6010 2205 6024 2257
rect 6076 2205 6090 2257
rect 6010 2191 6090 2205
rect 6160 2258 6240 2411
rect 6160 2224 6183 2258
rect 6217 2224 6240 2258
rect 6160 2178 6240 2224
rect 6010 2137 6090 2151
rect 6010 2085 6024 2137
rect 6076 2085 6090 2137
rect 6010 2071 6090 2085
rect 6160 2144 6183 2178
rect 6217 2144 6240 2178
rect 6160 2098 6240 2144
rect 6160 2064 6183 2098
rect 6217 2064 6240 2098
rect 6160 2041 6240 2064
rect 6460 2258 6540 2411
rect 6460 2224 6483 2258
rect 6517 2224 6540 2258
rect 6460 2178 6540 2224
rect 6460 2144 6483 2178
rect 6517 2144 6540 2178
rect 6460 2098 6540 2144
rect 6460 2064 6483 2098
rect 6517 2064 6540 2098
rect 6460 2041 6540 2064
rect 6760 2258 6840 2411
rect 6760 2224 6783 2258
rect 6817 2224 6840 2258
rect 6760 2178 6840 2224
rect 7140 2257 7220 2271
rect 7140 2205 7154 2257
rect 7206 2205 7220 2257
rect 7140 2191 7220 2205
rect 6760 2144 6783 2178
rect 6817 2144 6840 2178
rect 6760 2098 6840 2144
rect 6760 2064 6783 2098
rect 6817 2064 6840 2098
rect 6990 2137 7070 2151
rect 6990 2085 7004 2137
rect 7056 2085 7070 2137
rect 6990 2071 7070 2085
rect 6760 2041 6840 2064
rect 6510 1981 6590 2001
rect 6910 1981 6990 2001
rect 6510 1978 6990 1981
rect 6510 1944 6533 1978
rect 6567 1944 6933 1978
rect 6967 1944 6990 1978
rect 6510 1941 6990 1944
rect 6510 1921 6590 1941
rect 6910 1921 6990 1941
rect 7260 1731 7300 2411
rect 7340 1987 7420 2001
rect 7340 1935 7354 1987
rect 7406 1935 7420 1987
rect 7340 1921 7420 1935
rect 3401 1489 3620 1529
rect 3660 1698 3740 1731
rect 3660 1664 3683 1698
rect 3717 1664 3740 1698
rect 3660 1618 3740 1664
rect 3660 1584 3683 1618
rect 3717 1584 3740 1618
rect 3660 1538 3740 1584
rect 3660 1504 3683 1538
rect 3717 1504 3740 1538
rect 3401 1484 3415 1489
rect 1129 1427 1209 1441
rect 1129 1375 1143 1427
rect 1195 1375 1209 1427
rect 1129 1361 1209 1375
rect 1840 1331 1880 1481
rect 2140 1331 2180 1481
rect 2440 1331 2480 1481
rect 3335 1469 3415 1484
rect 3660 1481 3740 1504
rect 4140 1698 4220 1731
rect 4140 1664 4163 1698
rect 4197 1664 4220 1698
rect 4140 1618 4220 1664
rect 4140 1584 4163 1618
rect 4197 1584 4220 1618
rect 4140 1538 4220 1584
rect 4140 1504 4163 1538
rect 4197 1504 4220 1538
rect 4140 1481 4220 1504
rect 4440 1698 4520 1731
rect 4440 1664 4463 1698
rect 4497 1664 4520 1698
rect 4440 1618 4520 1664
rect 4440 1584 4463 1618
rect 4497 1584 4520 1618
rect 4440 1538 4520 1584
rect 4440 1504 4463 1538
rect 4497 1504 4520 1538
rect 4440 1481 4520 1504
rect 4740 1698 4820 1731
rect 4740 1664 4763 1698
rect 4797 1664 4820 1698
rect 4740 1618 4820 1664
rect 4740 1584 4763 1618
rect 4797 1584 4820 1618
rect 4740 1538 4820 1584
rect 4740 1504 4763 1538
rect 4797 1504 4820 1538
rect 4740 1481 4820 1504
rect 5070 1698 5150 1731
rect 5070 1664 5093 1698
rect 5127 1664 5150 1698
rect 5070 1618 5150 1664
rect 5070 1584 5093 1618
rect 5127 1584 5150 1618
rect 5070 1538 5150 1584
rect 5830 1698 5910 1731
rect 5830 1664 5853 1698
rect 5887 1664 5910 1698
rect 5830 1618 5910 1664
rect 5830 1584 5853 1618
rect 5887 1584 5910 1618
rect 5070 1504 5093 1538
rect 5127 1504 5150 1538
rect 5070 1481 5150 1504
rect 5328 1547 5408 1561
rect 5328 1495 5342 1547
rect 5394 1541 5408 1547
rect 5830 1541 5910 1584
rect 5394 1538 5910 1541
rect 5394 1504 5853 1538
rect 5887 1504 5910 1538
rect 5394 1501 5910 1504
rect 5394 1495 5408 1501
rect 5328 1481 5408 1495
rect 5830 1481 5910 1501
rect 6160 1698 6240 1731
rect 6160 1664 6183 1698
rect 6217 1664 6240 1698
rect 6160 1618 6240 1664
rect 6160 1584 6183 1618
rect 6217 1584 6240 1618
rect 6160 1538 6240 1584
rect 6160 1504 6183 1538
rect 6217 1504 6240 1538
rect 6160 1481 6240 1504
rect 6460 1698 6540 1731
rect 6460 1664 6483 1698
rect 6517 1664 6540 1698
rect 6460 1618 6540 1664
rect 6460 1584 6483 1618
rect 6517 1584 6540 1618
rect 6460 1538 6540 1584
rect 6460 1504 6483 1538
rect 6517 1504 6540 1538
rect 6460 1481 6540 1504
rect 6760 1698 6840 1731
rect 6760 1664 6783 1698
rect 6817 1664 6840 1698
rect 6760 1618 6840 1664
rect 6760 1584 6783 1618
rect 6817 1584 6840 1618
rect 6760 1538 6840 1584
rect 6760 1504 6783 1538
rect 6817 1504 6840 1538
rect 6760 1481 6840 1504
rect 7240 1698 7320 1731
rect 7240 1664 7263 1698
rect 7297 1664 7320 1698
rect 7240 1618 7320 1664
rect 7240 1584 7263 1618
rect 7297 1584 7320 1618
rect 7240 1538 7320 1584
rect 7240 1504 7263 1538
rect 7297 1504 7320 1538
rect 7240 1481 7320 1504
rect 4160 1331 4200 1481
rect 4460 1331 4500 1481
rect 4760 1331 4800 1481
rect 5742 1427 5822 1441
rect 5742 1375 5756 1427
rect 5808 1375 5822 1427
rect 5742 1361 5822 1375
rect 6180 1331 6220 1481
rect 6480 1331 6520 1481
rect 6780 1331 6820 1481
rect 912 1264 935 1298
rect 969 1264 992 1298
rect 912 -1522 992 1264
rect 1020 1298 7340 1331
rect 1020 1264 1103 1298
rect 1137 1264 1183 1298
rect 1217 1264 1263 1298
rect 1297 1264 1343 1298
rect 1377 1264 1423 1298
rect 1457 1264 1503 1298
rect 1537 1264 1583 1298
rect 1617 1264 1663 1298
rect 1697 1264 1743 1298
rect 1777 1264 1823 1298
rect 1857 1264 1903 1298
rect 1937 1264 1983 1298
rect 2017 1264 2063 1298
rect 2097 1264 2143 1298
rect 2177 1264 2223 1298
rect 2257 1264 2303 1298
rect 2337 1264 2383 1298
rect 2417 1264 2463 1298
rect 2497 1264 2543 1298
rect 2577 1264 2623 1298
rect 2657 1264 2703 1298
rect 2737 1264 2783 1298
rect 2817 1264 2863 1298
rect 2897 1264 2943 1298
rect 2977 1264 3023 1298
rect 3057 1264 3103 1298
rect 3137 1264 3183 1298
rect 3217 1264 3663 1298
rect 3697 1264 3743 1298
rect 3777 1264 3823 1298
rect 3857 1264 3903 1298
rect 3937 1264 3983 1298
rect 4017 1264 4063 1298
rect 4097 1264 4143 1298
rect 4177 1264 4223 1298
rect 4257 1264 4303 1298
rect 4337 1264 4383 1298
rect 4417 1264 4463 1298
rect 4497 1264 4543 1298
rect 4577 1264 4623 1298
rect 4657 1264 4703 1298
rect 4737 1264 4783 1298
rect 4817 1264 4863 1298
rect 4897 1264 4943 1298
rect 4977 1264 5023 1298
rect 5057 1264 5103 1298
rect 5137 1264 5183 1298
rect 5217 1264 5263 1298
rect 5297 1264 5683 1298
rect 5717 1264 5763 1298
rect 5797 1264 5843 1298
rect 5877 1264 5923 1298
rect 5957 1264 6003 1298
rect 6037 1264 6083 1298
rect 6117 1264 6163 1298
rect 6197 1264 6243 1298
rect 6277 1264 6323 1298
rect 6357 1264 6403 1298
rect 6437 1264 6483 1298
rect 6517 1264 6563 1298
rect 6597 1264 6643 1298
rect 6677 1264 6723 1298
rect 6757 1264 6803 1298
rect 6837 1264 6883 1298
rect 6917 1264 6963 1298
rect 6997 1264 7043 1298
rect 7077 1264 7123 1298
rect 7157 1264 7203 1298
rect 7237 1264 7283 1298
rect 7317 1264 7340 1298
rect 1020 1231 7340 1264
rect 1128 1187 1208 1201
rect 1128 1135 1142 1187
rect 1194 1135 1208 1187
rect 1128 1121 1208 1135
rect 1840 1081 1880 1231
rect 2140 1081 2180 1231
rect 2440 1081 2480 1231
rect 4160 1081 4200 1231
rect 4460 1081 4500 1231
rect 4760 1081 4800 1231
rect 5073 1188 5153 1202
rect 5073 1136 5087 1188
rect 5139 1136 5153 1188
rect 5922 1187 6002 1201
rect 5922 1181 5936 1187
rect 5073 1122 5153 1136
rect 5487 1141 5936 1181
rect 1490 1058 1570 1081
rect 1490 1024 1513 1058
rect 1547 1024 1570 1058
rect 1490 978 1570 1024
rect 1490 944 1513 978
rect 1547 944 1570 978
rect 1490 898 1570 944
rect 1490 864 1513 898
rect 1547 864 1570 898
rect 1490 831 1570 864
rect 1820 1058 1900 1081
rect 1820 1024 1843 1058
rect 1877 1024 1900 1058
rect 1820 978 1900 1024
rect 1820 944 1843 978
rect 1877 944 1900 978
rect 1820 898 1900 944
rect 1820 864 1843 898
rect 1877 864 1900 898
rect 1820 831 1900 864
rect 2120 1058 2200 1081
rect 2120 1024 2143 1058
rect 2177 1024 2200 1058
rect 2120 978 2200 1024
rect 2120 944 2143 978
rect 2177 944 2200 978
rect 2120 898 2200 944
rect 2120 864 2143 898
rect 2177 864 2200 898
rect 2120 831 2200 864
rect 2420 1058 2500 1081
rect 2420 1024 2443 1058
rect 2477 1024 2500 1058
rect 2420 978 2500 1024
rect 2420 944 2443 978
rect 2477 944 2500 978
rect 2420 898 2500 944
rect 2420 864 2443 898
rect 2477 864 2500 898
rect 2420 831 2500 864
rect 2900 1058 2980 1081
rect 2900 1024 2923 1058
rect 2957 1024 2980 1058
rect 2900 978 2980 1024
rect 2900 944 2923 978
rect 2957 944 2980 978
rect 2900 898 2980 944
rect 2900 864 2923 898
rect 2957 864 2980 898
rect 2900 831 2980 864
rect 3810 1058 3890 1081
rect 3810 1024 3833 1058
rect 3867 1024 3890 1058
rect 3810 978 3890 1024
rect 3810 944 3833 978
rect 3867 944 3890 978
rect 3810 898 3890 944
rect 3810 864 3833 898
rect 3867 864 3890 898
rect 3810 831 3890 864
rect 4140 1058 4220 1081
rect 4140 1024 4163 1058
rect 4197 1024 4220 1058
rect 4140 978 4220 1024
rect 4140 944 4163 978
rect 4197 944 4220 978
rect 4140 898 4220 944
rect 4140 864 4163 898
rect 4197 864 4220 898
rect 4140 831 4220 864
rect 4440 1058 4520 1081
rect 4440 1024 4463 1058
rect 4497 1024 4520 1058
rect 4440 978 4520 1024
rect 4440 944 4463 978
rect 4497 944 4520 978
rect 4440 898 4520 944
rect 4440 864 4463 898
rect 4497 864 4520 898
rect 4440 831 4520 864
rect 4740 1058 4820 1081
rect 4740 1024 4763 1058
rect 4797 1024 4820 1058
rect 4740 978 4820 1024
rect 4740 944 4763 978
rect 4797 944 4820 978
rect 4740 898 4820 944
rect 4740 864 4763 898
rect 4797 864 4820 898
rect 4740 831 4820 864
rect 5220 1067 5408 1081
rect 5220 1058 5342 1067
rect 5220 1024 5243 1058
rect 5277 1024 5342 1058
rect 5220 1015 5342 1024
rect 5394 1015 5408 1067
rect 5220 1001 5408 1015
rect 5220 978 5300 1001
rect 5220 944 5243 978
rect 5277 944 5300 978
rect 5487 973 5527 1141
rect 5922 1135 5936 1141
rect 5988 1135 6002 1187
rect 5922 1121 6002 1135
rect 6180 1081 6220 1231
rect 6480 1081 6520 1231
rect 6780 1081 6820 1231
rect 5220 898 5300 944
rect 5220 864 5243 898
rect 5277 864 5300 898
rect 5220 831 5300 864
rect 5402 933 5527 973
rect 5830 1058 5910 1081
rect 5830 1024 5853 1058
rect 5887 1024 5910 1058
rect 5830 978 5910 1024
rect 5830 944 5853 978
rect 5887 944 5910 978
rect 1510 151 1550 831
rect 2170 621 2250 641
rect 2570 621 2650 641
rect 2170 618 2650 621
rect 2170 584 2193 618
rect 2227 584 2593 618
rect 2627 584 2650 618
rect 2170 581 2650 584
rect 2170 561 2250 581
rect 2570 561 2650 581
rect 1820 498 1900 521
rect 1670 477 1750 491
rect 1670 425 1684 477
rect 1736 425 1750 477
rect 1670 411 1750 425
rect 1820 464 1843 498
rect 1877 464 1900 498
rect 1820 418 1900 464
rect 1820 384 1843 418
rect 1877 384 1900 418
rect 1670 357 1750 371
rect 1670 305 1684 357
rect 1736 305 1750 357
rect 1670 291 1750 305
rect 1820 338 1900 384
rect 1820 304 1843 338
rect 1877 304 1900 338
rect 1820 151 1900 304
rect 2120 498 2200 521
rect 2120 464 2143 498
rect 2177 464 2200 498
rect 2120 418 2200 464
rect 2120 384 2143 418
rect 2177 384 2200 418
rect 2120 338 2200 384
rect 2120 304 2143 338
rect 2177 304 2200 338
rect 2120 151 2200 304
rect 2420 498 2500 521
rect 2420 464 2443 498
rect 2477 464 2500 498
rect 2420 418 2500 464
rect 2420 384 2443 418
rect 2477 384 2500 418
rect 2650 477 2730 491
rect 2650 425 2664 477
rect 2716 425 2730 477
rect 2650 411 2730 425
rect 2420 338 2500 384
rect 2420 304 2443 338
rect 2477 304 2500 338
rect 2420 151 2500 304
rect 2800 357 2880 371
rect 2800 305 2814 357
rect 2866 305 2880 357
rect 2800 291 2880 305
rect 2920 151 2960 831
rect 3000 738 3080 761
rect 3000 704 3023 738
rect 3057 704 3080 738
rect 3000 681 3080 704
rect 3020 511 3060 681
rect 3560 577 3640 591
rect 3560 525 3574 577
rect 3626 525 3640 577
rect 3560 511 3640 525
rect 3000 488 3080 511
rect 3000 454 3023 488
rect 3057 454 3080 488
rect 3000 431 3080 454
rect 3054 357 3134 371
rect 3054 305 3068 357
rect 3120 305 3134 357
rect 3054 291 3134 305
rect 3830 151 3870 831
rect 4490 621 4570 641
rect 4890 621 4970 641
rect 4490 618 4970 621
rect 4490 584 4513 618
rect 4547 584 4913 618
rect 4947 584 4970 618
rect 4490 581 4970 584
rect 4490 561 4570 581
rect 4890 561 4970 581
rect 4140 498 4220 521
rect 3990 477 4070 491
rect 3990 425 4004 477
rect 4056 425 4070 477
rect 3990 411 4070 425
rect 4140 464 4163 498
rect 4197 464 4220 498
rect 4140 418 4220 464
rect 4140 384 4163 418
rect 4197 384 4220 418
rect 3990 357 4070 371
rect 3990 305 4004 357
rect 4056 305 4070 357
rect 3990 291 4070 305
rect 4140 338 4220 384
rect 4140 304 4163 338
rect 4197 304 4220 338
rect 4140 151 4220 304
rect 4440 498 4520 521
rect 4440 464 4463 498
rect 4497 464 4520 498
rect 4440 418 4520 464
rect 4440 384 4463 418
rect 4497 384 4520 418
rect 4440 338 4520 384
rect 4440 304 4463 338
rect 4497 304 4520 338
rect 4440 151 4520 304
rect 4740 498 4820 521
rect 4740 464 4763 498
rect 4797 464 4820 498
rect 4740 418 4820 464
rect 4740 384 4763 418
rect 4797 384 4820 418
rect 4970 477 5050 491
rect 4970 425 4984 477
rect 5036 425 5050 477
rect 4970 411 5050 425
rect 4740 338 4820 384
rect 4740 304 4763 338
rect 4797 304 4820 338
rect 4740 151 4820 304
rect 5120 357 5200 371
rect 5120 305 5134 357
rect 5186 305 5200 357
rect 5120 291 5200 305
rect 5240 151 5280 831
rect 1020 127 3000 151
rect 1020 75 1034 127
rect 1086 118 3000 127
rect 1086 84 1343 118
rect 1377 84 1423 118
rect 1457 84 1503 118
rect 1537 84 1583 118
rect 1617 84 1663 118
rect 1697 84 1743 118
rect 1777 84 1823 118
rect 1857 84 1903 118
rect 1937 84 1983 118
rect 2017 84 2063 118
rect 2097 84 2143 118
rect 2177 84 2223 118
rect 2257 84 2303 118
rect 2337 84 2383 118
rect 2417 84 2463 118
rect 2497 84 2543 118
rect 2577 84 2623 118
rect 2657 84 2703 118
rect 2737 84 2783 118
rect 2817 84 2863 118
rect 2897 84 2943 118
rect 2977 84 3000 118
rect 1086 75 3000 84
rect 1020 51 3000 75
rect 3640 118 5320 151
rect 3640 84 3663 118
rect 3697 84 3743 118
rect 3777 84 3823 118
rect 3857 84 3903 118
rect 3937 84 3983 118
rect 4017 84 4063 118
rect 4097 84 4143 118
rect 4177 84 4223 118
rect 4257 84 4303 118
rect 4337 84 4383 118
rect 4417 84 4463 118
rect 4497 84 4543 118
rect 4577 84 4623 118
rect 4657 84 4703 118
rect 4737 84 4783 118
rect 4817 84 4863 118
rect 4897 84 4943 118
rect 4977 84 5023 118
rect 5057 84 5103 118
rect 5137 84 5183 118
rect 5217 84 5263 118
rect 5297 84 5320 118
rect 3640 51 5320 84
rect 5136 -193 5216 -179
rect 5136 -245 5150 -193
rect 5202 -198 5216 -193
rect 5402 -198 5442 933
rect 5555 897 5635 911
rect 5555 891 5569 897
rect 5487 851 5569 891
rect 5487 641 5527 851
rect 5555 845 5569 851
rect 5621 845 5635 897
rect 5555 831 5635 845
rect 5830 898 5910 944
rect 5830 864 5853 898
rect 5887 864 5910 898
rect 5830 831 5910 864
rect 6160 1058 6240 1081
rect 6160 1024 6183 1058
rect 6217 1024 6240 1058
rect 6160 978 6240 1024
rect 6160 944 6183 978
rect 6217 944 6240 978
rect 6160 898 6240 944
rect 6160 864 6183 898
rect 6217 864 6240 898
rect 6160 831 6240 864
rect 6460 1058 6540 1081
rect 6460 1024 6483 1058
rect 6517 1024 6540 1058
rect 6460 978 6540 1024
rect 6460 944 6483 978
rect 6517 944 6540 978
rect 6460 898 6540 944
rect 6460 864 6483 898
rect 6517 864 6540 898
rect 6460 831 6540 864
rect 6760 1058 6840 1081
rect 6760 1024 6783 1058
rect 6817 1024 6840 1058
rect 6760 978 6840 1024
rect 6760 944 6783 978
rect 6817 944 6840 978
rect 6760 898 6840 944
rect 7240 1058 7320 1081
rect 7240 1024 7263 1058
rect 7297 1024 7320 1058
rect 7240 978 7320 1024
rect 7240 944 7263 978
rect 7297 944 7320 978
rect 6760 864 6783 898
rect 6817 864 6840 898
rect 6760 831 6840 864
rect 7090 897 7170 911
rect 7090 845 7104 897
rect 7156 845 7170 897
rect 7090 831 7170 845
rect 7240 898 7320 944
rect 7240 864 7263 898
rect 7297 864 7320 898
rect 7240 831 7320 864
rect 7348 897 7428 911
rect 7348 845 7362 897
rect 7414 845 7428 897
rect 7348 831 7428 845
rect 5660 747 5740 761
rect 5660 695 5674 747
rect 5726 695 5740 747
rect 5660 681 5740 695
rect 5471 618 5551 641
rect 5471 584 5494 618
rect 5528 584 5551 618
rect 5471 561 5551 584
rect 5660 627 5740 641
rect 5660 575 5674 627
rect 5726 575 5740 627
rect 5660 561 5740 575
rect 5730 387 5810 401
rect 5730 335 5744 387
rect 5796 335 5810 387
rect 5730 321 5810 335
rect 5850 151 5890 831
rect 6010 621 6090 641
rect 6410 621 6490 641
rect 6010 618 6490 621
rect 6010 584 6033 618
rect 6067 584 6433 618
rect 6467 584 6490 618
rect 6010 581 6490 584
rect 6010 561 6090 581
rect 6410 561 6490 581
rect 5930 507 6010 521
rect 5930 455 5944 507
rect 5996 455 6010 507
rect 5930 441 6010 455
rect 6160 498 6240 521
rect 6160 464 6183 498
rect 6217 464 6240 498
rect 6160 418 6240 464
rect 6160 384 6183 418
rect 6217 384 6240 418
rect 6160 338 6240 384
rect 6160 304 6183 338
rect 6217 304 6240 338
rect 6160 151 6240 304
rect 6460 498 6540 521
rect 6460 464 6483 498
rect 6517 464 6540 498
rect 6460 418 6540 464
rect 6460 384 6483 418
rect 6517 384 6540 418
rect 6460 338 6540 384
rect 6460 304 6483 338
rect 6517 304 6540 338
rect 6460 151 6540 304
rect 6760 498 6840 521
rect 6760 464 6783 498
rect 6817 464 6840 498
rect 6760 418 6840 464
rect 6910 507 6990 521
rect 6910 455 6924 507
rect 6976 455 6990 507
rect 6910 441 6990 455
rect 6760 384 6783 418
rect 6817 384 6840 418
rect 6760 338 6840 384
rect 6760 304 6783 338
rect 6817 304 6840 338
rect 6910 387 6990 401
rect 6910 335 6924 387
rect 6976 335 6990 387
rect 6910 321 6990 335
rect 6760 151 6840 304
rect 7260 151 7300 831
rect 7354 722 7394 831
rect 7334 699 7414 722
rect 7334 665 7357 699
rect 7391 665 7414 699
rect 7334 642 7414 665
rect 5478 127 7340 151
rect 5478 75 5492 127
rect 5544 118 5754 127
rect 5806 118 7340 127
rect 5544 84 5683 118
rect 5717 84 5754 118
rect 5806 84 5843 118
rect 5877 84 5923 118
rect 5957 84 6003 118
rect 6037 84 6083 118
rect 6117 84 6163 118
rect 6197 84 6243 118
rect 6277 84 6323 118
rect 6357 84 6403 118
rect 6437 84 6483 118
rect 6517 84 6563 118
rect 6597 84 6643 118
rect 6677 84 6723 118
rect 6757 84 6803 118
rect 6837 84 6883 118
rect 6917 84 6963 118
rect 6997 84 7043 118
rect 7077 84 7123 118
rect 7157 84 7203 118
rect 7237 84 7283 118
rect 7317 84 7340 118
rect 5544 75 5754 84
rect 5806 75 7340 84
rect 5478 51 7340 75
rect 5202 -238 5442 -198
rect 5202 -245 5216 -238
rect 5136 -259 5216 -245
rect 1020 -333 5040 -309
rect 1020 -385 1070 -333
rect 1122 -342 5040 -333
rect 1137 -376 1183 -342
rect 1217 -376 1263 -342
rect 1297 -376 1343 -342
rect 1377 -376 1423 -342
rect 1457 -376 1503 -342
rect 1537 -376 1583 -342
rect 1617 -376 1663 -342
rect 1697 -376 1743 -342
rect 1777 -376 1823 -342
rect 1857 -376 1903 -342
rect 1937 -376 1983 -342
rect 2017 -376 2063 -342
rect 2097 -376 2143 -342
rect 2177 -376 2223 -342
rect 2257 -376 2303 -342
rect 2337 -376 2383 -342
rect 2417 -376 2463 -342
rect 2497 -376 2543 -342
rect 2577 -376 2623 -342
rect 2657 -376 2703 -342
rect 2737 -376 2783 -342
rect 2817 -376 2863 -342
rect 2897 -376 2943 -342
rect 2977 -376 3023 -342
rect 3057 -376 3103 -342
rect 3137 -376 3183 -342
rect 3217 -376 3693 -342
rect 3727 -376 3773 -342
rect 3807 -376 3853 -342
rect 3887 -376 3933 -342
rect 3967 -376 4013 -342
rect 4047 -376 4093 -342
rect 4127 -376 4173 -342
rect 4207 -376 4253 -342
rect 4287 -376 4333 -342
rect 4367 -376 4413 -342
rect 4447 -376 4493 -342
rect 4527 -376 4573 -342
rect 4607 -376 4653 -342
rect 4687 -376 4733 -342
rect 4767 -376 4813 -342
rect 4847 -376 4893 -342
rect 4927 -376 4973 -342
rect 5007 -376 5040 -342
rect 1122 -385 5040 -376
rect 1020 -409 5040 -385
rect 5390 -333 7070 -309
rect 5390 -342 7004 -333
rect 5390 -376 5413 -342
rect 5447 -376 5493 -342
rect 5527 -376 5573 -342
rect 5607 -376 5653 -342
rect 5687 -376 5733 -342
rect 5767 -376 5813 -342
rect 5847 -376 5893 -342
rect 5927 -376 5973 -342
rect 6007 -376 6053 -342
rect 6087 -376 6133 -342
rect 6167 -376 6213 -342
rect 6247 -376 6293 -342
rect 6327 -376 6373 -342
rect 6407 -376 6453 -342
rect 6487 -376 6533 -342
rect 6567 -376 6613 -342
rect 6647 -376 6693 -342
rect 6727 -376 6773 -342
rect 6807 -376 6853 -342
rect 6887 -376 6933 -342
rect 6967 -376 7004 -342
rect 5390 -385 7004 -376
rect 7056 -385 7070 -333
rect 5390 -409 7070 -385
rect 1360 -1089 1400 -409
rect 1540 -463 1620 -449
rect 1540 -515 1554 -463
rect 1606 -515 1620 -463
rect 1540 -529 1620 -515
rect 1670 -563 1750 -549
rect 1670 -615 1684 -563
rect 1736 -615 1750 -563
rect 1670 -629 1750 -615
rect 1820 -562 1900 -409
rect 1820 -596 1843 -562
rect 1877 -596 1900 -562
rect 1820 -642 1900 -596
rect 1540 -663 1620 -649
rect 1540 -715 1554 -663
rect 1606 -715 1620 -663
rect 1540 -729 1620 -715
rect 1820 -676 1843 -642
rect 1877 -676 1900 -642
rect 1820 -722 1900 -676
rect 1670 -763 1750 -749
rect 1670 -815 1684 -763
rect 1736 -815 1750 -763
rect 1820 -756 1843 -722
rect 1877 -756 1900 -722
rect 1820 -779 1900 -756
rect 2120 -562 2200 -409
rect 2120 -596 2143 -562
rect 2177 -596 2200 -562
rect 2120 -642 2200 -596
rect 2120 -676 2143 -642
rect 2177 -676 2200 -642
rect 2120 -722 2200 -676
rect 2120 -756 2143 -722
rect 2177 -756 2200 -722
rect 2120 -779 2200 -756
rect 2420 -562 2500 -409
rect 2800 -463 2880 -449
rect 2800 -515 2814 -463
rect 2866 -515 2880 -463
rect 2800 -529 2880 -515
rect 2420 -596 2443 -562
rect 2477 -596 2500 -562
rect 2420 -642 2500 -596
rect 2420 -676 2443 -642
rect 2477 -676 2500 -642
rect 2420 -722 2500 -676
rect 2420 -756 2443 -722
rect 2477 -756 2500 -722
rect 2420 -779 2500 -756
rect 2700 -763 2780 -749
rect 1670 -829 1750 -815
rect 2700 -815 2714 -763
rect 2766 -815 2780 -763
rect 2170 -842 2250 -819
rect 2700 -829 2780 -815
rect 2170 -876 2193 -842
rect 2227 -859 2250 -842
rect 2540 -852 2620 -829
rect 2540 -859 2563 -852
rect 2227 -876 2563 -859
rect 2170 -886 2563 -876
rect 2597 -886 2620 -852
rect 2170 -899 2620 -886
rect 2540 -909 2620 -899
rect 2920 -1089 2960 -409
rect 3572 -529 3652 -515
rect 3000 -563 3080 -549
rect 3000 -615 3014 -563
rect 3066 -615 3080 -563
rect 3572 -581 3586 -529
rect 3638 -581 3652 -529
rect 3572 -595 3652 -581
rect 3000 -629 3080 -615
rect 3572 -640 3652 -626
rect 3150 -663 3230 -649
rect 3150 -715 3164 -663
rect 3216 -715 3230 -663
rect 3572 -692 3586 -640
rect 3638 -692 3652 -640
rect 3572 -706 3652 -692
rect 3150 -729 3230 -715
rect 3300 -964 3380 -943
rect 3591 -964 3631 -706
rect 3300 -966 3631 -964
rect 3300 -1000 3323 -966
rect 3357 -1000 3631 -966
rect 3300 -1004 3631 -1000
rect 3300 -1023 3380 -1004
rect 1340 -1122 1420 -1089
rect 1340 -1156 1363 -1122
rect 1397 -1156 1420 -1122
rect 1340 -1202 1420 -1156
rect 1340 -1236 1363 -1202
rect 1397 -1236 1420 -1202
rect 1340 -1282 1420 -1236
rect 1340 -1316 1363 -1282
rect 1397 -1316 1420 -1282
rect 1340 -1339 1420 -1316
rect 1820 -1122 1900 -1089
rect 1820 -1156 1843 -1122
rect 1877 -1156 1900 -1122
rect 1820 -1202 1900 -1156
rect 1820 -1236 1843 -1202
rect 1877 -1236 1900 -1202
rect 1820 -1282 1900 -1236
rect 1820 -1316 1843 -1282
rect 1877 -1316 1900 -1282
rect 1820 -1339 1900 -1316
rect 2120 -1122 2200 -1089
rect 2120 -1156 2143 -1122
rect 2177 -1156 2200 -1122
rect 2120 -1202 2200 -1156
rect 2120 -1236 2143 -1202
rect 2177 -1236 2200 -1202
rect 2120 -1282 2200 -1236
rect 2120 -1316 2143 -1282
rect 2177 -1316 2200 -1282
rect 2120 -1339 2200 -1316
rect 2420 -1122 2500 -1089
rect 2420 -1156 2443 -1122
rect 2477 -1156 2500 -1122
rect 2420 -1202 2500 -1156
rect 2420 -1236 2443 -1202
rect 2477 -1236 2500 -1202
rect 2420 -1282 2500 -1236
rect 2420 -1316 2443 -1282
rect 2477 -1316 2500 -1282
rect 2420 -1339 2500 -1316
rect 2900 -1122 2980 -1089
rect 2900 -1156 2923 -1122
rect 2957 -1156 2980 -1122
rect 3680 -1122 3760 -409
rect 3860 -460 3940 -447
rect 3860 -512 3874 -460
rect 3926 -512 3940 -460
rect 3860 -527 3940 -512
rect 3880 -699 3920 -527
rect 4010 -562 4090 -409
rect 4010 -596 4033 -562
rect 4067 -596 4090 -562
rect 4010 -642 4090 -596
rect 4010 -676 4033 -642
rect 4067 -676 4090 -642
rect 3860 -713 3940 -699
rect 3860 -765 3874 -713
rect 3926 -765 3940 -713
rect 3860 -779 3940 -765
rect 4010 -722 4090 -676
rect 4010 -756 4033 -722
rect 4067 -756 4090 -722
rect 4010 -779 4090 -756
rect 4310 -562 4390 -409
rect 4310 -596 4333 -562
rect 4367 -596 4390 -562
rect 4310 -642 4390 -596
rect 4310 -676 4333 -642
rect 4367 -676 4390 -642
rect 4310 -722 4390 -676
rect 4310 -756 4333 -722
rect 4367 -756 4390 -722
rect 4310 -779 4390 -756
rect 4610 -562 4690 -409
rect 4610 -596 4633 -562
rect 4667 -596 4690 -562
rect 4610 -642 4690 -596
rect 4610 -676 4633 -642
rect 4667 -676 4690 -642
rect 4610 -722 4690 -676
rect 4610 -756 4633 -722
rect 4667 -756 4690 -722
rect 4610 -779 4690 -756
rect 4760 -713 4840 -699
rect 4760 -765 4774 -713
rect 4826 -765 4840 -713
rect 4760 -779 4840 -765
rect 4360 -839 4440 -819
rect 4760 -839 4840 -819
rect 4360 -842 4840 -839
rect 4360 -876 4383 -842
rect 4417 -876 4783 -842
rect 4817 -876 4840 -842
rect 4360 -879 4840 -876
rect 4360 -899 4440 -879
rect 4760 -899 4840 -879
rect 2900 -1202 2980 -1156
rect 2900 -1236 2923 -1202
rect 2957 -1236 2980 -1202
rect 3314 -1161 3394 -1148
rect 3314 -1213 3328 -1161
rect 3380 -1213 3394 -1161
rect 3314 -1228 3394 -1213
rect 3680 -1156 3703 -1122
rect 3737 -1156 3760 -1122
rect 3680 -1202 3760 -1156
rect 2900 -1282 2980 -1236
rect 2900 -1316 2923 -1282
rect 2957 -1316 2980 -1282
rect 2900 -1339 2980 -1316
rect 3680 -1236 3703 -1202
rect 3737 -1236 3760 -1202
rect 3680 -1282 3760 -1236
rect 3680 -1316 3703 -1282
rect 3737 -1316 3760 -1282
rect 3680 -1339 3760 -1316
rect 4010 -1122 4090 -1089
rect 4010 -1156 4033 -1122
rect 4067 -1156 4090 -1122
rect 4010 -1202 4090 -1156
rect 4010 -1236 4033 -1202
rect 4067 -1236 4090 -1202
rect 4010 -1282 4090 -1236
rect 4010 -1316 4033 -1282
rect 4067 -1316 4090 -1282
rect 4010 -1339 4090 -1316
rect 4310 -1122 4390 -1089
rect 4310 -1156 4333 -1122
rect 4367 -1156 4390 -1122
rect 4310 -1202 4390 -1156
rect 4310 -1236 4333 -1202
rect 4367 -1236 4390 -1202
rect 4310 -1282 4390 -1236
rect 4310 -1316 4333 -1282
rect 4367 -1316 4390 -1282
rect 4310 -1339 4390 -1316
rect 4610 -1122 4690 -1089
rect 4610 -1156 4633 -1122
rect 4667 -1156 4690 -1122
rect 4610 -1202 4690 -1156
rect 4610 -1236 4633 -1202
rect 4667 -1236 4690 -1202
rect 4610 -1282 4690 -1236
rect 4610 -1316 4633 -1282
rect 4667 -1316 4690 -1282
rect 4610 -1339 4690 -1316
rect 4940 -1122 5020 -409
rect 5251 -449 5331 -435
rect 5251 -501 5265 -449
rect 5317 -501 5331 -449
rect 5251 -515 5331 -501
rect 5472 -451 5552 -437
rect 5472 -503 5486 -451
rect 5538 -503 5552 -451
rect 5472 -517 5552 -503
rect 5048 -550 5128 -536
rect 5048 -602 5062 -550
rect 5114 -564 5128 -550
rect 5310 -564 5390 -549
rect 5114 -572 5390 -564
rect 5114 -602 5333 -572
rect 5048 -604 5333 -602
rect 5048 -616 5128 -604
rect 5310 -606 5333 -604
rect 5367 -606 5390 -572
rect 5310 -629 5390 -606
rect 5048 -659 5128 -645
rect 5048 -711 5062 -659
rect 5114 -665 5128 -659
rect 5114 -705 5370 -665
rect 5114 -711 5128 -705
rect 5048 -725 5128 -711
rect 5330 -769 5370 -705
rect 5310 -792 5390 -769
rect 5048 -848 5128 -825
rect 5048 -882 5071 -848
rect 5105 -882 5128 -848
rect 5310 -826 5333 -792
rect 5367 -826 5390 -792
rect 5310 -849 5390 -826
rect 5048 -905 5128 -882
rect 5310 -905 5390 -889
rect 5048 -912 5390 -905
rect 5048 -945 5333 -912
rect 5310 -946 5333 -945
rect 5367 -946 5390 -912
rect 5310 -969 5390 -946
rect 5580 -1089 5620 -409
rect 5740 -563 5820 -549
rect 5740 -615 5754 -563
rect 5806 -615 5820 -563
rect 5740 -629 5820 -615
rect 5890 -562 5970 -409
rect 5890 -596 5913 -562
rect 5947 -596 5970 -562
rect 5890 -642 5970 -596
rect 5740 -683 5820 -669
rect 5740 -735 5754 -683
rect 5806 -735 5820 -683
rect 5740 -749 5820 -735
rect 5890 -676 5913 -642
rect 5947 -676 5970 -642
rect 5890 -722 5970 -676
rect 5890 -756 5913 -722
rect 5947 -756 5970 -722
rect 5890 -779 5970 -756
rect 6190 -562 6270 -409
rect 6190 -596 6213 -562
rect 6247 -596 6270 -562
rect 6190 -642 6270 -596
rect 6190 -676 6213 -642
rect 6247 -676 6270 -642
rect 6190 -722 6270 -676
rect 6190 -756 6213 -722
rect 6247 -756 6270 -722
rect 6190 -779 6270 -756
rect 6490 -562 6570 -409
rect 6490 -596 6513 -562
rect 6547 -596 6570 -562
rect 6490 -642 6570 -596
rect 6870 -563 6950 -549
rect 6870 -615 6884 -563
rect 6936 -615 6950 -563
rect 6870 -629 6950 -615
rect 6490 -676 6513 -642
rect 6547 -676 6570 -642
rect 6490 -722 6570 -676
rect 6490 -756 6513 -722
rect 6547 -756 6570 -722
rect 6720 -683 6800 -669
rect 6720 -735 6734 -683
rect 6786 -735 6800 -683
rect 6720 -749 6800 -735
rect 6490 -779 6570 -756
rect 6240 -839 6320 -819
rect 6640 -839 6720 -819
rect 6240 -842 6720 -839
rect 6240 -876 6263 -842
rect 6297 -876 6663 -842
rect 6697 -876 6720 -842
rect 6240 -879 6720 -876
rect 6240 -899 6320 -879
rect 6640 -899 6720 -879
rect 6990 -1089 7030 -409
rect 7073 -953 7153 -939
rect 7073 -1005 7087 -953
rect 7139 -1005 7153 -953
rect 7073 -1019 7153 -1005
rect 4940 -1156 4963 -1122
rect 4997 -1156 5020 -1122
rect 4940 -1202 5020 -1156
rect 4940 -1236 4963 -1202
rect 4997 -1236 5020 -1202
rect 4940 -1282 5020 -1236
rect 4940 -1316 4963 -1282
rect 4997 -1316 5020 -1282
rect 4940 -1339 5020 -1316
rect 5560 -1122 5640 -1089
rect 5560 -1156 5583 -1122
rect 5617 -1156 5640 -1122
rect 5560 -1202 5640 -1156
rect 5560 -1236 5583 -1202
rect 5617 -1236 5640 -1202
rect 5560 -1282 5640 -1236
rect 5560 -1316 5583 -1282
rect 5617 -1316 5640 -1282
rect 5560 -1339 5640 -1316
rect 5890 -1122 5970 -1089
rect 5890 -1156 5913 -1122
rect 5947 -1156 5970 -1122
rect 5890 -1202 5970 -1156
rect 5890 -1236 5913 -1202
rect 5947 -1236 5970 -1202
rect 5890 -1282 5970 -1236
rect 5890 -1316 5913 -1282
rect 5947 -1316 5970 -1282
rect 5890 -1339 5970 -1316
rect 6190 -1122 6270 -1089
rect 6190 -1156 6213 -1122
rect 6247 -1156 6270 -1122
rect 6190 -1202 6270 -1156
rect 6190 -1236 6213 -1202
rect 6247 -1236 6270 -1202
rect 6190 -1282 6270 -1236
rect 6190 -1316 6213 -1282
rect 6247 -1316 6270 -1282
rect 6190 -1339 6270 -1316
rect 6490 -1122 6570 -1089
rect 6490 -1156 6513 -1122
rect 6547 -1156 6570 -1122
rect 6490 -1202 6570 -1156
rect 6490 -1236 6513 -1202
rect 6547 -1236 6570 -1202
rect 6490 -1282 6570 -1236
rect 6490 -1316 6513 -1282
rect 6547 -1316 6570 -1282
rect 6490 -1339 6570 -1316
rect 6970 -1122 7050 -1089
rect 6970 -1156 6993 -1122
rect 7027 -1156 7050 -1122
rect 6970 -1202 7050 -1156
rect 6970 -1236 6993 -1202
rect 7027 -1236 7050 -1202
rect 6970 -1273 7050 -1236
rect 6970 -1325 6984 -1273
rect 7036 -1325 7050 -1273
rect 6970 -1339 7050 -1325
rect 1171 -1393 1251 -1379
rect 1171 -1445 1185 -1393
rect 1237 -1445 1251 -1393
rect 1171 -1459 1251 -1445
rect 1840 -1489 1880 -1339
rect 2140 -1489 2180 -1339
rect 2440 -1489 2480 -1339
rect 4030 -1489 4070 -1339
rect 4330 -1489 4370 -1339
rect 4630 -1489 4670 -1339
rect 5398 -1393 5478 -1379
rect 5398 -1445 5412 -1393
rect 5464 -1445 5478 -1393
rect 5398 -1459 5478 -1445
rect 5910 -1489 5950 -1339
rect 6210 -1489 6250 -1339
rect 6510 -1489 6550 -1339
rect 912 -1556 935 -1522
rect 969 -1556 992 -1522
rect 912 -4342 992 -1556
rect 1020 -1522 7070 -1489
rect 1020 -1556 1103 -1522
rect 1137 -1556 1183 -1522
rect 1217 -1556 1263 -1522
rect 1297 -1556 1343 -1522
rect 1377 -1556 1423 -1522
rect 1457 -1556 1503 -1522
rect 1537 -1556 1583 -1522
rect 1617 -1556 1663 -1522
rect 1697 -1556 1743 -1522
rect 1777 -1556 1823 -1522
rect 1857 -1556 1903 -1522
rect 1937 -1556 1983 -1522
rect 2017 -1556 2063 -1522
rect 2097 -1556 2143 -1522
rect 2177 -1556 2223 -1522
rect 2257 -1556 2303 -1522
rect 2337 -1556 2383 -1522
rect 2417 -1556 2463 -1522
rect 2497 -1556 2543 -1522
rect 2577 -1556 2623 -1522
rect 2657 -1556 2703 -1522
rect 2737 -1556 2783 -1522
rect 2817 -1556 2863 -1522
rect 2897 -1556 2943 -1522
rect 2977 -1556 3023 -1522
rect 3057 -1556 3103 -1522
rect 3137 -1556 3183 -1522
rect 3217 -1556 3693 -1522
rect 3727 -1556 3773 -1522
rect 3807 -1556 3853 -1522
rect 3887 -1556 3933 -1522
rect 3967 -1556 4013 -1522
rect 4047 -1556 4093 -1522
rect 4127 -1556 4173 -1522
rect 4207 -1556 4253 -1522
rect 4287 -1556 4333 -1522
rect 4367 -1556 4413 -1522
rect 4447 -1556 4493 -1522
rect 4527 -1556 4573 -1522
rect 4607 -1556 4653 -1522
rect 4687 -1556 4733 -1522
rect 4767 -1556 4813 -1522
rect 4847 -1556 4893 -1522
rect 4927 -1556 4973 -1522
rect 5007 -1556 5413 -1522
rect 5447 -1556 5493 -1522
rect 5527 -1556 5573 -1522
rect 5607 -1556 5653 -1522
rect 5687 -1556 5733 -1522
rect 5767 -1556 5813 -1522
rect 5847 -1556 5893 -1522
rect 5927 -1556 5973 -1522
rect 6007 -1556 6053 -1522
rect 6087 -1556 6133 -1522
rect 6167 -1556 6213 -1522
rect 6247 -1556 6293 -1522
rect 6327 -1556 6373 -1522
rect 6407 -1556 6453 -1522
rect 6487 -1556 6533 -1522
rect 6567 -1556 6613 -1522
rect 6647 -1556 6693 -1522
rect 6727 -1556 6773 -1522
rect 6807 -1556 6853 -1522
rect 6887 -1556 6933 -1522
rect 6967 -1556 7013 -1522
rect 7047 -1556 7070 -1522
rect 1020 -1589 7070 -1556
rect 1171 -1633 1251 -1619
rect 1171 -1685 1185 -1633
rect 1237 -1685 1251 -1633
rect 1171 -1699 1251 -1685
rect 1840 -1739 1880 -1589
rect 2140 -1739 2180 -1589
rect 2440 -1739 2480 -1589
rect 4030 -1739 4070 -1589
rect 4330 -1739 4370 -1589
rect 4630 -1739 4670 -1589
rect 5398 -1632 5478 -1618
rect 5398 -1684 5412 -1632
rect 5464 -1684 5478 -1632
rect 5398 -1698 5478 -1684
rect 5910 -1739 5950 -1589
rect 6210 -1739 6250 -1589
rect 6510 -1739 6550 -1589
rect 1340 -1762 1420 -1739
rect 1340 -1796 1363 -1762
rect 1397 -1796 1420 -1762
rect 1340 -1842 1420 -1796
rect 1340 -1876 1363 -1842
rect 1397 -1876 1420 -1842
rect 1340 -1922 1420 -1876
rect 1340 -1956 1363 -1922
rect 1397 -1956 1420 -1922
rect 1340 -1989 1420 -1956
rect 1820 -1762 1900 -1739
rect 1820 -1796 1843 -1762
rect 1877 -1796 1900 -1762
rect 1820 -1842 1900 -1796
rect 1820 -1876 1843 -1842
rect 1877 -1876 1900 -1842
rect 1820 -1922 1900 -1876
rect 1820 -1956 1843 -1922
rect 1877 -1956 1900 -1922
rect 1820 -1989 1900 -1956
rect 2120 -1762 2200 -1739
rect 2120 -1796 2143 -1762
rect 2177 -1796 2200 -1762
rect 2120 -1842 2200 -1796
rect 2120 -1876 2143 -1842
rect 2177 -1876 2200 -1842
rect 2120 -1922 2200 -1876
rect 2120 -1956 2143 -1922
rect 2177 -1956 2200 -1922
rect 2120 -1989 2200 -1956
rect 2420 -1762 2500 -1739
rect 2420 -1796 2443 -1762
rect 2477 -1796 2500 -1762
rect 2420 -1842 2500 -1796
rect 2420 -1876 2443 -1842
rect 2477 -1876 2500 -1842
rect 2420 -1922 2500 -1876
rect 2420 -1956 2443 -1922
rect 2477 -1956 2500 -1922
rect 2420 -1989 2500 -1956
rect 2900 -1762 2980 -1739
rect 2900 -1796 2923 -1762
rect 2957 -1796 2980 -1762
rect 2900 -1842 2980 -1796
rect 2900 -1876 2923 -1842
rect 2957 -1876 2980 -1842
rect 3680 -1762 3760 -1739
rect 3680 -1796 3703 -1762
rect 3737 -1796 3760 -1762
rect 3680 -1842 3760 -1796
rect 2900 -1922 2980 -1876
rect 2900 -1956 2923 -1922
rect 2957 -1956 2980 -1922
rect 3314 -1856 3394 -1843
rect 3314 -1908 3328 -1856
rect 3380 -1908 3394 -1856
rect 3314 -1923 3394 -1908
rect 3680 -1876 3703 -1842
rect 3737 -1876 3760 -1842
rect 3680 -1922 3760 -1876
rect 2900 -1989 2980 -1956
rect 3680 -1956 3703 -1922
rect 3737 -1956 3760 -1922
rect 1360 -2669 1400 -1989
rect 2540 -2179 2620 -2169
rect 2170 -2192 2620 -2179
rect 2170 -2202 2563 -2192
rect 2170 -2236 2193 -2202
rect 2227 -2219 2563 -2202
rect 2227 -2236 2250 -2219
rect 1670 -2263 1750 -2249
rect 2170 -2259 2250 -2236
rect 2540 -2226 2563 -2219
rect 2597 -2226 2620 -2192
rect 2540 -2249 2620 -2226
rect 1670 -2315 1684 -2263
rect 1736 -2315 1750 -2263
rect 2700 -2263 2780 -2249
rect 1670 -2329 1750 -2315
rect 1820 -2322 1900 -2299
rect 1540 -2363 1620 -2349
rect 1540 -2415 1554 -2363
rect 1606 -2415 1620 -2363
rect 1540 -2429 1620 -2415
rect 1820 -2356 1843 -2322
rect 1877 -2356 1900 -2322
rect 1820 -2402 1900 -2356
rect 1820 -2436 1843 -2402
rect 1877 -2436 1900 -2402
rect 1670 -2463 1750 -2449
rect 1670 -2515 1684 -2463
rect 1736 -2515 1750 -2463
rect 1670 -2529 1750 -2515
rect 1820 -2482 1900 -2436
rect 1820 -2516 1843 -2482
rect 1877 -2516 1900 -2482
rect 1540 -2563 1620 -2549
rect 1540 -2615 1554 -2563
rect 1606 -2615 1620 -2563
rect 1540 -2629 1620 -2615
rect 1820 -2669 1900 -2516
rect 2120 -2322 2200 -2299
rect 2120 -2356 2143 -2322
rect 2177 -2356 2200 -2322
rect 2120 -2402 2200 -2356
rect 2120 -2436 2143 -2402
rect 2177 -2436 2200 -2402
rect 2120 -2482 2200 -2436
rect 2120 -2516 2143 -2482
rect 2177 -2516 2200 -2482
rect 2120 -2669 2200 -2516
rect 2420 -2322 2500 -2299
rect 2420 -2356 2443 -2322
rect 2477 -2356 2500 -2322
rect 2700 -2315 2714 -2263
rect 2766 -2315 2780 -2263
rect 2700 -2329 2780 -2315
rect 2420 -2402 2500 -2356
rect 2420 -2436 2443 -2402
rect 2477 -2436 2500 -2402
rect 2420 -2482 2500 -2436
rect 2420 -2516 2443 -2482
rect 2477 -2516 2500 -2482
rect 2420 -2669 2500 -2516
rect 2800 -2563 2880 -2549
rect 2800 -2615 2814 -2563
rect 2866 -2615 2880 -2563
rect 2800 -2629 2880 -2615
rect 2920 -2669 2960 -1989
rect 3300 -2192 3631 -2169
rect 3300 -2226 3323 -2192
rect 3357 -2209 3631 -2192
rect 3357 -2226 3380 -2209
rect 3300 -2249 3380 -2226
rect 3150 -2363 3230 -2349
rect 3150 -2415 3164 -2363
rect 3216 -2415 3230 -2363
rect 3591 -2370 3631 -2209
rect 3150 -2429 3230 -2415
rect 3572 -2384 3652 -2370
rect 3572 -2436 3586 -2384
rect 3638 -2436 3652 -2384
rect 3000 -2463 3080 -2449
rect 3572 -2450 3652 -2436
rect 3000 -2515 3014 -2463
rect 3066 -2515 3080 -2463
rect 3000 -2529 3080 -2515
rect 3572 -2497 3652 -2483
rect 3572 -2549 3586 -2497
rect 3638 -2549 3652 -2497
rect 3572 -2563 3652 -2549
rect 3680 -2669 3760 -1956
rect 4010 -1762 4090 -1739
rect 4010 -1796 4033 -1762
rect 4067 -1796 4090 -1762
rect 4010 -1842 4090 -1796
rect 4010 -1876 4033 -1842
rect 4067 -1876 4090 -1842
rect 4010 -1922 4090 -1876
rect 4010 -1956 4033 -1922
rect 4067 -1956 4090 -1922
rect 4010 -1989 4090 -1956
rect 4310 -1762 4390 -1739
rect 4310 -1796 4333 -1762
rect 4367 -1796 4390 -1762
rect 4310 -1842 4390 -1796
rect 4310 -1876 4333 -1842
rect 4367 -1876 4390 -1842
rect 4310 -1922 4390 -1876
rect 4310 -1956 4333 -1922
rect 4367 -1956 4390 -1922
rect 4310 -1989 4390 -1956
rect 4610 -1762 4690 -1739
rect 4610 -1796 4633 -1762
rect 4667 -1796 4690 -1762
rect 4610 -1842 4690 -1796
rect 4610 -1876 4633 -1842
rect 4667 -1876 4690 -1842
rect 4610 -1922 4690 -1876
rect 4610 -1956 4633 -1922
rect 4667 -1956 4690 -1922
rect 4610 -1989 4690 -1956
rect 4940 -1762 5020 -1739
rect 4940 -1796 4963 -1762
rect 4997 -1796 5020 -1762
rect 4940 -1842 5020 -1796
rect 4940 -1876 4963 -1842
rect 4997 -1876 5020 -1842
rect 4940 -1922 5020 -1876
rect 4940 -1956 4963 -1922
rect 4997 -1956 5020 -1922
rect 4360 -2199 4440 -2179
rect 4760 -2199 4840 -2179
rect 4360 -2202 4840 -2199
rect 4360 -2236 4383 -2202
rect 4417 -2236 4783 -2202
rect 4817 -2236 4840 -2202
rect 4360 -2239 4840 -2236
rect 4360 -2259 4440 -2239
rect 4760 -2259 4840 -2239
rect 3860 -2313 3940 -2299
rect 3860 -2365 3874 -2313
rect 3926 -2365 3940 -2313
rect 3860 -2379 3940 -2365
rect 4010 -2322 4090 -2299
rect 4010 -2356 4033 -2322
rect 4067 -2356 4090 -2322
rect 3880 -2551 3920 -2379
rect 4010 -2402 4090 -2356
rect 4010 -2436 4033 -2402
rect 4067 -2436 4090 -2402
rect 4010 -2482 4090 -2436
rect 4010 -2516 4033 -2482
rect 4067 -2516 4090 -2482
rect 3860 -2564 3940 -2551
rect 3860 -2616 3874 -2564
rect 3926 -2616 3940 -2564
rect 3860 -2631 3940 -2616
rect 4010 -2669 4090 -2516
rect 4310 -2322 4390 -2299
rect 4310 -2356 4333 -2322
rect 4367 -2356 4390 -2322
rect 4310 -2402 4390 -2356
rect 4310 -2436 4333 -2402
rect 4367 -2436 4390 -2402
rect 4310 -2482 4390 -2436
rect 4310 -2516 4333 -2482
rect 4367 -2516 4390 -2482
rect 4310 -2669 4390 -2516
rect 4610 -2322 4690 -2299
rect 4610 -2356 4633 -2322
rect 4667 -2356 4690 -2322
rect 4610 -2402 4690 -2356
rect 4760 -2313 4840 -2299
rect 4760 -2365 4774 -2313
rect 4826 -2365 4840 -2313
rect 4760 -2379 4840 -2365
rect 4610 -2436 4633 -2402
rect 4667 -2436 4690 -2402
rect 4610 -2482 4690 -2436
rect 4610 -2516 4633 -2482
rect 4667 -2516 4690 -2482
rect 4610 -2669 4690 -2516
rect 4940 -2669 5020 -1956
rect 5560 -1762 5640 -1739
rect 5560 -1796 5583 -1762
rect 5617 -1796 5640 -1762
rect 5560 -1842 5640 -1796
rect 5560 -1876 5583 -1842
rect 5617 -1876 5640 -1842
rect 5560 -1922 5640 -1876
rect 5560 -1956 5583 -1922
rect 5617 -1956 5640 -1922
rect 5560 -1989 5640 -1956
rect 5890 -1762 5970 -1739
rect 5890 -1796 5913 -1762
rect 5947 -1796 5970 -1762
rect 5890 -1842 5970 -1796
rect 5890 -1876 5913 -1842
rect 5947 -1876 5970 -1842
rect 5890 -1922 5970 -1876
rect 5890 -1956 5913 -1922
rect 5947 -1956 5970 -1922
rect 5890 -1989 5970 -1956
rect 6190 -1762 6270 -1739
rect 6190 -1796 6213 -1762
rect 6247 -1796 6270 -1762
rect 6190 -1842 6270 -1796
rect 6190 -1876 6213 -1842
rect 6247 -1876 6270 -1842
rect 6190 -1922 6270 -1876
rect 6190 -1956 6213 -1922
rect 6247 -1956 6270 -1922
rect 6190 -1989 6270 -1956
rect 6490 -1762 6570 -1739
rect 6490 -1796 6513 -1762
rect 6547 -1796 6570 -1762
rect 6490 -1842 6570 -1796
rect 6490 -1876 6513 -1842
rect 6547 -1876 6570 -1842
rect 6490 -1922 6570 -1876
rect 6490 -1956 6513 -1922
rect 6547 -1956 6570 -1922
rect 6490 -1989 6570 -1956
rect 6970 -1753 7050 -1739
rect 6970 -1805 6984 -1753
rect 7036 -1805 7050 -1753
rect 6970 -1842 7050 -1805
rect 6970 -1876 6993 -1842
rect 7027 -1876 7050 -1842
rect 6970 -1922 7050 -1876
rect 6970 -1956 6993 -1922
rect 7027 -1956 7050 -1922
rect 6970 -1989 7050 -1956
rect 5310 -2252 5390 -2229
rect 5310 -2286 5333 -2252
rect 5367 -2286 5390 -2252
rect 5310 -2309 5390 -2286
rect 5048 -2351 5128 -2337
rect 5048 -2403 5062 -2351
rect 5114 -2357 5128 -2351
rect 5330 -2357 5370 -2309
rect 5114 -2397 5370 -2357
rect 5114 -2403 5128 -2397
rect 5048 -2417 5128 -2403
rect 5048 -2459 5128 -2445
rect 5048 -2511 5062 -2459
rect 5114 -2464 5128 -2459
rect 5310 -2464 5390 -2450
rect 5114 -2473 5390 -2464
rect 5114 -2504 5333 -2473
rect 5114 -2511 5128 -2504
rect 5048 -2525 5128 -2511
rect 5310 -2507 5333 -2504
rect 5367 -2507 5390 -2473
rect 5310 -2530 5390 -2507
rect 5580 -2669 5620 -1989
rect 6240 -2199 6320 -2179
rect 6640 -2199 6720 -2179
rect 6240 -2202 6720 -2199
rect 6240 -2236 6263 -2202
rect 6297 -2236 6663 -2202
rect 6697 -2236 6720 -2202
rect 6240 -2239 6720 -2236
rect 6240 -2259 6320 -2239
rect 6640 -2259 6720 -2239
rect 5890 -2322 5970 -2299
rect 5740 -2343 5820 -2329
rect 5740 -2395 5754 -2343
rect 5806 -2395 5820 -2343
rect 5740 -2409 5820 -2395
rect 5890 -2356 5913 -2322
rect 5947 -2356 5970 -2322
rect 5890 -2402 5970 -2356
rect 5890 -2436 5913 -2402
rect 5947 -2436 5970 -2402
rect 5740 -2463 5820 -2449
rect 5740 -2515 5754 -2463
rect 5806 -2515 5820 -2463
rect 5740 -2529 5820 -2515
rect 5890 -2482 5970 -2436
rect 5890 -2516 5913 -2482
rect 5947 -2516 5970 -2482
rect 5890 -2669 5970 -2516
rect 6190 -2322 6270 -2299
rect 6190 -2356 6213 -2322
rect 6247 -2356 6270 -2322
rect 6190 -2402 6270 -2356
rect 6190 -2436 6213 -2402
rect 6247 -2436 6270 -2402
rect 6190 -2482 6270 -2436
rect 6190 -2516 6213 -2482
rect 6247 -2516 6270 -2482
rect 6190 -2669 6270 -2516
rect 6490 -2322 6570 -2299
rect 6490 -2356 6513 -2322
rect 6547 -2356 6570 -2322
rect 6490 -2402 6570 -2356
rect 6490 -2436 6513 -2402
rect 6547 -2436 6570 -2402
rect 6720 -2343 6800 -2329
rect 6720 -2395 6734 -2343
rect 6786 -2395 6800 -2343
rect 6720 -2409 6800 -2395
rect 6490 -2482 6570 -2436
rect 6490 -2516 6513 -2482
rect 6547 -2516 6570 -2482
rect 6490 -2669 6570 -2516
rect 6870 -2463 6950 -2449
rect 6870 -2515 6884 -2463
rect 6936 -2515 6950 -2463
rect 6870 -2529 6950 -2515
rect 6990 -2669 7030 -1989
rect 7073 -2073 7153 -2059
rect 7073 -2125 7087 -2073
rect 7139 -2125 7153 -2073
rect 7073 -2139 7153 -2125
rect 1020 -2693 5040 -2669
rect 1020 -2745 1069 -2693
rect 1121 -2702 5040 -2693
rect 1137 -2736 1183 -2702
rect 1217 -2736 1263 -2702
rect 1297 -2736 1343 -2702
rect 1377 -2736 1423 -2702
rect 1457 -2736 1503 -2702
rect 1537 -2736 1583 -2702
rect 1617 -2736 1663 -2702
rect 1697 -2736 1743 -2702
rect 1777 -2736 1823 -2702
rect 1857 -2736 1903 -2702
rect 1937 -2736 1983 -2702
rect 2017 -2736 2063 -2702
rect 2097 -2736 2143 -2702
rect 2177 -2736 2223 -2702
rect 2257 -2736 2303 -2702
rect 2337 -2736 2383 -2702
rect 2417 -2736 2463 -2702
rect 2497 -2736 2543 -2702
rect 2577 -2736 2623 -2702
rect 2657 -2736 2703 -2702
rect 2737 -2736 2783 -2702
rect 2817 -2736 2863 -2702
rect 2897 -2736 2943 -2702
rect 2977 -2736 3023 -2702
rect 3057 -2736 3103 -2702
rect 3137 -2736 3183 -2702
rect 3217 -2736 3693 -2702
rect 3727 -2736 3773 -2702
rect 3807 -2736 3853 -2702
rect 3887 -2736 3933 -2702
rect 3967 -2736 4013 -2702
rect 4047 -2736 4093 -2702
rect 4127 -2736 4173 -2702
rect 4207 -2736 4253 -2702
rect 4287 -2736 4333 -2702
rect 4367 -2736 4413 -2702
rect 4447 -2736 4493 -2702
rect 4527 -2736 4573 -2702
rect 4607 -2736 4653 -2702
rect 4687 -2736 4733 -2702
rect 4767 -2736 4813 -2702
rect 4847 -2736 4893 -2702
rect 4927 -2736 4973 -2702
rect 5007 -2736 5040 -2702
rect 1121 -2745 5040 -2736
rect 1020 -2769 5040 -2745
rect 5170 -2702 7070 -2669
rect 5170 -2736 5413 -2702
rect 5447 -2736 5493 -2702
rect 5527 -2736 5573 -2702
rect 5607 -2736 5653 -2702
rect 5687 -2736 5733 -2702
rect 5767 -2736 5813 -2702
rect 5847 -2736 5893 -2702
rect 5927 -2736 5973 -2702
rect 6007 -2736 6053 -2702
rect 6087 -2736 6133 -2702
rect 6167 -2736 6213 -2702
rect 6247 -2736 6293 -2702
rect 6327 -2736 6373 -2702
rect 6407 -2736 6453 -2702
rect 6487 -2736 6533 -2702
rect 6567 -2736 6613 -2702
rect 6647 -2736 6693 -2702
rect 6727 -2736 6773 -2702
rect 6807 -2736 6853 -2702
rect 6887 -2736 6933 -2702
rect 6967 -2736 7013 -2702
rect 7047 -2736 7070 -2702
rect 5170 -2769 7070 -2736
rect 5170 -2899 5270 -2769
rect 4801 -2999 5270 -2899
rect 5398 -2927 5478 -2913
rect 5398 -2979 5412 -2927
rect 5464 -2979 5478 -2927
rect 5398 -2993 5478 -2979
rect 7343 -2960 7423 -2946
rect 4801 -3129 4901 -2999
rect 7343 -3012 7357 -2960
rect 7409 -3012 7423 -2960
rect 7343 -3026 7423 -3012
rect 1055 -3154 3161 -3129
rect 1055 -3206 1069 -3154
rect 1121 -3162 3161 -3154
rect 1121 -3196 1184 -3162
rect 1218 -3196 1264 -3162
rect 1298 -3196 1344 -3162
rect 1378 -3196 1424 -3162
rect 1458 -3196 1504 -3162
rect 1538 -3196 1584 -3162
rect 1618 -3196 1664 -3162
rect 1698 -3196 1744 -3162
rect 1778 -3196 1824 -3162
rect 1858 -3196 1904 -3162
rect 1938 -3196 1984 -3162
rect 2018 -3196 2064 -3162
rect 2098 -3196 2144 -3162
rect 2178 -3196 2224 -3162
rect 2258 -3196 2304 -3162
rect 2338 -3196 2384 -3162
rect 2418 -3196 2464 -3162
rect 2498 -3196 2544 -3162
rect 2578 -3196 2624 -3162
rect 2658 -3196 2704 -3162
rect 2738 -3196 2784 -3162
rect 2818 -3196 2864 -3162
rect 2898 -3196 2944 -3162
rect 2978 -3196 3024 -3162
rect 3058 -3196 3104 -3162
rect 3138 -3196 3161 -3162
rect 1121 -3206 3161 -3196
rect 1055 -3229 3161 -3206
rect 3521 -3162 4901 -3129
rect 3521 -3196 3554 -3162
rect 3588 -3196 3634 -3162
rect 3668 -3196 3714 -3162
rect 3748 -3196 3794 -3162
rect 3828 -3196 3874 -3162
rect 3908 -3196 3954 -3162
rect 3988 -3196 4034 -3162
rect 4068 -3196 4114 -3162
rect 4148 -3196 4194 -3162
rect 4228 -3196 4274 -3162
rect 4308 -3196 4354 -3162
rect 4388 -3196 4434 -3162
rect 4468 -3196 4514 -3162
rect 4548 -3196 4594 -3162
rect 4628 -3196 4674 -3162
rect 4708 -3196 4754 -3162
rect 4788 -3196 4834 -3162
rect 4868 -3196 4901 -3162
rect 3521 -3229 4901 -3196
rect 5251 -3154 7251 -3130
rect 5251 -3206 5265 -3154
rect 5317 -3163 7251 -3154
rect 5317 -3197 5354 -3163
rect 5388 -3197 5434 -3163
rect 5468 -3197 5514 -3163
rect 5548 -3197 5594 -3163
rect 5628 -3197 5674 -3163
rect 5708 -3197 5754 -3163
rect 5788 -3197 5834 -3163
rect 5868 -3197 5914 -3163
rect 5948 -3197 5994 -3163
rect 6028 -3197 6074 -3163
rect 6108 -3197 6154 -3163
rect 6188 -3197 6234 -3163
rect 6268 -3197 6314 -3163
rect 6348 -3197 6394 -3163
rect 6428 -3197 6474 -3163
rect 6508 -3197 6554 -3163
rect 6588 -3197 6634 -3163
rect 6668 -3197 6714 -3163
rect 6748 -3197 6794 -3163
rect 6828 -3197 6874 -3163
rect 6908 -3197 6954 -3163
rect 6988 -3197 7034 -3163
rect 7068 -3197 7114 -3163
rect 7148 -3197 7194 -3163
rect 7228 -3197 7251 -3163
rect 5317 -3206 7251 -3197
rect 1211 -3909 1251 -3229
rect 1511 -3909 1551 -3229
rect 1581 -3273 1661 -3259
rect 1581 -3325 1595 -3273
rect 1647 -3325 1661 -3273
rect 1581 -3339 1661 -3325
rect 1671 -3393 1751 -3379
rect 1671 -3445 1685 -3393
rect 1737 -3445 1751 -3393
rect 1671 -3459 1751 -3445
rect 1821 -3382 1901 -3229
rect 1821 -3416 1844 -3382
rect 1878 -3416 1901 -3382
rect 1821 -3462 1901 -3416
rect 1821 -3496 1844 -3462
rect 1878 -3496 1901 -3462
rect 1641 -3513 1721 -3499
rect 1641 -3565 1655 -3513
rect 1707 -3565 1721 -3513
rect 1641 -3579 1721 -3565
rect 1821 -3542 1901 -3496
rect 1821 -3576 1844 -3542
rect 1878 -3576 1901 -3542
rect 1821 -3599 1901 -3576
rect 2121 -3382 2201 -3229
rect 2121 -3416 2144 -3382
rect 2178 -3416 2201 -3382
rect 2121 -3462 2201 -3416
rect 2121 -3496 2144 -3462
rect 2178 -3496 2201 -3462
rect 2121 -3542 2201 -3496
rect 2121 -3576 2144 -3542
rect 2178 -3576 2201 -3542
rect 2121 -3599 2201 -3576
rect 2421 -3382 2501 -3229
rect 2951 -3273 3031 -3259
rect 2951 -3325 2965 -3273
rect 3017 -3325 3031 -3273
rect 2951 -3339 3031 -3325
rect 2421 -3416 2444 -3382
rect 2478 -3416 2501 -3382
rect 2421 -3462 2501 -3416
rect 2801 -3393 2881 -3379
rect 2801 -3445 2815 -3393
rect 2867 -3445 2881 -3393
rect 2801 -3459 2881 -3445
rect 2421 -3496 2444 -3462
rect 2478 -3496 2501 -3462
rect 2421 -3542 2501 -3496
rect 2421 -3576 2444 -3542
rect 2478 -3576 2501 -3542
rect 2421 -3599 2501 -3576
rect 2671 -3513 2751 -3499
rect 2671 -3565 2685 -3513
rect 2737 -3565 2751 -3513
rect 2671 -3579 2751 -3565
rect 2171 -3659 2251 -3639
rect 2571 -3659 2651 -3639
rect 2171 -3662 2651 -3659
rect 2171 -3696 2194 -3662
rect 2228 -3696 2594 -3662
rect 2628 -3696 2651 -3662
rect 2171 -3699 2651 -3696
rect 2171 -3719 2251 -3699
rect 2571 -3719 2651 -3699
rect 3071 -3909 3111 -3229
rect 3433 -3539 3513 -3519
rect 3172 -3542 3513 -3539
rect 3172 -3576 3456 -3542
rect 3490 -3576 3513 -3542
rect 3172 -3579 3513 -3576
rect 3172 -3758 3212 -3579
rect 3433 -3599 3513 -3579
rect 3151 -3781 3231 -3758
rect 3151 -3815 3174 -3781
rect 3208 -3815 3231 -3781
rect 3151 -3838 3231 -3815
rect 1191 -3942 1271 -3909
rect 1191 -3976 1214 -3942
rect 1248 -3976 1271 -3942
rect 1191 -4022 1271 -3976
rect 1191 -4056 1214 -4022
rect 1248 -4056 1271 -4022
rect 1191 -4102 1271 -4056
rect 1191 -4136 1214 -4102
rect 1248 -4136 1271 -4102
rect 1191 -4159 1271 -4136
rect 1491 -3942 1571 -3909
rect 1491 -3976 1514 -3942
rect 1548 -3976 1571 -3942
rect 1491 -4022 1571 -3976
rect 1491 -4056 1514 -4022
rect 1548 -4056 1571 -4022
rect 1491 -4102 1571 -4056
rect 1491 -4136 1514 -4102
rect 1548 -4136 1571 -4102
rect 1491 -4159 1571 -4136
rect 1821 -3942 1901 -3909
rect 1821 -3976 1844 -3942
rect 1878 -3976 1901 -3942
rect 1821 -4022 1901 -3976
rect 1821 -4056 1844 -4022
rect 1878 -4056 1901 -4022
rect 1821 -4102 1901 -4056
rect 1821 -4136 1844 -4102
rect 1878 -4136 1901 -4102
rect 1821 -4159 1901 -4136
rect 2121 -3942 2201 -3909
rect 2121 -3976 2144 -3942
rect 2178 -3976 2201 -3942
rect 2121 -4022 2201 -3976
rect 2121 -4056 2144 -4022
rect 2178 -4056 2201 -4022
rect 2121 -4102 2201 -4056
rect 2121 -4136 2144 -4102
rect 2178 -4136 2201 -4102
rect 2121 -4159 2201 -4136
rect 2421 -3942 2501 -3909
rect 2421 -3976 2444 -3942
rect 2478 -3976 2501 -3942
rect 2421 -4022 2501 -3976
rect 2421 -4056 2444 -4022
rect 2478 -4056 2501 -4022
rect 2421 -4102 2501 -4056
rect 2421 -4136 2444 -4102
rect 2478 -4136 2501 -4102
rect 2421 -4159 2501 -4136
rect 3051 -3942 3131 -3909
rect 3051 -3976 3074 -3942
rect 3108 -3976 3131 -3942
rect 3051 -4022 3131 -3976
rect 3051 -4056 3074 -4022
rect 3108 -4056 3131 -4022
rect 3051 -4093 3131 -4056
rect 3051 -4145 3065 -4093
rect 3117 -4145 3131 -4093
rect 3051 -4159 3131 -4145
rect 3541 -3942 3621 -3229
rect 3871 -3382 3951 -3229
rect 3871 -3416 3894 -3382
rect 3928 -3416 3951 -3382
rect 3871 -3462 3951 -3416
rect 3871 -3496 3894 -3462
rect 3928 -3496 3951 -3462
rect 3721 -3533 3801 -3519
rect 3721 -3585 3735 -3533
rect 3787 -3585 3801 -3533
rect 3721 -3599 3801 -3585
rect 3871 -3542 3951 -3496
rect 3871 -3576 3894 -3542
rect 3928 -3576 3951 -3542
rect 3871 -3599 3951 -3576
rect 4171 -3382 4251 -3229
rect 4171 -3416 4194 -3382
rect 4228 -3416 4251 -3382
rect 4171 -3462 4251 -3416
rect 4171 -3496 4194 -3462
rect 4228 -3496 4251 -3462
rect 4171 -3542 4251 -3496
rect 4171 -3576 4194 -3542
rect 4228 -3576 4251 -3542
rect 4171 -3599 4251 -3576
rect 4471 -3382 4551 -3229
rect 4471 -3416 4494 -3382
rect 4528 -3416 4551 -3382
rect 4471 -3462 4551 -3416
rect 4471 -3496 4494 -3462
rect 4528 -3496 4551 -3462
rect 4471 -3542 4551 -3496
rect 4471 -3576 4494 -3542
rect 4528 -3576 4551 -3542
rect 4471 -3599 4551 -3576
rect 4621 -3533 4701 -3519
rect 4621 -3585 4635 -3533
rect 4687 -3585 4701 -3533
rect 4621 -3599 4701 -3585
rect 4221 -3659 4301 -3639
rect 4621 -3659 4701 -3639
rect 4221 -3662 4701 -3659
rect 4221 -3696 4244 -3662
rect 4278 -3696 4644 -3662
rect 4678 -3696 4701 -3662
rect 4221 -3699 4701 -3696
rect 4221 -3719 4301 -3699
rect 4621 -3719 4701 -3699
rect 3541 -3976 3564 -3942
rect 3598 -3976 3621 -3942
rect 3541 -4022 3621 -3976
rect 3541 -4056 3564 -4022
rect 3598 -4056 3621 -4022
rect 3541 -4102 3621 -4056
rect 3541 -4136 3564 -4102
rect 3598 -4136 3621 -4102
rect 3541 -4159 3621 -4136
rect 3871 -3942 3951 -3909
rect 3871 -3976 3894 -3942
rect 3928 -3976 3951 -3942
rect 3871 -4022 3951 -3976
rect 3871 -4056 3894 -4022
rect 3928 -4056 3951 -4022
rect 3871 -4102 3951 -4056
rect 3871 -4136 3894 -4102
rect 3928 -4136 3951 -4102
rect 3871 -4159 3951 -4136
rect 4171 -3942 4251 -3909
rect 4171 -3976 4194 -3942
rect 4228 -3976 4251 -3942
rect 4171 -4022 4251 -3976
rect 4171 -4056 4194 -4022
rect 4228 -4056 4251 -4022
rect 4171 -4102 4251 -4056
rect 4171 -4136 4194 -4102
rect 4228 -4136 4251 -4102
rect 4171 -4159 4251 -4136
rect 4471 -3942 4551 -3909
rect 4471 -3976 4494 -3942
rect 4528 -3976 4551 -3942
rect 4471 -4022 4551 -3976
rect 4471 -4056 4494 -4022
rect 4528 -4056 4551 -4022
rect 4471 -4102 4551 -4056
rect 4471 -4136 4494 -4102
rect 4528 -4136 4551 -4102
rect 4471 -4159 4551 -4136
rect 4801 -3942 4881 -3229
rect 5251 -3230 7251 -3206
rect 5004 -3360 5084 -3346
rect 5004 -3412 5018 -3360
rect 5070 -3412 5084 -3360
rect 5004 -3426 5084 -3412
rect 5180 -3446 5260 -3432
rect 5180 -3454 5194 -3446
rect 4935 -3494 5194 -3454
rect 4935 -3809 4975 -3494
rect 5180 -3498 5194 -3494
rect 5246 -3498 5260 -3446
rect 5180 -3512 5260 -3498
rect 5180 -3556 5260 -3542
rect 5180 -3608 5194 -3556
rect 5246 -3608 5260 -3556
rect 5180 -3622 5260 -3608
rect 5181 -3670 5261 -3656
rect 5181 -3722 5195 -3670
rect 5247 -3722 5261 -3670
rect 5181 -3736 5261 -3722
rect 5181 -3784 5261 -3770
rect 4915 -3832 4995 -3809
rect 4915 -3866 4938 -3832
rect 4972 -3866 4995 -3832
rect 5181 -3836 5195 -3784
rect 5247 -3836 5261 -3784
rect 5181 -3850 5261 -3836
rect 4915 -3889 4995 -3866
rect 5301 -3910 5341 -3230
rect 5381 -3279 5461 -3265
rect 5381 -3331 5395 -3279
rect 5447 -3331 5461 -3279
rect 5381 -3345 5461 -3331
rect 5481 -3404 5561 -3390
rect 5481 -3456 5495 -3404
rect 5547 -3456 5561 -3404
rect 5481 -3470 5561 -3456
rect 5601 -3910 5641 -3230
rect 5911 -3383 5991 -3230
rect 5911 -3417 5934 -3383
rect 5968 -3417 5991 -3383
rect 5911 -3463 5991 -3417
rect 5681 -3494 5761 -3480
rect 5681 -3546 5695 -3494
rect 5747 -3546 5761 -3494
rect 5681 -3560 5761 -3546
rect 5911 -3497 5934 -3463
rect 5968 -3497 5991 -3463
rect 5911 -3543 5991 -3497
rect 5911 -3577 5934 -3543
rect 5968 -3577 5991 -3543
rect 5911 -3600 5991 -3577
rect 6211 -3383 6291 -3230
rect 6211 -3417 6234 -3383
rect 6268 -3417 6291 -3383
rect 6211 -3463 6291 -3417
rect 6211 -3497 6234 -3463
rect 6268 -3497 6291 -3463
rect 6211 -3543 6291 -3497
rect 6211 -3577 6234 -3543
rect 6268 -3577 6291 -3543
rect 6211 -3600 6291 -3577
rect 6511 -3383 6591 -3230
rect 6661 -3284 6741 -3270
rect 6661 -3336 6675 -3284
rect 6727 -3336 6741 -3284
rect 6661 -3350 6741 -3336
rect 6511 -3417 6534 -3383
rect 6568 -3417 6591 -3383
rect 6511 -3463 6591 -3417
rect 6781 -3394 6861 -3380
rect 6781 -3446 6795 -3394
rect 6847 -3446 6861 -3394
rect 6781 -3460 6861 -3446
rect 7033 -3394 7113 -3380
rect 7033 -3446 7047 -3394
rect 7099 -3446 7113 -3394
rect 7033 -3460 7113 -3446
rect 6511 -3497 6534 -3463
rect 6568 -3497 6591 -3463
rect 6511 -3543 6591 -3497
rect 6511 -3577 6534 -3543
rect 6568 -3577 6591 -3543
rect 6661 -3494 6741 -3480
rect 6661 -3546 6675 -3494
rect 6727 -3546 6741 -3494
rect 6661 -3560 6741 -3546
rect 6511 -3600 6591 -3577
rect 6791 -3582 6871 -3568
rect 6791 -3634 6805 -3582
rect 6857 -3634 6871 -3582
rect 5761 -3660 5841 -3640
rect 6161 -3660 6241 -3640
rect 6791 -3648 6871 -3634
rect 5761 -3663 6241 -3660
rect 5761 -3697 5784 -3663
rect 5818 -3697 6184 -3663
rect 6218 -3697 6241 -3663
rect 5761 -3700 6241 -3697
rect 5761 -3720 5841 -3700
rect 6161 -3720 6241 -3700
rect 6811 -3770 6851 -3648
rect 6791 -3793 6871 -3770
rect 6791 -3827 6814 -3793
rect 6848 -3827 6871 -3793
rect 6791 -3850 6871 -3827
rect 7161 -3910 7201 -3230
rect 7229 -3284 7309 -3270
rect 7229 -3336 7243 -3284
rect 7295 -3336 7309 -3284
rect 7229 -3350 7309 -3336
rect 7275 -3582 7355 -3568
rect 7275 -3634 7289 -3582
rect 7341 -3634 7355 -3582
rect 7275 -3648 7355 -3634
rect 4801 -3976 4824 -3942
rect 4858 -3976 4881 -3942
rect 4801 -4022 4881 -3976
rect 4998 -3937 5078 -3923
rect 4998 -3989 5012 -3937
rect 5064 -3989 5078 -3937
rect 4998 -4003 5078 -3989
rect 5281 -3943 5361 -3910
rect 5281 -3977 5304 -3943
rect 5338 -3977 5361 -3943
rect 4801 -4056 4824 -4022
rect 4858 -4056 4881 -4022
rect 4801 -4093 4881 -4056
rect 4801 -4145 4815 -4093
rect 4867 -4145 4881 -4093
rect 4801 -4159 4881 -4145
rect 5281 -4023 5361 -3977
rect 5281 -4057 5304 -4023
rect 5338 -4057 5361 -4023
rect 5281 -4103 5361 -4057
rect 5281 -4137 5304 -4103
rect 5338 -4137 5361 -4103
rect 1171 -4213 1251 -4199
rect 1171 -4265 1185 -4213
rect 1237 -4265 1251 -4213
rect 1171 -4279 1251 -4265
rect 1841 -4309 1881 -4159
rect 2141 -4309 2181 -4159
rect 2441 -4309 2481 -4159
rect 3891 -4309 3931 -4159
rect 4191 -4309 4231 -4159
rect 4491 -4309 4531 -4159
rect 5281 -4160 5361 -4137
rect 5581 -3943 5661 -3910
rect 5581 -3977 5604 -3943
rect 5638 -3977 5661 -3943
rect 5581 -4023 5661 -3977
rect 5581 -4057 5604 -4023
rect 5638 -4057 5661 -4023
rect 5581 -4103 5661 -4057
rect 5581 -4137 5604 -4103
rect 5638 -4137 5661 -4103
rect 5581 -4160 5661 -4137
rect 5911 -3943 5991 -3910
rect 5911 -3977 5934 -3943
rect 5968 -3977 5991 -3943
rect 5911 -4023 5991 -3977
rect 5911 -4057 5934 -4023
rect 5968 -4057 5991 -4023
rect 5911 -4103 5991 -4057
rect 5911 -4137 5934 -4103
rect 5968 -4137 5991 -4103
rect 5911 -4160 5991 -4137
rect 6211 -3943 6291 -3910
rect 6211 -3977 6234 -3943
rect 6268 -3977 6291 -3943
rect 6211 -4023 6291 -3977
rect 6211 -4057 6234 -4023
rect 6268 -4057 6291 -4023
rect 6211 -4103 6291 -4057
rect 6211 -4137 6234 -4103
rect 6268 -4137 6291 -4103
rect 6211 -4160 6291 -4137
rect 6511 -3943 6591 -3910
rect 6511 -3977 6534 -3943
rect 6568 -3977 6591 -3943
rect 6511 -4023 6591 -3977
rect 6511 -4057 6534 -4023
rect 6568 -4057 6591 -4023
rect 6511 -4103 6591 -4057
rect 6511 -4137 6534 -4103
rect 6568 -4137 6591 -4103
rect 6511 -4160 6591 -4137
rect 7141 -3943 7221 -3910
rect 7141 -3977 7164 -3943
rect 7198 -3977 7221 -3943
rect 7141 -4023 7221 -3977
rect 7141 -4057 7164 -4023
rect 7198 -4057 7221 -4023
rect 7141 -4093 7221 -4057
rect 7141 -4145 7155 -4093
rect 7207 -4145 7221 -4093
rect 7141 -4160 7221 -4145
rect 5092 -4215 5172 -4201
rect 5092 -4267 5106 -4215
rect 5158 -4267 5172 -4215
rect 5092 -4281 5172 -4267
rect 912 -4376 935 -4342
rect 969 -4376 992 -4342
rect 912 -4399 992 -4376
rect 1040 -4310 5251 -4309
rect 5931 -4310 5971 -4160
rect 6231 -4310 6271 -4160
rect 6531 -4310 6571 -4160
rect 7251 -4310 7470 -4309
rect 1040 -4342 7470 -4310
rect 1040 -4376 1184 -4342
rect 1218 -4376 1264 -4342
rect 1298 -4376 1344 -4342
rect 1378 -4376 1424 -4342
rect 1458 -4376 1504 -4342
rect 1538 -4376 1584 -4342
rect 1618 -4376 1664 -4342
rect 1698 -4376 1744 -4342
rect 1778 -4376 1824 -4342
rect 1858 -4376 1904 -4342
rect 1938 -4376 1984 -4342
rect 2018 -4376 2064 -4342
rect 2098 -4376 2144 -4342
rect 2178 -4376 2224 -4342
rect 2258 -4376 2304 -4342
rect 2338 -4376 2384 -4342
rect 2418 -4376 2464 -4342
rect 2498 -4376 2544 -4342
rect 2578 -4376 2624 -4342
rect 2658 -4376 2704 -4342
rect 2738 -4376 2784 -4342
rect 2818 -4376 2864 -4342
rect 2898 -4376 2944 -4342
rect 2978 -4376 3024 -4342
rect 3058 -4376 3104 -4342
rect 3138 -4376 3184 -4342
rect 3218 -4376 3264 -4342
rect 3298 -4376 3554 -4342
rect 3588 -4376 3634 -4342
rect 3668 -4376 3714 -4342
rect 3748 -4376 3794 -4342
rect 3828 -4376 3874 -4342
rect 3908 -4376 3954 -4342
rect 3988 -4376 4034 -4342
rect 4068 -4376 4114 -4342
rect 4148 -4376 4194 -4342
rect 4228 -4376 4274 -4342
rect 4308 -4376 4354 -4342
rect 4388 -4376 4434 -4342
rect 4468 -4376 4514 -4342
rect 4548 -4376 4594 -4342
rect 4628 -4376 4674 -4342
rect 4708 -4376 4754 -4342
rect 4788 -4376 4834 -4342
rect 4868 -4376 4914 -4342
rect 4948 -4376 4994 -4342
rect 5028 -4343 7274 -4342
rect 5028 -4376 5274 -4343
rect 1040 -4377 5274 -4376
rect 5308 -4377 5354 -4343
rect 5388 -4377 5434 -4343
rect 5468 -4377 5514 -4343
rect 5548 -4377 5594 -4343
rect 5628 -4377 5674 -4343
rect 5708 -4377 5754 -4343
rect 5788 -4377 5834 -4343
rect 5868 -4377 5914 -4343
rect 5948 -4377 5994 -4343
rect 6028 -4377 6074 -4343
rect 6108 -4377 6154 -4343
rect 6188 -4377 6234 -4343
rect 6268 -4377 6314 -4343
rect 6348 -4377 6394 -4343
rect 6428 -4377 6474 -4343
rect 6508 -4377 6554 -4343
rect 6588 -4377 6634 -4343
rect 6668 -4377 6714 -4343
rect 6748 -4377 6794 -4343
rect 6828 -4377 6874 -4343
rect 6908 -4377 6954 -4343
rect 6988 -4377 7034 -4343
rect 7068 -4377 7114 -4343
rect 7148 -4377 7194 -4343
rect 7228 -4376 7274 -4343
rect 7308 -4376 7354 -4342
rect 7388 -4376 7470 -4342
rect 7228 -4377 7470 -4376
rect 912 -4422 993 -4399
rect 912 -4456 936 -4422
rect 970 -4456 993 -4422
rect 912 -4479 993 -4456
rect 1040 -4422 7470 -4377
rect 1040 -4456 1063 -4422
rect 1097 -4456 1143 -4422
rect 1177 -4456 1223 -4422
rect 1257 -4456 1303 -4422
rect 1337 -4456 1383 -4422
rect 1417 -4456 1463 -4422
rect 1497 -4456 1543 -4422
rect 1577 -4456 1623 -4422
rect 1657 -4456 1703 -4422
rect 1737 -4456 1783 -4422
rect 1817 -4456 1863 -4422
rect 1897 -4456 1943 -4422
rect 1977 -4456 2023 -4422
rect 2057 -4456 2103 -4422
rect 2137 -4456 2183 -4422
rect 2217 -4456 2263 -4422
rect 2297 -4456 2343 -4422
rect 2377 -4456 2423 -4422
rect 2457 -4456 2503 -4422
rect 2537 -4456 2583 -4422
rect 2617 -4456 2663 -4422
rect 2697 -4456 2743 -4422
rect 2777 -4456 2823 -4422
rect 2857 -4456 2903 -4422
rect 2937 -4456 2983 -4422
rect 3017 -4456 3063 -4422
rect 3097 -4456 3143 -4422
rect 3177 -4456 3223 -4422
rect 3257 -4456 3303 -4422
rect 3337 -4423 7470 -4422
rect 3337 -4456 3594 -4423
rect 1040 -4457 3594 -4456
rect 3628 -4457 3674 -4423
rect 3708 -4457 3754 -4423
rect 3788 -4457 3834 -4423
rect 3868 -4457 3914 -4423
rect 3948 -4457 3994 -4423
rect 4028 -4457 4074 -4423
rect 4108 -4457 4154 -4423
rect 4188 -4457 4234 -4423
rect 4268 -4457 4314 -4423
rect 4348 -4457 4394 -4423
rect 4428 -4457 4474 -4423
rect 4508 -4457 4554 -4423
rect 4588 -4457 4634 -4423
rect 4668 -4457 4714 -4423
rect 4748 -4457 4794 -4423
rect 4828 -4457 4874 -4423
rect 4908 -4457 4954 -4423
rect 4988 -4457 5034 -4423
rect 5068 -4457 5333 -4423
rect 5367 -4457 5413 -4423
rect 5447 -4457 5493 -4423
rect 5527 -4457 5573 -4423
rect 5607 -4457 5653 -4423
rect 5687 -4457 5733 -4423
rect 5767 -4457 5813 -4423
rect 5847 -4457 5893 -4423
rect 5927 -4457 5973 -4423
rect 6007 -4457 6053 -4423
rect 6087 -4457 6133 -4423
rect 6167 -4457 6213 -4423
rect 6247 -4457 6293 -4423
rect 6327 -4457 6373 -4423
rect 6407 -4457 6453 -4423
rect 6487 -4457 6533 -4423
rect 6567 -4457 6613 -4423
rect 6647 -4457 6693 -4423
rect 6727 -4457 6773 -4423
rect 6807 -4457 6853 -4423
rect 6887 -4457 6933 -4423
rect 6967 -4457 7013 -4423
rect 7047 -4457 7093 -4423
rect 7127 -4457 7173 -4423
rect 7207 -4457 7253 -4423
rect 7287 -4457 7333 -4423
rect 7367 -4457 7413 -4423
rect 7447 -4457 7470 -4423
rect 912 -7243 992 -4479
rect 1040 -4489 7470 -4457
rect 1041 -4536 1121 -4522
rect 1041 -4588 1055 -4536
rect 1107 -4588 1121 -4536
rect 1041 -4602 1121 -4588
rect 1880 -4639 1920 -4489
rect 2180 -4639 2220 -4489
rect 2480 -4639 2520 -4489
rect 3360 -4490 7470 -4489
rect 1230 -4662 1310 -4639
rect 1230 -4696 1253 -4662
rect 1287 -4696 1310 -4662
rect 1230 -4742 1310 -4696
rect 1230 -4776 1253 -4742
rect 1287 -4776 1310 -4742
rect 1230 -4822 1310 -4776
rect 1230 -4856 1253 -4822
rect 1287 -4856 1310 -4822
rect 1230 -4889 1310 -4856
rect 1530 -4662 1610 -4639
rect 1530 -4696 1553 -4662
rect 1587 -4696 1610 -4662
rect 1530 -4742 1610 -4696
rect 1530 -4776 1553 -4742
rect 1587 -4776 1610 -4742
rect 1530 -4822 1610 -4776
rect 1530 -4856 1553 -4822
rect 1587 -4856 1610 -4822
rect 1530 -4889 1610 -4856
rect 1860 -4662 1940 -4639
rect 1860 -4696 1883 -4662
rect 1917 -4696 1940 -4662
rect 1860 -4742 1940 -4696
rect 1860 -4776 1883 -4742
rect 1917 -4776 1940 -4742
rect 1860 -4822 1940 -4776
rect 1860 -4856 1883 -4822
rect 1917 -4856 1940 -4822
rect 1860 -4889 1940 -4856
rect 2160 -4662 2240 -4639
rect 2160 -4696 2183 -4662
rect 2217 -4696 2240 -4662
rect 2160 -4742 2240 -4696
rect 2160 -4776 2183 -4742
rect 2217 -4776 2240 -4742
rect 2160 -4822 2240 -4776
rect 2160 -4856 2183 -4822
rect 2217 -4856 2240 -4822
rect 2160 -4889 2240 -4856
rect 2460 -4662 2540 -4639
rect 2460 -4696 2483 -4662
rect 2517 -4696 2540 -4662
rect 2460 -4742 2540 -4696
rect 2460 -4776 2483 -4742
rect 2517 -4776 2540 -4742
rect 2460 -4822 2540 -4776
rect 2460 -4856 2483 -4822
rect 2517 -4856 2540 -4822
rect 2460 -4889 2540 -4856
rect 3240 -4654 3320 -4639
rect 4091 -4640 4131 -4490
rect 4391 -4640 4431 -4490
rect 4691 -4640 4731 -4490
rect 5115 -4534 5195 -4520
rect 5115 -4586 5129 -4534
rect 5181 -4586 5195 -4534
rect 5115 -4600 5195 -4586
rect 5312 -4534 5392 -4520
rect 5312 -4586 5326 -4534
rect 5378 -4586 5392 -4534
rect 5312 -4600 5392 -4586
rect 6150 -4640 6190 -4490
rect 6450 -4640 6490 -4490
rect 6750 -4640 6790 -4490
rect 3240 -4706 3254 -4654
rect 3306 -4706 3320 -4654
rect 3240 -4742 3320 -4706
rect 3240 -4776 3263 -4742
rect 3297 -4776 3320 -4742
rect 3240 -4822 3320 -4776
rect 3240 -4856 3263 -4822
rect 3297 -4856 3320 -4822
rect 3240 -4889 3320 -4856
rect 3741 -4663 3821 -4640
rect 3741 -4697 3764 -4663
rect 3798 -4697 3821 -4663
rect 3741 -4743 3821 -4697
rect 3741 -4777 3764 -4743
rect 3798 -4777 3821 -4743
rect 3741 -4823 3821 -4777
rect 3741 -4857 3764 -4823
rect 3798 -4857 3821 -4823
rect 1130 -5423 1210 -5409
rect 1130 -5475 1144 -5423
rect 1196 -5475 1210 -5423
rect 1130 -5489 1210 -5475
rect 1130 -5543 1210 -5529
rect 1130 -5595 1144 -5543
rect 1196 -5595 1210 -5543
rect 1130 -5609 1210 -5595
rect 1130 -5663 1210 -5649
rect 1130 -5715 1144 -5663
rect 1196 -5715 1210 -5663
rect 1130 -5729 1210 -5715
rect 1130 -5783 1210 -5769
rect 1130 -5835 1144 -5783
rect 1196 -5835 1210 -5783
rect 1130 -5849 1210 -5835
rect 1250 -5889 1290 -4889
rect 1550 -5889 1590 -4889
rect 2690 -5032 2770 -5009
rect 2690 -5066 2713 -5032
rect 2747 -5066 2770 -5032
rect 2690 -5089 2770 -5066
rect 2840 -5032 2920 -5009
rect 2840 -5066 2863 -5032
rect 2897 -5066 2920 -5032
rect 2840 -5089 2920 -5066
rect 2990 -5032 3070 -5009
rect 2990 -5066 3013 -5032
rect 3047 -5066 3070 -5032
rect 2990 -5089 3070 -5066
rect 3140 -5032 3220 -5009
rect 3140 -5066 3163 -5032
rect 3197 -5066 3220 -5032
rect 3140 -5089 3220 -5066
rect 2210 -5329 2290 -5309
rect 2410 -5329 2490 -5309
rect 2210 -5332 2490 -5329
rect 2210 -5366 2233 -5332
rect 2267 -5366 2433 -5332
rect 2467 -5366 2490 -5332
rect 2210 -5369 2490 -5366
rect 2210 -5389 2290 -5369
rect 2410 -5389 2490 -5369
rect 2710 -5409 2750 -5089
rect 2690 -5423 2770 -5409
rect 2690 -5475 2704 -5423
rect 2756 -5475 2770 -5423
rect 2690 -5489 2770 -5475
rect 1860 -5542 1940 -5519
rect 1860 -5576 1883 -5542
rect 1917 -5576 1940 -5542
rect 1860 -5622 1940 -5576
rect 1860 -5656 1883 -5622
rect 1917 -5656 1940 -5622
rect 1860 -5702 1940 -5656
rect 1860 -5736 1883 -5702
rect 1917 -5736 1940 -5702
rect 1860 -5889 1940 -5736
rect 2160 -5542 2240 -5519
rect 2160 -5576 2183 -5542
rect 2217 -5576 2240 -5542
rect 2160 -5622 2240 -5576
rect 2160 -5656 2183 -5622
rect 2217 -5656 2240 -5622
rect 2160 -5702 2240 -5656
rect 2160 -5736 2183 -5702
rect 2217 -5736 2240 -5702
rect 2160 -5889 2240 -5736
rect 2460 -5542 2540 -5519
rect 2860 -5529 2900 -5089
rect 2460 -5576 2483 -5542
rect 2517 -5576 2540 -5542
rect 2460 -5622 2540 -5576
rect 2840 -5543 2920 -5529
rect 2840 -5595 2854 -5543
rect 2906 -5595 2920 -5543
rect 2840 -5609 2920 -5595
rect 2460 -5656 2483 -5622
rect 2517 -5656 2540 -5622
rect 3010 -5649 3050 -5089
rect 2460 -5702 2540 -5656
rect 2460 -5736 2483 -5702
rect 2517 -5736 2540 -5702
rect 2990 -5663 3070 -5649
rect 2990 -5715 3004 -5663
rect 3056 -5715 3070 -5663
rect 2990 -5729 3070 -5715
rect 2460 -5889 2540 -5736
rect 3160 -5769 3200 -5089
rect 3140 -5783 3220 -5769
rect 3140 -5835 3154 -5783
rect 3206 -5835 3220 -5783
rect 3140 -5849 3220 -5835
rect 3260 -5889 3300 -4889
rect 3633 -4980 3713 -4960
rect 3360 -4983 3713 -4980
rect 3360 -5017 3656 -4983
rect 3690 -5017 3713 -4983
rect 3360 -5020 3713 -5017
rect 3360 -5310 3400 -5020
rect 3633 -5040 3713 -5020
rect 3340 -5333 3420 -5310
rect 3340 -5367 3363 -5333
rect 3397 -5367 3420 -5333
rect 3340 -5390 3420 -5367
rect 3741 -5570 3821 -4857
rect 4071 -4663 4151 -4640
rect 4071 -4697 4094 -4663
rect 4128 -4697 4151 -4663
rect 4071 -4743 4151 -4697
rect 4071 -4777 4094 -4743
rect 4128 -4777 4151 -4743
rect 4071 -4823 4151 -4777
rect 4071 -4857 4094 -4823
rect 4128 -4857 4151 -4823
rect 4071 -4890 4151 -4857
rect 4371 -4663 4451 -4640
rect 4371 -4697 4394 -4663
rect 4428 -4697 4451 -4663
rect 4371 -4743 4451 -4697
rect 4371 -4777 4394 -4743
rect 4428 -4777 4451 -4743
rect 4371 -4823 4451 -4777
rect 4371 -4857 4394 -4823
rect 4428 -4857 4451 -4823
rect 4371 -4890 4451 -4857
rect 4671 -4663 4751 -4640
rect 4671 -4697 4694 -4663
rect 4728 -4697 4751 -4663
rect 4671 -4743 4751 -4697
rect 4671 -4777 4694 -4743
rect 4728 -4777 4751 -4743
rect 4671 -4823 4751 -4777
rect 4671 -4857 4694 -4823
rect 4728 -4857 4751 -4823
rect 4671 -4890 4751 -4857
rect 5001 -4654 5081 -4640
rect 5001 -4706 5015 -4654
rect 5067 -4706 5081 -4654
rect 5001 -4743 5081 -4706
rect 5001 -4777 5024 -4743
rect 5058 -4777 5081 -4743
rect 5001 -4823 5081 -4777
rect 5001 -4857 5024 -4823
rect 5058 -4857 5081 -4823
rect 4421 -5100 4501 -5080
rect 4821 -5100 4901 -5080
rect 4421 -5103 4901 -5100
rect 4421 -5137 4444 -5103
rect 4478 -5137 4844 -5103
rect 4878 -5137 4901 -5103
rect 4421 -5140 4901 -5137
rect 4421 -5160 4501 -5140
rect 4821 -5160 4901 -5140
rect 3921 -5214 4001 -5200
rect 3921 -5266 3935 -5214
rect 3987 -5266 4001 -5214
rect 3921 -5280 4001 -5266
rect 4071 -5223 4151 -5200
rect 4071 -5257 4094 -5223
rect 4128 -5257 4151 -5223
rect 4071 -5303 4151 -5257
rect 4071 -5337 4094 -5303
rect 4128 -5337 4151 -5303
rect 4071 -5383 4151 -5337
rect 4071 -5417 4094 -5383
rect 4128 -5417 4151 -5383
rect 4071 -5570 4151 -5417
rect 4371 -5223 4451 -5200
rect 4371 -5257 4394 -5223
rect 4428 -5257 4451 -5223
rect 4371 -5303 4451 -5257
rect 4371 -5337 4394 -5303
rect 4428 -5337 4451 -5303
rect 4371 -5383 4451 -5337
rect 4371 -5417 4394 -5383
rect 4428 -5417 4451 -5383
rect 4371 -5570 4451 -5417
rect 4671 -5223 4751 -5200
rect 4671 -5257 4694 -5223
rect 4728 -5257 4751 -5223
rect 4671 -5303 4751 -5257
rect 4821 -5214 4901 -5200
rect 4821 -5266 4835 -5214
rect 4887 -5266 4901 -5214
rect 4821 -5280 4901 -5266
rect 4671 -5337 4694 -5303
rect 4728 -5337 4751 -5303
rect 4671 -5383 4751 -5337
rect 4671 -5417 4694 -5383
rect 4728 -5417 4751 -5383
rect 4671 -5570 4751 -5417
rect 5001 -5570 5081 -4857
rect 5500 -4663 5580 -4640
rect 5500 -4697 5523 -4663
rect 5557 -4697 5580 -4663
rect 5500 -4743 5580 -4697
rect 5500 -4777 5523 -4743
rect 5557 -4777 5580 -4743
rect 5500 -4823 5580 -4777
rect 5500 -4857 5523 -4823
rect 5557 -4857 5580 -4823
rect 5500 -4890 5580 -4857
rect 5800 -4663 5880 -4640
rect 5800 -4697 5823 -4663
rect 5857 -4697 5880 -4663
rect 5800 -4743 5880 -4697
rect 5800 -4777 5823 -4743
rect 5857 -4777 5880 -4743
rect 5800 -4823 5880 -4777
rect 5800 -4857 5823 -4823
rect 5857 -4857 5880 -4823
rect 5800 -4890 5880 -4857
rect 6130 -4663 6210 -4640
rect 6130 -4697 6153 -4663
rect 6187 -4697 6210 -4663
rect 6130 -4743 6210 -4697
rect 6130 -4777 6153 -4743
rect 6187 -4777 6210 -4743
rect 6130 -4823 6210 -4777
rect 6130 -4857 6153 -4823
rect 6187 -4857 6210 -4823
rect 6130 -4890 6210 -4857
rect 6430 -4663 6510 -4640
rect 6430 -4697 6453 -4663
rect 6487 -4697 6510 -4663
rect 6430 -4743 6510 -4697
rect 6430 -4777 6453 -4743
rect 6487 -4777 6510 -4743
rect 6430 -4823 6510 -4777
rect 6430 -4857 6453 -4823
rect 6487 -4857 6510 -4823
rect 6430 -4890 6510 -4857
rect 6730 -4663 6810 -4640
rect 6730 -4697 6753 -4663
rect 6787 -4697 6810 -4663
rect 6730 -4743 6810 -4697
rect 6730 -4777 6753 -4743
rect 6787 -4777 6810 -4743
rect 6730 -4823 6810 -4777
rect 6730 -4857 6753 -4823
rect 6787 -4857 6810 -4823
rect 6730 -4890 6810 -4857
rect 7360 -4654 7440 -4640
rect 7360 -4706 7374 -4654
rect 7426 -4706 7440 -4654
rect 7360 -4743 7440 -4706
rect 7360 -4777 7383 -4743
rect 7417 -4777 7440 -4743
rect 7360 -4823 7440 -4777
rect 7360 -4857 7383 -4823
rect 7417 -4857 7440 -4823
rect 7360 -4890 7440 -4857
rect 5115 -4933 5195 -4910
rect 5115 -4967 5138 -4933
rect 5172 -4967 5195 -4933
rect 5115 -4990 5195 -4967
rect 5400 -4954 5480 -4940
rect 5135 -5303 5175 -4990
rect 5400 -5006 5414 -4954
rect 5466 -5006 5480 -4954
rect 5400 -5020 5480 -5006
rect 5400 -5074 5480 -5060
rect 5400 -5126 5414 -5074
rect 5466 -5126 5480 -5074
rect 5400 -5140 5480 -5126
rect 5400 -5202 5480 -5188
rect 5400 -5254 5414 -5202
rect 5466 -5254 5480 -5202
rect 5400 -5268 5480 -5254
rect 5135 -5317 5480 -5303
rect 5135 -5343 5414 -5317
rect 5400 -5369 5414 -5343
rect 5466 -5369 5480 -5317
rect 5115 -5387 5195 -5373
rect 5400 -5383 5480 -5369
rect 5115 -5439 5129 -5387
rect 5181 -5439 5195 -5387
rect 5115 -5453 5195 -5439
rect 5520 -5570 5560 -4890
rect 5700 -5344 5780 -5330
rect 5700 -5396 5714 -5344
rect 5766 -5396 5780 -5344
rect 5700 -5410 5780 -5396
rect 5600 -5469 5680 -5455
rect 5600 -5521 5614 -5469
rect 5666 -5521 5680 -5469
rect 5600 -5535 5680 -5521
rect 5820 -5570 5860 -4890
rect 7010 -4973 7090 -4950
rect 7010 -5007 7033 -4973
rect 7067 -5007 7090 -4973
rect 7010 -5030 7090 -5007
rect 5980 -5100 6060 -5080
rect 6380 -5100 6460 -5080
rect 5980 -5103 6460 -5100
rect 5980 -5137 6003 -5103
rect 6037 -5137 6403 -5103
rect 6437 -5137 6460 -5103
rect 5980 -5140 6460 -5137
rect 5980 -5160 6060 -5140
rect 6380 -5160 6460 -5140
rect 7030 -5153 7070 -5030
rect 7010 -5167 7090 -5153
rect 6130 -5223 6210 -5200
rect 5900 -5254 5980 -5240
rect 5900 -5306 5914 -5254
rect 5966 -5306 5980 -5254
rect 5900 -5320 5980 -5306
rect 6130 -5257 6153 -5223
rect 6187 -5257 6210 -5223
rect 6130 -5303 6210 -5257
rect 6130 -5337 6153 -5303
rect 6187 -5337 6210 -5303
rect 6130 -5383 6210 -5337
rect 6130 -5417 6153 -5383
rect 6187 -5417 6210 -5383
rect 6130 -5570 6210 -5417
rect 6430 -5223 6510 -5200
rect 6430 -5257 6453 -5223
rect 6487 -5257 6510 -5223
rect 6430 -5303 6510 -5257
rect 6430 -5337 6453 -5303
rect 6487 -5337 6510 -5303
rect 6430 -5383 6510 -5337
rect 6430 -5417 6453 -5383
rect 6487 -5417 6510 -5383
rect 6430 -5570 6510 -5417
rect 6730 -5223 6810 -5200
rect 6730 -5257 6753 -5223
rect 6787 -5257 6810 -5223
rect 7010 -5219 7024 -5167
rect 7076 -5219 7090 -5167
rect 7010 -5233 7090 -5219
rect 6730 -5303 6810 -5257
rect 6730 -5337 6753 -5303
rect 6787 -5337 6810 -5303
rect 6880 -5254 6960 -5240
rect 6880 -5306 6894 -5254
rect 6946 -5306 6960 -5254
rect 6880 -5320 6960 -5306
rect 6730 -5383 6810 -5337
rect 6730 -5417 6753 -5383
rect 6787 -5417 6810 -5383
rect 6730 -5570 6810 -5417
rect 7000 -5354 7080 -5340
rect 7000 -5406 7014 -5354
rect 7066 -5406 7080 -5354
rect 7000 -5420 7080 -5406
rect 7132 -5353 7212 -5339
rect 7132 -5405 7146 -5353
rect 7198 -5405 7212 -5353
rect 7132 -5419 7212 -5405
rect 6880 -5464 6960 -5450
rect 6880 -5516 6894 -5464
rect 6946 -5516 6960 -5464
rect 6880 -5530 6960 -5516
rect 7270 -5464 7350 -5450
rect 7270 -5516 7284 -5464
rect 7336 -5516 7350 -5464
rect 7270 -5530 7350 -5516
rect 7380 -5570 7420 -4890
rect 7494 -5167 7574 -5153
rect 7494 -5219 7508 -5167
rect 7560 -5219 7574 -5167
rect 7494 -5233 7574 -5219
rect 3721 -5603 5101 -5570
rect 3721 -5637 3754 -5603
rect 3788 -5637 3834 -5603
rect 3868 -5637 3914 -5603
rect 3948 -5637 3994 -5603
rect 4028 -5637 4074 -5603
rect 4108 -5637 4154 -5603
rect 4188 -5637 4234 -5603
rect 4268 -5637 4314 -5603
rect 4348 -5637 4394 -5603
rect 4428 -5637 4474 -5603
rect 4508 -5637 4554 -5603
rect 4588 -5637 4634 -5603
rect 4668 -5637 4714 -5603
rect 4748 -5637 4794 -5603
rect 4828 -5637 4874 -5603
rect 4908 -5637 4954 -5603
rect 4988 -5637 5034 -5603
rect 5068 -5637 5101 -5603
rect 3721 -5670 5101 -5637
rect 5470 -5594 7470 -5570
rect 5470 -5603 5580 -5594
rect 5632 -5603 7470 -5594
rect 5470 -5637 5493 -5603
rect 5527 -5637 5573 -5603
rect 5632 -5637 5653 -5603
rect 5687 -5637 5733 -5603
rect 5767 -5637 5813 -5603
rect 5847 -5637 5893 -5603
rect 5927 -5637 5973 -5603
rect 6007 -5637 6053 -5603
rect 6087 -5637 6133 -5603
rect 6167 -5637 6213 -5603
rect 6247 -5637 6293 -5603
rect 6327 -5637 6373 -5603
rect 6407 -5637 6453 -5603
rect 6487 -5637 6533 -5603
rect 6567 -5637 6613 -5603
rect 6647 -5637 6693 -5603
rect 6727 -5637 6773 -5603
rect 6807 -5637 6853 -5603
rect 6887 -5637 6933 -5603
rect 6967 -5637 7013 -5603
rect 7047 -5637 7093 -5603
rect 7127 -5637 7173 -5603
rect 7207 -5637 7253 -5603
rect 7287 -5637 7333 -5603
rect 7367 -5637 7413 -5603
rect 7447 -5637 7470 -5603
rect 5470 -5646 5580 -5637
rect 5632 -5646 7470 -5637
rect 5470 -5670 7470 -5646
rect 4861 -5800 4961 -5670
rect 7494 -5788 7574 -5774
rect 1040 -5922 3360 -5889
rect 4861 -5900 5330 -5800
rect 5458 -5820 5538 -5806
rect 5458 -5872 5472 -5820
rect 5524 -5872 5538 -5820
rect 7494 -5840 7508 -5788
rect 7560 -5840 7574 -5788
rect 7494 -5854 7574 -5840
rect 5458 -5886 5538 -5872
rect 1040 -5956 1063 -5922
rect 1097 -5956 1143 -5922
rect 1177 -5956 1223 -5922
rect 1257 -5956 1303 -5922
rect 1337 -5956 1383 -5922
rect 1417 -5956 1463 -5922
rect 1497 -5956 1543 -5922
rect 1577 -5956 1623 -5922
rect 1657 -5956 1703 -5922
rect 1737 -5956 1783 -5922
rect 1817 -5956 1863 -5922
rect 1897 -5956 1943 -5922
rect 1977 -5956 2023 -5922
rect 2057 -5956 2103 -5922
rect 2137 -5956 2183 -5922
rect 2217 -5956 2263 -5922
rect 2297 -5956 2343 -5922
rect 2377 -5956 2423 -5922
rect 2457 -5956 2503 -5922
rect 2537 -5956 2583 -5922
rect 2617 -5956 2663 -5922
rect 2697 -5956 2743 -5922
rect 2777 -5956 2823 -5922
rect 2857 -5956 2903 -5922
rect 2937 -5956 2983 -5922
rect 3017 -5956 3063 -5922
rect 3097 -5956 3143 -5922
rect 3177 -5956 3223 -5922
rect 3257 -5956 3303 -5922
rect 3337 -5956 3360 -5922
rect 1040 -6030 3360 -5956
rect 5230 -6030 5330 -5900
rect 1040 -6063 5100 -6030
rect 1040 -6097 1063 -6063
rect 1097 -6097 1143 -6063
rect 1177 -6097 1223 -6063
rect 1257 -6097 1303 -6063
rect 1337 -6097 1383 -6063
rect 1417 -6097 1463 -6063
rect 1497 -6097 1543 -6063
rect 1577 -6097 1623 -6063
rect 1657 -6097 1703 -6063
rect 1737 -6097 1783 -6063
rect 1817 -6097 1863 -6063
rect 1897 -6097 1943 -6063
rect 1977 -6097 2023 -6063
rect 2057 -6097 2103 -6063
rect 2137 -6097 2183 -6063
rect 2217 -6097 2263 -6063
rect 2297 -6097 2343 -6063
rect 2377 -6097 2423 -6063
rect 2457 -6097 2503 -6063
rect 2537 -6097 2583 -6063
rect 2617 -6097 2663 -6063
rect 2697 -6097 2743 -6063
rect 2777 -6097 2823 -6063
rect 2857 -6097 2903 -6063
rect 2937 -6097 2983 -6063
rect 3017 -6097 3063 -6063
rect 3097 -6097 3143 -6063
rect 3177 -6097 3223 -6063
rect 3257 -6097 3303 -6063
rect 3337 -6097 3753 -6063
rect 3787 -6097 3833 -6063
rect 3867 -6097 3913 -6063
rect 3947 -6097 3993 -6063
rect 4027 -6097 4073 -6063
rect 4107 -6097 4153 -6063
rect 4187 -6097 4233 -6063
rect 4267 -6097 4313 -6063
rect 4347 -6097 4393 -6063
rect 4427 -6097 4473 -6063
rect 4507 -6097 4553 -6063
rect 4587 -6097 4633 -6063
rect 4667 -6097 4713 -6063
rect 4747 -6097 4793 -6063
rect 4827 -6097 4873 -6063
rect 4907 -6097 4953 -6063
rect 4987 -6097 5033 -6063
rect 5067 -6097 5100 -6063
rect 1040 -6130 5100 -6097
rect 5230 -6063 7129 -6030
rect 5230 -6097 5472 -6063
rect 5506 -6097 5552 -6063
rect 5586 -6097 5632 -6063
rect 5666 -6097 5712 -6063
rect 5746 -6097 5792 -6063
rect 5826 -6097 5872 -6063
rect 5906 -6097 5952 -6063
rect 5986 -6097 6032 -6063
rect 6066 -6097 6112 -6063
rect 6146 -6097 6192 -6063
rect 6226 -6097 6272 -6063
rect 6306 -6097 6352 -6063
rect 6386 -6097 6432 -6063
rect 6466 -6097 6512 -6063
rect 6546 -6097 6592 -6063
rect 6626 -6097 6672 -6063
rect 6706 -6097 6752 -6063
rect 6786 -6097 6832 -6063
rect 6866 -6097 6912 -6063
rect 6946 -6097 6992 -6063
rect 7026 -6097 7072 -6063
rect 7106 -6097 7129 -6063
rect 5230 -6130 7129 -6097
rect 1400 -6810 1440 -6130
rect 1580 -6184 1660 -6170
rect 1580 -6236 1594 -6184
rect 1646 -6236 1660 -6184
rect 1580 -6250 1660 -6236
rect 1710 -6284 1790 -6270
rect 1710 -6336 1724 -6284
rect 1776 -6336 1790 -6284
rect 1710 -6350 1790 -6336
rect 1860 -6283 1940 -6130
rect 1860 -6317 1883 -6283
rect 1917 -6317 1940 -6283
rect 1860 -6363 1940 -6317
rect 1580 -6384 1660 -6370
rect 1580 -6436 1594 -6384
rect 1646 -6436 1660 -6384
rect 1580 -6450 1660 -6436
rect 1860 -6397 1883 -6363
rect 1917 -6397 1940 -6363
rect 1860 -6443 1940 -6397
rect 1710 -6484 1790 -6470
rect 1710 -6536 1724 -6484
rect 1776 -6536 1790 -6484
rect 1860 -6477 1883 -6443
rect 1917 -6477 1940 -6443
rect 1860 -6500 1940 -6477
rect 2160 -6283 2240 -6130
rect 2160 -6317 2183 -6283
rect 2217 -6317 2240 -6283
rect 2160 -6363 2240 -6317
rect 2160 -6397 2183 -6363
rect 2217 -6397 2240 -6363
rect 2160 -6443 2240 -6397
rect 2160 -6477 2183 -6443
rect 2217 -6477 2240 -6443
rect 2160 -6500 2240 -6477
rect 2460 -6283 2540 -6130
rect 2840 -6184 2920 -6170
rect 2840 -6236 2854 -6184
rect 2906 -6236 2920 -6184
rect 2840 -6250 2920 -6236
rect 2460 -6317 2483 -6283
rect 2517 -6317 2540 -6283
rect 2460 -6363 2540 -6317
rect 2460 -6397 2483 -6363
rect 2517 -6397 2540 -6363
rect 2460 -6443 2540 -6397
rect 2460 -6477 2483 -6443
rect 2517 -6477 2540 -6443
rect 2460 -6500 2540 -6477
rect 2740 -6484 2820 -6470
rect 1710 -6550 1790 -6536
rect 2740 -6536 2754 -6484
rect 2806 -6536 2820 -6484
rect 2210 -6563 2290 -6540
rect 2740 -6550 2820 -6536
rect 2210 -6597 2233 -6563
rect 2267 -6580 2290 -6563
rect 2580 -6573 2660 -6550
rect 2580 -6580 2603 -6573
rect 2267 -6597 2603 -6580
rect 2210 -6607 2603 -6597
rect 2637 -6607 2660 -6573
rect 2210 -6620 2660 -6607
rect 2580 -6630 2660 -6620
rect 2960 -6810 3000 -6130
rect 3040 -6284 3120 -6270
rect 3040 -6336 3054 -6284
rect 3106 -6336 3120 -6284
rect 3040 -6350 3120 -6336
rect 3632 -6284 3712 -6270
rect 3632 -6336 3646 -6284
rect 3698 -6336 3712 -6284
rect 3632 -6350 3712 -6336
rect 3190 -6384 3270 -6370
rect 3190 -6436 3204 -6384
rect 3256 -6436 3270 -6384
rect 3190 -6450 3270 -6436
rect 3340 -6573 3692 -6550
rect 3340 -6607 3363 -6573
rect 3397 -6590 3692 -6573
rect 3397 -6607 3420 -6590
rect 3340 -6630 3420 -6607
rect 1380 -6843 1460 -6810
rect 1380 -6877 1403 -6843
rect 1437 -6877 1460 -6843
rect 1380 -6923 1460 -6877
rect 1380 -6957 1403 -6923
rect 1437 -6957 1460 -6923
rect 1380 -7003 1460 -6957
rect 1380 -7037 1403 -7003
rect 1437 -7037 1460 -7003
rect 1380 -7060 1460 -7037
rect 1860 -6843 1940 -6810
rect 1860 -6877 1883 -6843
rect 1917 -6877 1940 -6843
rect 1860 -6923 1940 -6877
rect 1860 -6957 1883 -6923
rect 1917 -6957 1940 -6923
rect 1860 -7003 1940 -6957
rect 1860 -7037 1883 -7003
rect 1917 -7037 1940 -7003
rect 1860 -7060 1940 -7037
rect 2160 -6843 2240 -6810
rect 2160 -6877 2183 -6843
rect 2217 -6877 2240 -6843
rect 2160 -6923 2240 -6877
rect 2160 -6957 2183 -6923
rect 2217 -6957 2240 -6923
rect 2160 -7003 2240 -6957
rect 2160 -7037 2183 -7003
rect 2217 -7037 2240 -7003
rect 2160 -7060 2240 -7037
rect 2460 -6843 2540 -6810
rect 2460 -6877 2483 -6843
rect 2517 -6877 2540 -6843
rect 2460 -6923 2540 -6877
rect 2460 -6957 2483 -6923
rect 2517 -6957 2540 -6923
rect 2460 -7003 2540 -6957
rect 2460 -7037 2483 -7003
rect 2517 -7037 2540 -7003
rect 2460 -7060 2540 -7037
rect 2940 -6843 3020 -6810
rect 3652 -6829 3692 -6590
rect 2940 -6877 2963 -6843
rect 2997 -6877 3020 -6843
rect 2940 -6923 3020 -6877
rect 3631 -6843 3711 -6829
rect 3631 -6895 3645 -6843
rect 3697 -6895 3711 -6843
rect 2940 -6957 2963 -6923
rect 2997 -6957 3020 -6923
rect 2940 -6994 3020 -6957
rect 3354 -6914 3434 -6899
rect 3631 -6909 3711 -6895
rect 3740 -6843 3820 -6130
rect 3920 -6183 4000 -6168
rect 3920 -6235 3934 -6183
rect 3986 -6235 4000 -6183
rect 3920 -6248 4000 -6235
rect 3940 -6420 3980 -6248
rect 4070 -6283 4150 -6130
rect 4070 -6317 4093 -6283
rect 4127 -6317 4150 -6283
rect 4070 -6363 4150 -6317
rect 4070 -6397 4093 -6363
rect 4127 -6397 4150 -6363
rect 3920 -6434 4000 -6420
rect 3920 -6486 3934 -6434
rect 3986 -6486 4000 -6434
rect 3920 -6500 4000 -6486
rect 4070 -6443 4150 -6397
rect 4070 -6477 4093 -6443
rect 4127 -6477 4150 -6443
rect 4070 -6500 4150 -6477
rect 4370 -6283 4450 -6130
rect 4370 -6317 4393 -6283
rect 4427 -6317 4450 -6283
rect 4370 -6363 4450 -6317
rect 4370 -6397 4393 -6363
rect 4427 -6397 4450 -6363
rect 4370 -6443 4450 -6397
rect 4370 -6477 4393 -6443
rect 4427 -6477 4450 -6443
rect 4370 -6500 4450 -6477
rect 4670 -6283 4750 -6130
rect 4670 -6317 4693 -6283
rect 4727 -6317 4750 -6283
rect 4670 -6363 4750 -6317
rect 4820 -6284 4900 -6270
rect 4820 -6336 4834 -6284
rect 4886 -6336 4900 -6284
rect 4820 -6350 4900 -6336
rect 4670 -6397 4693 -6363
rect 4727 -6397 4750 -6363
rect 4670 -6443 4750 -6397
rect 4670 -6477 4693 -6443
rect 4727 -6477 4750 -6443
rect 4670 -6500 4750 -6477
rect 4820 -6434 4900 -6420
rect 4820 -6486 4834 -6434
rect 4886 -6486 4900 -6434
rect 4820 -6500 4900 -6486
rect 4420 -6560 4500 -6540
rect 4820 -6560 4900 -6540
rect 4420 -6563 4900 -6560
rect 4420 -6597 4443 -6563
rect 4477 -6597 4843 -6563
rect 4877 -6597 4900 -6563
rect 4420 -6600 4900 -6597
rect 4420 -6620 4500 -6600
rect 4820 -6620 4900 -6600
rect 3740 -6877 3763 -6843
rect 3797 -6877 3820 -6843
rect 3354 -6966 3368 -6914
rect 3420 -6966 3434 -6914
rect 3354 -6979 3434 -6966
rect 3740 -6923 3820 -6877
rect 3740 -6957 3763 -6923
rect 3797 -6957 3820 -6923
rect 2940 -7046 2954 -6994
rect 3006 -7046 3020 -6994
rect 2940 -7060 3020 -7046
rect 3740 -7003 3820 -6957
rect 3740 -7037 3763 -7003
rect 3797 -7037 3820 -7003
rect 3740 -7060 3820 -7037
rect 4070 -6843 4150 -6810
rect 4070 -6877 4093 -6843
rect 4127 -6877 4150 -6843
rect 4070 -6923 4150 -6877
rect 4070 -6957 4093 -6923
rect 4127 -6957 4150 -6923
rect 4070 -7003 4150 -6957
rect 4070 -7037 4093 -7003
rect 4127 -7037 4150 -7003
rect 4070 -7060 4150 -7037
rect 4370 -6843 4450 -6810
rect 4370 -6877 4393 -6843
rect 4427 -6877 4450 -6843
rect 4370 -6923 4450 -6877
rect 4370 -6957 4393 -6923
rect 4427 -6957 4450 -6923
rect 4370 -7003 4450 -6957
rect 4370 -7037 4393 -7003
rect 4427 -7037 4450 -7003
rect 4370 -7060 4450 -7037
rect 4670 -6843 4750 -6810
rect 4670 -6877 4693 -6843
rect 4727 -6877 4750 -6843
rect 4670 -6923 4750 -6877
rect 4670 -6957 4693 -6923
rect 4727 -6957 4750 -6923
rect 4670 -7003 4750 -6957
rect 4670 -7037 4693 -7003
rect 4727 -7037 4750 -7003
rect 4670 -7060 4750 -7037
rect 5000 -6843 5080 -6130
rect 5370 -6390 5450 -6370
rect 5128 -6393 5450 -6390
rect 5128 -6427 5393 -6393
rect 5427 -6427 5450 -6393
rect 5128 -6430 5450 -6427
rect 5128 -6710 5168 -6430
rect 5370 -6450 5450 -6430
rect 5370 -6510 5450 -6490
rect 5216 -6513 5450 -6510
rect 5216 -6547 5393 -6513
rect 5427 -6547 5450 -6513
rect 5216 -6550 5450 -6547
rect 5108 -6733 5188 -6710
rect 5108 -6767 5131 -6733
rect 5165 -6767 5188 -6733
rect 5108 -6790 5188 -6767
rect 5000 -6877 5023 -6843
rect 5057 -6877 5080 -6843
rect 5000 -6923 5080 -6877
rect 5108 -6844 5188 -6830
rect 5108 -6896 5122 -6844
rect 5174 -6850 5188 -6844
rect 5216 -6850 5256 -6550
rect 5370 -6570 5450 -6550
rect 5639 -6810 5679 -6130
rect 5799 -6284 5879 -6270
rect 5799 -6336 5813 -6284
rect 5865 -6336 5879 -6284
rect 5799 -6350 5879 -6336
rect 5949 -6283 6029 -6130
rect 5949 -6317 5972 -6283
rect 6006 -6317 6029 -6283
rect 5949 -6363 6029 -6317
rect 5799 -6404 5879 -6390
rect 5799 -6456 5813 -6404
rect 5865 -6456 5879 -6404
rect 5799 -6470 5879 -6456
rect 5949 -6397 5972 -6363
rect 6006 -6397 6029 -6363
rect 5949 -6443 6029 -6397
rect 5949 -6477 5972 -6443
rect 6006 -6477 6029 -6443
rect 5949 -6500 6029 -6477
rect 6249 -6283 6329 -6130
rect 6249 -6317 6272 -6283
rect 6306 -6317 6329 -6283
rect 6249 -6363 6329 -6317
rect 6249 -6397 6272 -6363
rect 6306 -6397 6329 -6363
rect 6249 -6443 6329 -6397
rect 6249 -6477 6272 -6443
rect 6306 -6477 6329 -6443
rect 6249 -6500 6329 -6477
rect 6549 -6283 6629 -6130
rect 6549 -6317 6572 -6283
rect 6606 -6317 6629 -6283
rect 6549 -6363 6629 -6317
rect 6929 -6284 7009 -6270
rect 6929 -6336 6943 -6284
rect 6995 -6336 7009 -6284
rect 6929 -6350 7009 -6336
rect 6549 -6397 6572 -6363
rect 6606 -6397 6629 -6363
rect 6549 -6443 6629 -6397
rect 6549 -6477 6572 -6443
rect 6606 -6477 6629 -6443
rect 6779 -6404 6859 -6390
rect 6779 -6456 6793 -6404
rect 6845 -6456 6859 -6404
rect 6779 -6470 6859 -6456
rect 6549 -6500 6629 -6477
rect 6299 -6560 6379 -6540
rect 6699 -6560 6779 -6540
rect 6299 -6563 6779 -6560
rect 6299 -6597 6322 -6563
rect 6356 -6597 6722 -6563
rect 6756 -6597 6779 -6563
rect 6299 -6600 6779 -6597
rect 6299 -6620 6379 -6600
rect 6699 -6620 6779 -6600
rect 7049 -6810 7089 -6130
rect 7129 -6674 7209 -6660
rect 7129 -6726 7143 -6674
rect 7195 -6726 7209 -6674
rect 7129 -6740 7209 -6726
rect 5174 -6890 5256 -6850
rect 5619 -6843 5699 -6810
rect 5619 -6877 5642 -6843
rect 5676 -6877 5699 -6843
rect 5174 -6896 5188 -6890
rect 5108 -6910 5188 -6896
rect 5000 -6957 5023 -6923
rect 5057 -6957 5080 -6923
rect 5000 -7003 5080 -6957
rect 5000 -7037 5023 -7003
rect 5057 -7037 5080 -7003
rect 5000 -7060 5080 -7037
rect 5619 -6923 5699 -6877
rect 5619 -6957 5642 -6923
rect 5676 -6957 5699 -6923
rect 5619 -7003 5699 -6957
rect 5619 -7037 5642 -7003
rect 5676 -7037 5699 -7003
rect 5619 -7060 5699 -7037
rect 5949 -6843 6029 -6810
rect 5949 -6877 5972 -6843
rect 6006 -6877 6029 -6843
rect 5949 -6923 6029 -6877
rect 5949 -6957 5972 -6923
rect 6006 -6957 6029 -6923
rect 5949 -7003 6029 -6957
rect 5949 -7037 5972 -7003
rect 6006 -7037 6029 -7003
rect 5949 -7060 6029 -7037
rect 6249 -6843 6329 -6810
rect 6249 -6877 6272 -6843
rect 6306 -6877 6329 -6843
rect 6249 -6923 6329 -6877
rect 6249 -6957 6272 -6923
rect 6306 -6957 6329 -6923
rect 6249 -7003 6329 -6957
rect 6249 -7037 6272 -7003
rect 6306 -7037 6329 -7003
rect 6249 -7060 6329 -7037
rect 6549 -6843 6629 -6810
rect 6549 -6877 6572 -6843
rect 6606 -6877 6629 -6843
rect 6549 -6923 6629 -6877
rect 6549 -6957 6572 -6923
rect 6606 -6957 6629 -6923
rect 6549 -7003 6629 -6957
rect 6549 -7037 6572 -7003
rect 6606 -7037 6629 -7003
rect 6549 -7060 6629 -7037
rect 7029 -6843 7109 -6810
rect 7029 -6877 7052 -6843
rect 7086 -6877 7109 -6843
rect 7029 -6923 7109 -6877
rect 7029 -6957 7052 -6923
rect 7086 -6957 7109 -6923
rect 7029 -6980 7109 -6957
rect 7029 -6994 7110 -6980
rect 7029 -7046 7044 -6994
rect 7096 -7046 7110 -6994
rect 7029 -7060 7110 -7046
rect 1492 -7114 1572 -7100
rect 1492 -7166 1506 -7114
rect 1558 -7166 1572 -7114
rect 1492 -7180 1572 -7166
rect 1880 -7210 1920 -7060
rect 2180 -7210 2220 -7060
rect 2480 -7210 2520 -7060
rect 4090 -7210 4130 -7060
rect 4390 -7210 4430 -7060
rect 4690 -7210 4730 -7060
rect 5456 -7114 5536 -7100
rect 5456 -7166 5470 -7114
rect 5522 -7166 5536 -7114
rect 5456 -7180 5536 -7166
rect 5969 -7210 6009 -7060
rect 6269 -7210 6309 -7060
rect 6569 -7210 6609 -7060
rect 912 -7277 935 -7243
rect 969 -7277 992 -7243
rect 912 -10063 992 -7277
rect 1060 -7243 7129 -7210
rect 1060 -7277 1143 -7243
rect 1177 -7277 1223 -7243
rect 1257 -7277 1303 -7243
rect 1337 -7277 1383 -7243
rect 1417 -7277 1463 -7243
rect 1497 -7277 1543 -7243
rect 1577 -7277 1623 -7243
rect 1657 -7277 1703 -7243
rect 1737 -7277 1783 -7243
rect 1817 -7277 1863 -7243
rect 1897 -7277 1943 -7243
rect 1977 -7277 2023 -7243
rect 2057 -7277 2103 -7243
rect 2137 -7277 2183 -7243
rect 2217 -7277 2263 -7243
rect 2297 -7277 2343 -7243
rect 2377 -7277 2423 -7243
rect 2457 -7277 2503 -7243
rect 2537 -7277 2583 -7243
rect 2617 -7277 2663 -7243
rect 2697 -7277 2743 -7243
rect 2777 -7277 2823 -7243
rect 2857 -7277 2903 -7243
rect 2937 -7277 2983 -7243
rect 3017 -7277 3063 -7243
rect 3097 -7277 3143 -7243
rect 3177 -7277 3223 -7243
rect 3257 -7277 3753 -7243
rect 3787 -7277 3833 -7243
rect 3867 -7277 3913 -7243
rect 3947 -7277 3993 -7243
rect 4027 -7277 4073 -7243
rect 4107 -7277 4153 -7243
rect 4187 -7277 4233 -7243
rect 4267 -7277 4313 -7243
rect 4347 -7277 4393 -7243
rect 4427 -7277 4473 -7243
rect 4507 -7277 4553 -7243
rect 4587 -7277 4633 -7243
rect 4667 -7277 4713 -7243
rect 4747 -7277 4793 -7243
rect 4827 -7277 4873 -7243
rect 4907 -7277 4953 -7243
rect 4987 -7277 5033 -7243
rect 5067 -7277 5472 -7243
rect 5506 -7277 5552 -7243
rect 5586 -7277 5632 -7243
rect 5666 -7277 5712 -7243
rect 5746 -7277 5792 -7243
rect 5826 -7277 5872 -7243
rect 5906 -7277 5952 -7243
rect 5986 -7277 6032 -7243
rect 6066 -7277 6112 -7243
rect 6146 -7277 6192 -7243
rect 6226 -7277 6272 -7243
rect 6306 -7277 6352 -7243
rect 6386 -7277 6432 -7243
rect 6466 -7277 6512 -7243
rect 6546 -7277 6592 -7243
rect 6626 -7277 6672 -7243
rect 6706 -7277 6752 -7243
rect 6786 -7277 6832 -7243
rect 6866 -7277 6912 -7243
rect 6946 -7277 6992 -7243
rect 7026 -7277 7072 -7243
rect 7106 -7277 7129 -7243
rect 1060 -7310 7129 -7277
rect 1492 -7354 1572 -7340
rect 1492 -7406 1506 -7354
rect 1558 -7406 1572 -7354
rect 1492 -7420 1572 -7406
rect 1880 -7460 1920 -7310
rect 2180 -7460 2220 -7310
rect 2480 -7460 2520 -7310
rect 4090 -7460 4130 -7310
rect 4390 -7460 4430 -7310
rect 4690 -7460 4730 -7310
rect 5458 -7354 5538 -7340
rect 5458 -7406 5472 -7354
rect 5524 -7406 5538 -7354
rect 5458 -7420 5538 -7406
rect 5969 -7460 6009 -7310
rect 6269 -7460 6309 -7310
rect 6569 -7460 6609 -7310
rect 1380 -7483 1460 -7460
rect 1380 -7517 1403 -7483
rect 1437 -7517 1460 -7483
rect 1380 -7563 1460 -7517
rect 1380 -7597 1403 -7563
rect 1437 -7597 1460 -7563
rect 1380 -7643 1460 -7597
rect 1380 -7677 1403 -7643
rect 1437 -7677 1460 -7643
rect 1380 -7710 1460 -7677
rect 1860 -7483 1940 -7460
rect 1860 -7517 1883 -7483
rect 1917 -7517 1940 -7483
rect 1860 -7563 1940 -7517
rect 1860 -7597 1883 -7563
rect 1917 -7597 1940 -7563
rect 1860 -7643 1940 -7597
rect 1860 -7677 1883 -7643
rect 1917 -7677 1940 -7643
rect 1860 -7710 1940 -7677
rect 2160 -7483 2240 -7460
rect 2160 -7517 2183 -7483
rect 2217 -7517 2240 -7483
rect 2160 -7563 2240 -7517
rect 2160 -7597 2183 -7563
rect 2217 -7597 2240 -7563
rect 2160 -7643 2240 -7597
rect 2160 -7677 2183 -7643
rect 2217 -7677 2240 -7643
rect 2160 -7710 2240 -7677
rect 2460 -7483 2540 -7460
rect 2460 -7517 2483 -7483
rect 2517 -7517 2540 -7483
rect 2460 -7563 2540 -7517
rect 2460 -7597 2483 -7563
rect 2517 -7597 2540 -7563
rect 2460 -7643 2540 -7597
rect 2460 -7677 2483 -7643
rect 2517 -7677 2540 -7643
rect 2460 -7710 2540 -7677
rect 2940 -7474 3020 -7460
rect 2940 -7526 2954 -7474
rect 3006 -7526 3020 -7474
rect 2940 -7563 3020 -7526
rect 3740 -7483 3820 -7460
rect 3740 -7517 3763 -7483
rect 3797 -7517 3820 -7483
rect 2940 -7597 2963 -7563
rect 2997 -7597 3020 -7563
rect 2940 -7643 3020 -7597
rect 3354 -7552 3434 -7537
rect 3354 -7604 3368 -7552
rect 3420 -7604 3434 -7552
rect 3354 -7617 3434 -7604
rect 3740 -7563 3820 -7517
rect 3740 -7597 3763 -7563
rect 3797 -7597 3820 -7563
rect 2940 -7677 2963 -7643
rect 2997 -7677 3020 -7643
rect 2940 -7710 3020 -7677
rect 3740 -7643 3820 -7597
rect 3740 -7677 3763 -7643
rect 3797 -7677 3820 -7643
rect 1400 -8390 1440 -7710
rect 2580 -7900 2660 -7890
rect 2210 -7913 2660 -7900
rect 2210 -7923 2603 -7913
rect 2210 -7957 2233 -7923
rect 2267 -7940 2603 -7923
rect 2267 -7957 2290 -7940
rect 1710 -7984 1790 -7970
rect 2210 -7980 2290 -7957
rect 2580 -7947 2603 -7940
rect 2637 -7947 2660 -7913
rect 2580 -7970 2660 -7947
rect 1710 -8036 1724 -7984
rect 1776 -8036 1790 -7984
rect 2740 -7984 2820 -7970
rect 1710 -8050 1790 -8036
rect 1860 -8043 1940 -8020
rect 1580 -8084 1660 -8070
rect 1580 -8136 1594 -8084
rect 1646 -8136 1660 -8084
rect 1580 -8150 1660 -8136
rect 1860 -8077 1883 -8043
rect 1917 -8077 1940 -8043
rect 1860 -8123 1940 -8077
rect 1860 -8157 1883 -8123
rect 1917 -8157 1940 -8123
rect 1710 -8184 1790 -8170
rect 1710 -8236 1724 -8184
rect 1776 -8236 1790 -8184
rect 1710 -8250 1790 -8236
rect 1860 -8203 1940 -8157
rect 1860 -8237 1883 -8203
rect 1917 -8237 1940 -8203
rect 1580 -8284 1660 -8270
rect 1580 -8336 1594 -8284
rect 1646 -8336 1660 -8284
rect 1580 -8350 1660 -8336
rect 1860 -8390 1940 -8237
rect 2160 -8043 2240 -8020
rect 2160 -8077 2183 -8043
rect 2217 -8077 2240 -8043
rect 2160 -8123 2240 -8077
rect 2160 -8157 2183 -8123
rect 2217 -8157 2240 -8123
rect 2160 -8203 2240 -8157
rect 2160 -8237 2183 -8203
rect 2217 -8237 2240 -8203
rect 2160 -8390 2240 -8237
rect 2460 -8043 2540 -8020
rect 2460 -8077 2483 -8043
rect 2517 -8077 2540 -8043
rect 2740 -8036 2754 -7984
rect 2806 -8036 2820 -7984
rect 2740 -8050 2820 -8036
rect 2460 -8123 2540 -8077
rect 2460 -8157 2483 -8123
rect 2517 -8157 2540 -8123
rect 2460 -8203 2540 -8157
rect 2460 -8237 2483 -8203
rect 2517 -8237 2540 -8203
rect 2460 -8390 2540 -8237
rect 2840 -8284 2920 -8270
rect 2840 -8336 2854 -8284
rect 2906 -8336 2920 -8284
rect 2840 -8350 2920 -8336
rect 2960 -8390 3000 -7710
rect 3340 -7795 3420 -7776
rect 3340 -7799 3692 -7795
rect 3340 -7833 3363 -7799
rect 3397 -7833 3692 -7799
rect 3340 -7835 3692 -7833
rect 3340 -7856 3420 -7835
rect 3190 -8084 3270 -8070
rect 3190 -8136 3204 -8084
rect 3256 -8136 3270 -8084
rect 3652 -8096 3692 -7835
rect 3190 -8150 3270 -8136
rect 3632 -8110 3712 -8096
rect 3632 -8162 3646 -8110
rect 3698 -8162 3712 -8110
rect 3040 -8184 3120 -8170
rect 3632 -8176 3712 -8162
rect 3040 -8236 3054 -8184
rect 3106 -8236 3120 -8184
rect 3040 -8250 3120 -8236
rect 3632 -8218 3712 -8204
rect 3632 -8270 3646 -8218
rect 3698 -8270 3712 -8218
rect 3632 -8284 3712 -8270
rect 3740 -8390 3820 -7677
rect 4070 -7483 4150 -7460
rect 4070 -7517 4093 -7483
rect 4127 -7517 4150 -7483
rect 4070 -7563 4150 -7517
rect 4070 -7597 4093 -7563
rect 4127 -7597 4150 -7563
rect 4070 -7643 4150 -7597
rect 4070 -7677 4093 -7643
rect 4127 -7677 4150 -7643
rect 4070 -7710 4150 -7677
rect 4370 -7483 4450 -7460
rect 4370 -7517 4393 -7483
rect 4427 -7517 4450 -7483
rect 4370 -7563 4450 -7517
rect 4370 -7597 4393 -7563
rect 4427 -7597 4450 -7563
rect 4370 -7643 4450 -7597
rect 4370 -7677 4393 -7643
rect 4427 -7677 4450 -7643
rect 4370 -7710 4450 -7677
rect 4670 -7483 4750 -7460
rect 4670 -7517 4693 -7483
rect 4727 -7517 4750 -7483
rect 4670 -7563 4750 -7517
rect 4670 -7597 4693 -7563
rect 4727 -7597 4750 -7563
rect 4670 -7643 4750 -7597
rect 4670 -7677 4693 -7643
rect 4727 -7677 4750 -7643
rect 4670 -7710 4750 -7677
rect 5000 -7483 5080 -7460
rect 5000 -7517 5023 -7483
rect 5057 -7517 5080 -7483
rect 5000 -7563 5080 -7517
rect 5000 -7597 5023 -7563
rect 5057 -7597 5080 -7563
rect 5000 -7643 5080 -7597
rect 5000 -7677 5023 -7643
rect 5057 -7677 5080 -7643
rect 4420 -7920 4500 -7900
rect 4820 -7920 4900 -7900
rect 4420 -7923 4900 -7920
rect 4420 -7957 4443 -7923
rect 4477 -7957 4843 -7923
rect 4877 -7957 4900 -7923
rect 4420 -7960 4900 -7957
rect 4420 -7980 4500 -7960
rect 4820 -7980 4900 -7960
rect 3920 -8034 4000 -8020
rect 3920 -8086 3934 -8034
rect 3986 -8086 4000 -8034
rect 3920 -8100 4000 -8086
rect 4070 -8043 4150 -8020
rect 4070 -8077 4093 -8043
rect 4127 -8077 4150 -8043
rect 3940 -8272 3980 -8100
rect 4070 -8123 4150 -8077
rect 4070 -8157 4093 -8123
rect 4127 -8157 4150 -8123
rect 4070 -8203 4150 -8157
rect 4070 -8237 4093 -8203
rect 4127 -8237 4150 -8203
rect 3920 -8287 4000 -8272
rect 3920 -8339 3934 -8287
rect 3986 -8339 4000 -8287
rect 3920 -8352 4000 -8339
rect 4070 -8390 4150 -8237
rect 4370 -8043 4450 -8020
rect 4370 -8077 4393 -8043
rect 4427 -8077 4450 -8043
rect 4370 -8123 4450 -8077
rect 4370 -8157 4393 -8123
rect 4427 -8157 4450 -8123
rect 4370 -8203 4450 -8157
rect 4370 -8237 4393 -8203
rect 4427 -8237 4450 -8203
rect 4370 -8390 4450 -8237
rect 4670 -8043 4750 -8020
rect 4670 -8077 4693 -8043
rect 4727 -8077 4750 -8043
rect 4670 -8123 4750 -8077
rect 4820 -8034 4900 -8020
rect 4820 -8086 4834 -8034
rect 4886 -8086 4900 -8034
rect 4820 -8100 4900 -8086
rect 4670 -8157 4693 -8123
rect 4727 -8157 4750 -8123
rect 4670 -8203 4750 -8157
rect 4670 -8237 4693 -8203
rect 4727 -8237 4750 -8203
rect 4670 -8390 4750 -8237
rect 5000 -8390 5080 -7677
rect 5619 -7483 5699 -7460
rect 5619 -7517 5642 -7483
rect 5676 -7517 5699 -7483
rect 5619 -7563 5699 -7517
rect 5619 -7597 5642 -7563
rect 5676 -7597 5699 -7563
rect 5619 -7643 5699 -7597
rect 5619 -7677 5642 -7643
rect 5676 -7677 5699 -7643
rect 5619 -7710 5699 -7677
rect 5949 -7483 6029 -7460
rect 5949 -7517 5972 -7483
rect 6006 -7517 6029 -7483
rect 5949 -7563 6029 -7517
rect 5949 -7597 5972 -7563
rect 6006 -7597 6029 -7563
rect 5949 -7643 6029 -7597
rect 5949 -7677 5972 -7643
rect 6006 -7677 6029 -7643
rect 5949 -7710 6029 -7677
rect 6249 -7483 6329 -7460
rect 6249 -7517 6272 -7483
rect 6306 -7517 6329 -7483
rect 6249 -7563 6329 -7517
rect 6249 -7597 6272 -7563
rect 6306 -7597 6329 -7563
rect 6249 -7643 6329 -7597
rect 6249 -7677 6272 -7643
rect 6306 -7677 6329 -7643
rect 6249 -7710 6329 -7677
rect 6549 -7483 6629 -7460
rect 6549 -7517 6572 -7483
rect 6606 -7517 6629 -7483
rect 6549 -7563 6629 -7517
rect 6549 -7597 6572 -7563
rect 6606 -7597 6629 -7563
rect 6549 -7643 6629 -7597
rect 6549 -7677 6572 -7643
rect 6606 -7677 6629 -7643
rect 6549 -7710 6629 -7677
rect 7029 -7474 7110 -7460
rect 7029 -7526 7044 -7474
rect 7096 -7526 7110 -7474
rect 7029 -7540 7110 -7526
rect 7029 -7563 7109 -7540
rect 7029 -7597 7052 -7563
rect 7086 -7597 7109 -7563
rect 7029 -7643 7109 -7597
rect 7029 -7677 7052 -7643
rect 7086 -7677 7109 -7643
rect 7029 -7710 7109 -7677
rect 5108 -7770 5188 -7750
rect 5108 -7773 5430 -7770
rect 5108 -7807 5131 -7773
rect 5165 -7807 5430 -7773
rect 5108 -7810 5430 -7807
rect 5108 -7830 5188 -7810
rect 5390 -8070 5430 -7810
rect 5108 -8103 5188 -8089
rect 5108 -8155 5122 -8103
rect 5174 -8155 5188 -8103
rect 5370 -8093 5450 -8070
rect 5370 -8127 5393 -8093
rect 5427 -8127 5450 -8093
rect 5370 -8150 5450 -8127
rect 5108 -8169 5188 -8155
rect 5108 -8218 5188 -8204
rect 5108 -8270 5122 -8218
rect 5174 -8270 5188 -8218
rect 5108 -8284 5188 -8270
rect 5639 -8390 5679 -7710
rect 6299 -7920 6379 -7900
rect 6699 -7920 6779 -7900
rect 6299 -7923 6779 -7920
rect 6299 -7957 6322 -7923
rect 6356 -7957 6722 -7923
rect 6756 -7957 6779 -7923
rect 6299 -7960 6779 -7957
rect 6299 -7980 6379 -7960
rect 6699 -7980 6779 -7960
rect 5949 -8043 6029 -8020
rect 5799 -8064 5879 -8050
rect 5799 -8116 5813 -8064
rect 5865 -8116 5879 -8064
rect 5799 -8130 5879 -8116
rect 5949 -8077 5972 -8043
rect 6006 -8077 6029 -8043
rect 5949 -8123 6029 -8077
rect 5949 -8157 5972 -8123
rect 6006 -8157 6029 -8123
rect 5799 -8184 5879 -8170
rect 5799 -8236 5813 -8184
rect 5865 -8236 5879 -8184
rect 5799 -8250 5879 -8236
rect 5949 -8203 6029 -8157
rect 5949 -8237 5972 -8203
rect 6006 -8237 6029 -8203
rect 5949 -8390 6029 -8237
rect 6249 -8043 6329 -8020
rect 6249 -8077 6272 -8043
rect 6306 -8077 6329 -8043
rect 6249 -8123 6329 -8077
rect 6249 -8157 6272 -8123
rect 6306 -8157 6329 -8123
rect 6249 -8203 6329 -8157
rect 6249 -8237 6272 -8203
rect 6306 -8237 6329 -8203
rect 6249 -8390 6329 -8237
rect 6549 -8043 6629 -8020
rect 6549 -8077 6572 -8043
rect 6606 -8077 6629 -8043
rect 6549 -8123 6629 -8077
rect 6549 -8157 6572 -8123
rect 6606 -8157 6629 -8123
rect 6779 -8064 6859 -8050
rect 6779 -8116 6793 -8064
rect 6845 -8116 6859 -8064
rect 6779 -8130 6859 -8116
rect 6549 -8203 6629 -8157
rect 6549 -8237 6572 -8203
rect 6606 -8237 6629 -8203
rect 6549 -8390 6629 -8237
rect 6929 -8184 7009 -8170
rect 6929 -8236 6943 -8184
rect 6995 -8236 7009 -8184
rect 6929 -8250 7009 -8236
rect 7049 -8390 7089 -7710
rect 7133 -7795 7213 -7781
rect 7133 -7847 7147 -7795
rect 7199 -7847 7213 -7795
rect 7133 -7861 7213 -7847
rect 1060 -8414 5100 -8390
rect 1060 -8466 1134 -8414
rect 1186 -8423 5100 -8414
rect 1186 -8457 1223 -8423
rect 1257 -8457 1303 -8423
rect 1337 -8457 1383 -8423
rect 1417 -8457 1463 -8423
rect 1497 -8457 1543 -8423
rect 1577 -8457 1623 -8423
rect 1657 -8457 1703 -8423
rect 1737 -8457 1783 -8423
rect 1817 -8457 1863 -8423
rect 1897 -8457 1943 -8423
rect 1977 -8457 2023 -8423
rect 2057 -8457 2103 -8423
rect 2137 -8457 2183 -8423
rect 2217 -8457 2263 -8423
rect 2297 -8457 2343 -8423
rect 2377 -8457 2423 -8423
rect 2457 -8457 2503 -8423
rect 2537 -8457 2583 -8423
rect 2617 -8457 2663 -8423
rect 2697 -8457 2743 -8423
rect 2777 -8457 2823 -8423
rect 2857 -8457 2903 -8423
rect 2937 -8457 2983 -8423
rect 3017 -8457 3063 -8423
rect 3097 -8457 3143 -8423
rect 3177 -8457 3223 -8423
rect 3257 -8457 3753 -8423
rect 3787 -8457 3833 -8423
rect 3867 -8457 3913 -8423
rect 3947 -8457 3993 -8423
rect 4027 -8457 4073 -8423
rect 4107 -8457 4153 -8423
rect 4187 -8457 4233 -8423
rect 4267 -8457 4313 -8423
rect 4347 -8457 4393 -8423
rect 4427 -8457 4473 -8423
rect 4507 -8457 4553 -8423
rect 4587 -8457 4633 -8423
rect 4667 -8457 4713 -8423
rect 4747 -8457 4793 -8423
rect 4827 -8457 4873 -8423
rect 4907 -8457 4953 -8423
rect 4987 -8457 5033 -8423
rect 5067 -8457 5100 -8423
rect 1186 -8466 5100 -8457
rect 1060 -8490 5100 -8466
rect 5449 -8414 7129 -8390
rect 5449 -8423 5704 -8414
rect 5756 -8423 7129 -8414
rect 5449 -8457 5472 -8423
rect 5506 -8457 5552 -8423
rect 5586 -8457 5632 -8423
rect 5666 -8457 5704 -8423
rect 5756 -8457 5792 -8423
rect 5826 -8457 5872 -8423
rect 5906 -8457 5952 -8423
rect 5986 -8457 6032 -8423
rect 6066 -8457 6112 -8423
rect 6146 -8457 6192 -8423
rect 6226 -8457 6272 -8423
rect 6306 -8457 6352 -8423
rect 6386 -8457 6432 -8423
rect 6466 -8457 6512 -8423
rect 6546 -8457 6592 -8423
rect 6626 -8457 6672 -8423
rect 6706 -8457 6752 -8423
rect 6786 -8457 6832 -8423
rect 6866 -8457 6912 -8423
rect 6946 -8457 6992 -8423
rect 7026 -8457 7072 -8423
rect 7106 -8457 7129 -8423
rect 5449 -8466 5704 -8457
rect 5756 -8466 7129 -8457
rect 5449 -8490 7129 -8466
rect 5418 -8532 5538 -8518
rect 5418 -8584 5472 -8532
rect 5524 -8584 5538 -8532
rect 5418 -8598 5538 -8584
rect 5418 -8742 5458 -8598
rect 5398 -8756 5478 -8742
rect 5398 -8808 5412 -8756
rect 5464 -8808 5478 -8756
rect 5398 -8822 5478 -8808
rect 1020 -8874 5040 -8850
rect 1020 -8926 1070 -8874
rect 1122 -8883 5040 -8874
rect 1137 -8917 1183 -8883
rect 1217 -8917 1263 -8883
rect 1297 -8917 1343 -8883
rect 1377 -8917 1423 -8883
rect 1457 -8917 1503 -8883
rect 1537 -8917 1583 -8883
rect 1617 -8917 1663 -8883
rect 1697 -8917 1743 -8883
rect 1777 -8917 1823 -8883
rect 1857 -8917 1903 -8883
rect 1937 -8917 1983 -8883
rect 2017 -8917 2063 -8883
rect 2097 -8917 2143 -8883
rect 2177 -8917 2223 -8883
rect 2257 -8917 2303 -8883
rect 2337 -8917 2383 -8883
rect 2417 -8917 2463 -8883
rect 2497 -8917 2543 -8883
rect 2577 -8917 2623 -8883
rect 2657 -8917 2703 -8883
rect 2737 -8917 2783 -8883
rect 2817 -8917 2863 -8883
rect 2897 -8917 2943 -8883
rect 2977 -8917 3023 -8883
rect 3057 -8917 3103 -8883
rect 3137 -8917 3183 -8883
rect 3217 -8917 3693 -8883
rect 3727 -8917 3773 -8883
rect 3807 -8917 3853 -8883
rect 3887 -8917 3933 -8883
rect 3967 -8917 4013 -8883
rect 4047 -8917 4093 -8883
rect 4127 -8917 4173 -8883
rect 4207 -8917 4253 -8883
rect 4287 -8917 4333 -8883
rect 4367 -8917 4413 -8883
rect 4447 -8917 4493 -8883
rect 4527 -8917 4573 -8883
rect 4607 -8917 4653 -8883
rect 4687 -8917 4733 -8883
rect 4767 -8917 4813 -8883
rect 4847 -8917 4893 -8883
rect 4927 -8917 4973 -8883
rect 5007 -8917 5040 -8883
rect 1122 -8926 5040 -8917
rect 1020 -8950 5040 -8926
rect 5390 -8874 7070 -8850
rect 5390 -8883 5704 -8874
rect 5756 -8883 7004 -8874
rect 5390 -8917 5413 -8883
rect 5447 -8917 5493 -8883
rect 5527 -8917 5573 -8883
rect 5607 -8917 5653 -8883
rect 5687 -8917 5704 -8883
rect 5767 -8917 5813 -8883
rect 5847 -8917 5893 -8883
rect 5927 -8917 5973 -8883
rect 6007 -8917 6053 -8883
rect 6087 -8917 6133 -8883
rect 6167 -8917 6213 -8883
rect 6247 -8917 6293 -8883
rect 6327 -8917 6373 -8883
rect 6407 -8917 6453 -8883
rect 6487 -8917 6533 -8883
rect 6567 -8917 6613 -8883
rect 6647 -8917 6693 -8883
rect 6727 -8917 6773 -8883
rect 6807 -8917 6853 -8883
rect 6887 -8917 6933 -8883
rect 6967 -8917 7004 -8883
rect 5390 -8926 5704 -8917
rect 5756 -8926 7004 -8917
rect 7056 -8926 7070 -8874
rect 5390 -8950 7070 -8926
rect 1360 -9630 1400 -8950
rect 1540 -9004 1620 -8990
rect 1540 -9056 1554 -9004
rect 1606 -9056 1620 -9004
rect 1540 -9070 1620 -9056
rect 1670 -9104 1750 -9090
rect 1670 -9156 1684 -9104
rect 1736 -9156 1750 -9104
rect 1670 -9170 1750 -9156
rect 1820 -9103 1900 -8950
rect 1820 -9137 1843 -9103
rect 1877 -9137 1900 -9103
rect 1820 -9183 1900 -9137
rect 1540 -9204 1620 -9190
rect 1540 -9256 1554 -9204
rect 1606 -9256 1620 -9204
rect 1540 -9270 1620 -9256
rect 1820 -9217 1843 -9183
rect 1877 -9217 1900 -9183
rect 1820 -9263 1900 -9217
rect 1670 -9304 1750 -9290
rect 1670 -9356 1684 -9304
rect 1736 -9356 1750 -9304
rect 1820 -9297 1843 -9263
rect 1877 -9297 1900 -9263
rect 1820 -9320 1900 -9297
rect 2120 -9103 2200 -8950
rect 2120 -9137 2143 -9103
rect 2177 -9137 2200 -9103
rect 2120 -9183 2200 -9137
rect 2120 -9217 2143 -9183
rect 2177 -9217 2200 -9183
rect 2120 -9263 2200 -9217
rect 2120 -9297 2143 -9263
rect 2177 -9297 2200 -9263
rect 2120 -9320 2200 -9297
rect 2420 -9103 2500 -8950
rect 2800 -9004 2880 -8990
rect 2800 -9056 2814 -9004
rect 2866 -9056 2880 -9004
rect 2800 -9070 2880 -9056
rect 2420 -9137 2443 -9103
rect 2477 -9137 2500 -9103
rect 2420 -9183 2500 -9137
rect 2420 -9217 2443 -9183
rect 2477 -9217 2500 -9183
rect 2420 -9263 2500 -9217
rect 2420 -9297 2443 -9263
rect 2477 -9297 2500 -9263
rect 2420 -9320 2500 -9297
rect 2700 -9304 2780 -9290
rect 1670 -9370 1750 -9356
rect 2700 -9356 2714 -9304
rect 2766 -9356 2780 -9304
rect 2170 -9383 2250 -9360
rect 2700 -9370 2780 -9356
rect 2170 -9417 2193 -9383
rect 2227 -9400 2250 -9383
rect 2540 -9393 2620 -9370
rect 2540 -9400 2563 -9393
rect 2227 -9417 2563 -9400
rect 2170 -9427 2563 -9417
rect 2597 -9427 2620 -9393
rect 2170 -9440 2620 -9427
rect 2540 -9450 2620 -9440
rect 2920 -9630 2960 -8950
rect 3572 -9070 3652 -9056
rect 3000 -9104 3080 -9090
rect 3000 -9156 3014 -9104
rect 3066 -9156 3080 -9104
rect 3572 -9122 3586 -9070
rect 3638 -9122 3652 -9070
rect 3572 -9136 3652 -9122
rect 3000 -9170 3080 -9156
rect 3572 -9181 3652 -9167
rect 3150 -9204 3230 -9190
rect 3150 -9256 3164 -9204
rect 3216 -9256 3230 -9204
rect 3572 -9233 3586 -9181
rect 3638 -9233 3652 -9181
rect 3572 -9247 3652 -9233
rect 3150 -9270 3230 -9256
rect 3300 -9505 3380 -9484
rect 3591 -9505 3631 -9247
rect 3300 -9507 3631 -9505
rect 3300 -9541 3323 -9507
rect 3357 -9541 3631 -9507
rect 3300 -9545 3631 -9541
rect 3300 -9564 3380 -9545
rect 1340 -9663 1420 -9630
rect 1340 -9697 1363 -9663
rect 1397 -9697 1420 -9663
rect 1340 -9743 1420 -9697
rect 1340 -9777 1363 -9743
rect 1397 -9777 1420 -9743
rect 1340 -9823 1420 -9777
rect 1340 -9857 1363 -9823
rect 1397 -9857 1420 -9823
rect 1340 -9880 1420 -9857
rect 1820 -9663 1900 -9630
rect 1820 -9697 1843 -9663
rect 1877 -9697 1900 -9663
rect 1820 -9743 1900 -9697
rect 1820 -9777 1843 -9743
rect 1877 -9777 1900 -9743
rect 1820 -9823 1900 -9777
rect 1820 -9857 1843 -9823
rect 1877 -9857 1900 -9823
rect 1820 -9880 1900 -9857
rect 2120 -9663 2200 -9630
rect 2120 -9697 2143 -9663
rect 2177 -9697 2200 -9663
rect 2120 -9743 2200 -9697
rect 2120 -9777 2143 -9743
rect 2177 -9777 2200 -9743
rect 2120 -9823 2200 -9777
rect 2120 -9857 2143 -9823
rect 2177 -9857 2200 -9823
rect 2120 -9880 2200 -9857
rect 2420 -9663 2500 -9630
rect 2420 -9697 2443 -9663
rect 2477 -9697 2500 -9663
rect 2420 -9743 2500 -9697
rect 2420 -9777 2443 -9743
rect 2477 -9777 2500 -9743
rect 2420 -9823 2500 -9777
rect 2420 -9857 2443 -9823
rect 2477 -9857 2500 -9823
rect 2420 -9880 2500 -9857
rect 2900 -9663 2980 -9630
rect 2900 -9697 2923 -9663
rect 2957 -9697 2980 -9663
rect 3680 -9663 3760 -8950
rect 3860 -9001 3940 -8988
rect 3860 -9053 3874 -9001
rect 3926 -9053 3940 -9001
rect 3860 -9068 3940 -9053
rect 3880 -9240 3920 -9068
rect 4010 -9103 4090 -8950
rect 4010 -9137 4033 -9103
rect 4067 -9137 4090 -9103
rect 4010 -9183 4090 -9137
rect 4010 -9217 4033 -9183
rect 4067 -9217 4090 -9183
rect 3860 -9254 3940 -9240
rect 3860 -9306 3874 -9254
rect 3926 -9306 3940 -9254
rect 3860 -9320 3940 -9306
rect 4010 -9263 4090 -9217
rect 4010 -9297 4033 -9263
rect 4067 -9297 4090 -9263
rect 4010 -9320 4090 -9297
rect 4310 -9103 4390 -8950
rect 4310 -9137 4333 -9103
rect 4367 -9137 4390 -9103
rect 4310 -9183 4390 -9137
rect 4310 -9217 4333 -9183
rect 4367 -9217 4390 -9183
rect 4310 -9263 4390 -9217
rect 4310 -9297 4333 -9263
rect 4367 -9297 4390 -9263
rect 4310 -9320 4390 -9297
rect 4610 -9103 4690 -8950
rect 4610 -9137 4633 -9103
rect 4667 -9137 4690 -9103
rect 4610 -9183 4690 -9137
rect 4610 -9217 4633 -9183
rect 4667 -9217 4690 -9183
rect 4610 -9263 4690 -9217
rect 4610 -9297 4633 -9263
rect 4667 -9297 4690 -9263
rect 4610 -9320 4690 -9297
rect 4760 -9254 4840 -9240
rect 4760 -9306 4774 -9254
rect 4826 -9306 4840 -9254
rect 4760 -9320 4840 -9306
rect 4360 -9380 4440 -9360
rect 4760 -9380 4840 -9360
rect 4360 -9383 4840 -9380
rect 4360 -9417 4383 -9383
rect 4417 -9417 4783 -9383
rect 4817 -9417 4840 -9383
rect 4360 -9420 4840 -9417
rect 4360 -9440 4440 -9420
rect 4760 -9440 4840 -9420
rect 2900 -9743 2980 -9697
rect 2900 -9777 2923 -9743
rect 2957 -9777 2980 -9743
rect 3314 -9702 3394 -9689
rect 3314 -9754 3328 -9702
rect 3380 -9754 3394 -9702
rect 3314 -9769 3394 -9754
rect 3680 -9697 3703 -9663
rect 3737 -9697 3760 -9663
rect 3680 -9743 3760 -9697
rect 2900 -9823 2980 -9777
rect 2900 -9857 2923 -9823
rect 2957 -9857 2980 -9823
rect 2900 -9880 2980 -9857
rect 3680 -9777 3703 -9743
rect 3737 -9777 3760 -9743
rect 3680 -9823 3760 -9777
rect 3680 -9857 3703 -9823
rect 3737 -9857 3760 -9823
rect 3680 -9880 3760 -9857
rect 4010 -9663 4090 -9630
rect 4010 -9697 4033 -9663
rect 4067 -9697 4090 -9663
rect 4010 -9743 4090 -9697
rect 4010 -9777 4033 -9743
rect 4067 -9777 4090 -9743
rect 4010 -9823 4090 -9777
rect 4010 -9857 4033 -9823
rect 4067 -9857 4090 -9823
rect 4010 -9880 4090 -9857
rect 4310 -9663 4390 -9630
rect 4310 -9697 4333 -9663
rect 4367 -9697 4390 -9663
rect 4310 -9743 4390 -9697
rect 4310 -9777 4333 -9743
rect 4367 -9777 4390 -9743
rect 4310 -9823 4390 -9777
rect 4310 -9857 4333 -9823
rect 4367 -9857 4390 -9823
rect 4310 -9880 4390 -9857
rect 4610 -9663 4690 -9630
rect 4610 -9697 4633 -9663
rect 4667 -9697 4690 -9663
rect 4610 -9743 4690 -9697
rect 4610 -9777 4633 -9743
rect 4667 -9777 4690 -9743
rect 4610 -9823 4690 -9777
rect 4610 -9857 4633 -9823
rect 4667 -9857 4690 -9823
rect 4610 -9880 4690 -9857
rect 4940 -9663 5020 -8950
rect 5048 -9091 5128 -9077
rect 5048 -9143 5062 -9091
rect 5114 -9105 5128 -9091
rect 5310 -9105 5390 -9090
rect 5114 -9113 5390 -9105
rect 5114 -9143 5333 -9113
rect 5048 -9145 5333 -9143
rect 5048 -9157 5128 -9145
rect 5310 -9147 5333 -9145
rect 5367 -9147 5390 -9113
rect 5310 -9170 5390 -9147
rect 5048 -9200 5128 -9186
rect 5048 -9252 5062 -9200
rect 5114 -9206 5128 -9200
rect 5114 -9246 5370 -9206
rect 5114 -9252 5128 -9246
rect 5048 -9266 5128 -9252
rect 5330 -9310 5370 -9246
rect 5310 -9333 5390 -9310
rect 5048 -9389 5128 -9366
rect 5048 -9423 5071 -9389
rect 5105 -9423 5128 -9389
rect 5310 -9367 5333 -9333
rect 5367 -9367 5390 -9333
rect 5310 -9390 5390 -9367
rect 5048 -9446 5128 -9423
rect 5310 -9446 5390 -9430
rect 5048 -9453 5390 -9446
rect 5048 -9486 5333 -9453
rect 5310 -9487 5333 -9486
rect 5367 -9487 5390 -9453
rect 5310 -9510 5390 -9487
rect 5580 -9630 5620 -8950
rect 5740 -9104 5820 -9090
rect 5740 -9156 5754 -9104
rect 5806 -9156 5820 -9104
rect 5740 -9170 5820 -9156
rect 5890 -9103 5970 -8950
rect 5890 -9137 5913 -9103
rect 5947 -9137 5970 -9103
rect 5890 -9183 5970 -9137
rect 5740 -9224 5820 -9210
rect 5740 -9276 5754 -9224
rect 5806 -9276 5820 -9224
rect 5740 -9290 5820 -9276
rect 5890 -9217 5913 -9183
rect 5947 -9217 5970 -9183
rect 5890 -9263 5970 -9217
rect 5890 -9297 5913 -9263
rect 5947 -9297 5970 -9263
rect 5890 -9320 5970 -9297
rect 6190 -9103 6270 -8950
rect 6190 -9137 6213 -9103
rect 6247 -9137 6270 -9103
rect 6190 -9183 6270 -9137
rect 6190 -9217 6213 -9183
rect 6247 -9217 6270 -9183
rect 6190 -9263 6270 -9217
rect 6190 -9297 6213 -9263
rect 6247 -9297 6270 -9263
rect 6190 -9320 6270 -9297
rect 6490 -9103 6570 -8950
rect 6490 -9137 6513 -9103
rect 6547 -9137 6570 -9103
rect 6490 -9183 6570 -9137
rect 6870 -9104 6950 -9090
rect 6870 -9156 6884 -9104
rect 6936 -9156 6950 -9104
rect 6870 -9170 6950 -9156
rect 6490 -9217 6513 -9183
rect 6547 -9217 6570 -9183
rect 6490 -9263 6570 -9217
rect 6490 -9297 6513 -9263
rect 6547 -9297 6570 -9263
rect 6720 -9224 6800 -9210
rect 6720 -9276 6734 -9224
rect 6786 -9276 6800 -9224
rect 6720 -9290 6800 -9276
rect 6490 -9320 6570 -9297
rect 6240 -9380 6320 -9360
rect 6640 -9380 6720 -9360
rect 6240 -9383 6720 -9380
rect 6240 -9417 6263 -9383
rect 6297 -9417 6663 -9383
rect 6697 -9417 6720 -9383
rect 6240 -9420 6720 -9417
rect 6240 -9440 6320 -9420
rect 6640 -9440 6720 -9420
rect 6990 -9630 7030 -8950
rect 7073 -9494 7153 -9480
rect 7073 -9546 7087 -9494
rect 7139 -9546 7153 -9494
rect 7073 -9560 7153 -9546
rect 4940 -9697 4963 -9663
rect 4997 -9697 5020 -9663
rect 4940 -9743 5020 -9697
rect 4940 -9777 4963 -9743
rect 4997 -9777 5020 -9743
rect 4940 -9823 5020 -9777
rect 4940 -9857 4963 -9823
rect 4997 -9857 5020 -9823
rect 4940 -9880 5020 -9857
rect 5560 -9663 5640 -9630
rect 5560 -9697 5583 -9663
rect 5617 -9697 5640 -9663
rect 5560 -9743 5640 -9697
rect 5560 -9777 5583 -9743
rect 5617 -9777 5640 -9743
rect 5560 -9823 5640 -9777
rect 5560 -9857 5583 -9823
rect 5617 -9857 5640 -9823
rect 5560 -9880 5640 -9857
rect 5890 -9663 5970 -9630
rect 5890 -9697 5913 -9663
rect 5947 -9697 5970 -9663
rect 5890 -9743 5970 -9697
rect 5890 -9777 5913 -9743
rect 5947 -9777 5970 -9743
rect 5890 -9823 5970 -9777
rect 5890 -9857 5913 -9823
rect 5947 -9857 5970 -9823
rect 5890 -9880 5970 -9857
rect 6190 -9663 6270 -9630
rect 6190 -9697 6213 -9663
rect 6247 -9697 6270 -9663
rect 6190 -9743 6270 -9697
rect 6190 -9777 6213 -9743
rect 6247 -9777 6270 -9743
rect 6190 -9823 6270 -9777
rect 6190 -9857 6213 -9823
rect 6247 -9857 6270 -9823
rect 6190 -9880 6270 -9857
rect 6490 -9663 6570 -9630
rect 6490 -9697 6513 -9663
rect 6547 -9697 6570 -9663
rect 6490 -9743 6570 -9697
rect 6490 -9777 6513 -9743
rect 6547 -9777 6570 -9743
rect 6490 -9823 6570 -9777
rect 6490 -9857 6513 -9823
rect 6547 -9857 6570 -9823
rect 6490 -9880 6570 -9857
rect 6970 -9663 7050 -9630
rect 6970 -9697 6993 -9663
rect 7027 -9697 7050 -9663
rect 6970 -9743 7050 -9697
rect 6970 -9777 6993 -9743
rect 7027 -9777 7050 -9743
rect 6970 -9814 7050 -9777
rect 6970 -9866 6984 -9814
rect 7036 -9866 7050 -9814
rect 6970 -9880 7050 -9866
rect 1171 -9934 1251 -9920
rect 1171 -9986 1185 -9934
rect 1237 -9986 1251 -9934
rect 1171 -10000 1251 -9986
rect 1840 -10030 1880 -9880
rect 2140 -10030 2180 -9880
rect 2440 -10030 2480 -9880
rect 4030 -10030 4070 -9880
rect 4330 -10030 4370 -9880
rect 4630 -10030 4670 -9880
rect 5398 -9934 5478 -9920
rect 5398 -9986 5412 -9934
rect 5464 -9986 5478 -9934
rect 5398 -10000 5478 -9986
rect 5910 -10030 5950 -9880
rect 6210 -10030 6250 -9880
rect 6510 -10030 6550 -9880
rect 912 -10097 935 -10063
rect 969 -10097 992 -10063
rect 912 -12883 992 -10097
rect 1020 -10063 7070 -10030
rect 1020 -10097 1103 -10063
rect 1137 -10097 1183 -10063
rect 1217 -10097 1263 -10063
rect 1297 -10097 1343 -10063
rect 1377 -10097 1423 -10063
rect 1457 -10097 1503 -10063
rect 1537 -10097 1583 -10063
rect 1617 -10097 1663 -10063
rect 1697 -10097 1743 -10063
rect 1777 -10097 1823 -10063
rect 1857 -10097 1903 -10063
rect 1937 -10097 1983 -10063
rect 2017 -10097 2063 -10063
rect 2097 -10097 2143 -10063
rect 2177 -10097 2223 -10063
rect 2257 -10097 2303 -10063
rect 2337 -10097 2383 -10063
rect 2417 -10097 2463 -10063
rect 2497 -10097 2543 -10063
rect 2577 -10097 2623 -10063
rect 2657 -10097 2703 -10063
rect 2737 -10097 2783 -10063
rect 2817 -10097 2863 -10063
rect 2897 -10097 2943 -10063
rect 2977 -10097 3023 -10063
rect 3057 -10097 3103 -10063
rect 3137 -10097 3183 -10063
rect 3217 -10097 3693 -10063
rect 3727 -10097 3773 -10063
rect 3807 -10097 3853 -10063
rect 3887 -10097 3933 -10063
rect 3967 -10097 4013 -10063
rect 4047 -10097 4093 -10063
rect 4127 -10097 4173 -10063
rect 4207 -10097 4253 -10063
rect 4287 -10097 4333 -10063
rect 4367 -10097 4413 -10063
rect 4447 -10097 4493 -10063
rect 4527 -10097 4573 -10063
rect 4607 -10097 4653 -10063
rect 4687 -10097 4733 -10063
rect 4767 -10097 4813 -10063
rect 4847 -10097 4893 -10063
rect 4927 -10097 4973 -10063
rect 5007 -10097 5413 -10063
rect 5447 -10097 5493 -10063
rect 5527 -10097 5573 -10063
rect 5607 -10097 5653 -10063
rect 5687 -10097 5733 -10063
rect 5767 -10097 5813 -10063
rect 5847 -10097 5893 -10063
rect 5927 -10097 5973 -10063
rect 6007 -10097 6053 -10063
rect 6087 -10097 6133 -10063
rect 6167 -10097 6213 -10063
rect 6247 -10097 6293 -10063
rect 6327 -10097 6373 -10063
rect 6407 -10097 6453 -10063
rect 6487 -10097 6533 -10063
rect 6567 -10097 6613 -10063
rect 6647 -10097 6693 -10063
rect 6727 -10097 6773 -10063
rect 6807 -10097 6853 -10063
rect 6887 -10097 6933 -10063
rect 6967 -10097 7013 -10063
rect 7047 -10097 7070 -10063
rect 1020 -10130 7070 -10097
rect 1171 -10174 1251 -10160
rect 1171 -10226 1185 -10174
rect 1237 -10226 1251 -10174
rect 1171 -10240 1251 -10226
rect 1840 -10280 1880 -10130
rect 2140 -10280 2180 -10130
rect 2440 -10280 2480 -10130
rect 4030 -10280 4070 -10130
rect 4330 -10280 4370 -10130
rect 4630 -10280 4670 -10130
rect 5398 -10173 5478 -10159
rect 5398 -10225 5412 -10173
rect 5464 -10225 5478 -10173
rect 5398 -10239 5478 -10225
rect 5910 -10280 5950 -10130
rect 6210 -10280 6250 -10130
rect 6510 -10280 6550 -10130
rect 1340 -10303 1420 -10280
rect 1340 -10337 1363 -10303
rect 1397 -10337 1420 -10303
rect 1340 -10383 1420 -10337
rect 1340 -10417 1363 -10383
rect 1397 -10417 1420 -10383
rect 1340 -10463 1420 -10417
rect 1340 -10497 1363 -10463
rect 1397 -10497 1420 -10463
rect 1340 -10530 1420 -10497
rect 1820 -10303 1900 -10280
rect 1820 -10337 1843 -10303
rect 1877 -10337 1900 -10303
rect 1820 -10383 1900 -10337
rect 1820 -10417 1843 -10383
rect 1877 -10417 1900 -10383
rect 1820 -10463 1900 -10417
rect 1820 -10497 1843 -10463
rect 1877 -10497 1900 -10463
rect 1820 -10530 1900 -10497
rect 2120 -10303 2200 -10280
rect 2120 -10337 2143 -10303
rect 2177 -10337 2200 -10303
rect 2120 -10383 2200 -10337
rect 2120 -10417 2143 -10383
rect 2177 -10417 2200 -10383
rect 2120 -10463 2200 -10417
rect 2120 -10497 2143 -10463
rect 2177 -10497 2200 -10463
rect 2120 -10530 2200 -10497
rect 2420 -10303 2500 -10280
rect 2420 -10337 2443 -10303
rect 2477 -10337 2500 -10303
rect 2420 -10383 2500 -10337
rect 2420 -10417 2443 -10383
rect 2477 -10417 2500 -10383
rect 2420 -10463 2500 -10417
rect 2420 -10497 2443 -10463
rect 2477 -10497 2500 -10463
rect 2420 -10530 2500 -10497
rect 2900 -10303 2980 -10280
rect 2900 -10337 2923 -10303
rect 2957 -10337 2980 -10303
rect 2900 -10383 2980 -10337
rect 2900 -10417 2923 -10383
rect 2957 -10417 2980 -10383
rect 3680 -10303 3760 -10280
rect 3680 -10337 3703 -10303
rect 3737 -10337 3760 -10303
rect 3680 -10383 3760 -10337
rect 2900 -10463 2980 -10417
rect 2900 -10497 2923 -10463
rect 2957 -10497 2980 -10463
rect 3314 -10397 3394 -10384
rect 3314 -10449 3328 -10397
rect 3380 -10449 3394 -10397
rect 3314 -10464 3394 -10449
rect 3680 -10417 3703 -10383
rect 3737 -10417 3760 -10383
rect 3680 -10463 3760 -10417
rect 2900 -10530 2980 -10497
rect 3680 -10497 3703 -10463
rect 3737 -10497 3760 -10463
rect 1360 -11210 1400 -10530
rect 2540 -10720 2620 -10710
rect 2170 -10733 2620 -10720
rect 2170 -10743 2563 -10733
rect 2170 -10777 2193 -10743
rect 2227 -10760 2563 -10743
rect 2227 -10777 2250 -10760
rect 1670 -10804 1750 -10790
rect 2170 -10800 2250 -10777
rect 2540 -10767 2563 -10760
rect 2597 -10767 2620 -10733
rect 2540 -10790 2620 -10767
rect 1670 -10856 1684 -10804
rect 1736 -10856 1750 -10804
rect 2700 -10804 2780 -10790
rect 1670 -10870 1750 -10856
rect 1820 -10863 1900 -10840
rect 1540 -10904 1620 -10890
rect 1540 -10956 1554 -10904
rect 1606 -10956 1620 -10904
rect 1540 -10970 1620 -10956
rect 1820 -10897 1843 -10863
rect 1877 -10897 1900 -10863
rect 1820 -10943 1900 -10897
rect 1820 -10977 1843 -10943
rect 1877 -10977 1900 -10943
rect 1670 -11004 1750 -10990
rect 1670 -11056 1684 -11004
rect 1736 -11056 1750 -11004
rect 1670 -11070 1750 -11056
rect 1820 -11023 1900 -10977
rect 1820 -11057 1843 -11023
rect 1877 -11057 1900 -11023
rect 1540 -11104 1620 -11090
rect 1540 -11156 1554 -11104
rect 1606 -11156 1620 -11104
rect 1540 -11170 1620 -11156
rect 1820 -11210 1900 -11057
rect 2120 -10863 2200 -10840
rect 2120 -10897 2143 -10863
rect 2177 -10897 2200 -10863
rect 2120 -10943 2200 -10897
rect 2120 -10977 2143 -10943
rect 2177 -10977 2200 -10943
rect 2120 -11023 2200 -10977
rect 2120 -11057 2143 -11023
rect 2177 -11057 2200 -11023
rect 2120 -11210 2200 -11057
rect 2420 -10863 2500 -10840
rect 2420 -10897 2443 -10863
rect 2477 -10897 2500 -10863
rect 2700 -10856 2714 -10804
rect 2766 -10856 2780 -10804
rect 2700 -10870 2780 -10856
rect 2420 -10943 2500 -10897
rect 2420 -10977 2443 -10943
rect 2477 -10977 2500 -10943
rect 2420 -11023 2500 -10977
rect 2420 -11057 2443 -11023
rect 2477 -11057 2500 -11023
rect 2420 -11210 2500 -11057
rect 2800 -11104 2880 -11090
rect 2800 -11156 2814 -11104
rect 2866 -11156 2880 -11104
rect 2800 -11170 2880 -11156
rect 2920 -11210 2960 -10530
rect 3300 -10733 3631 -10710
rect 3300 -10767 3323 -10733
rect 3357 -10750 3631 -10733
rect 3357 -10767 3380 -10750
rect 3300 -10790 3380 -10767
rect 3150 -10904 3230 -10890
rect 3150 -10956 3164 -10904
rect 3216 -10956 3230 -10904
rect 3591 -10911 3631 -10750
rect 3150 -10970 3230 -10956
rect 3572 -10925 3652 -10911
rect 3572 -10977 3586 -10925
rect 3638 -10977 3652 -10925
rect 3000 -11004 3080 -10990
rect 3572 -10991 3652 -10977
rect 3000 -11056 3014 -11004
rect 3066 -11056 3080 -11004
rect 3000 -11070 3080 -11056
rect 3572 -11038 3652 -11024
rect 3572 -11090 3586 -11038
rect 3638 -11090 3652 -11038
rect 3572 -11104 3652 -11090
rect 3680 -11210 3760 -10497
rect 4010 -10303 4090 -10280
rect 4010 -10337 4033 -10303
rect 4067 -10337 4090 -10303
rect 4010 -10383 4090 -10337
rect 4010 -10417 4033 -10383
rect 4067 -10417 4090 -10383
rect 4010 -10463 4090 -10417
rect 4010 -10497 4033 -10463
rect 4067 -10497 4090 -10463
rect 4010 -10530 4090 -10497
rect 4310 -10303 4390 -10280
rect 4310 -10337 4333 -10303
rect 4367 -10337 4390 -10303
rect 4310 -10383 4390 -10337
rect 4310 -10417 4333 -10383
rect 4367 -10417 4390 -10383
rect 4310 -10463 4390 -10417
rect 4310 -10497 4333 -10463
rect 4367 -10497 4390 -10463
rect 4310 -10530 4390 -10497
rect 4610 -10303 4690 -10280
rect 4610 -10337 4633 -10303
rect 4667 -10337 4690 -10303
rect 4610 -10383 4690 -10337
rect 4610 -10417 4633 -10383
rect 4667 -10417 4690 -10383
rect 4610 -10463 4690 -10417
rect 4610 -10497 4633 -10463
rect 4667 -10497 4690 -10463
rect 4610 -10530 4690 -10497
rect 4940 -10303 5020 -10280
rect 4940 -10337 4963 -10303
rect 4997 -10337 5020 -10303
rect 4940 -10383 5020 -10337
rect 4940 -10417 4963 -10383
rect 4997 -10417 5020 -10383
rect 4940 -10463 5020 -10417
rect 4940 -10497 4963 -10463
rect 4997 -10497 5020 -10463
rect 4360 -10740 4440 -10720
rect 4760 -10740 4840 -10720
rect 4360 -10743 4840 -10740
rect 4360 -10777 4383 -10743
rect 4417 -10777 4783 -10743
rect 4817 -10777 4840 -10743
rect 4360 -10780 4840 -10777
rect 4360 -10800 4440 -10780
rect 4760 -10800 4840 -10780
rect 3860 -10854 3940 -10840
rect 3860 -10906 3874 -10854
rect 3926 -10906 3940 -10854
rect 3860 -10920 3940 -10906
rect 4010 -10863 4090 -10840
rect 4010 -10897 4033 -10863
rect 4067 -10897 4090 -10863
rect 3880 -11092 3920 -10920
rect 4010 -10943 4090 -10897
rect 4010 -10977 4033 -10943
rect 4067 -10977 4090 -10943
rect 4010 -11023 4090 -10977
rect 4010 -11057 4033 -11023
rect 4067 -11057 4090 -11023
rect 3860 -11105 3940 -11092
rect 3860 -11157 3874 -11105
rect 3926 -11157 3940 -11105
rect 3860 -11172 3940 -11157
rect 4010 -11210 4090 -11057
rect 4310 -10863 4390 -10840
rect 4310 -10897 4333 -10863
rect 4367 -10897 4390 -10863
rect 4310 -10943 4390 -10897
rect 4310 -10977 4333 -10943
rect 4367 -10977 4390 -10943
rect 4310 -11023 4390 -10977
rect 4310 -11057 4333 -11023
rect 4367 -11057 4390 -11023
rect 4310 -11210 4390 -11057
rect 4610 -10863 4690 -10840
rect 4610 -10897 4633 -10863
rect 4667 -10897 4690 -10863
rect 4610 -10943 4690 -10897
rect 4760 -10854 4840 -10840
rect 4760 -10906 4774 -10854
rect 4826 -10906 4840 -10854
rect 4760 -10920 4840 -10906
rect 4610 -10977 4633 -10943
rect 4667 -10977 4690 -10943
rect 4610 -11023 4690 -10977
rect 4610 -11057 4633 -11023
rect 4667 -11057 4690 -11023
rect 4610 -11210 4690 -11057
rect 4940 -11210 5020 -10497
rect 5560 -10303 5640 -10280
rect 5560 -10337 5583 -10303
rect 5617 -10337 5640 -10303
rect 5560 -10383 5640 -10337
rect 5560 -10417 5583 -10383
rect 5617 -10417 5640 -10383
rect 5560 -10463 5640 -10417
rect 5560 -10497 5583 -10463
rect 5617 -10497 5640 -10463
rect 5560 -10530 5640 -10497
rect 5890 -10303 5970 -10280
rect 5890 -10337 5913 -10303
rect 5947 -10337 5970 -10303
rect 5890 -10383 5970 -10337
rect 5890 -10417 5913 -10383
rect 5947 -10417 5970 -10383
rect 5890 -10463 5970 -10417
rect 5890 -10497 5913 -10463
rect 5947 -10497 5970 -10463
rect 5890 -10530 5970 -10497
rect 6190 -10303 6270 -10280
rect 6190 -10337 6213 -10303
rect 6247 -10337 6270 -10303
rect 6190 -10383 6270 -10337
rect 6190 -10417 6213 -10383
rect 6247 -10417 6270 -10383
rect 6190 -10463 6270 -10417
rect 6190 -10497 6213 -10463
rect 6247 -10497 6270 -10463
rect 6190 -10530 6270 -10497
rect 6490 -10303 6570 -10280
rect 6490 -10337 6513 -10303
rect 6547 -10337 6570 -10303
rect 6490 -10383 6570 -10337
rect 6490 -10417 6513 -10383
rect 6547 -10417 6570 -10383
rect 6490 -10463 6570 -10417
rect 6490 -10497 6513 -10463
rect 6547 -10497 6570 -10463
rect 6490 -10530 6570 -10497
rect 6970 -10294 7050 -10280
rect 6970 -10346 6984 -10294
rect 7036 -10346 7050 -10294
rect 6970 -10383 7050 -10346
rect 6970 -10417 6993 -10383
rect 7027 -10417 7050 -10383
rect 6970 -10463 7050 -10417
rect 6970 -10497 6993 -10463
rect 7027 -10497 7050 -10463
rect 6970 -10530 7050 -10497
rect 5048 -10570 5128 -10550
rect 5048 -10573 5370 -10570
rect 5048 -10607 5071 -10573
rect 5105 -10607 5370 -10573
rect 5048 -10610 5370 -10607
rect 5048 -10630 5128 -10610
rect 5330 -10870 5370 -10610
rect 5048 -10892 5128 -10878
rect 5048 -10944 5062 -10892
rect 5114 -10944 5128 -10892
rect 5048 -10958 5128 -10944
rect 5310 -10893 5390 -10870
rect 5310 -10927 5333 -10893
rect 5367 -10927 5390 -10893
rect 5310 -10950 5390 -10927
rect 5048 -11000 5128 -10986
rect 5048 -11052 5062 -11000
rect 5114 -11005 5128 -11000
rect 5310 -11005 5390 -10991
rect 5114 -11014 5390 -11005
rect 5114 -11045 5333 -11014
rect 5114 -11052 5128 -11045
rect 5048 -11066 5128 -11052
rect 5310 -11048 5333 -11045
rect 5367 -11048 5390 -11014
rect 5310 -11071 5390 -11048
rect 5580 -11210 5620 -10530
rect 6240 -10740 6320 -10720
rect 6640 -10740 6720 -10720
rect 6240 -10743 6720 -10740
rect 6240 -10777 6263 -10743
rect 6297 -10777 6663 -10743
rect 6697 -10777 6720 -10743
rect 6240 -10780 6720 -10777
rect 6240 -10800 6320 -10780
rect 6640 -10800 6720 -10780
rect 5890 -10863 5970 -10840
rect 5740 -10884 5820 -10870
rect 5740 -10936 5754 -10884
rect 5806 -10936 5820 -10884
rect 5740 -10950 5820 -10936
rect 5890 -10897 5913 -10863
rect 5947 -10897 5970 -10863
rect 5890 -10943 5970 -10897
rect 5890 -10977 5913 -10943
rect 5947 -10977 5970 -10943
rect 5740 -11004 5820 -10990
rect 5740 -11056 5754 -11004
rect 5806 -11056 5820 -11004
rect 5740 -11070 5820 -11056
rect 5890 -11023 5970 -10977
rect 5890 -11057 5913 -11023
rect 5947 -11057 5970 -11023
rect 5890 -11210 5970 -11057
rect 6190 -10863 6270 -10840
rect 6190 -10897 6213 -10863
rect 6247 -10897 6270 -10863
rect 6190 -10943 6270 -10897
rect 6190 -10977 6213 -10943
rect 6247 -10977 6270 -10943
rect 6190 -11023 6270 -10977
rect 6190 -11057 6213 -11023
rect 6247 -11057 6270 -11023
rect 6190 -11210 6270 -11057
rect 6490 -10863 6570 -10840
rect 6490 -10897 6513 -10863
rect 6547 -10897 6570 -10863
rect 6490 -10943 6570 -10897
rect 6490 -10977 6513 -10943
rect 6547 -10977 6570 -10943
rect 6720 -10884 6800 -10870
rect 6720 -10936 6734 -10884
rect 6786 -10936 6800 -10884
rect 6720 -10950 6800 -10936
rect 6490 -11023 6570 -10977
rect 6490 -11057 6513 -11023
rect 6547 -11057 6570 -11023
rect 6490 -11210 6570 -11057
rect 6870 -11004 6950 -10990
rect 6870 -11056 6884 -11004
rect 6936 -11056 6950 -11004
rect 6870 -11070 6950 -11056
rect 6990 -11210 7030 -10530
rect 7073 -10614 7153 -10600
rect 7073 -10666 7087 -10614
rect 7139 -10666 7153 -10614
rect 7073 -10680 7153 -10666
rect 1020 -11234 5040 -11210
rect 1020 -11286 1069 -11234
rect 1121 -11243 5040 -11234
rect 1137 -11277 1183 -11243
rect 1217 -11277 1263 -11243
rect 1297 -11277 1343 -11243
rect 1377 -11277 1423 -11243
rect 1457 -11277 1503 -11243
rect 1537 -11277 1583 -11243
rect 1617 -11277 1663 -11243
rect 1697 -11277 1743 -11243
rect 1777 -11277 1823 -11243
rect 1857 -11277 1903 -11243
rect 1937 -11277 1983 -11243
rect 2017 -11277 2063 -11243
rect 2097 -11277 2143 -11243
rect 2177 -11277 2223 -11243
rect 2257 -11277 2303 -11243
rect 2337 -11277 2383 -11243
rect 2417 -11277 2463 -11243
rect 2497 -11277 2543 -11243
rect 2577 -11277 2623 -11243
rect 2657 -11277 2703 -11243
rect 2737 -11277 2783 -11243
rect 2817 -11277 2863 -11243
rect 2897 -11277 2943 -11243
rect 2977 -11277 3023 -11243
rect 3057 -11277 3103 -11243
rect 3137 -11277 3183 -11243
rect 3217 -11277 3693 -11243
rect 3727 -11277 3773 -11243
rect 3807 -11277 3853 -11243
rect 3887 -11277 3933 -11243
rect 3967 -11277 4013 -11243
rect 4047 -11277 4093 -11243
rect 4127 -11277 4173 -11243
rect 4207 -11277 4253 -11243
rect 4287 -11277 4333 -11243
rect 4367 -11277 4413 -11243
rect 4447 -11277 4493 -11243
rect 4527 -11277 4573 -11243
rect 4607 -11277 4653 -11243
rect 4687 -11277 4733 -11243
rect 4767 -11277 4813 -11243
rect 4847 -11277 4893 -11243
rect 4927 -11277 4973 -11243
rect 5007 -11277 5040 -11243
rect 1121 -11286 5040 -11277
rect 1020 -11310 5040 -11286
rect 5170 -11243 7070 -11210
rect 5170 -11277 5413 -11243
rect 5447 -11277 5493 -11243
rect 5527 -11277 5573 -11243
rect 5607 -11277 5653 -11243
rect 5687 -11277 5733 -11243
rect 5767 -11277 5813 -11243
rect 5847 -11277 5893 -11243
rect 5927 -11277 5973 -11243
rect 6007 -11277 6053 -11243
rect 6087 -11277 6133 -11243
rect 6167 -11277 6213 -11243
rect 6247 -11277 6293 -11243
rect 6327 -11277 6373 -11243
rect 6407 -11277 6453 -11243
rect 6487 -11277 6533 -11243
rect 6567 -11277 6613 -11243
rect 6647 -11277 6693 -11243
rect 6727 -11277 6773 -11243
rect 6807 -11277 6853 -11243
rect 6887 -11277 6933 -11243
rect 6967 -11277 7013 -11243
rect 7047 -11277 7070 -11243
rect 5170 -11310 7070 -11277
rect 5170 -11440 5270 -11310
rect 4801 -11540 5270 -11440
rect 5398 -11468 5478 -11454
rect 5398 -11520 5412 -11468
rect 5464 -11520 5478 -11468
rect 5398 -11534 5478 -11520
rect 7343 -11501 7423 -11487
rect 4801 -11670 4901 -11540
rect 7343 -11553 7357 -11501
rect 7409 -11553 7423 -11501
rect 7343 -11567 7423 -11553
rect 1055 -11695 3161 -11670
rect 1055 -11747 1069 -11695
rect 1121 -11703 3161 -11695
rect 1121 -11737 1184 -11703
rect 1218 -11737 1264 -11703
rect 1298 -11737 1344 -11703
rect 1378 -11737 1424 -11703
rect 1458 -11737 1504 -11703
rect 1538 -11737 1584 -11703
rect 1618 -11737 1664 -11703
rect 1698 -11737 1744 -11703
rect 1778 -11737 1824 -11703
rect 1858 -11737 1904 -11703
rect 1938 -11737 1984 -11703
rect 2018 -11737 2064 -11703
rect 2098 -11737 2144 -11703
rect 2178 -11737 2224 -11703
rect 2258 -11737 2304 -11703
rect 2338 -11737 2384 -11703
rect 2418 -11737 2464 -11703
rect 2498 -11737 2544 -11703
rect 2578 -11737 2624 -11703
rect 2658 -11737 2704 -11703
rect 2738 -11737 2784 -11703
rect 2818 -11737 2864 -11703
rect 2898 -11737 2944 -11703
rect 2978 -11737 3024 -11703
rect 3058 -11737 3104 -11703
rect 3138 -11737 3161 -11703
rect 1121 -11747 3161 -11737
rect 1055 -11770 3161 -11747
rect 3521 -11703 4901 -11670
rect 3521 -11737 3554 -11703
rect 3588 -11737 3634 -11703
rect 3668 -11737 3714 -11703
rect 3748 -11737 3794 -11703
rect 3828 -11737 3874 -11703
rect 3908 -11737 3954 -11703
rect 3988 -11737 4034 -11703
rect 4068 -11737 4114 -11703
rect 4148 -11737 4194 -11703
rect 4228 -11737 4274 -11703
rect 4308 -11737 4354 -11703
rect 4388 -11737 4434 -11703
rect 4468 -11737 4514 -11703
rect 4548 -11737 4594 -11703
rect 4628 -11737 4674 -11703
rect 4708 -11737 4754 -11703
rect 4788 -11737 4834 -11703
rect 4868 -11737 4901 -11703
rect 3521 -11770 4901 -11737
rect 5251 -11695 7251 -11671
rect 5251 -11747 5265 -11695
rect 5317 -11704 7251 -11695
rect 5317 -11738 5354 -11704
rect 5388 -11738 5434 -11704
rect 5468 -11738 5514 -11704
rect 5548 -11738 5594 -11704
rect 5628 -11738 5674 -11704
rect 5708 -11738 5754 -11704
rect 5788 -11738 5834 -11704
rect 5868 -11738 5914 -11704
rect 5948 -11738 5994 -11704
rect 6028 -11738 6074 -11704
rect 6108 -11738 6154 -11704
rect 6188 -11738 6234 -11704
rect 6268 -11738 6314 -11704
rect 6348 -11738 6394 -11704
rect 6428 -11738 6474 -11704
rect 6508 -11738 6554 -11704
rect 6588 -11738 6634 -11704
rect 6668 -11738 6714 -11704
rect 6748 -11738 6794 -11704
rect 6828 -11738 6874 -11704
rect 6908 -11738 6954 -11704
rect 6988 -11738 7034 -11704
rect 7068 -11738 7114 -11704
rect 7148 -11738 7194 -11704
rect 7228 -11738 7251 -11704
rect 5317 -11747 7251 -11738
rect 1211 -12450 1251 -11770
rect 1511 -12450 1551 -11770
rect 1581 -11814 1661 -11800
rect 1581 -11866 1595 -11814
rect 1647 -11866 1661 -11814
rect 1581 -11880 1661 -11866
rect 1671 -11934 1751 -11920
rect 1671 -11986 1685 -11934
rect 1737 -11986 1751 -11934
rect 1671 -12000 1751 -11986
rect 1821 -11923 1901 -11770
rect 1821 -11957 1844 -11923
rect 1878 -11957 1901 -11923
rect 1821 -12003 1901 -11957
rect 1821 -12037 1844 -12003
rect 1878 -12037 1901 -12003
rect 1641 -12054 1721 -12040
rect 1641 -12106 1655 -12054
rect 1707 -12106 1721 -12054
rect 1641 -12120 1721 -12106
rect 1821 -12083 1901 -12037
rect 1821 -12117 1844 -12083
rect 1878 -12117 1901 -12083
rect 1821 -12140 1901 -12117
rect 2121 -11923 2201 -11770
rect 2121 -11957 2144 -11923
rect 2178 -11957 2201 -11923
rect 2121 -12003 2201 -11957
rect 2121 -12037 2144 -12003
rect 2178 -12037 2201 -12003
rect 2121 -12083 2201 -12037
rect 2121 -12117 2144 -12083
rect 2178 -12117 2201 -12083
rect 2121 -12140 2201 -12117
rect 2421 -11923 2501 -11770
rect 2951 -11814 3031 -11800
rect 2951 -11866 2965 -11814
rect 3017 -11866 3031 -11814
rect 2951 -11880 3031 -11866
rect 2421 -11957 2444 -11923
rect 2478 -11957 2501 -11923
rect 2421 -12003 2501 -11957
rect 2801 -11934 2881 -11920
rect 2801 -11986 2815 -11934
rect 2867 -11986 2881 -11934
rect 2801 -12000 2881 -11986
rect 2421 -12037 2444 -12003
rect 2478 -12037 2501 -12003
rect 2421 -12083 2501 -12037
rect 2421 -12117 2444 -12083
rect 2478 -12117 2501 -12083
rect 2421 -12140 2501 -12117
rect 2671 -12054 2751 -12040
rect 2671 -12106 2685 -12054
rect 2737 -12106 2751 -12054
rect 2671 -12120 2751 -12106
rect 2171 -12200 2251 -12180
rect 2571 -12200 2651 -12180
rect 2171 -12203 2651 -12200
rect 2171 -12237 2194 -12203
rect 2228 -12237 2594 -12203
rect 2628 -12237 2651 -12203
rect 2171 -12240 2651 -12237
rect 2171 -12260 2251 -12240
rect 2571 -12260 2651 -12240
rect 3071 -12450 3111 -11770
rect 3433 -12080 3513 -12060
rect 3172 -12083 3513 -12080
rect 3172 -12117 3456 -12083
rect 3490 -12117 3513 -12083
rect 3172 -12120 3513 -12117
rect 3172 -12299 3212 -12120
rect 3433 -12140 3513 -12120
rect 3151 -12322 3231 -12299
rect 3151 -12356 3174 -12322
rect 3208 -12356 3231 -12322
rect 3151 -12379 3231 -12356
rect 1191 -12483 1271 -12450
rect 1191 -12517 1214 -12483
rect 1248 -12517 1271 -12483
rect 1191 -12563 1271 -12517
rect 1191 -12597 1214 -12563
rect 1248 -12597 1271 -12563
rect 1191 -12643 1271 -12597
rect 1191 -12677 1214 -12643
rect 1248 -12677 1271 -12643
rect 1191 -12700 1271 -12677
rect 1491 -12483 1571 -12450
rect 1491 -12517 1514 -12483
rect 1548 -12517 1571 -12483
rect 1491 -12563 1571 -12517
rect 1491 -12597 1514 -12563
rect 1548 -12597 1571 -12563
rect 1491 -12643 1571 -12597
rect 1491 -12677 1514 -12643
rect 1548 -12677 1571 -12643
rect 1491 -12700 1571 -12677
rect 1821 -12483 1901 -12450
rect 1821 -12517 1844 -12483
rect 1878 -12517 1901 -12483
rect 1821 -12563 1901 -12517
rect 1821 -12597 1844 -12563
rect 1878 -12597 1901 -12563
rect 1821 -12643 1901 -12597
rect 1821 -12677 1844 -12643
rect 1878 -12677 1901 -12643
rect 1821 -12700 1901 -12677
rect 2121 -12483 2201 -12450
rect 2121 -12517 2144 -12483
rect 2178 -12517 2201 -12483
rect 2121 -12563 2201 -12517
rect 2121 -12597 2144 -12563
rect 2178 -12597 2201 -12563
rect 2121 -12643 2201 -12597
rect 2121 -12677 2144 -12643
rect 2178 -12677 2201 -12643
rect 2121 -12700 2201 -12677
rect 2421 -12483 2501 -12450
rect 2421 -12517 2444 -12483
rect 2478 -12517 2501 -12483
rect 2421 -12563 2501 -12517
rect 2421 -12597 2444 -12563
rect 2478 -12597 2501 -12563
rect 2421 -12643 2501 -12597
rect 2421 -12677 2444 -12643
rect 2478 -12677 2501 -12643
rect 2421 -12700 2501 -12677
rect 3051 -12483 3131 -12450
rect 3051 -12517 3074 -12483
rect 3108 -12517 3131 -12483
rect 3051 -12563 3131 -12517
rect 3051 -12597 3074 -12563
rect 3108 -12597 3131 -12563
rect 3051 -12643 3131 -12597
rect 3051 -12677 3074 -12643
rect 3108 -12677 3131 -12643
rect 3051 -12700 3131 -12677
rect 3541 -12483 3621 -11770
rect 3871 -11923 3951 -11770
rect 3871 -11957 3894 -11923
rect 3928 -11957 3951 -11923
rect 3871 -12003 3951 -11957
rect 3871 -12037 3894 -12003
rect 3928 -12037 3951 -12003
rect 3721 -12074 3801 -12060
rect 3721 -12126 3735 -12074
rect 3787 -12126 3801 -12074
rect 3721 -12140 3801 -12126
rect 3871 -12083 3951 -12037
rect 3871 -12117 3894 -12083
rect 3928 -12117 3951 -12083
rect 3871 -12140 3951 -12117
rect 4171 -11923 4251 -11770
rect 4171 -11957 4194 -11923
rect 4228 -11957 4251 -11923
rect 4171 -12003 4251 -11957
rect 4171 -12037 4194 -12003
rect 4228 -12037 4251 -12003
rect 4171 -12083 4251 -12037
rect 4171 -12117 4194 -12083
rect 4228 -12117 4251 -12083
rect 4171 -12140 4251 -12117
rect 4471 -11923 4551 -11770
rect 4471 -11957 4494 -11923
rect 4528 -11957 4551 -11923
rect 4471 -12003 4551 -11957
rect 4471 -12037 4494 -12003
rect 4528 -12037 4551 -12003
rect 4471 -12083 4551 -12037
rect 4471 -12117 4494 -12083
rect 4528 -12117 4551 -12083
rect 4471 -12140 4551 -12117
rect 4621 -12074 4701 -12060
rect 4621 -12126 4635 -12074
rect 4687 -12126 4701 -12074
rect 4621 -12140 4701 -12126
rect 4221 -12200 4301 -12180
rect 4621 -12200 4701 -12180
rect 4221 -12203 4701 -12200
rect 4221 -12237 4244 -12203
rect 4278 -12237 4644 -12203
rect 4678 -12237 4701 -12203
rect 4221 -12240 4701 -12237
rect 4221 -12260 4301 -12240
rect 4621 -12260 4701 -12240
rect 3541 -12517 3564 -12483
rect 3598 -12517 3621 -12483
rect 3541 -12563 3621 -12517
rect 3541 -12597 3564 -12563
rect 3598 -12597 3621 -12563
rect 3541 -12643 3621 -12597
rect 3541 -12677 3564 -12643
rect 3598 -12677 3621 -12643
rect 3541 -12700 3621 -12677
rect 3871 -12483 3951 -12450
rect 3871 -12517 3894 -12483
rect 3928 -12517 3951 -12483
rect 3871 -12563 3951 -12517
rect 3871 -12597 3894 -12563
rect 3928 -12597 3951 -12563
rect 3871 -12643 3951 -12597
rect 3871 -12677 3894 -12643
rect 3928 -12677 3951 -12643
rect 3871 -12700 3951 -12677
rect 4171 -12483 4251 -12450
rect 4171 -12517 4194 -12483
rect 4228 -12517 4251 -12483
rect 4171 -12563 4251 -12517
rect 4171 -12597 4194 -12563
rect 4228 -12597 4251 -12563
rect 4171 -12643 4251 -12597
rect 4171 -12677 4194 -12643
rect 4228 -12677 4251 -12643
rect 4171 -12700 4251 -12677
rect 4471 -12483 4551 -12450
rect 4471 -12517 4494 -12483
rect 4528 -12517 4551 -12483
rect 4471 -12563 4551 -12517
rect 4471 -12597 4494 -12563
rect 4528 -12597 4551 -12563
rect 4471 -12643 4551 -12597
rect 4471 -12677 4494 -12643
rect 4528 -12677 4551 -12643
rect 4471 -12700 4551 -12677
rect 4801 -12483 4881 -11770
rect 5251 -11771 7251 -11747
rect 5004 -11901 5084 -11887
rect 5004 -11953 5018 -11901
rect 5070 -11953 5084 -11901
rect 5004 -11967 5084 -11953
rect 5180 -11987 5260 -11973
rect 5180 -11995 5194 -11987
rect 4935 -12035 5194 -11995
rect 4935 -12350 4975 -12035
rect 5180 -12039 5194 -12035
rect 5246 -12039 5260 -11987
rect 5180 -12053 5260 -12039
rect 5180 -12097 5260 -12083
rect 5180 -12149 5194 -12097
rect 5246 -12149 5260 -12097
rect 5180 -12163 5260 -12149
rect 5181 -12211 5261 -12197
rect 5181 -12263 5195 -12211
rect 5247 -12263 5261 -12211
rect 5181 -12277 5261 -12263
rect 5181 -12325 5261 -12311
rect 4915 -12373 4995 -12350
rect 4915 -12407 4938 -12373
rect 4972 -12407 4995 -12373
rect 5181 -12377 5195 -12325
rect 5247 -12377 5261 -12325
rect 5181 -12391 5261 -12377
rect 4915 -12430 4995 -12407
rect 5301 -12451 5341 -11771
rect 5381 -11820 5461 -11806
rect 5381 -11872 5395 -11820
rect 5447 -11872 5461 -11820
rect 5381 -11886 5461 -11872
rect 5481 -11945 5561 -11931
rect 5481 -11997 5495 -11945
rect 5547 -11997 5561 -11945
rect 5481 -12011 5561 -11997
rect 5601 -12451 5641 -11771
rect 5911 -11924 5991 -11771
rect 5911 -11958 5934 -11924
rect 5968 -11958 5991 -11924
rect 5911 -12004 5991 -11958
rect 5681 -12035 5761 -12021
rect 5681 -12087 5695 -12035
rect 5747 -12087 5761 -12035
rect 5681 -12101 5761 -12087
rect 5911 -12038 5934 -12004
rect 5968 -12038 5991 -12004
rect 5911 -12084 5991 -12038
rect 5911 -12118 5934 -12084
rect 5968 -12118 5991 -12084
rect 5911 -12141 5991 -12118
rect 6211 -11924 6291 -11771
rect 6211 -11958 6234 -11924
rect 6268 -11958 6291 -11924
rect 6211 -12004 6291 -11958
rect 6211 -12038 6234 -12004
rect 6268 -12038 6291 -12004
rect 6211 -12084 6291 -12038
rect 6211 -12118 6234 -12084
rect 6268 -12118 6291 -12084
rect 6211 -12141 6291 -12118
rect 6511 -11924 6591 -11771
rect 6661 -11825 6741 -11811
rect 6661 -11877 6675 -11825
rect 6727 -11877 6741 -11825
rect 6661 -11891 6741 -11877
rect 6511 -11958 6534 -11924
rect 6568 -11958 6591 -11924
rect 6511 -12004 6591 -11958
rect 6781 -11935 6861 -11921
rect 6781 -11987 6795 -11935
rect 6847 -11987 6861 -11935
rect 6781 -12001 6861 -11987
rect 7033 -11935 7113 -11921
rect 7033 -11987 7047 -11935
rect 7099 -11987 7113 -11935
rect 7033 -12001 7113 -11987
rect 6511 -12038 6534 -12004
rect 6568 -12038 6591 -12004
rect 6511 -12084 6591 -12038
rect 6511 -12118 6534 -12084
rect 6568 -12118 6591 -12084
rect 6661 -12035 6741 -12021
rect 6661 -12087 6675 -12035
rect 6727 -12087 6741 -12035
rect 6661 -12101 6741 -12087
rect 6511 -12141 6591 -12118
rect 6791 -12123 6871 -12109
rect 6791 -12175 6805 -12123
rect 6857 -12175 6871 -12123
rect 5761 -12201 5841 -12181
rect 6161 -12201 6241 -12181
rect 6791 -12189 6871 -12175
rect 5761 -12204 6241 -12201
rect 5761 -12238 5784 -12204
rect 5818 -12238 6184 -12204
rect 6218 -12238 6241 -12204
rect 5761 -12241 6241 -12238
rect 5761 -12261 5841 -12241
rect 6161 -12261 6241 -12241
rect 6811 -12311 6851 -12189
rect 6791 -12334 6871 -12311
rect 6791 -12368 6814 -12334
rect 6848 -12368 6871 -12334
rect 6791 -12391 6871 -12368
rect 7161 -12451 7201 -11771
rect 7229 -11825 7309 -11811
rect 7229 -11877 7243 -11825
rect 7295 -11877 7309 -11825
rect 7229 -11891 7309 -11877
rect 7275 -12123 7355 -12109
rect 7275 -12175 7289 -12123
rect 7341 -12175 7355 -12123
rect 7275 -12189 7355 -12175
rect 4801 -12517 4824 -12483
rect 4858 -12517 4881 -12483
rect 4801 -12563 4881 -12517
rect 4998 -12478 5078 -12464
rect 4998 -12530 5012 -12478
rect 5064 -12530 5078 -12478
rect 4998 -12544 5078 -12530
rect 5281 -12484 5361 -12451
rect 5281 -12518 5304 -12484
rect 5338 -12518 5361 -12484
rect 4801 -12597 4824 -12563
rect 4858 -12597 4881 -12563
rect 4801 -12643 4881 -12597
rect 4801 -12677 4824 -12643
rect 4858 -12677 4881 -12643
rect 4801 -12700 4881 -12677
rect 5281 -12564 5361 -12518
rect 5281 -12598 5304 -12564
rect 5338 -12598 5361 -12564
rect 5281 -12644 5361 -12598
rect 5281 -12678 5304 -12644
rect 5338 -12678 5361 -12644
rect 1171 -12754 1251 -12740
rect 1171 -12806 1185 -12754
rect 1237 -12806 1251 -12754
rect 1171 -12820 1251 -12806
rect 1841 -12850 1881 -12700
rect 2141 -12850 2181 -12700
rect 2441 -12850 2481 -12700
rect 3891 -12850 3931 -12700
rect 4191 -12850 4231 -12700
rect 4491 -12850 4531 -12700
rect 5281 -12701 5361 -12678
rect 5581 -12484 5661 -12451
rect 5581 -12518 5604 -12484
rect 5638 -12518 5661 -12484
rect 5581 -12564 5661 -12518
rect 5581 -12598 5604 -12564
rect 5638 -12598 5661 -12564
rect 5581 -12644 5661 -12598
rect 5581 -12678 5604 -12644
rect 5638 -12678 5661 -12644
rect 5581 -12701 5661 -12678
rect 5911 -12484 5991 -12451
rect 5911 -12518 5934 -12484
rect 5968 -12518 5991 -12484
rect 5911 -12564 5991 -12518
rect 5911 -12598 5934 -12564
rect 5968 -12598 5991 -12564
rect 5911 -12644 5991 -12598
rect 5911 -12678 5934 -12644
rect 5968 -12678 5991 -12644
rect 5911 -12701 5991 -12678
rect 6211 -12484 6291 -12451
rect 6211 -12518 6234 -12484
rect 6268 -12518 6291 -12484
rect 6211 -12564 6291 -12518
rect 6211 -12598 6234 -12564
rect 6268 -12598 6291 -12564
rect 6211 -12644 6291 -12598
rect 6211 -12678 6234 -12644
rect 6268 -12678 6291 -12644
rect 6211 -12701 6291 -12678
rect 6511 -12484 6591 -12451
rect 6511 -12518 6534 -12484
rect 6568 -12518 6591 -12484
rect 6511 -12564 6591 -12518
rect 6511 -12598 6534 -12564
rect 6568 -12598 6591 -12564
rect 6511 -12644 6591 -12598
rect 6511 -12678 6534 -12644
rect 6568 -12678 6591 -12644
rect 6511 -12701 6591 -12678
rect 7141 -12484 7221 -12451
rect 7141 -12518 7164 -12484
rect 7198 -12518 7221 -12484
rect 7141 -12564 7221 -12518
rect 7141 -12598 7164 -12564
rect 7198 -12598 7221 -12564
rect 7141 -12644 7221 -12598
rect 7141 -12678 7164 -12644
rect 7198 -12678 7221 -12644
rect 7141 -12701 7221 -12678
rect 5092 -12756 5172 -12742
rect 5092 -12808 5106 -12756
rect 5158 -12808 5172 -12756
rect 5092 -12822 5172 -12808
rect 912 -12917 935 -12883
rect 969 -12917 992 -12883
rect 912 -12940 992 -12917
rect 1161 -12851 5251 -12850
rect 5931 -12851 5971 -12701
rect 6231 -12851 6271 -12701
rect 6531 -12851 6571 -12701
rect 1161 -12883 7251 -12851
rect 1161 -12917 1184 -12883
rect 1218 -12917 1264 -12883
rect 1298 -12917 1344 -12883
rect 1378 -12917 1424 -12883
rect 1458 -12917 1504 -12883
rect 1538 -12917 1584 -12883
rect 1618 -12917 1664 -12883
rect 1698 -12917 1744 -12883
rect 1778 -12917 1824 -12883
rect 1858 -12917 1904 -12883
rect 1938 -12917 1984 -12883
rect 2018 -12917 2064 -12883
rect 2098 -12917 2144 -12883
rect 2178 -12917 2224 -12883
rect 2258 -12917 2304 -12883
rect 2338 -12917 2384 -12883
rect 2418 -12917 2464 -12883
rect 2498 -12917 2544 -12883
rect 2578 -12917 2624 -12883
rect 2658 -12917 2704 -12883
rect 2738 -12917 2784 -12883
rect 2818 -12917 2864 -12883
rect 2898 -12917 2944 -12883
rect 2978 -12917 3024 -12883
rect 3058 -12917 3104 -12883
rect 3138 -12917 3554 -12883
rect 3588 -12917 3634 -12883
rect 3668 -12917 3714 -12883
rect 3748 -12917 3794 -12883
rect 3828 -12917 3874 -12883
rect 3908 -12917 3954 -12883
rect 3988 -12917 4034 -12883
rect 4068 -12917 4114 -12883
rect 4148 -12917 4194 -12883
rect 4228 -12917 4274 -12883
rect 4308 -12917 4354 -12883
rect 4388 -12917 4434 -12883
rect 4468 -12917 4514 -12883
rect 4548 -12917 4594 -12883
rect 4628 -12917 4674 -12883
rect 4708 -12917 4754 -12883
rect 4788 -12917 4834 -12883
rect 4868 -12884 7251 -12883
rect 4868 -12917 5274 -12884
rect 1161 -12918 5274 -12917
rect 5308 -12918 5354 -12884
rect 5388 -12918 5434 -12884
rect 5468 -12918 5514 -12884
rect 5548 -12918 5594 -12884
rect 5628 -12918 5674 -12884
rect 5708 -12918 5754 -12884
rect 5788 -12918 5834 -12884
rect 5868 -12918 5914 -12884
rect 5948 -12918 5994 -12884
rect 6028 -12918 6074 -12884
rect 6108 -12918 6154 -12884
rect 6188 -12918 6234 -12884
rect 6268 -12918 6314 -12884
rect 6348 -12918 6394 -12884
rect 6428 -12918 6474 -12884
rect 6508 -12918 6554 -12884
rect 6588 -12918 6634 -12884
rect 6668 -12918 6714 -12884
rect 6748 -12918 6794 -12884
rect 6828 -12918 6874 -12884
rect 6908 -12918 6954 -12884
rect 6988 -12918 7034 -12884
rect 7068 -12918 7114 -12884
rect 7148 -12918 7194 -12884
rect 7228 -12918 7251 -12884
rect 1161 -12950 7251 -12918
rect 5251 -12951 7251 -12950
<< via1 >>
rect 1034 2435 1086 2487
rect 5844 2478 5896 2487
rect 5844 2444 5877 2478
rect 5877 2444 5896 2478
rect 5844 2435 5896 2444
rect 242 2318 294 2370
rect 242 -7604 294 -7552
rect 242 -11157 294 -11105
rect 356 1484 408 1536
rect 356 -8339 408 -8287
rect 356 -10450 408 -10398
rect 470 1644 522 1696
rect 584 2175 636 2227
rect 582 -1909 634 -1857
rect 470 -2616 522 -2564
rect 470 -6966 522 -6914
rect 584 -6235 636 -6183
rect 698 -512 750 -460
rect 698 -9754 750 -9702
rect 812 -1213 864 -1161
rect 812 -9054 864 -9002
rect 1554 2348 1606 2357
rect 1554 2314 1563 2348
rect 1563 2314 1597 2348
rect 1597 2314 1606 2348
rect 1554 2305 1606 2314
rect 1684 2248 1736 2257
rect 1684 2214 1693 2248
rect 1693 2214 1727 2248
rect 1727 2214 1736 2248
rect 1684 2205 1736 2214
rect 1554 2148 1606 2157
rect 1554 2114 1563 2148
rect 1563 2114 1597 2148
rect 1597 2114 1606 2148
rect 1554 2105 1606 2114
rect 1684 2048 1736 2057
rect 1684 2014 1693 2048
rect 1693 2014 1727 2048
rect 1727 2014 1736 2048
rect 1684 2005 1736 2014
rect 2814 2348 2866 2357
rect 2814 2314 2823 2348
rect 2823 2314 2857 2348
rect 2857 2314 2866 2348
rect 2814 2305 2866 2314
rect 2714 2048 2766 2057
rect 2714 2014 2723 2048
rect 2723 2014 2757 2048
rect 2757 2014 2766 2048
rect 2714 2005 2766 2014
rect 3002 2318 3054 2370
rect 3014 2248 3066 2257
rect 3014 2214 3023 2248
rect 3023 2214 3057 2248
rect 3057 2214 3066 2248
rect 3014 2205 3066 2214
rect 3282 2178 3334 2230
rect 3164 2148 3216 2157
rect 3164 2114 3173 2148
rect 3173 2114 3207 2148
rect 3207 2114 3216 2148
rect 3164 2105 3216 2114
rect 3314 2056 3366 2065
rect 3314 2022 3323 2056
rect 3323 2022 3357 2056
rect 3357 2022 3366 2056
rect 3314 2013 3366 2022
rect 3068 1968 3120 1977
rect 3068 1934 3077 1968
rect 3077 1934 3111 1968
rect 3111 1934 3120 1968
rect 3068 1925 3120 1934
rect 3314 1854 3366 1863
rect 3314 1820 3323 1854
rect 3323 1820 3357 1854
rect 3357 1820 3366 1854
rect 3314 1811 3366 1820
rect 3349 1644 3401 1696
rect 3349 1484 3401 1536
rect 4004 2218 4056 2227
rect 4004 2184 4013 2218
rect 4013 2184 4047 2218
rect 4047 2184 4056 2218
rect 4004 2175 4056 2184
rect 4004 2098 4056 2107
rect 4004 2064 4013 2098
rect 4013 2064 4047 2098
rect 4047 2064 4056 2098
rect 4004 2055 4056 2064
rect 4984 2098 5036 2107
rect 4984 2064 4993 2098
rect 4993 2064 5027 2098
rect 5027 2064 5036 2098
rect 4984 2055 5036 2064
rect 5298 2283 5350 2335
rect 5184 2218 5236 2227
rect 5184 2184 5193 2218
rect 5193 2184 5227 2218
rect 5227 2184 5236 2218
rect 5184 2175 5236 2184
rect 5384 1944 5436 1996
rect 6024 2248 6076 2257
rect 6024 2214 6033 2248
rect 6033 2214 6067 2248
rect 6067 2214 6076 2248
rect 6024 2205 6076 2214
rect 6024 2128 6076 2137
rect 6024 2094 6033 2128
rect 6033 2094 6067 2128
rect 6067 2094 6076 2128
rect 6024 2085 6076 2094
rect 7154 2248 7206 2257
rect 7154 2214 7163 2248
rect 7163 2214 7197 2248
rect 7197 2214 7206 2248
rect 7154 2205 7206 2214
rect 7004 2128 7056 2137
rect 7004 2094 7013 2128
rect 7013 2094 7047 2128
rect 7047 2094 7056 2128
rect 7004 2085 7056 2094
rect 7354 1978 7406 1987
rect 7354 1944 7363 1978
rect 7363 1944 7397 1978
rect 7397 1944 7406 1978
rect 7354 1935 7406 1944
rect 1143 1418 1195 1427
rect 1143 1384 1152 1418
rect 1152 1384 1186 1418
rect 1186 1384 1195 1418
rect 1143 1375 1195 1384
rect 5342 1495 5394 1547
rect 5756 1418 5808 1427
rect 5756 1384 5765 1418
rect 5765 1384 5799 1418
rect 5799 1384 5808 1418
rect 5756 1375 5808 1384
rect 1142 1178 1194 1187
rect 1142 1144 1151 1178
rect 1151 1144 1185 1178
rect 1185 1144 1194 1178
rect 1142 1135 1194 1144
rect 5087 1179 5139 1188
rect 5087 1145 5096 1179
rect 5096 1145 5130 1179
rect 5130 1145 5139 1179
rect 5087 1136 5139 1145
rect 5936 1178 5988 1187
rect 5936 1144 5945 1178
rect 5945 1144 5979 1178
rect 5979 1144 5988 1178
rect 5342 1015 5394 1067
rect 5936 1135 5988 1144
rect 1684 468 1736 477
rect 1684 434 1693 468
rect 1693 434 1727 468
rect 1727 434 1736 468
rect 1684 425 1736 434
rect 1684 348 1736 357
rect 1684 314 1693 348
rect 1693 314 1727 348
rect 1727 314 1736 348
rect 1684 305 1736 314
rect 2664 468 2716 477
rect 2664 434 2673 468
rect 2673 434 2707 468
rect 2707 434 2716 468
rect 2664 425 2716 434
rect 2814 348 2866 357
rect 2814 314 2823 348
rect 2823 314 2857 348
rect 2857 314 2866 348
rect 2814 305 2866 314
rect 3574 568 3626 577
rect 3574 534 3583 568
rect 3583 534 3617 568
rect 3617 534 3626 568
rect 3574 525 3626 534
rect 3068 348 3120 357
rect 3068 314 3077 348
rect 3077 314 3111 348
rect 3111 314 3120 348
rect 3068 305 3120 314
rect 4004 468 4056 477
rect 4004 434 4013 468
rect 4013 434 4047 468
rect 4047 434 4056 468
rect 4004 425 4056 434
rect 4004 348 4056 357
rect 4004 314 4013 348
rect 4013 314 4047 348
rect 4047 314 4056 348
rect 4004 305 4056 314
rect 4984 468 5036 477
rect 4984 434 4993 468
rect 4993 434 5027 468
rect 5027 434 5036 468
rect 4984 425 5036 434
rect 5134 348 5186 357
rect 5134 314 5143 348
rect 5143 314 5177 348
rect 5177 314 5186 348
rect 5134 305 5186 314
rect 1034 75 1086 127
rect 5150 -245 5202 -193
rect 5569 845 5621 897
rect 7104 888 7156 897
rect 7104 854 7113 888
rect 7113 854 7147 888
rect 7147 854 7156 888
rect 7104 845 7156 854
rect 7362 845 7414 897
rect 5674 738 5726 747
rect 5674 704 5683 738
rect 5683 704 5717 738
rect 5717 704 5726 738
rect 5674 695 5726 704
rect 5674 618 5726 627
rect 5674 584 5683 618
rect 5683 584 5717 618
rect 5717 584 5726 618
rect 5674 575 5726 584
rect 5744 378 5796 387
rect 5744 344 5753 378
rect 5753 344 5787 378
rect 5787 344 5796 378
rect 5744 335 5796 344
rect 5944 498 5996 507
rect 5944 464 5953 498
rect 5953 464 5987 498
rect 5987 464 5996 498
rect 5944 455 5996 464
rect 6924 498 6976 507
rect 6924 464 6933 498
rect 6933 464 6967 498
rect 6967 464 6976 498
rect 6924 455 6976 464
rect 6924 378 6976 387
rect 6924 344 6933 378
rect 6933 344 6967 378
rect 6967 344 6976 378
rect 6924 335 6976 344
rect 5492 75 5544 127
rect 5754 118 5806 127
rect 5754 84 5763 118
rect 5763 84 5797 118
rect 5797 84 5806 118
rect 5754 75 5806 84
rect 1070 -342 1122 -333
rect 1070 -376 1103 -342
rect 1103 -376 1122 -342
rect 1070 -385 1122 -376
rect 7004 -342 7056 -333
rect 7004 -376 7013 -342
rect 7013 -376 7047 -342
rect 7047 -376 7056 -342
rect 7004 -385 7056 -376
rect 1554 -472 1606 -463
rect 1554 -506 1563 -472
rect 1563 -506 1597 -472
rect 1597 -506 1606 -472
rect 1554 -515 1606 -506
rect 1684 -572 1736 -563
rect 1684 -606 1693 -572
rect 1693 -606 1727 -572
rect 1727 -606 1736 -572
rect 1684 -615 1736 -606
rect 1554 -672 1606 -663
rect 1554 -706 1563 -672
rect 1563 -706 1597 -672
rect 1597 -706 1606 -672
rect 1554 -715 1606 -706
rect 1684 -772 1736 -763
rect 1684 -806 1693 -772
rect 1693 -806 1727 -772
rect 1727 -806 1736 -772
rect 1684 -815 1736 -806
rect 2814 -472 2866 -463
rect 2814 -506 2823 -472
rect 2823 -506 2857 -472
rect 2857 -506 2866 -472
rect 2814 -515 2866 -506
rect 2714 -772 2766 -763
rect 2714 -806 2723 -772
rect 2723 -806 2757 -772
rect 2757 -806 2766 -772
rect 2714 -815 2766 -806
rect 3014 -572 3066 -563
rect 3014 -606 3023 -572
rect 3023 -606 3057 -572
rect 3057 -606 3066 -572
rect 3014 -615 3066 -606
rect 3586 -538 3638 -529
rect 3586 -572 3595 -538
rect 3595 -572 3629 -538
rect 3629 -572 3638 -538
rect 3586 -581 3638 -572
rect 3164 -672 3216 -663
rect 3164 -706 3173 -672
rect 3173 -706 3207 -672
rect 3207 -706 3216 -672
rect 3164 -715 3216 -706
rect 3586 -692 3638 -640
rect 3874 -512 3926 -460
rect 3874 -722 3926 -713
rect 3874 -756 3883 -722
rect 3883 -756 3917 -722
rect 3917 -756 3926 -722
rect 3874 -765 3926 -756
rect 4774 -722 4826 -713
rect 4774 -756 4783 -722
rect 4783 -756 4817 -722
rect 4817 -756 4826 -722
rect 4774 -765 4826 -756
rect 3328 -1170 3380 -1161
rect 3328 -1204 3337 -1170
rect 3337 -1204 3371 -1170
rect 3371 -1204 3380 -1170
rect 3328 -1213 3380 -1204
rect 5265 -458 5317 -449
rect 5265 -492 5274 -458
rect 5274 -492 5308 -458
rect 5308 -492 5317 -458
rect 5265 -501 5317 -492
rect 5486 -460 5538 -451
rect 5486 -494 5495 -460
rect 5495 -494 5529 -460
rect 5529 -494 5538 -460
rect 5486 -503 5538 -494
rect 5062 -602 5114 -550
rect 5062 -711 5114 -659
rect 5754 -572 5806 -563
rect 5754 -606 5763 -572
rect 5763 -606 5797 -572
rect 5797 -606 5806 -572
rect 5754 -615 5806 -606
rect 5754 -692 5806 -683
rect 5754 -726 5763 -692
rect 5763 -726 5797 -692
rect 5797 -726 5806 -692
rect 5754 -735 5806 -726
rect 6884 -572 6936 -563
rect 6884 -606 6893 -572
rect 6893 -606 6927 -572
rect 6927 -606 6936 -572
rect 6884 -615 6936 -606
rect 6734 -692 6786 -683
rect 6734 -726 6743 -692
rect 6743 -726 6777 -692
rect 6777 -726 6786 -692
rect 6734 -735 6786 -726
rect 7087 -962 7139 -953
rect 7087 -996 7096 -962
rect 7096 -996 7130 -962
rect 7130 -996 7139 -962
rect 7087 -1005 7139 -996
rect 6984 -1282 7036 -1273
rect 6984 -1316 6993 -1282
rect 6993 -1316 7027 -1282
rect 7027 -1316 7036 -1282
rect 6984 -1325 7036 -1316
rect 1185 -1402 1237 -1393
rect 1185 -1436 1194 -1402
rect 1194 -1436 1228 -1402
rect 1228 -1436 1237 -1402
rect 1185 -1445 1237 -1436
rect 5412 -1402 5464 -1393
rect 5412 -1436 5421 -1402
rect 5421 -1436 5455 -1402
rect 5455 -1436 5464 -1402
rect 5412 -1445 5464 -1436
rect 1185 -1642 1237 -1633
rect 1185 -1676 1194 -1642
rect 1194 -1676 1228 -1642
rect 1228 -1676 1237 -1642
rect 1185 -1685 1237 -1676
rect 5412 -1641 5464 -1632
rect 5412 -1675 5421 -1641
rect 5421 -1675 5455 -1641
rect 5455 -1675 5464 -1641
rect 5412 -1684 5464 -1675
rect 3328 -1865 3380 -1856
rect 3328 -1899 3337 -1865
rect 3337 -1899 3371 -1865
rect 3371 -1899 3380 -1865
rect 3328 -1908 3380 -1899
rect 1684 -2272 1736 -2263
rect 1684 -2306 1693 -2272
rect 1693 -2306 1727 -2272
rect 1727 -2306 1736 -2272
rect 1684 -2315 1736 -2306
rect 1554 -2372 1606 -2363
rect 1554 -2406 1563 -2372
rect 1563 -2406 1597 -2372
rect 1597 -2406 1606 -2372
rect 1554 -2415 1606 -2406
rect 1684 -2472 1736 -2463
rect 1684 -2506 1693 -2472
rect 1693 -2506 1727 -2472
rect 1727 -2506 1736 -2472
rect 1684 -2515 1736 -2506
rect 1554 -2572 1606 -2563
rect 1554 -2606 1563 -2572
rect 1563 -2606 1597 -2572
rect 1597 -2606 1606 -2572
rect 1554 -2615 1606 -2606
rect 2714 -2272 2766 -2263
rect 2714 -2306 2723 -2272
rect 2723 -2306 2757 -2272
rect 2757 -2306 2766 -2272
rect 2714 -2315 2766 -2306
rect 2814 -2572 2866 -2563
rect 2814 -2606 2823 -2572
rect 2823 -2606 2857 -2572
rect 2857 -2606 2866 -2572
rect 2814 -2615 2866 -2606
rect 3164 -2372 3216 -2363
rect 3164 -2406 3173 -2372
rect 3173 -2406 3207 -2372
rect 3207 -2406 3216 -2372
rect 3164 -2415 3216 -2406
rect 3586 -2436 3638 -2384
rect 3014 -2472 3066 -2463
rect 3014 -2506 3023 -2472
rect 3023 -2506 3057 -2472
rect 3057 -2506 3066 -2472
rect 3014 -2515 3066 -2506
rect 3586 -2506 3638 -2497
rect 3586 -2540 3595 -2506
rect 3595 -2540 3629 -2506
rect 3629 -2540 3638 -2506
rect 3586 -2549 3638 -2540
rect 3874 -2322 3926 -2313
rect 3874 -2356 3883 -2322
rect 3883 -2356 3917 -2322
rect 3917 -2356 3926 -2322
rect 3874 -2365 3926 -2356
rect 3874 -2616 3926 -2564
rect 4774 -2322 4826 -2313
rect 4774 -2356 4783 -2322
rect 4783 -2356 4817 -2322
rect 4817 -2356 4826 -2322
rect 4774 -2365 4826 -2356
rect 6984 -1762 7036 -1753
rect 6984 -1796 6993 -1762
rect 6993 -1796 7027 -1762
rect 7027 -1796 7036 -1762
rect 6984 -1805 7036 -1796
rect 5062 -2403 5114 -2351
rect 5062 -2511 5114 -2459
rect 5754 -2352 5806 -2343
rect 5754 -2386 5763 -2352
rect 5763 -2386 5797 -2352
rect 5797 -2386 5806 -2352
rect 5754 -2395 5806 -2386
rect 5754 -2472 5806 -2463
rect 5754 -2506 5763 -2472
rect 5763 -2506 5797 -2472
rect 5797 -2506 5806 -2472
rect 5754 -2515 5806 -2506
rect 6734 -2352 6786 -2343
rect 6734 -2386 6743 -2352
rect 6743 -2386 6777 -2352
rect 6777 -2386 6786 -2352
rect 6734 -2395 6786 -2386
rect 6884 -2472 6936 -2463
rect 6884 -2506 6893 -2472
rect 6893 -2506 6927 -2472
rect 6927 -2506 6936 -2472
rect 6884 -2515 6936 -2506
rect 7087 -2082 7139 -2073
rect 7087 -2116 7096 -2082
rect 7096 -2116 7130 -2082
rect 7130 -2116 7139 -2082
rect 7087 -2125 7139 -2116
rect 1069 -2702 1121 -2693
rect 1069 -2736 1103 -2702
rect 1103 -2736 1121 -2702
rect 1069 -2745 1121 -2736
rect 5412 -2936 5464 -2927
rect 5412 -2970 5421 -2936
rect 5421 -2970 5455 -2936
rect 5455 -2970 5464 -2936
rect 5412 -2979 5464 -2970
rect 7357 -2969 7409 -2960
rect 7357 -3003 7366 -2969
rect 7366 -3003 7400 -2969
rect 7400 -3003 7409 -2969
rect 7357 -3012 7409 -3003
rect 1069 -3206 1121 -3154
rect 5265 -3163 5317 -3154
rect 5265 -3197 5274 -3163
rect 5274 -3197 5308 -3163
rect 5308 -3197 5317 -3163
rect 5265 -3206 5317 -3197
rect 1595 -3282 1647 -3273
rect 1595 -3316 1604 -3282
rect 1604 -3316 1638 -3282
rect 1638 -3316 1647 -3282
rect 1595 -3325 1647 -3316
rect 1685 -3402 1737 -3393
rect 1685 -3436 1694 -3402
rect 1694 -3436 1728 -3402
rect 1728 -3436 1737 -3402
rect 1685 -3445 1737 -3436
rect 1655 -3522 1707 -3513
rect 1655 -3556 1664 -3522
rect 1664 -3556 1698 -3522
rect 1698 -3556 1707 -3522
rect 1655 -3565 1707 -3556
rect 2965 -3282 3017 -3273
rect 2965 -3316 2974 -3282
rect 2974 -3316 3008 -3282
rect 3008 -3316 3017 -3282
rect 2965 -3325 3017 -3316
rect 2815 -3402 2867 -3393
rect 2815 -3436 2824 -3402
rect 2824 -3436 2858 -3402
rect 2858 -3436 2867 -3402
rect 2815 -3445 2867 -3436
rect 2685 -3522 2737 -3513
rect 2685 -3556 2694 -3522
rect 2694 -3556 2728 -3522
rect 2728 -3556 2737 -3522
rect 2685 -3565 2737 -3556
rect 3065 -4102 3117 -4093
rect 3065 -4136 3074 -4102
rect 3074 -4136 3108 -4102
rect 3108 -4136 3117 -4102
rect 3065 -4145 3117 -4136
rect 3735 -3542 3787 -3533
rect 3735 -3576 3744 -3542
rect 3744 -3576 3778 -3542
rect 3778 -3576 3787 -3542
rect 3735 -3585 3787 -3576
rect 4635 -3542 4687 -3533
rect 4635 -3576 4644 -3542
rect 4644 -3576 4678 -3542
rect 4678 -3576 4687 -3542
rect 4635 -3585 4687 -3576
rect 5018 -3369 5070 -3360
rect 5018 -3403 5027 -3369
rect 5027 -3403 5061 -3369
rect 5061 -3403 5070 -3369
rect 5018 -3412 5070 -3403
rect 5194 -3498 5246 -3446
rect 5194 -3565 5246 -3556
rect 5194 -3599 5203 -3565
rect 5203 -3599 5237 -3565
rect 5237 -3599 5246 -3565
rect 5194 -3608 5246 -3599
rect 5195 -3679 5247 -3670
rect 5195 -3713 5204 -3679
rect 5204 -3713 5238 -3679
rect 5238 -3713 5247 -3679
rect 5195 -3722 5247 -3713
rect 5195 -3793 5247 -3784
rect 5195 -3827 5204 -3793
rect 5204 -3827 5238 -3793
rect 5238 -3827 5247 -3793
rect 5195 -3836 5247 -3827
rect 5395 -3288 5447 -3279
rect 5395 -3322 5404 -3288
rect 5404 -3322 5438 -3288
rect 5438 -3322 5447 -3288
rect 5395 -3331 5447 -3322
rect 5495 -3413 5547 -3404
rect 5495 -3447 5504 -3413
rect 5504 -3447 5538 -3413
rect 5538 -3447 5547 -3413
rect 5495 -3456 5547 -3447
rect 5695 -3503 5747 -3494
rect 5695 -3537 5704 -3503
rect 5704 -3537 5738 -3503
rect 5738 -3537 5747 -3503
rect 5695 -3546 5747 -3537
rect 6675 -3293 6727 -3284
rect 6675 -3327 6684 -3293
rect 6684 -3327 6718 -3293
rect 6718 -3327 6727 -3293
rect 6675 -3336 6727 -3327
rect 6795 -3403 6847 -3394
rect 6795 -3437 6804 -3403
rect 6804 -3437 6838 -3403
rect 6838 -3437 6847 -3403
rect 6795 -3446 6847 -3437
rect 7047 -3403 7099 -3394
rect 7047 -3437 7056 -3403
rect 7056 -3437 7090 -3403
rect 7090 -3437 7099 -3403
rect 7047 -3446 7099 -3437
rect 6675 -3503 6727 -3494
rect 6675 -3537 6684 -3503
rect 6684 -3537 6718 -3503
rect 6718 -3537 6727 -3503
rect 6675 -3546 6727 -3537
rect 6805 -3634 6857 -3582
rect 7243 -3293 7295 -3284
rect 7243 -3327 7252 -3293
rect 7252 -3327 7286 -3293
rect 7286 -3327 7295 -3293
rect 7243 -3336 7295 -3327
rect 7289 -3591 7341 -3582
rect 7289 -3625 7298 -3591
rect 7298 -3625 7332 -3591
rect 7332 -3625 7341 -3591
rect 7289 -3634 7341 -3625
rect 5012 -3946 5064 -3937
rect 5012 -3980 5021 -3946
rect 5021 -3980 5055 -3946
rect 5055 -3980 5064 -3946
rect 5012 -3989 5064 -3980
rect 4815 -4102 4867 -4093
rect 4815 -4136 4824 -4102
rect 4824 -4136 4858 -4102
rect 4858 -4136 4867 -4102
rect 4815 -4145 4867 -4136
rect 1185 -4222 1237 -4213
rect 1185 -4256 1194 -4222
rect 1194 -4256 1228 -4222
rect 1228 -4256 1237 -4222
rect 1185 -4265 1237 -4256
rect 7155 -4103 7207 -4093
rect 7155 -4137 7164 -4103
rect 7164 -4137 7198 -4103
rect 7198 -4137 7207 -4103
rect 7155 -4145 7207 -4137
rect 5106 -4224 5158 -4215
rect 5106 -4258 5115 -4224
rect 5115 -4258 5149 -4224
rect 5149 -4258 5158 -4224
rect 5106 -4267 5158 -4258
rect 1055 -4545 1107 -4536
rect 1055 -4579 1064 -4545
rect 1064 -4579 1098 -4545
rect 1098 -4579 1107 -4545
rect 1055 -4588 1107 -4579
rect 5129 -4543 5181 -4534
rect 5129 -4577 5138 -4543
rect 5138 -4577 5172 -4543
rect 5172 -4577 5181 -4543
rect 5129 -4586 5181 -4577
rect 5326 -4543 5378 -4534
rect 5326 -4577 5335 -4543
rect 5335 -4577 5369 -4543
rect 5369 -4577 5378 -4543
rect 5326 -4586 5378 -4577
rect 3254 -4662 3306 -4654
rect 3254 -4696 3263 -4662
rect 3263 -4696 3297 -4662
rect 3297 -4696 3306 -4662
rect 3254 -4706 3306 -4696
rect 1144 -5432 1196 -5423
rect 1144 -5466 1153 -5432
rect 1153 -5466 1187 -5432
rect 1187 -5466 1196 -5432
rect 1144 -5475 1196 -5466
rect 1144 -5552 1196 -5543
rect 1144 -5586 1153 -5552
rect 1153 -5586 1187 -5552
rect 1187 -5586 1196 -5552
rect 1144 -5595 1196 -5586
rect 1144 -5672 1196 -5663
rect 1144 -5706 1153 -5672
rect 1153 -5706 1187 -5672
rect 1187 -5706 1196 -5672
rect 1144 -5715 1196 -5706
rect 1144 -5792 1196 -5783
rect 1144 -5826 1153 -5792
rect 1153 -5826 1187 -5792
rect 1187 -5826 1196 -5792
rect 1144 -5835 1196 -5826
rect 2704 -5475 2756 -5423
rect 2854 -5595 2906 -5543
rect 3004 -5715 3056 -5663
rect 3154 -5835 3206 -5783
rect 5015 -4663 5067 -4654
rect 5015 -4697 5024 -4663
rect 5024 -4697 5058 -4663
rect 5058 -4697 5067 -4663
rect 5015 -4706 5067 -4697
rect 3935 -5223 3987 -5214
rect 3935 -5257 3944 -5223
rect 3944 -5257 3978 -5223
rect 3978 -5257 3987 -5223
rect 3935 -5266 3987 -5257
rect 4835 -5223 4887 -5214
rect 4835 -5257 4844 -5223
rect 4844 -5257 4878 -5223
rect 4878 -5257 4887 -5223
rect 4835 -5266 4887 -5257
rect 7374 -4663 7426 -4654
rect 7374 -4697 7383 -4663
rect 7383 -4697 7417 -4663
rect 7417 -4697 7426 -4663
rect 7374 -4706 7426 -4697
rect 5414 -4963 5466 -4954
rect 5414 -4997 5423 -4963
rect 5423 -4997 5457 -4963
rect 5457 -4997 5466 -4963
rect 5414 -5006 5466 -4997
rect 5414 -5083 5466 -5074
rect 5414 -5117 5423 -5083
rect 5423 -5117 5457 -5083
rect 5457 -5117 5466 -5083
rect 5414 -5126 5466 -5117
rect 5414 -5211 5466 -5202
rect 5414 -5245 5423 -5211
rect 5423 -5245 5457 -5211
rect 5457 -5245 5466 -5211
rect 5414 -5254 5466 -5245
rect 5414 -5369 5466 -5317
rect 5129 -5396 5181 -5387
rect 5129 -5430 5138 -5396
rect 5138 -5430 5172 -5396
rect 5172 -5430 5181 -5396
rect 5129 -5439 5181 -5430
rect 5714 -5353 5766 -5344
rect 5714 -5387 5723 -5353
rect 5723 -5387 5757 -5353
rect 5757 -5387 5766 -5353
rect 5714 -5396 5766 -5387
rect 5614 -5478 5666 -5469
rect 5614 -5512 5623 -5478
rect 5623 -5512 5657 -5478
rect 5657 -5512 5666 -5478
rect 5614 -5521 5666 -5512
rect 5914 -5263 5966 -5254
rect 5914 -5297 5923 -5263
rect 5923 -5297 5957 -5263
rect 5957 -5297 5966 -5263
rect 5914 -5306 5966 -5297
rect 7024 -5219 7076 -5167
rect 6894 -5263 6946 -5254
rect 6894 -5297 6903 -5263
rect 6903 -5297 6937 -5263
rect 6937 -5297 6946 -5263
rect 6894 -5306 6946 -5297
rect 7014 -5363 7066 -5354
rect 7014 -5397 7023 -5363
rect 7023 -5397 7057 -5363
rect 7057 -5397 7066 -5363
rect 7014 -5406 7066 -5397
rect 7146 -5362 7198 -5353
rect 7146 -5396 7155 -5362
rect 7155 -5396 7189 -5362
rect 7189 -5396 7198 -5362
rect 7146 -5405 7198 -5396
rect 6894 -5473 6946 -5464
rect 6894 -5507 6903 -5473
rect 6903 -5507 6937 -5473
rect 6937 -5507 6946 -5473
rect 6894 -5516 6946 -5507
rect 7284 -5473 7336 -5464
rect 7284 -5507 7293 -5473
rect 7293 -5507 7327 -5473
rect 7327 -5507 7336 -5473
rect 7284 -5516 7336 -5507
rect 7508 -5176 7560 -5167
rect 7508 -5210 7517 -5176
rect 7517 -5210 7551 -5176
rect 7551 -5210 7560 -5176
rect 7508 -5219 7560 -5210
rect 5580 -5603 5632 -5594
rect 5580 -5637 5607 -5603
rect 5607 -5637 5632 -5603
rect 5580 -5646 5632 -5637
rect 5472 -5829 5524 -5820
rect 5472 -5863 5481 -5829
rect 5481 -5863 5515 -5829
rect 5515 -5863 5524 -5829
rect 5472 -5872 5524 -5863
rect 7508 -5797 7560 -5788
rect 7508 -5831 7517 -5797
rect 7517 -5831 7551 -5797
rect 7551 -5831 7560 -5797
rect 7508 -5840 7560 -5831
rect 1594 -6193 1646 -6184
rect 1594 -6227 1603 -6193
rect 1603 -6227 1637 -6193
rect 1637 -6227 1646 -6193
rect 1594 -6236 1646 -6227
rect 1724 -6293 1776 -6284
rect 1724 -6327 1733 -6293
rect 1733 -6327 1767 -6293
rect 1767 -6327 1776 -6293
rect 1724 -6336 1776 -6327
rect 1594 -6393 1646 -6384
rect 1594 -6427 1603 -6393
rect 1603 -6427 1637 -6393
rect 1637 -6427 1646 -6393
rect 1594 -6436 1646 -6427
rect 1724 -6493 1776 -6484
rect 1724 -6527 1733 -6493
rect 1733 -6527 1767 -6493
rect 1767 -6527 1776 -6493
rect 1724 -6536 1776 -6527
rect 2854 -6193 2906 -6184
rect 2854 -6227 2863 -6193
rect 2863 -6227 2897 -6193
rect 2897 -6227 2906 -6193
rect 2854 -6236 2906 -6227
rect 2754 -6493 2806 -6484
rect 2754 -6527 2763 -6493
rect 2763 -6527 2797 -6493
rect 2797 -6527 2806 -6493
rect 2754 -6536 2806 -6527
rect 3054 -6293 3106 -6284
rect 3054 -6327 3063 -6293
rect 3063 -6327 3097 -6293
rect 3097 -6327 3106 -6293
rect 3054 -6336 3106 -6327
rect 3646 -6293 3698 -6284
rect 3646 -6327 3655 -6293
rect 3655 -6327 3689 -6293
rect 3689 -6327 3698 -6293
rect 3646 -6336 3698 -6327
rect 3204 -6393 3256 -6384
rect 3204 -6427 3213 -6393
rect 3213 -6427 3247 -6393
rect 3247 -6427 3256 -6393
rect 3204 -6436 3256 -6427
rect 3645 -6895 3697 -6843
rect 3934 -6235 3986 -6183
rect 3934 -6443 3986 -6434
rect 3934 -6477 3943 -6443
rect 3943 -6477 3977 -6443
rect 3977 -6477 3986 -6443
rect 3934 -6486 3986 -6477
rect 4834 -6293 4886 -6284
rect 4834 -6327 4843 -6293
rect 4843 -6327 4877 -6293
rect 4877 -6327 4886 -6293
rect 4834 -6336 4886 -6327
rect 4834 -6443 4886 -6434
rect 4834 -6477 4843 -6443
rect 4843 -6477 4877 -6443
rect 4877 -6477 4886 -6443
rect 4834 -6486 4886 -6477
rect 3368 -6923 3420 -6914
rect 3368 -6957 3377 -6923
rect 3377 -6957 3411 -6923
rect 3411 -6957 3420 -6923
rect 3368 -6966 3420 -6957
rect 2954 -7003 3006 -6994
rect 2954 -7037 2963 -7003
rect 2963 -7037 2997 -7003
rect 2997 -7037 3006 -7003
rect 2954 -7046 3006 -7037
rect 5122 -6896 5174 -6844
rect 5813 -6293 5865 -6284
rect 5813 -6327 5822 -6293
rect 5822 -6327 5856 -6293
rect 5856 -6327 5865 -6293
rect 5813 -6336 5865 -6327
rect 5813 -6413 5865 -6404
rect 5813 -6447 5822 -6413
rect 5822 -6447 5856 -6413
rect 5856 -6447 5865 -6413
rect 5813 -6456 5865 -6447
rect 6943 -6293 6995 -6284
rect 6943 -6327 6952 -6293
rect 6952 -6327 6986 -6293
rect 6986 -6327 6995 -6293
rect 6943 -6336 6995 -6327
rect 6793 -6413 6845 -6404
rect 6793 -6447 6802 -6413
rect 6802 -6447 6836 -6413
rect 6836 -6447 6845 -6413
rect 6793 -6456 6845 -6447
rect 7143 -6683 7195 -6674
rect 7143 -6717 7152 -6683
rect 7152 -6717 7186 -6683
rect 7186 -6717 7195 -6683
rect 7143 -6726 7195 -6717
rect 7044 -7003 7096 -6994
rect 7044 -7037 7052 -7003
rect 7052 -7037 7086 -7003
rect 7086 -7037 7096 -7003
rect 7044 -7046 7096 -7037
rect 1506 -7123 1558 -7114
rect 1506 -7157 1515 -7123
rect 1515 -7157 1549 -7123
rect 1549 -7157 1558 -7123
rect 1506 -7166 1558 -7157
rect 5470 -7123 5522 -7114
rect 5470 -7157 5479 -7123
rect 5479 -7157 5513 -7123
rect 5513 -7157 5522 -7123
rect 5470 -7166 5522 -7157
rect 1506 -7363 1558 -7354
rect 1506 -7397 1515 -7363
rect 1515 -7397 1549 -7363
rect 1549 -7397 1558 -7363
rect 1506 -7406 1558 -7397
rect 5472 -7363 5524 -7354
rect 5472 -7397 5481 -7363
rect 5481 -7397 5515 -7363
rect 5515 -7397 5524 -7363
rect 5472 -7406 5524 -7397
rect 2954 -7483 3006 -7474
rect 2954 -7517 2963 -7483
rect 2963 -7517 2997 -7483
rect 2997 -7517 3006 -7483
rect 2954 -7526 3006 -7517
rect 3368 -7561 3420 -7552
rect 3368 -7595 3377 -7561
rect 3377 -7595 3411 -7561
rect 3411 -7595 3420 -7561
rect 3368 -7604 3420 -7595
rect 1724 -7993 1776 -7984
rect 1724 -8027 1733 -7993
rect 1733 -8027 1767 -7993
rect 1767 -8027 1776 -7993
rect 1724 -8036 1776 -8027
rect 1594 -8093 1646 -8084
rect 1594 -8127 1603 -8093
rect 1603 -8127 1637 -8093
rect 1637 -8127 1646 -8093
rect 1594 -8136 1646 -8127
rect 1724 -8193 1776 -8184
rect 1724 -8227 1733 -8193
rect 1733 -8227 1767 -8193
rect 1767 -8227 1776 -8193
rect 1724 -8236 1776 -8227
rect 1594 -8293 1646 -8284
rect 1594 -8327 1603 -8293
rect 1603 -8327 1637 -8293
rect 1637 -8327 1646 -8293
rect 1594 -8336 1646 -8327
rect 2754 -7993 2806 -7984
rect 2754 -8027 2763 -7993
rect 2763 -8027 2797 -7993
rect 2797 -8027 2806 -7993
rect 2754 -8036 2806 -8027
rect 2854 -8293 2906 -8284
rect 2854 -8327 2863 -8293
rect 2863 -8327 2897 -8293
rect 2897 -8327 2906 -8293
rect 2854 -8336 2906 -8327
rect 3204 -8093 3256 -8084
rect 3204 -8127 3213 -8093
rect 3213 -8127 3247 -8093
rect 3247 -8127 3256 -8093
rect 3204 -8136 3256 -8127
rect 3646 -8162 3698 -8110
rect 3054 -8193 3106 -8184
rect 3054 -8227 3063 -8193
rect 3063 -8227 3097 -8193
rect 3097 -8227 3106 -8193
rect 3054 -8236 3106 -8227
rect 3646 -8227 3698 -8218
rect 3646 -8261 3655 -8227
rect 3655 -8261 3689 -8227
rect 3689 -8261 3698 -8227
rect 3646 -8270 3698 -8261
rect 3934 -8043 3986 -8034
rect 3934 -8077 3943 -8043
rect 3943 -8077 3977 -8043
rect 3977 -8077 3986 -8043
rect 3934 -8086 3986 -8077
rect 3934 -8339 3986 -8287
rect 4834 -8043 4886 -8034
rect 4834 -8077 4843 -8043
rect 4843 -8077 4877 -8043
rect 4877 -8077 4886 -8043
rect 4834 -8086 4886 -8077
rect 7044 -7483 7096 -7474
rect 7044 -7517 7052 -7483
rect 7052 -7517 7086 -7483
rect 7086 -7517 7096 -7483
rect 7044 -7526 7096 -7517
rect 5122 -8112 5174 -8103
rect 5122 -8146 5131 -8112
rect 5131 -8146 5165 -8112
rect 5165 -8146 5174 -8112
rect 5122 -8155 5174 -8146
rect 5122 -8227 5174 -8218
rect 5122 -8261 5131 -8227
rect 5131 -8261 5165 -8227
rect 5165 -8261 5174 -8227
rect 5122 -8270 5174 -8261
rect 5813 -8073 5865 -8064
rect 5813 -8107 5822 -8073
rect 5822 -8107 5856 -8073
rect 5856 -8107 5865 -8073
rect 5813 -8116 5865 -8107
rect 5813 -8193 5865 -8184
rect 5813 -8227 5822 -8193
rect 5822 -8227 5856 -8193
rect 5856 -8227 5865 -8193
rect 5813 -8236 5865 -8227
rect 6793 -8073 6845 -8064
rect 6793 -8107 6802 -8073
rect 6802 -8107 6836 -8073
rect 6836 -8107 6845 -8073
rect 6793 -8116 6845 -8107
rect 6943 -8193 6995 -8184
rect 6943 -8227 6952 -8193
rect 6952 -8227 6986 -8193
rect 6986 -8227 6995 -8193
rect 6943 -8236 6995 -8227
rect 7147 -7804 7199 -7795
rect 7147 -7838 7156 -7804
rect 7156 -7838 7190 -7804
rect 7190 -7838 7199 -7804
rect 7147 -7847 7199 -7838
rect 1134 -8423 1186 -8414
rect 1134 -8457 1143 -8423
rect 1143 -8457 1177 -8423
rect 1177 -8457 1186 -8423
rect 1134 -8466 1186 -8457
rect 5704 -8423 5756 -8414
rect 5704 -8457 5712 -8423
rect 5712 -8457 5746 -8423
rect 5746 -8457 5756 -8423
rect 5704 -8466 5756 -8457
rect 5472 -8584 5524 -8532
rect 5412 -8808 5464 -8756
rect 1070 -8883 1122 -8874
rect 1070 -8917 1103 -8883
rect 1103 -8917 1122 -8883
rect 1070 -8926 1122 -8917
rect 5704 -8883 5756 -8874
rect 7004 -8883 7056 -8874
rect 5704 -8917 5733 -8883
rect 5733 -8917 5756 -8883
rect 7004 -8917 7013 -8883
rect 7013 -8917 7047 -8883
rect 7047 -8917 7056 -8883
rect 5704 -8926 5756 -8917
rect 7004 -8926 7056 -8917
rect 1554 -9013 1606 -9004
rect 1554 -9047 1563 -9013
rect 1563 -9047 1597 -9013
rect 1597 -9047 1606 -9013
rect 1554 -9056 1606 -9047
rect 1684 -9113 1736 -9104
rect 1684 -9147 1693 -9113
rect 1693 -9147 1727 -9113
rect 1727 -9147 1736 -9113
rect 1684 -9156 1736 -9147
rect 1554 -9213 1606 -9204
rect 1554 -9247 1563 -9213
rect 1563 -9247 1597 -9213
rect 1597 -9247 1606 -9213
rect 1554 -9256 1606 -9247
rect 1684 -9313 1736 -9304
rect 1684 -9347 1693 -9313
rect 1693 -9347 1727 -9313
rect 1727 -9347 1736 -9313
rect 1684 -9356 1736 -9347
rect 2814 -9013 2866 -9004
rect 2814 -9047 2823 -9013
rect 2823 -9047 2857 -9013
rect 2857 -9047 2866 -9013
rect 2814 -9056 2866 -9047
rect 2714 -9313 2766 -9304
rect 2714 -9347 2723 -9313
rect 2723 -9347 2757 -9313
rect 2757 -9347 2766 -9313
rect 2714 -9356 2766 -9347
rect 3014 -9113 3066 -9104
rect 3014 -9147 3023 -9113
rect 3023 -9147 3057 -9113
rect 3057 -9147 3066 -9113
rect 3014 -9156 3066 -9147
rect 3586 -9079 3638 -9070
rect 3586 -9113 3595 -9079
rect 3595 -9113 3629 -9079
rect 3629 -9113 3638 -9079
rect 3586 -9122 3638 -9113
rect 3164 -9213 3216 -9204
rect 3164 -9247 3173 -9213
rect 3173 -9247 3207 -9213
rect 3207 -9247 3216 -9213
rect 3164 -9256 3216 -9247
rect 3586 -9233 3638 -9181
rect 3874 -9053 3926 -9001
rect 3874 -9263 3926 -9254
rect 3874 -9297 3883 -9263
rect 3883 -9297 3917 -9263
rect 3917 -9297 3926 -9263
rect 3874 -9306 3926 -9297
rect 4774 -9263 4826 -9254
rect 4774 -9297 4783 -9263
rect 4783 -9297 4817 -9263
rect 4817 -9297 4826 -9263
rect 4774 -9306 4826 -9297
rect 3328 -9711 3380 -9702
rect 3328 -9745 3337 -9711
rect 3337 -9745 3371 -9711
rect 3371 -9745 3380 -9711
rect 3328 -9754 3380 -9745
rect 5062 -9143 5114 -9091
rect 5062 -9252 5114 -9200
rect 5754 -9113 5806 -9104
rect 5754 -9147 5763 -9113
rect 5763 -9147 5797 -9113
rect 5797 -9147 5806 -9113
rect 5754 -9156 5806 -9147
rect 5754 -9233 5806 -9224
rect 5754 -9267 5763 -9233
rect 5763 -9267 5797 -9233
rect 5797 -9267 5806 -9233
rect 5754 -9276 5806 -9267
rect 6884 -9113 6936 -9104
rect 6884 -9147 6893 -9113
rect 6893 -9147 6927 -9113
rect 6927 -9147 6936 -9113
rect 6884 -9156 6936 -9147
rect 6734 -9233 6786 -9224
rect 6734 -9267 6743 -9233
rect 6743 -9267 6777 -9233
rect 6777 -9267 6786 -9233
rect 6734 -9276 6786 -9267
rect 7087 -9503 7139 -9494
rect 7087 -9537 7096 -9503
rect 7096 -9537 7130 -9503
rect 7130 -9537 7139 -9503
rect 7087 -9546 7139 -9537
rect 6984 -9823 7036 -9814
rect 6984 -9857 6993 -9823
rect 6993 -9857 7027 -9823
rect 7027 -9857 7036 -9823
rect 6984 -9866 7036 -9857
rect 1185 -9943 1237 -9934
rect 1185 -9977 1194 -9943
rect 1194 -9977 1228 -9943
rect 1228 -9977 1237 -9943
rect 1185 -9986 1237 -9977
rect 5412 -9943 5464 -9934
rect 5412 -9977 5421 -9943
rect 5421 -9977 5455 -9943
rect 5455 -9977 5464 -9943
rect 5412 -9986 5464 -9977
rect 1185 -10183 1237 -10174
rect 1185 -10217 1194 -10183
rect 1194 -10217 1228 -10183
rect 1228 -10217 1237 -10183
rect 1185 -10226 1237 -10217
rect 5412 -10182 5464 -10173
rect 5412 -10216 5421 -10182
rect 5421 -10216 5455 -10182
rect 5455 -10216 5464 -10182
rect 5412 -10225 5464 -10216
rect 3328 -10406 3380 -10397
rect 3328 -10440 3337 -10406
rect 3337 -10440 3371 -10406
rect 3371 -10440 3380 -10406
rect 3328 -10449 3380 -10440
rect 1684 -10813 1736 -10804
rect 1684 -10847 1693 -10813
rect 1693 -10847 1727 -10813
rect 1727 -10847 1736 -10813
rect 1684 -10856 1736 -10847
rect 1554 -10913 1606 -10904
rect 1554 -10947 1563 -10913
rect 1563 -10947 1597 -10913
rect 1597 -10947 1606 -10913
rect 1554 -10956 1606 -10947
rect 1684 -11013 1736 -11004
rect 1684 -11047 1693 -11013
rect 1693 -11047 1727 -11013
rect 1727 -11047 1736 -11013
rect 1684 -11056 1736 -11047
rect 1554 -11113 1606 -11104
rect 1554 -11147 1563 -11113
rect 1563 -11147 1597 -11113
rect 1597 -11147 1606 -11113
rect 1554 -11156 1606 -11147
rect 2714 -10813 2766 -10804
rect 2714 -10847 2723 -10813
rect 2723 -10847 2757 -10813
rect 2757 -10847 2766 -10813
rect 2714 -10856 2766 -10847
rect 2814 -11113 2866 -11104
rect 2814 -11147 2823 -11113
rect 2823 -11147 2857 -11113
rect 2857 -11147 2866 -11113
rect 2814 -11156 2866 -11147
rect 3164 -10913 3216 -10904
rect 3164 -10947 3173 -10913
rect 3173 -10947 3207 -10913
rect 3207 -10947 3216 -10913
rect 3164 -10956 3216 -10947
rect 3586 -10977 3638 -10925
rect 3014 -11013 3066 -11004
rect 3014 -11047 3023 -11013
rect 3023 -11047 3057 -11013
rect 3057 -11047 3066 -11013
rect 3014 -11056 3066 -11047
rect 3586 -11047 3638 -11038
rect 3586 -11081 3595 -11047
rect 3595 -11081 3629 -11047
rect 3629 -11081 3638 -11047
rect 3586 -11090 3638 -11081
rect 3874 -10863 3926 -10854
rect 3874 -10897 3883 -10863
rect 3883 -10897 3917 -10863
rect 3917 -10897 3926 -10863
rect 3874 -10906 3926 -10897
rect 3874 -11157 3926 -11105
rect 4774 -10863 4826 -10854
rect 4774 -10897 4783 -10863
rect 4783 -10897 4817 -10863
rect 4817 -10897 4826 -10863
rect 4774 -10906 4826 -10897
rect 6984 -10303 7036 -10294
rect 6984 -10337 6993 -10303
rect 6993 -10337 7027 -10303
rect 7027 -10337 7036 -10303
rect 6984 -10346 7036 -10337
rect 5062 -10901 5114 -10892
rect 5062 -10935 5071 -10901
rect 5071 -10935 5105 -10901
rect 5105 -10935 5114 -10901
rect 5062 -10944 5114 -10935
rect 5062 -11052 5114 -11000
rect 5754 -10893 5806 -10884
rect 5754 -10927 5763 -10893
rect 5763 -10927 5797 -10893
rect 5797 -10927 5806 -10893
rect 5754 -10936 5806 -10927
rect 5754 -11013 5806 -11004
rect 5754 -11047 5763 -11013
rect 5763 -11047 5797 -11013
rect 5797 -11047 5806 -11013
rect 5754 -11056 5806 -11047
rect 6734 -10893 6786 -10884
rect 6734 -10927 6743 -10893
rect 6743 -10927 6777 -10893
rect 6777 -10927 6786 -10893
rect 6734 -10936 6786 -10927
rect 6884 -11013 6936 -11004
rect 6884 -11047 6893 -11013
rect 6893 -11047 6927 -11013
rect 6927 -11047 6936 -11013
rect 6884 -11056 6936 -11047
rect 7087 -10623 7139 -10614
rect 7087 -10657 7096 -10623
rect 7096 -10657 7130 -10623
rect 7130 -10657 7139 -10623
rect 7087 -10666 7139 -10657
rect 1069 -11243 1121 -11234
rect 1069 -11277 1103 -11243
rect 1103 -11277 1121 -11243
rect 1069 -11286 1121 -11277
rect 5412 -11477 5464 -11468
rect 5412 -11511 5421 -11477
rect 5421 -11511 5455 -11477
rect 5455 -11511 5464 -11477
rect 5412 -11520 5464 -11511
rect 7357 -11510 7409 -11501
rect 7357 -11544 7366 -11510
rect 7366 -11544 7400 -11510
rect 7400 -11544 7409 -11510
rect 7357 -11553 7409 -11544
rect 1069 -11747 1121 -11695
rect 5265 -11704 5317 -11695
rect 5265 -11738 5274 -11704
rect 5274 -11738 5308 -11704
rect 5308 -11738 5317 -11704
rect 5265 -11747 5317 -11738
rect 1595 -11823 1647 -11814
rect 1595 -11857 1604 -11823
rect 1604 -11857 1638 -11823
rect 1638 -11857 1647 -11823
rect 1595 -11866 1647 -11857
rect 1685 -11943 1737 -11934
rect 1685 -11977 1694 -11943
rect 1694 -11977 1728 -11943
rect 1728 -11977 1737 -11943
rect 1685 -11986 1737 -11977
rect 1655 -12063 1707 -12054
rect 1655 -12097 1664 -12063
rect 1664 -12097 1698 -12063
rect 1698 -12097 1707 -12063
rect 1655 -12106 1707 -12097
rect 2965 -11823 3017 -11814
rect 2965 -11857 2974 -11823
rect 2974 -11857 3008 -11823
rect 3008 -11857 3017 -11823
rect 2965 -11866 3017 -11857
rect 2815 -11943 2867 -11934
rect 2815 -11977 2824 -11943
rect 2824 -11977 2858 -11943
rect 2858 -11977 2867 -11943
rect 2815 -11986 2867 -11977
rect 2685 -12063 2737 -12054
rect 2685 -12097 2694 -12063
rect 2694 -12097 2728 -12063
rect 2728 -12097 2737 -12063
rect 2685 -12106 2737 -12097
rect 3735 -12083 3787 -12074
rect 3735 -12117 3744 -12083
rect 3744 -12117 3778 -12083
rect 3778 -12117 3787 -12083
rect 3735 -12126 3787 -12117
rect 4635 -12083 4687 -12074
rect 4635 -12117 4644 -12083
rect 4644 -12117 4678 -12083
rect 4678 -12117 4687 -12083
rect 4635 -12126 4687 -12117
rect 5018 -11910 5070 -11901
rect 5018 -11944 5027 -11910
rect 5027 -11944 5061 -11910
rect 5061 -11944 5070 -11910
rect 5018 -11953 5070 -11944
rect 5194 -12039 5246 -11987
rect 5194 -12106 5246 -12097
rect 5194 -12140 5203 -12106
rect 5203 -12140 5237 -12106
rect 5237 -12140 5246 -12106
rect 5194 -12149 5246 -12140
rect 5195 -12220 5247 -12211
rect 5195 -12254 5204 -12220
rect 5204 -12254 5238 -12220
rect 5238 -12254 5247 -12220
rect 5195 -12263 5247 -12254
rect 5195 -12334 5247 -12325
rect 5195 -12368 5204 -12334
rect 5204 -12368 5238 -12334
rect 5238 -12368 5247 -12334
rect 5195 -12377 5247 -12368
rect 5395 -11829 5447 -11820
rect 5395 -11863 5404 -11829
rect 5404 -11863 5438 -11829
rect 5438 -11863 5447 -11829
rect 5395 -11872 5447 -11863
rect 5495 -11954 5547 -11945
rect 5495 -11988 5504 -11954
rect 5504 -11988 5538 -11954
rect 5538 -11988 5547 -11954
rect 5495 -11997 5547 -11988
rect 5695 -12044 5747 -12035
rect 5695 -12078 5704 -12044
rect 5704 -12078 5738 -12044
rect 5738 -12078 5747 -12044
rect 5695 -12087 5747 -12078
rect 6675 -11834 6727 -11825
rect 6675 -11868 6684 -11834
rect 6684 -11868 6718 -11834
rect 6718 -11868 6727 -11834
rect 6675 -11877 6727 -11868
rect 6795 -11944 6847 -11935
rect 6795 -11978 6804 -11944
rect 6804 -11978 6838 -11944
rect 6838 -11978 6847 -11944
rect 6795 -11987 6847 -11978
rect 7047 -11944 7099 -11935
rect 7047 -11978 7056 -11944
rect 7056 -11978 7090 -11944
rect 7090 -11978 7099 -11944
rect 7047 -11987 7099 -11978
rect 6675 -12044 6727 -12035
rect 6675 -12078 6684 -12044
rect 6684 -12078 6718 -12044
rect 6718 -12078 6727 -12044
rect 6675 -12087 6727 -12078
rect 6805 -12175 6857 -12123
rect 7243 -11834 7295 -11825
rect 7243 -11868 7252 -11834
rect 7252 -11868 7286 -11834
rect 7286 -11868 7295 -11834
rect 7243 -11877 7295 -11868
rect 7289 -12132 7341 -12123
rect 7289 -12166 7298 -12132
rect 7298 -12166 7332 -12132
rect 7332 -12166 7341 -12132
rect 7289 -12175 7341 -12166
rect 5012 -12487 5064 -12478
rect 5012 -12521 5021 -12487
rect 5021 -12521 5055 -12487
rect 5055 -12521 5064 -12487
rect 5012 -12530 5064 -12521
rect 1185 -12763 1237 -12754
rect 1185 -12797 1194 -12763
rect 1194 -12797 1228 -12763
rect 1228 -12797 1237 -12763
rect 1185 -12806 1237 -12797
rect 5106 -12765 5158 -12756
rect 5106 -12799 5115 -12765
rect 5115 -12799 5149 -12765
rect 5149 -12799 5158 -12765
rect 5106 -12808 5158 -12799
<< metal2 >>
rect 1020 2487 1100 2501
rect 1020 2435 1034 2487
rect 1086 2435 1100 2487
rect 228 2372 308 2383
rect 228 2316 240 2372
rect 296 2316 308 2372
rect 228 2303 308 2316
rect 570 2229 650 2240
rect 570 2173 582 2229
rect 638 2173 650 2229
rect 570 2160 650 2173
rect 456 1698 536 1709
rect 456 1642 468 1698
rect 524 1642 536 1698
rect 456 1629 536 1642
rect 342 1538 422 1549
rect 342 1482 354 1538
rect 410 1482 422 1538
rect 342 1469 422 1482
rect 1020 127 1100 2435
rect 1149 1441 1189 2501
rect 2988 2372 3068 2383
rect 1540 2357 1620 2371
rect 1540 2305 1554 2357
rect 1606 2351 1620 2357
rect 2800 2357 2880 2371
rect 2800 2351 2814 2357
rect 1606 2311 2814 2351
rect 1606 2305 1620 2311
rect 1540 2291 1620 2305
rect 2800 2305 2814 2311
rect 2866 2305 2880 2357
rect 2800 2291 2880 2305
rect 2988 2316 3000 2372
rect 3056 2316 3068 2372
rect 5284 2335 5364 2349
rect 5284 2329 5298 2335
rect 2988 2303 3068 2316
rect 3410 2289 5298 2329
rect 1670 2257 1750 2271
rect 1670 2205 1684 2257
rect 1736 2251 1750 2257
rect 3000 2257 3080 2271
rect 3000 2251 3014 2257
rect 1736 2211 3014 2251
rect 1736 2205 1750 2211
rect 1670 2191 1750 2205
rect 3000 2205 3014 2211
rect 3066 2205 3080 2257
rect 3000 2191 3080 2205
rect 3268 2232 3348 2243
rect 3268 2176 3280 2232
rect 3336 2176 3348 2232
rect 1540 2157 1620 2171
rect 1540 2105 1554 2157
rect 1606 2151 1620 2157
rect 3150 2157 3230 2171
rect 3268 2163 3348 2176
rect 3150 2151 3164 2157
rect 1606 2111 3164 2151
rect 1606 2105 1620 2111
rect 1540 2091 1620 2105
rect 3150 2105 3164 2111
rect 3216 2105 3230 2157
rect 3150 2091 3230 2105
rect 1670 2057 1750 2071
rect 1670 2005 1684 2057
rect 1736 2051 1750 2057
rect 2700 2057 2780 2071
rect 2700 2051 2714 2057
rect 1736 2011 2714 2051
rect 1736 2005 1750 2011
rect 1670 1991 1750 2005
rect 2700 2005 2714 2011
rect 2766 2005 2780 2057
rect 2700 1991 2780 2005
rect 3300 2065 3380 2079
rect 3300 2013 3314 2065
rect 3366 2059 3380 2065
rect 3410 2059 3450 2289
rect 5284 2283 5298 2289
rect 5350 2283 5364 2335
rect 5284 2269 5364 2283
rect 3990 2227 4070 2241
rect 3990 2175 4004 2227
rect 4056 2221 4070 2227
rect 5170 2227 5250 2241
rect 5170 2221 5184 2227
rect 4056 2181 5184 2221
rect 4056 2175 4070 2181
rect 3990 2161 4070 2175
rect 5170 2175 5184 2181
rect 5236 2175 5250 2227
rect 5170 2161 5250 2175
rect 3366 2019 3450 2059
rect 3990 2107 4070 2121
rect 3990 2055 4004 2107
rect 4056 2101 4070 2107
rect 4970 2107 5050 2121
rect 4970 2101 4984 2107
rect 4056 2061 4984 2101
rect 4056 2055 4070 2061
rect 3990 2041 4070 2055
rect 4970 2055 4984 2061
rect 5036 2055 5050 2107
rect 4970 2041 5050 2055
rect 3366 2013 3380 2019
rect 3300 1999 3380 2013
rect 5370 1996 5450 2010
rect 3054 1977 3134 1991
rect 3054 1925 3068 1977
rect 3120 1970 3134 1977
rect 5370 1970 5384 1996
rect 3120 1944 5384 1970
rect 5436 1944 5450 1996
rect 3120 1930 5450 1944
rect 3120 1925 3134 1930
rect 3054 1911 3134 1925
rect 1129 1427 1209 1441
rect 1129 1375 1143 1427
rect 1195 1375 1209 1427
rect 1129 1361 1209 1375
rect 1149 1201 1189 1361
rect 1128 1187 1208 1201
rect 1128 1135 1142 1187
rect 1194 1135 1208 1187
rect 1128 1121 1208 1135
rect 1148 189 1188 1121
rect 1670 477 1750 491
rect 1670 425 1684 477
rect 1736 471 1750 477
rect 2650 477 2730 491
rect 2650 471 2664 477
rect 1736 431 2664 471
rect 1736 425 1750 431
rect 1670 411 1750 425
rect 2650 425 2664 431
rect 2716 425 2730 477
rect 2650 411 2730 425
rect 3074 371 3114 1911
rect 3300 1863 3380 1877
rect 3300 1811 3314 1863
rect 3366 1857 3380 1863
rect 3366 1817 3532 1857
rect 3366 1811 3380 1817
rect 3300 1797 3380 1811
rect 3335 1698 3415 1709
rect 3335 1642 3347 1698
rect 3403 1642 3415 1698
rect 3335 1629 3415 1642
rect 3335 1538 3415 1549
rect 3335 1482 3347 1538
rect 3403 1482 3415 1538
rect 3335 1469 3415 1482
rect 3492 571 3532 1817
rect 5328 1547 5408 1561
rect 5328 1495 5342 1547
rect 5394 1495 5408 1547
rect 5328 1481 5408 1495
rect 5073 1188 5153 1202
rect 5073 1136 5087 1188
rect 5139 1136 5153 1188
rect 5073 1122 5153 1136
rect 5093 973 5133 1122
rect 5348 1081 5388 1481
rect 5328 1067 5408 1081
rect 5328 1015 5342 1067
rect 5394 1015 5408 1067
rect 5328 1001 5408 1015
rect 5093 933 5438 973
rect 3560 577 3640 591
rect 3560 571 3574 577
rect 3492 531 3574 571
rect 3560 525 3574 531
rect 3626 525 3640 577
rect 3560 511 3640 525
rect 3990 477 4070 491
rect 3990 425 4004 477
rect 4056 471 4070 477
rect 4970 477 5050 491
rect 4970 471 4984 477
rect 4056 431 4984 471
rect 4056 425 4070 431
rect 3990 411 4070 425
rect 4970 425 4984 431
rect 5036 425 5050 477
rect 4970 411 5050 425
rect 1670 357 1750 371
rect 1670 305 1684 357
rect 1736 351 1750 357
rect 2800 357 2880 371
rect 2800 351 2814 357
rect 1736 311 2814 351
rect 1736 305 1750 311
rect 1670 291 1750 305
rect 2800 305 2814 311
rect 2866 305 2880 357
rect 2800 291 2880 305
rect 3054 357 3134 371
rect 3054 305 3068 357
rect 3120 305 3134 357
rect 3054 291 3134 305
rect 3990 357 4070 371
rect 3990 305 4004 357
rect 4056 351 4070 357
rect 5120 357 5200 371
rect 5120 351 5134 357
rect 4056 311 5134 351
rect 4056 305 4070 311
rect 3990 291 4070 305
rect 5120 305 5134 311
rect 5186 305 5200 357
rect 5120 291 5200 305
rect 1148 149 1231 189
rect 1020 75 1034 127
rect 1086 75 1100 127
rect 1020 61 1100 75
rect 1055 -319 1135 61
rect 1055 -333 1136 -319
rect 1055 -385 1070 -333
rect 1122 -385 1136 -333
rect 1055 -399 1136 -385
rect 684 -458 764 -447
rect 684 -514 696 -458
rect 752 -514 764 -458
rect 684 -527 764 -514
rect 798 -1159 878 -1148
rect 798 -1215 810 -1159
rect 866 -1215 878 -1159
rect 798 -1228 878 -1215
rect 568 -1855 648 -1844
rect 568 -1911 580 -1855
rect 636 -1911 648 -1855
rect 568 -1924 648 -1911
rect 456 -2562 536 -2551
rect 456 -2618 468 -2562
rect 524 -2618 536 -2562
rect 456 -2631 536 -2618
rect 1055 -2693 1135 -399
rect 1191 -1379 1231 149
rect 5136 -193 5216 -179
rect 5136 -245 5150 -193
rect 5202 -245 5216 -193
rect 5136 -259 5216 -245
rect 1540 -463 1620 -449
rect 1540 -515 1554 -463
rect 1606 -469 1620 -463
rect 2800 -463 2880 -449
rect 2800 -469 2814 -463
rect 1606 -509 2814 -469
rect 1606 -515 1620 -509
rect 1540 -529 1620 -515
rect 2800 -515 2814 -509
rect 2866 -515 2880 -463
rect 3860 -458 3940 -447
rect 3860 -514 3872 -458
rect 3928 -514 3940 -458
rect 2800 -529 2880 -515
rect 3572 -529 3652 -515
rect 3860 -527 3940 -514
rect 1670 -563 1750 -549
rect 1670 -615 1684 -563
rect 1736 -569 1750 -563
rect 3000 -563 3080 -549
rect 3000 -569 3014 -563
rect 1736 -609 3014 -569
rect 1736 -615 1750 -609
rect 1670 -629 1750 -615
rect 3000 -615 3014 -609
rect 3066 -615 3080 -563
rect 3572 -581 3586 -529
rect 3638 -555 3652 -529
rect 5048 -550 5128 -536
rect 5048 -555 5062 -550
rect 3638 -581 5062 -555
rect 3572 -595 5062 -581
rect 3000 -629 3080 -615
rect 5048 -602 5062 -595
rect 5114 -602 5128 -550
rect 5048 -616 5128 -602
rect 3572 -640 4996 -626
rect 1540 -663 1620 -649
rect 1540 -715 1554 -663
rect 1606 -669 1620 -663
rect 3150 -663 3230 -649
rect 3150 -669 3164 -663
rect 1606 -709 3164 -669
rect 1606 -715 1620 -709
rect 1540 -729 1620 -715
rect 3150 -715 3164 -709
rect 3216 -715 3230 -663
rect 3572 -692 3586 -640
rect 3638 -666 4996 -640
rect 3638 -692 3652 -666
rect 3572 -706 3652 -692
rect 4956 -667 4996 -666
rect 5048 -659 5128 -645
rect 5048 -667 5062 -659
rect 3150 -729 3230 -715
rect 3860 -713 3940 -699
rect 1670 -763 1750 -749
rect 1670 -815 1684 -763
rect 1736 -769 1750 -763
rect 2700 -763 2780 -749
rect 2700 -769 2714 -763
rect 1736 -809 2714 -769
rect 1736 -815 1750 -809
rect 1670 -829 1750 -815
rect 2700 -815 2714 -809
rect 2766 -815 2780 -763
rect 3860 -765 3874 -713
rect 3926 -719 3940 -713
rect 4760 -713 4840 -699
rect 4956 -707 5062 -667
rect 4760 -719 4774 -713
rect 3926 -759 4774 -719
rect 3926 -765 3940 -759
rect 3860 -779 3940 -765
rect 4760 -765 4774 -759
rect 4826 -765 4840 -713
rect 5048 -711 5062 -707
rect 5114 -711 5128 -659
rect 5048 -725 5128 -711
rect 4760 -779 4840 -765
rect 2700 -829 2780 -815
rect 3314 -1159 3394 -1148
rect 3314 -1215 3326 -1159
rect 3382 -1215 3394 -1159
rect 3314 -1228 3394 -1215
rect 1171 -1393 1251 -1379
rect 1171 -1445 1185 -1393
rect 1237 -1445 1251 -1393
rect 1171 -1459 1251 -1445
rect 1191 -1619 1231 -1459
rect 1171 -1633 1251 -1619
rect 1171 -1685 1185 -1633
rect 1237 -1685 1251 -1633
rect 1171 -1699 1251 -1685
rect 1055 -2745 1069 -2693
rect 1121 -2745 1135 -2693
rect 1055 -3154 1135 -2745
rect 1055 -3206 1069 -3154
rect 1121 -3206 1135 -3154
rect 1055 -3220 1135 -3206
rect 1191 -4199 1231 -1699
rect 3314 -1854 3394 -1843
rect 3314 -1910 3326 -1854
rect 3382 -1910 3394 -1854
rect 3314 -1923 3394 -1910
rect 1670 -2263 1750 -2249
rect 1670 -2315 1684 -2263
rect 1736 -2269 1750 -2263
rect 2700 -2263 2780 -2249
rect 2700 -2269 2714 -2263
rect 1736 -2309 2714 -2269
rect 1736 -2315 1750 -2309
rect 1670 -2329 1750 -2315
rect 2700 -2315 2714 -2309
rect 2766 -2315 2780 -2263
rect 2700 -2329 2780 -2315
rect 3860 -2313 3940 -2299
rect 1540 -2363 1620 -2349
rect 1540 -2415 1554 -2363
rect 1606 -2369 1620 -2363
rect 3150 -2363 3230 -2349
rect 3150 -2369 3164 -2363
rect 1606 -2409 3164 -2369
rect 1606 -2415 1620 -2409
rect 1540 -2429 1620 -2415
rect 3150 -2415 3164 -2409
rect 3216 -2415 3230 -2363
rect 3860 -2365 3874 -2313
rect 3926 -2319 3940 -2313
rect 4760 -2313 4840 -2299
rect 4760 -2319 4774 -2313
rect 3926 -2359 4774 -2319
rect 3926 -2365 3940 -2359
rect 3150 -2429 3230 -2415
rect 3572 -2384 3652 -2370
rect 3860 -2379 3940 -2365
rect 4760 -2365 4774 -2359
rect 4826 -2365 4840 -2313
rect 5048 -2351 5128 -2337
rect 5048 -2358 5062 -2351
rect 4760 -2379 4840 -2365
rect 3572 -2436 3586 -2384
rect 3638 -2410 3652 -2384
rect 4900 -2398 5062 -2358
rect 4900 -2410 4940 -2398
rect 3638 -2436 4940 -2410
rect 5048 -2403 5062 -2398
rect 5114 -2403 5128 -2351
rect 5048 -2417 5128 -2403
rect 1670 -2463 1750 -2449
rect 1670 -2515 1684 -2463
rect 1736 -2469 1750 -2463
rect 3000 -2463 3080 -2449
rect 3572 -2450 4940 -2436
rect 3000 -2469 3014 -2463
rect 1736 -2509 3014 -2469
rect 1736 -2515 1750 -2509
rect 1670 -2529 1750 -2515
rect 3000 -2515 3014 -2509
rect 3066 -2515 3080 -2463
rect 5048 -2459 5128 -2445
rect 5048 -2483 5062 -2459
rect 3000 -2529 3080 -2515
rect 3572 -2497 5062 -2483
rect 3572 -2549 3586 -2497
rect 3638 -2511 5062 -2497
rect 5114 -2511 5128 -2459
rect 3638 -2523 5128 -2511
rect 3638 -2549 3652 -2523
rect 5048 -2525 5128 -2523
rect 1540 -2563 1620 -2549
rect 1540 -2615 1554 -2563
rect 1606 -2569 1620 -2563
rect 2800 -2563 2880 -2549
rect 3572 -2563 3652 -2549
rect 3860 -2562 3940 -2551
rect 2800 -2569 2814 -2563
rect 1606 -2609 2814 -2569
rect 1606 -2615 1620 -2609
rect 1540 -2629 1620 -2615
rect 2800 -2615 2814 -2609
rect 2866 -2615 2880 -2563
rect 2800 -2629 2880 -2615
rect 3860 -2618 3872 -2562
rect 3928 -2618 3940 -2562
rect 5156 -2576 5196 -259
rect 3860 -2631 3940 -2618
rect 5112 -2616 5196 -2576
rect 5251 -449 5331 -319
rect 5251 -501 5265 -449
rect 5317 -501 5331 -449
rect 1581 -3273 1661 -3259
rect 1581 -3325 1595 -3273
rect 1647 -3279 1661 -3273
rect 2951 -3273 3031 -3259
rect 2951 -3279 2965 -3273
rect 1647 -3319 2965 -3279
rect 1647 -3325 1661 -3319
rect 1581 -3339 1661 -3325
rect 2951 -3325 2965 -3319
rect 3017 -3325 3031 -3273
rect 2951 -3339 3031 -3325
rect 5004 -3360 5084 -3346
rect 1671 -3393 1751 -3379
rect 1671 -3445 1685 -3393
rect 1737 -3399 1751 -3393
rect 2801 -3393 2881 -3379
rect 2801 -3399 2815 -3393
rect 1737 -3439 2815 -3399
rect 1737 -3445 1751 -3439
rect 1671 -3459 1751 -3445
rect 2801 -3445 2815 -3439
rect 2867 -3445 2881 -3393
rect 5004 -3412 5018 -3360
rect 5070 -3412 5084 -3360
rect 5004 -3426 5084 -3412
rect 2801 -3459 2881 -3445
rect 1641 -3513 1721 -3499
rect 1641 -3565 1655 -3513
rect 1707 -3519 1721 -3513
rect 2671 -3513 2751 -3499
rect 2671 -3519 2685 -3513
rect 1707 -3559 2685 -3519
rect 1707 -3565 1721 -3559
rect 1641 -3579 1721 -3565
rect 2671 -3565 2685 -3559
rect 2737 -3565 2751 -3513
rect 2671 -3579 2751 -3565
rect 3721 -3533 3801 -3519
rect 3721 -3585 3735 -3533
rect 3787 -3539 3801 -3533
rect 4621 -3533 4701 -3519
rect 4621 -3539 4635 -3533
rect 3787 -3579 4635 -3539
rect 3787 -3585 3801 -3579
rect 3721 -3599 3801 -3585
rect 4621 -3585 4635 -3579
rect 4687 -3585 4701 -3533
rect 4621 -3599 4701 -3585
rect 5023 -3923 5063 -3426
rect 4998 -3937 5078 -3923
rect 4998 -3989 5012 -3937
rect 5064 -3989 5078 -3937
rect 4998 -4003 5078 -3989
rect 3051 -4093 3131 -4079
rect 3051 -4145 3065 -4093
rect 3117 -4097 3131 -4093
rect 4801 -4093 4881 -4079
rect 3117 -4137 3300 -4097
rect 3117 -4145 3131 -4137
rect 3051 -4159 3131 -4145
rect 1171 -4213 1251 -4199
rect 1171 -4219 1185 -4213
rect 1060 -4259 1185 -4219
rect 1060 -4522 1100 -4259
rect 1171 -4265 1185 -4259
rect 1237 -4265 1251 -4213
rect 1171 -4279 1251 -4265
rect 1041 -4536 1121 -4522
rect 1041 -4588 1055 -4536
rect 1107 -4588 1121 -4536
rect 1041 -4602 1121 -4588
rect 1062 -5920 1102 -4602
rect 3260 -4640 3300 -4137
rect 4801 -4145 4815 -4093
rect 4867 -4145 4881 -4093
rect 4801 -4640 4881 -4145
rect 5018 -4540 5058 -4003
rect 5112 -4201 5152 -2616
rect 5251 -3154 5331 -501
rect 5398 -1379 5438 933
rect 5478 141 5518 2501
rect 5762 1441 5802 2501
rect 5830 2487 5910 2501
rect 5830 2435 5844 2487
rect 5896 2435 5910 2487
rect 5830 2421 5910 2435
rect 5742 1427 5822 1441
rect 5742 1375 5756 1427
rect 5808 1375 5822 1427
rect 5742 1361 5822 1375
rect 5942 1201 5982 2501
rect 6010 2257 6090 2271
rect 6010 2205 6024 2257
rect 6076 2251 6090 2257
rect 7140 2257 7220 2271
rect 7140 2251 7154 2257
rect 6076 2211 7154 2251
rect 6076 2205 6090 2211
rect 6010 2191 6090 2205
rect 7140 2205 7154 2211
rect 7206 2205 7220 2257
rect 7140 2191 7220 2205
rect 6010 2137 6090 2151
rect 6010 2085 6024 2137
rect 6076 2131 6090 2137
rect 6990 2137 7070 2151
rect 6990 2131 7004 2137
rect 6076 2091 7004 2131
rect 6076 2085 6090 2091
rect 6010 2071 6090 2085
rect 6990 2085 7004 2091
rect 7056 2085 7070 2137
rect 6990 2071 7070 2085
rect 7340 1987 7420 2001
rect 7340 1935 7354 1987
rect 7406 1935 7420 1987
rect 7340 1921 7420 1935
rect 5922 1187 6002 1201
rect 5922 1135 5936 1187
rect 5988 1135 6002 1187
rect 5922 1121 6002 1135
rect 7366 911 7406 1921
rect 5555 897 5635 911
rect 5555 845 5569 897
rect 5621 891 5635 897
rect 7090 897 7170 911
rect 7090 891 7104 897
rect 5621 851 7104 891
rect 5621 845 5635 851
rect 5555 831 5635 845
rect 7090 845 7104 851
rect 7156 845 7170 897
rect 7090 831 7170 845
rect 7348 897 7428 911
rect 7348 845 7362 897
rect 7414 845 7428 897
rect 7348 831 7428 845
rect 5660 747 5740 761
rect 5660 695 5674 747
rect 5726 741 5740 747
rect 5726 701 7511 741
rect 5726 695 5740 701
rect 5660 681 5740 695
rect 5660 627 5740 641
rect 5660 575 5674 627
rect 5726 621 5740 627
rect 5726 581 7511 621
rect 5726 575 5740 581
rect 5660 561 5740 575
rect 5930 507 6010 521
rect 5930 455 5944 507
rect 5996 501 6010 507
rect 6910 507 6990 521
rect 6910 501 6924 507
rect 5996 461 6924 501
rect 5996 455 6010 461
rect 5930 441 6010 455
rect 6910 455 6924 461
rect 6976 455 6990 507
rect 6910 441 6990 455
rect 5730 387 5810 401
rect 5730 335 5744 387
rect 5796 381 5810 387
rect 6910 387 6990 401
rect 6910 381 6924 387
rect 5796 341 6924 381
rect 5796 335 5810 341
rect 5730 321 5810 335
rect 6910 335 6924 341
rect 6976 335 6990 387
rect 6910 321 6990 335
rect 5478 127 5558 141
rect 5478 75 5492 127
rect 5544 75 5558 127
rect 5478 61 5558 75
rect 5740 127 5820 141
rect 5740 75 5754 127
rect 5806 75 5820 127
rect 5740 -437 5820 75
rect 6990 -333 7070 -319
rect 6990 -385 7004 -333
rect 7056 -385 7070 -333
rect 6990 -399 7070 -385
rect 5472 -451 5820 -437
rect 5472 -503 5486 -451
rect 5538 -503 5820 -451
rect 5472 -517 5820 -503
rect 5740 -563 5820 -549
rect 5740 -615 5754 -563
rect 5806 -569 5820 -563
rect 6870 -563 6950 -549
rect 6870 -569 6884 -563
rect 5806 -609 6884 -569
rect 5806 -615 5820 -609
rect 5740 -629 5820 -615
rect 6870 -615 6884 -609
rect 6936 -615 6950 -563
rect 6870 -629 6950 -615
rect 5740 -683 5820 -669
rect 5740 -735 5754 -683
rect 5806 -689 5820 -683
rect 6720 -683 6800 -669
rect 6720 -689 6734 -683
rect 5806 -729 6734 -689
rect 5806 -735 5820 -729
rect 5740 -749 5820 -735
rect 6720 -735 6734 -729
rect 6786 -735 6800 -683
rect 6720 -749 6800 -735
rect 7073 -953 7153 -939
rect 7073 -1005 7087 -953
rect 7139 -959 7153 -953
rect 7139 -999 7269 -959
rect 7139 -1005 7153 -999
rect 7073 -1019 7153 -1005
rect 6970 -1273 7050 -1259
rect 6970 -1325 6984 -1273
rect 7036 -1325 7050 -1273
rect 5398 -1393 5478 -1379
rect 5398 -1445 5412 -1393
rect 5464 -1445 5478 -1393
rect 5398 -1459 5478 -1445
rect 5418 -1618 5458 -1459
rect 5398 -1632 5478 -1618
rect 5398 -1684 5412 -1632
rect 5464 -1684 5478 -1632
rect 5398 -1698 5478 -1684
rect 5418 -2913 5458 -1698
rect 6970 -1753 7050 -1325
rect 6970 -1805 6984 -1753
rect 7036 -1805 7050 -1753
rect 6970 -1819 7050 -1805
rect 7073 -2073 7153 -2059
rect 7073 -2125 7087 -2073
rect 7139 -2125 7153 -2073
rect 7073 -2139 7153 -2125
rect 5740 -2343 5820 -2329
rect 5740 -2395 5754 -2343
rect 5806 -2349 5820 -2343
rect 6720 -2343 6800 -2329
rect 6720 -2349 6734 -2343
rect 5806 -2389 6734 -2349
rect 5806 -2395 5820 -2389
rect 5740 -2409 5820 -2395
rect 6720 -2395 6734 -2389
rect 6786 -2395 6800 -2343
rect 6720 -2409 6800 -2395
rect 5740 -2463 5820 -2449
rect 5740 -2515 5754 -2463
rect 5806 -2469 5820 -2463
rect 6870 -2463 6950 -2449
rect 6870 -2469 6884 -2463
rect 5806 -2509 6884 -2469
rect 5806 -2515 5820 -2509
rect 5740 -2529 5820 -2515
rect 6870 -2515 6884 -2509
rect 6936 -2515 6950 -2463
rect 6870 -2529 6950 -2515
rect 5398 -2927 5478 -2913
rect 5398 -2979 5412 -2927
rect 5464 -2979 5478 -2927
rect 5398 -2993 5478 -2979
rect 5251 -3206 5265 -3154
rect 5317 -3206 5331 -3154
rect 5251 -3220 5331 -3206
rect 5381 -3279 5461 -3265
rect 5381 -3331 5395 -3279
rect 5447 -3290 5461 -3279
rect 6661 -3284 6741 -3270
rect 6661 -3290 6675 -3284
rect 5447 -3330 6675 -3290
rect 5447 -3331 5461 -3330
rect 5381 -3345 5461 -3331
rect 6661 -3336 6675 -3330
rect 6727 -3336 6741 -3284
rect 6661 -3350 6741 -3336
rect 7073 -3380 7113 -2139
rect 7229 -3270 7269 -999
rect 7343 -2960 7423 -2946
rect 7343 -3012 7357 -2960
rect 7409 -3012 7423 -2960
rect 7343 -3026 7423 -3012
rect 7229 -3284 7309 -3270
rect 7229 -3336 7243 -3284
rect 7295 -3336 7309 -3284
rect 7229 -3350 7309 -3336
rect 5481 -3400 5561 -3390
rect 6781 -3394 6861 -3380
rect 6781 -3400 6795 -3394
rect 5481 -3404 6795 -3400
rect 5180 -3446 5260 -3432
rect 5180 -3498 5194 -3446
rect 5246 -3452 5260 -3446
rect 5246 -3492 5353 -3452
rect 5481 -3456 5495 -3404
rect 5547 -3440 6795 -3404
rect 5547 -3456 5561 -3440
rect 5481 -3470 5561 -3456
rect 6781 -3446 6795 -3440
rect 6847 -3446 6861 -3394
rect 6781 -3460 6861 -3446
rect 7033 -3394 7113 -3380
rect 7033 -3446 7047 -3394
rect 7099 -3446 7113 -3394
rect 7033 -3460 7113 -3446
rect 5246 -3498 5260 -3492
rect 5180 -3512 5260 -3498
rect 5313 -3500 5353 -3492
rect 5681 -3494 5761 -3480
rect 5681 -3500 5695 -3494
rect 5313 -3540 5695 -3500
rect 5180 -3556 5260 -3542
rect 5180 -3608 5194 -3556
rect 5246 -3588 5260 -3556
rect 5681 -3546 5695 -3540
rect 5747 -3500 5761 -3494
rect 6661 -3494 6741 -3480
rect 6661 -3500 6675 -3494
rect 5747 -3540 6675 -3500
rect 5747 -3546 5761 -3540
rect 5681 -3560 5761 -3546
rect 6661 -3546 6675 -3540
rect 6727 -3546 6741 -3494
rect 6661 -3560 6741 -3546
rect 6791 -3582 6871 -3568
rect 6791 -3588 6805 -3582
rect 5246 -3608 6805 -3588
rect 5180 -3628 6805 -3608
rect 6791 -3634 6805 -3628
rect 6857 -3634 6871 -3582
rect 6791 -3648 6871 -3634
rect 7275 -3582 7355 -3568
rect 7275 -3634 7289 -3582
rect 7341 -3590 7355 -3582
rect 7383 -3590 7423 -3026
rect 7341 -3630 7423 -3590
rect 7341 -3634 7355 -3630
rect 7275 -3648 7355 -3634
rect 5181 -3670 5261 -3656
rect 5181 -3722 5195 -3670
rect 5247 -3676 5261 -3670
rect 5247 -3716 7291 -3676
rect 5247 -3722 5261 -3716
rect 5181 -3736 5261 -3722
rect 5181 -3780 5261 -3770
rect 5181 -3784 7291 -3780
rect 5181 -3836 5195 -3784
rect 5247 -3820 7291 -3784
rect 5247 -3836 5261 -3820
rect 5181 -3850 5261 -3836
rect 7141 -4093 7221 -4079
rect 7141 -4145 7155 -4093
rect 7207 -4099 7221 -4093
rect 7207 -4139 7420 -4099
rect 7207 -4145 7221 -4139
rect 7141 -4159 7221 -4145
rect 5092 -4215 5172 -4201
rect 5092 -4267 5106 -4215
rect 5158 -4219 5172 -4215
rect 5158 -4259 5372 -4219
rect 5158 -4267 5172 -4259
rect 5092 -4281 5172 -4267
rect 5332 -4520 5372 -4259
rect 5115 -4534 5195 -4520
rect 5115 -4540 5129 -4534
rect 5018 -4580 5129 -4540
rect 5115 -4586 5129 -4580
rect 5181 -4586 5195 -4534
rect 5115 -4600 5195 -4586
rect 5312 -4534 5392 -4520
rect 5312 -4586 5326 -4534
rect 5378 -4586 5392 -4534
rect 5312 -4600 5392 -4586
rect 3240 -4654 3320 -4640
rect 3240 -4706 3254 -4654
rect 3306 -4706 3320 -4654
rect 3240 -4720 3320 -4706
rect 4801 -4654 5081 -4640
rect 4801 -4706 5015 -4654
rect 5067 -4706 5081 -4654
rect 4801 -4720 5081 -4706
rect 3921 -5214 4001 -5200
rect 3921 -5266 3935 -5214
rect 3987 -5220 4001 -5214
rect 4821 -5214 4901 -5200
rect 4821 -5220 4835 -5214
rect 3987 -5260 4835 -5220
rect 3987 -5266 4001 -5260
rect 3921 -5280 4001 -5266
rect 4821 -5266 4835 -5260
rect 4887 -5266 4901 -5214
rect 4821 -5280 4901 -5266
rect 5135 -5373 5175 -4600
rect 5115 -5387 5195 -5373
rect 1130 -5423 1210 -5409
rect 1130 -5475 1144 -5423
rect 1196 -5429 1210 -5423
rect 2690 -5423 2770 -5409
rect 2690 -5429 2704 -5423
rect 1196 -5469 2704 -5429
rect 1196 -5475 1210 -5469
rect 1130 -5489 1210 -5475
rect 2690 -5475 2704 -5469
rect 2756 -5475 2770 -5423
rect 5115 -5439 5129 -5387
rect 5181 -5439 5195 -5387
rect 5115 -5453 5195 -5439
rect 2690 -5489 2770 -5475
rect 1130 -5543 1210 -5529
rect 1130 -5595 1144 -5543
rect 1196 -5549 1210 -5543
rect 2840 -5543 2920 -5529
rect 2840 -5549 2854 -5543
rect 1196 -5589 2854 -5549
rect 1196 -5595 1210 -5589
rect 1130 -5609 1210 -5595
rect 2840 -5595 2854 -5589
rect 2906 -5595 2920 -5543
rect 2840 -5609 2920 -5595
rect 1130 -5663 1210 -5649
rect 1130 -5715 1144 -5663
rect 1196 -5669 1210 -5663
rect 2990 -5663 3070 -5649
rect 2990 -5669 3004 -5663
rect 1196 -5709 3004 -5669
rect 1196 -5715 1210 -5709
rect 1130 -5729 1210 -5715
rect 2990 -5715 3004 -5709
rect 3056 -5715 3070 -5663
rect 2990 -5729 3070 -5715
rect 1130 -5783 1210 -5769
rect 1130 -5835 1144 -5783
rect 1196 -5789 1210 -5783
rect 3140 -5783 3220 -5769
rect 3140 -5789 3154 -5783
rect 1196 -5829 3154 -5789
rect 1196 -5835 1210 -5829
rect 1130 -5849 1210 -5835
rect 3140 -5835 3154 -5829
rect 3206 -5835 3220 -5783
rect 3140 -5849 3220 -5835
rect 1062 -5960 1552 -5920
rect 570 -6181 650 -6168
rect 570 -6237 582 -6181
rect 638 -6237 650 -6181
rect 570 -6248 650 -6237
rect 456 -6912 536 -6899
rect 456 -6968 468 -6912
rect 524 -6968 536 -6912
rect 456 -6979 536 -6968
rect 1512 -7100 1552 -5960
rect 1580 -6184 1660 -6170
rect 1580 -6236 1594 -6184
rect 1646 -6190 1660 -6184
rect 2840 -6184 2920 -6170
rect 2840 -6190 2854 -6184
rect 1646 -6230 2854 -6190
rect 1646 -6236 1660 -6230
rect 1580 -6250 1660 -6236
rect 2840 -6236 2854 -6230
rect 2906 -6236 2920 -6184
rect 2840 -6250 2920 -6236
rect 3920 -6181 4000 -6168
rect 3920 -6237 3932 -6181
rect 3988 -6237 4000 -6181
rect 3920 -6248 4000 -6237
rect 1710 -6284 1790 -6270
rect 1710 -6336 1724 -6284
rect 1776 -6290 1790 -6284
rect 3040 -6284 3120 -6270
rect 3040 -6290 3054 -6284
rect 1776 -6330 3054 -6290
rect 1776 -6336 1790 -6330
rect 1710 -6350 1790 -6336
rect 3040 -6336 3054 -6330
rect 3106 -6336 3120 -6284
rect 3040 -6350 3120 -6336
rect 3632 -6284 3712 -6270
rect 3632 -6336 3646 -6284
rect 3698 -6290 3712 -6284
rect 4820 -6284 4900 -6270
rect 4820 -6290 4834 -6284
rect 3698 -6330 4834 -6290
rect 3698 -6336 3712 -6330
rect 3632 -6350 3712 -6336
rect 4820 -6336 4834 -6330
rect 4886 -6336 4900 -6284
rect 4820 -6350 4900 -6336
rect 1580 -6384 1660 -6370
rect 1580 -6436 1594 -6384
rect 1646 -6390 1660 -6384
rect 3190 -6384 3270 -6370
rect 3190 -6390 3204 -6384
rect 1646 -6430 3204 -6390
rect 1646 -6436 1660 -6430
rect 1580 -6450 1660 -6436
rect 3190 -6436 3204 -6430
rect 3256 -6436 3270 -6384
rect 3190 -6450 3270 -6436
rect 3920 -6434 4000 -6420
rect 1710 -6484 1790 -6470
rect 1710 -6536 1724 -6484
rect 1776 -6490 1790 -6484
rect 2740 -6484 2820 -6470
rect 2740 -6490 2754 -6484
rect 1776 -6530 2754 -6490
rect 1776 -6536 1790 -6530
rect 1710 -6550 1790 -6536
rect 2740 -6536 2754 -6530
rect 2806 -6536 2820 -6484
rect 3920 -6486 3934 -6434
rect 3986 -6440 4000 -6434
rect 4820 -6434 4900 -6420
rect 4820 -6440 4834 -6434
rect 3986 -6480 4834 -6440
rect 3986 -6486 4000 -6480
rect 3920 -6500 4000 -6486
rect 4820 -6486 4834 -6480
rect 4886 -6486 4900 -6434
rect 4820 -6500 4900 -6486
rect 2740 -6550 2820 -6536
rect 3631 -6843 3711 -6829
rect 3631 -6895 3645 -6843
rect 3697 -6850 3711 -6843
rect 5108 -6844 5188 -6830
rect 5108 -6850 5122 -6844
rect 3697 -6890 5122 -6850
rect 3697 -6895 3711 -6890
rect 3354 -6912 3434 -6899
rect 3631 -6909 3711 -6895
rect 5108 -6896 5122 -6890
rect 5174 -6896 5188 -6844
rect 5108 -6910 5188 -6896
rect 3354 -6968 3366 -6912
rect 3422 -6968 3434 -6912
rect 3354 -6979 3434 -6968
rect 2940 -6994 3020 -6980
rect 2940 -7046 2954 -6994
rect 3006 -7046 3020 -6994
rect 2940 -7060 3020 -7046
rect 1492 -7114 1572 -7100
rect 1492 -7166 1506 -7114
rect 1558 -7166 1572 -7114
rect 1492 -7180 1572 -7166
rect 1512 -7340 1552 -7180
rect 1492 -7354 1572 -7340
rect 1492 -7406 1506 -7354
rect 1558 -7406 1572 -7354
rect 1492 -7420 1572 -7406
rect 228 -7550 308 -7537
rect 228 -7606 240 -7550
rect 296 -7606 308 -7550
rect 228 -7617 308 -7606
rect 342 -8285 422 -8272
rect 342 -8341 354 -8285
rect 410 -8341 422 -8285
rect 342 -8352 422 -8341
rect 1055 -8414 1200 -8400
rect 1055 -8466 1134 -8414
rect 1186 -8466 1200 -8414
rect 1055 -8480 1200 -8466
rect 1055 -8860 1135 -8480
rect 1512 -8642 1552 -7420
rect 2960 -7460 3000 -7060
rect 2940 -7474 3020 -7460
rect 2940 -7526 2954 -7474
rect 3006 -7526 3020 -7474
rect 2940 -7540 3020 -7526
rect 3354 -7550 3434 -7537
rect 3354 -7606 3366 -7550
rect 3422 -7606 3434 -7550
rect 3354 -7617 3434 -7606
rect 1710 -7984 1790 -7970
rect 1710 -8036 1724 -7984
rect 1776 -7990 1790 -7984
rect 2740 -7984 2820 -7970
rect 2740 -7990 2754 -7984
rect 1776 -8030 2754 -7990
rect 1776 -8036 1790 -8030
rect 1710 -8050 1790 -8036
rect 2740 -8036 2754 -8030
rect 2806 -8036 2820 -7984
rect 2740 -8050 2820 -8036
rect 3920 -8034 4000 -8020
rect 1580 -8084 1660 -8070
rect 1580 -8136 1594 -8084
rect 1646 -8090 1660 -8084
rect 3190 -8084 3270 -8070
rect 3190 -8090 3204 -8084
rect 1646 -8130 3204 -8090
rect 1646 -8136 1660 -8130
rect 1580 -8150 1660 -8136
rect 3190 -8136 3204 -8130
rect 3256 -8136 3270 -8084
rect 3920 -8086 3934 -8034
rect 3986 -8040 4000 -8034
rect 4820 -8034 4900 -8020
rect 4820 -8040 4834 -8034
rect 3986 -8080 4834 -8040
rect 3986 -8086 4000 -8080
rect 3190 -8150 3270 -8136
rect 3632 -8110 3712 -8096
rect 3920 -8100 4000 -8086
rect 4820 -8086 4834 -8080
rect 4886 -8086 4900 -8034
rect 4820 -8100 4900 -8086
rect 3632 -8162 3646 -8110
rect 3698 -8129 3712 -8110
rect 5108 -8103 5188 -8089
rect 5108 -8129 5122 -8103
rect 3698 -8155 5122 -8129
rect 5174 -8155 5188 -8103
rect 3698 -8162 5188 -8155
rect 3632 -8169 5188 -8162
rect 1710 -8184 1790 -8170
rect 1710 -8236 1724 -8184
rect 1776 -8190 1790 -8184
rect 3040 -8184 3120 -8170
rect 3632 -8176 3712 -8169
rect 3040 -8190 3054 -8184
rect 1776 -8230 3054 -8190
rect 1776 -8236 1790 -8230
rect 1710 -8250 1790 -8236
rect 3040 -8236 3054 -8230
rect 3106 -8236 3120 -8184
rect 3040 -8250 3120 -8236
rect 3632 -8218 5188 -8204
rect 3632 -8270 3646 -8218
rect 3698 -8244 5122 -8218
rect 3698 -8270 3712 -8244
rect 1580 -8284 1660 -8270
rect 1580 -8336 1594 -8284
rect 1646 -8290 1660 -8284
rect 2840 -8284 2920 -8270
rect 3632 -8284 3712 -8270
rect 5108 -8270 5122 -8244
rect 5174 -8270 5188 -8218
rect 2840 -8290 2854 -8284
rect 1646 -8330 2854 -8290
rect 1646 -8336 1660 -8330
rect 1580 -8350 1660 -8336
rect 2840 -8336 2854 -8330
rect 2906 -8336 2920 -8284
rect 2840 -8350 2920 -8336
rect 3920 -8285 4000 -8272
rect 5108 -8284 5188 -8270
rect 3920 -8341 3932 -8285
rect 3988 -8341 4000 -8285
rect 3920 -8352 4000 -8341
rect 5332 -8460 5372 -4600
rect 7380 -4640 7420 -4139
rect 7360 -4654 7440 -4640
rect 7360 -4706 7374 -4654
rect 7426 -4706 7440 -4654
rect 7360 -4720 7440 -4706
rect 5400 -4954 5480 -4940
rect 5400 -5006 5414 -4954
rect 5466 -4960 5480 -4954
rect 5466 -5000 7551 -4960
rect 5466 -5006 5480 -5000
rect 5400 -5020 5480 -5006
rect 5400 -5074 5480 -5060
rect 5400 -5126 5414 -5074
rect 5466 -5085 5480 -5074
rect 5466 -5125 7551 -5085
rect 5466 -5126 5480 -5125
rect 5400 -5140 5480 -5126
rect 7010 -5167 7090 -5153
rect 7010 -5172 7024 -5167
rect 5508 -5188 7024 -5172
rect 5400 -5202 7024 -5188
rect 5400 -5254 5414 -5202
rect 5466 -5212 7024 -5202
rect 5466 -5228 5548 -5212
rect 7010 -5219 7024 -5212
rect 7076 -5219 7090 -5167
rect 5466 -5254 5480 -5228
rect 7010 -5233 7090 -5219
rect 7494 -5167 7574 -5153
rect 7494 -5219 7508 -5167
rect 7560 -5219 7574 -5167
rect 7494 -5233 7574 -5219
rect 5400 -5268 5480 -5254
rect 5900 -5254 5980 -5240
rect 5900 -5260 5914 -5254
rect 5508 -5300 5914 -5260
rect 5508 -5303 5548 -5300
rect 5400 -5317 5548 -5303
rect 5400 -5369 5414 -5317
rect 5466 -5343 5548 -5317
rect 5900 -5306 5914 -5300
rect 5966 -5260 5980 -5254
rect 6880 -5254 6960 -5240
rect 6880 -5260 6894 -5254
rect 5966 -5300 6894 -5260
rect 5966 -5306 5980 -5300
rect 5900 -5320 5980 -5306
rect 6880 -5306 6894 -5300
rect 6946 -5306 6960 -5254
rect 6880 -5320 6960 -5306
rect 5466 -5369 5480 -5343
rect 5400 -5383 5480 -5369
rect 5700 -5344 5780 -5330
rect 5700 -5396 5714 -5344
rect 5766 -5360 5780 -5344
rect 7000 -5354 7080 -5340
rect 7000 -5360 7014 -5354
rect 5766 -5396 7014 -5360
rect 5700 -5400 7014 -5396
rect 5700 -5410 5780 -5400
rect 7000 -5406 7014 -5400
rect 7066 -5406 7080 -5354
rect 7000 -5420 7080 -5406
rect 7132 -5353 7212 -5339
rect 7132 -5405 7146 -5353
rect 7198 -5405 7212 -5353
rect 7132 -5419 7212 -5405
rect 5600 -5469 5680 -5455
rect 5600 -5521 5614 -5469
rect 5666 -5470 5680 -5469
rect 6880 -5464 6960 -5450
rect 6880 -5470 6894 -5464
rect 5666 -5510 6894 -5470
rect 5666 -5521 5680 -5510
rect 5600 -5535 5680 -5521
rect 6880 -5516 6894 -5510
rect 6946 -5516 6960 -5464
rect 6880 -5530 6960 -5516
rect 5566 -5594 5646 -5580
rect 5566 -5646 5580 -5594
rect 5632 -5646 5646 -5594
rect 5458 -5820 5538 -5806
rect 5458 -5872 5472 -5820
rect 5524 -5872 5538 -5820
rect 5458 -5886 5538 -5872
rect 5478 -7100 5518 -5886
rect 5456 -7114 5536 -7100
rect 5456 -7166 5470 -7114
rect 5522 -7166 5536 -7114
rect 5456 -7180 5536 -7166
rect 5478 -7340 5518 -7180
rect 5458 -7354 5538 -7340
rect 5458 -7406 5472 -7354
rect 5524 -7406 5538 -7354
rect 5458 -7420 5538 -7406
rect 1191 -8682 1552 -8642
rect 5156 -8500 5372 -8460
rect 1055 -8874 1136 -8860
rect 1055 -8926 1070 -8874
rect 1122 -8926 1136 -8874
rect 1055 -8940 1136 -8926
rect 798 -9000 878 -8989
rect 798 -9056 810 -9000
rect 866 -9056 878 -9000
rect 798 -9069 878 -9056
rect 684 -9700 764 -9689
rect 684 -9756 696 -9700
rect 752 -9756 764 -9700
rect 684 -9769 764 -9756
rect 342 -10396 422 -10385
rect 342 -10452 354 -10396
rect 410 -10452 422 -10396
rect 342 -10465 422 -10452
rect 228 -11103 308 -11092
rect 228 -11159 240 -11103
rect 296 -11159 308 -11103
rect 228 -11172 308 -11159
rect 1055 -11234 1135 -8940
rect 1191 -9920 1231 -8682
rect 1540 -9004 1620 -8990
rect 1540 -9056 1554 -9004
rect 1606 -9010 1620 -9004
rect 2800 -9004 2880 -8990
rect 2800 -9010 2814 -9004
rect 1606 -9050 2814 -9010
rect 1606 -9056 1620 -9050
rect 1540 -9070 1620 -9056
rect 2800 -9056 2814 -9050
rect 2866 -9056 2880 -9004
rect 3860 -8999 3940 -8988
rect 3860 -9055 3872 -8999
rect 3928 -9055 3940 -8999
rect 2800 -9070 2880 -9056
rect 3572 -9070 3652 -9056
rect 3860 -9068 3940 -9055
rect 1670 -9104 1750 -9090
rect 1670 -9156 1684 -9104
rect 1736 -9110 1750 -9104
rect 3000 -9104 3080 -9090
rect 3000 -9110 3014 -9104
rect 1736 -9150 3014 -9110
rect 1736 -9156 1750 -9150
rect 1670 -9170 1750 -9156
rect 3000 -9156 3014 -9150
rect 3066 -9156 3080 -9104
rect 3572 -9122 3586 -9070
rect 3638 -9096 3652 -9070
rect 5048 -9091 5128 -9077
rect 5048 -9096 5062 -9091
rect 3638 -9122 5062 -9096
rect 3572 -9136 5062 -9122
rect 3000 -9170 3080 -9156
rect 5048 -9143 5062 -9136
rect 5114 -9143 5128 -9091
rect 5048 -9157 5128 -9143
rect 3572 -9181 4996 -9167
rect 1540 -9204 1620 -9190
rect 1540 -9256 1554 -9204
rect 1606 -9210 1620 -9204
rect 3150 -9204 3230 -9190
rect 3150 -9210 3164 -9204
rect 1606 -9250 3164 -9210
rect 1606 -9256 1620 -9250
rect 1540 -9270 1620 -9256
rect 3150 -9256 3164 -9250
rect 3216 -9256 3230 -9204
rect 3572 -9233 3586 -9181
rect 3638 -9207 4996 -9181
rect 3638 -9233 3652 -9207
rect 3572 -9247 3652 -9233
rect 4956 -9208 4996 -9207
rect 5048 -9200 5128 -9186
rect 5048 -9208 5062 -9200
rect 3150 -9270 3230 -9256
rect 3860 -9254 3940 -9240
rect 1670 -9304 1750 -9290
rect 1670 -9356 1684 -9304
rect 1736 -9310 1750 -9304
rect 2700 -9304 2780 -9290
rect 2700 -9310 2714 -9304
rect 1736 -9350 2714 -9310
rect 1736 -9356 1750 -9350
rect 1670 -9370 1750 -9356
rect 2700 -9356 2714 -9350
rect 2766 -9356 2780 -9304
rect 3860 -9306 3874 -9254
rect 3926 -9260 3940 -9254
rect 4760 -9254 4840 -9240
rect 4956 -9248 5062 -9208
rect 4760 -9260 4774 -9254
rect 3926 -9300 4774 -9260
rect 3926 -9306 3940 -9300
rect 3860 -9320 3940 -9306
rect 4760 -9306 4774 -9300
rect 4826 -9306 4840 -9254
rect 5048 -9252 5062 -9248
rect 5114 -9252 5128 -9200
rect 5048 -9266 5128 -9252
rect 4760 -9320 4840 -9306
rect 2700 -9370 2780 -9356
rect 3314 -9700 3394 -9689
rect 3314 -9756 3326 -9700
rect 3382 -9756 3394 -9700
rect 3314 -9769 3394 -9756
rect 1171 -9934 1251 -9920
rect 1171 -9986 1185 -9934
rect 1237 -9986 1251 -9934
rect 1171 -10000 1251 -9986
rect 1191 -10160 1231 -10000
rect 1171 -10174 1251 -10160
rect 1171 -10226 1185 -10174
rect 1237 -10226 1251 -10174
rect 1171 -10240 1251 -10226
rect 1055 -11286 1069 -11234
rect 1121 -11286 1135 -11234
rect 1055 -11695 1135 -11286
rect 1055 -11747 1069 -11695
rect 1121 -11747 1135 -11695
rect 1055 -11761 1135 -11747
rect 1191 -12740 1231 -10240
rect 3314 -10395 3394 -10384
rect 3314 -10451 3326 -10395
rect 3382 -10451 3394 -10395
rect 3314 -10464 3394 -10451
rect 1670 -10804 1750 -10790
rect 1670 -10856 1684 -10804
rect 1736 -10810 1750 -10804
rect 2700 -10804 2780 -10790
rect 2700 -10810 2714 -10804
rect 1736 -10850 2714 -10810
rect 1736 -10856 1750 -10850
rect 1670 -10870 1750 -10856
rect 2700 -10856 2714 -10850
rect 2766 -10856 2780 -10804
rect 2700 -10870 2780 -10856
rect 3860 -10854 3940 -10840
rect 1540 -10904 1620 -10890
rect 1540 -10956 1554 -10904
rect 1606 -10910 1620 -10904
rect 3150 -10904 3230 -10890
rect 3150 -10910 3164 -10904
rect 1606 -10950 3164 -10910
rect 1606 -10956 1620 -10950
rect 1540 -10970 1620 -10956
rect 3150 -10956 3164 -10950
rect 3216 -10956 3230 -10904
rect 3860 -10906 3874 -10854
rect 3926 -10860 3940 -10854
rect 4760 -10854 4840 -10840
rect 4760 -10860 4774 -10854
rect 3926 -10900 4774 -10860
rect 3926 -10906 3940 -10900
rect 3150 -10970 3230 -10956
rect 3572 -10925 3652 -10911
rect 3860 -10920 3940 -10906
rect 4760 -10906 4774 -10900
rect 4826 -10906 4840 -10854
rect 5048 -10892 5128 -10878
rect 5048 -10898 5062 -10892
rect 4760 -10920 4840 -10906
rect 3572 -10977 3586 -10925
rect 3638 -10951 3652 -10925
rect 4900 -10938 5062 -10898
rect 4900 -10951 4940 -10938
rect 3638 -10977 4940 -10951
rect 5048 -10944 5062 -10938
rect 5114 -10944 5128 -10892
rect 5048 -10958 5128 -10944
rect 1670 -11004 1750 -10990
rect 1670 -11056 1684 -11004
rect 1736 -11010 1750 -11004
rect 3000 -11004 3080 -10990
rect 3572 -10991 4940 -10977
rect 3000 -11010 3014 -11004
rect 1736 -11050 3014 -11010
rect 1736 -11056 1750 -11050
rect 1670 -11070 1750 -11056
rect 3000 -11056 3014 -11050
rect 3066 -11056 3080 -11004
rect 5048 -11000 5128 -10986
rect 5048 -11024 5062 -11000
rect 3000 -11070 3080 -11056
rect 3572 -11038 5062 -11024
rect 3572 -11090 3586 -11038
rect 3638 -11052 5062 -11038
rect 5114 -11052 5128 -11000
rect 3638 -11064 5128 -11052
rect 3638 -11090 3652 -11064
rect 5048 -11066 5128 -11064
rect 1540 -11104 1620 -11090
rect 1540 -11156 1554 -11104
rect 1606 -11110 1620 -11104
rect 2800 -11104 2880 -11090
rect 3572 -11104 3652 -11090
rect 3860 -11103 3940 -11092
rect 2800 -11110 2814 -11104
rect 1606 -11150 2814 -11110
rect 1606 -11156 1620 -11150
rect 1540 -11170 1620 -11156
rect 2800 -11156 2814 -11150
rect 2866 -11156 2880 -11104
rect 2800 -11170 2880 -11156
rect 3860 -11159 3872 -11103
rect 3928 -11159 3940 -11103
rect 5156 -11117 5196 -8500
rect 5478 -8518 5518 -7420
rect 5458 -8532 5538 -8518
rect 5458 -8584 5472 -8532
rect 5524 -8584 5538 -8532
rect 5458 -8598 5538 -8584
rect 5566 -8626 5646 -5646
rect 5799 -6284 5879 -6270
rect 5799 -6336 5813 -6284
rect 5865 -6290 5879 -6284
rect 6929 -6284 7009 -6270
rect 6929 -6290 6943 -6284
rect 5865 -6330 6943 -6290
rect 5865 -6336 5879 -6330
rect 5799 -6350 5879 -6336
rect 6929 -6336 6943 -6330
rect 6995 -6336 7009 -6284
rect 6929 -6350 7009 -6336
rect 5799 -6404 5879 -6390
rect 5799 -6456 5813 -6404
rect 5865 -6410 5879 -6404
rect 6779 -6404 6859 -6390
rect 6779 -6410 6793 -6404
rect 5865 -6450 6793 -6410
rect 5865 -6456 5879 -6450
rect 5799 -6470 5879 -6456
rect 6779 -6456 6793 -6450
rect 6845 -6456 6859 -6404
rect 6779 -6470 6859 -6456
rect 7153 -6660 7193 -5419
rect 7270 -5464 7350 -5450
rect 7270 -5516 7284 -5464
rect 7336 -5516 7350 -5464
rect 7270 -5530 7350 -5516
rect 7129 -6674 7209 -6660
rect 7129 -6726 7143 -6674
rect 7195 -6726 7209 -6674
rect 7129 -6740 7209 -6726
rect 7030 -6994 7110 -6980
rect 7030 -7046 7044 -6994
rect 7096 -7046 7110 -6994
rect 7030 -7474 7110 -7046
rect 7030 -7526 7044 -7474
rect 7096 -7526 7110 -7474
rect 7030 -7540 7110 -7526
rect 7133 -7795 7213 -7781
rect 7133 -7847 7147 -7795
rect 7199 -7800 7213 -7795
rect 7291 -7800 7331 -5530
rect 7514 -5774 7554 -5233
rect 7494 -5788 7574 -5774
rect 7494 -5840 7508 -5788
rect 7560 -5840 7574 -5788
rect 7494 -5854 7574 -5840
rect 7199 -7840 7331 -7800
rect 7199 -7847 7213 -7840
rect 7133 -7861 7213 -7847
rect 5799 -8064 5879 -8050
rect 5799 -8116 5813 -8064
rect 5865 -8070 5879 -8064
rect 6779 -8064 6859 -8050
rect 6779 -8070 6793 -8064
rect 5865 -8110 6793 -8070
rect 5865 -8116 5879 -8110
rect 5799 -8130 5879 -8116
rect 6779 -8116 6793 -8110
rect 6845 -8116 6859 -8064
rect 6779 -8130 6859 -8116
rect 5799 -8184 5879 -8170
rect 5799 -8236 5813 -8184
rect 5865 -8190 5879 -8184
rect 6929 -8184 7009 -8170
rect 6929 -8190 6943 -8184
rect 5865 -8230 6943 -8190
rect 5865 -8236 5879 -8230
rect 5799 -8250 5879 -8236
rect 6929 -8236 6943 -8230
rect 6995 -8236 7009 -8184
rect 6929 -8250 7009 -8236
rect 3860 -11172 3940 -11159
rect 5112 -11157 5196 -11117
rect 5251 -8706 5646 -8626
rect 5690 -8414 5770 -8400
rect 5690 -8466 5704 -8414
rect 5756 -8466 5770 -8414
rect 1581 -11814 1661 -11800
rect 1581 -11866 1595 -11814
rect 1647 -11820 1661 -11814
rect 2951 -11814 3031 -11800
rect 2951 -11820 2965 -11814
rect 1647 -11860 2965 -11820
rect 1647 -11866 1661 -11860
rect 1581 -11880 1661 -11866
rect 2951 -11866 2965 -11860
rect 3017 -11866 3031 -11814
rect 2951 -11880 3031 -11866
rect 5004 -11901 5084 -11887
rect 1671 -11934 1751 -11920
rect 1671 -11986 1685 -11934
rect 1737 -11940 1751 -11934
rect 2801 -11934 2881 -11920
rect 2801 -11940 2815 -11934
rect 1737 -11980 2815 -11940
rect 1737 -11986 1751 -11980
rect 1671 -12000 1751 -11986
rect 2801 -11986 2815 -11980
rect 2867 -11986 2881 -11934
rect 5004 -11953 5018 -11901
rect 5070 -11953 5084 -11901
rect 5004 -11967 5084 -11953
rect 2801 -12000 2881 -11986
rect 1641 -12054 1721 -12040
rect 1641 -12106 1655 -12054
rect 1707 -12060 1721 -12054
rect 2671 -12054 2751 -12040
rect 2671 -12060 2685 -12054
rect 1707 -12100 2685 -12060
rect 1707 -12106 1721 -12100
rect 1641 -12120 1721 -12106
rect 2671 -12106 2685 -12100
rect 2737 -12106 2751 -12054
rect 2671 -12120 2751 -12106
rect 3721 -12074 3801 -12060
rect 3721 -12126 3735 -12074
rect 3787 -12080 3801 -12074
rect 4621 -12074 4701 -12060
rect 4621 -12080 4635 -12074
rect 3787 -12120 4635 -12080
rect 3787 -12126 3801 -12120
rect 3721 -12140 3801 -12126
rect 4621 -12126 4635 -12120
rect 4687 -12126 4701 -12074
rect 4621 -12140 4701 -12126
rect 5023 -12464 5063 -11967
rect 4998 -12478 5078 -12464
rect 4998 -12530 5012 -12478
rect 5064 -12530 5078 -12478
rect 4998 -12544 5078 -12530
rect 1171 -12754 1251 -12740
rect 5112 -12742 5152 -11157
rect 5251 -11695 5331 -8706
rect 5398 -8756 5478 -8742
rect 5398 -8808 5412 -8756
rect 5464 -8808 5478 -8756
rect 5398 -8822 5478 -8808
rect 5418 -9920 5458 -8822
rect 5690 -8874 5770 -8466
rect 5690 -8926 5704 -8874
rect 5756 -8926 5770 -8874
rect 5690 -8940 5770 -8926
rect 6990 -8874 7070 -8860
rect 6990 -8926 7004 -8874
rect 7056 -8926 7070 -8874
rect 6990 -8940 7070 -8926
rect 5740 -9104 5820 -9090
rect 5740 -9156 5754 -9104
rect 5806 -9110 5820 -9104
rect 6870 -9104 6950 -9090
rect 6870 -9110 6884 -9104
rect 5806 -9150 6884 -9110
rect 5806 -9156 5820 -9150
rect 5740 -9170 5820 -9156
rect 6870 -9156 6884 -9150
rect 6936 -9156 6950 -9104
rect 6870 -9170 6950 -9156
rect 5740 -9224 5820 -9210
rect 5740 -9276 5754 -9224
rect 5806 -9230 5820 -9224
rect 6720 -9224 6800 -9210
rect 6720 -9230 6734 -9224
rect 5806 -9270 6734 -9230
rect 5806 -9276 5820 -9270
rect 5740 -9290 5820 -9276
rect 6720 -9276 6734 -9270
rect 6786 -9276 6800 -9224
rect 6720 -9290 6800 -9276
rect 7073 -9494 7153 -9480
rect 7073 -9546 7087 -9494
rect 7139 -9500 7153 -9494
rect 7139 -9540 7269 -9500
rect 7139 -9546 7153 -9540
rect 7073 -9560 7153 -9546
rect 6970 -9814 7050 -9800
rect 6970 -9866 6984 -9814
rect 7036 -9866 7050 -9814
rect 5398 -9934 5478 -9920
rect 5398 -9986 5412 -9934
rect 5464 -9986 5478 -9934
rect 5398 -10000 5478 -9986
rect 5418 -10159 5458 -10000
rect 5398 -10173 5478 -10159
rect 5398 -10225 5412 -10173
rect 5464 -10225 5478 -10173
rect 5398 -10239 5478 -10225
rect 5418 -11454 5458 -10239
rect 6970 -10294 7050 -9866
rect 6970 -10346 6984 -10294
rect 7036 -10346 7050 -10294
rect 6970 -10360 7050 -10346
rect 7073 -10614 7153 -10600
rect 7073 -10666 7087 -10614
rect 7139 -10666 7153 -10614
rect 7073 -10680 7153 -10666
rect 5740 -10884 5820 -10870
rect 5740 -10936 5754 -10884
rect 5806 -10890 5820 -10884
rect 6720 -10884 6800 -10870
rect 6720 -10890 6734 -10884
rect 5806 -10930 6734 -10890
rect 5806 -10936 5820 -10930
rect 5740 -10950 5820 -10936
rect 6720 -10936 6734 -10930
rect 6786 -10936 6800 -10884
rect 6720 -10950 6800 -10936
rect 5740 -11004 5820 -10990
rect 5740 -11056 5754 -11004
rect 5806 -11010 5820 -11004
rect 6870 -11004 6950 -10990
rect 6870 -11010 6884 -11004
rect 5806 -11050 6884 -11010
rect 5806 -11056 5820 -11050
rect 5740 -11070 5820 -11056
rect 6870 -11056 6884 -11050
rect 6936 -11056 6950 -11004
rect 6870 -11070 6950 -11056
rect 5398 -11468 5478 -11454
rect 5398 -11520 5412 -11468
rect 5464 -11520 5478 -11468
rect 5398 -11534 5478 -11520
rect 5251 -11747 5265 -11695
rect 5317 -11747 5331 -11695
rect 5251 -11761 5331 -11747
rect 5381 -11820 5461 -11806
rect 5381 -11872 5395 -11820
rect 5447 -11831 5461 -11820
rect 6661 -11825 6741 -11811
rect 6661 -11831 6675 -11825
rect 5447 -11871 6675 -11831
rect 5447 -11872 5461 -11871
rect 5381 -11886 5461 -11872
rect 6661 -11877 6675 -11871
rect 6727 -11877 6741 -11825
rect 6661 -11891 6741 -11877
rect 7073 -11921 7113 -10680
rect 7229 -11811 7269 -9540
rect 7343 -11501 7423 -11487
rect 7343 -11553 7357 -11501
rect 7409 -11553 7423 -11501
rect 7343 -11567 7423 -11553
rect 7229 -11825 7309 -11811
rect 7229 -11877 7243 -11825
rect 7295 -11877 7309 -11825
rect 7229 -11891 7309 -11877
rect 5481 -11941 5561 -11931
rect 6781 -11935 6861 -11921
rect 6781 -11941 6795 -11935
rect 5481 -11945 6795 -11941
rect 5180 -11987 5260 -11973
rect 5180 -12039 5194 -11987
rect 5246 -11993 5260 -11987
rect 5246 -12033 5353 -11993
rect 5481 -11997 5495 -11945
rect 5547 -11981 6795 -11945
rect 5547 -11997 5561 -11981
rect 5481 -12011 5561 -11997
rect 6781 -11987 6795 -11981
rect 6847 -11987 6861 -11935
rect 6781 -12001 6861 -11987
rect 7033 -11935 7113 -11921
rect 7033 -11987 7047 -11935
rect 7099 -11987 7113 -11935
rect 7033 -12001 7113 -11987
rect 5246 -12039 5260 -12033
rect 5180 -12053 5260 -12039
rect 5313 -12041 5353 -12033
rect 5681 -12035 5761 -12021
rect 5681 -12041 5695 -12035
rect 5313 -12081 5695 -12041
rect 5180 -12097 5260 -12083
rect 5180 -12149 5194 -12097
rect 5246 -12129 5260 -12097
rect 5681 -12087 5695 -12081
rect 5747 -12041 5761 -12035
rect 6661 -12035 6741 -12021
rect 6661 -12041 6675 -12035
rect 5747 -12081 6675 -12041
rect 5747 -12087 5761 -12081
rect 5681 -12101 5761 -12087
rect 6661 -12087 6675 -12081
rect 6727 -12087 6741 -12035
rect 6661 -12101 6741 -12087
rect 6791 -12123 6871 -12109
rect 6791 -12129 6805 -12123
rect 5246 -12149 6805 -12129
rect 5180 -12169 6805 -12149
rect 6791 -12175 6805 -12169
rect 6857 -12175 6871 -12123
rect 6791 -12189 6871 -12175
rect 7275 -12123 7355 -12109
rect 7275 -12175 7289 -12123
rect 7341 -12131 7355 -12123
rect 7383 -12131 7423 -11567
rect 7341 -12171 7423 -12131
rect 7341 -12175 7355 -12171
rect 7275 -12189 7355 -12175
rect 5181 -12211 5261 -12197
rect 5181 -12263 5195 -12211
rect 5247 -12217 5261 -12211
rect 5247 -12257 7291 -12217
rect 5247 -12263 5261 -12257
rect 5181 -12277 5261 -12263
rect 5181 -12321 5261 -12311
rect 5181 -12325 7291 -12321
rect 5181 -12377 5195 -12325
rect 5247 -12361 7291 -12325
rect 5247 -12377 5261 -12361
rect 5181 -12391 5261 -12377
rect 1171 -12806 1185 -12754
rect 1237 -12806 1251 -12754
rect 1171 -12820 1251 -12806
rect 5092 -12756 5172 -12742
rect 5092 -12808 5106 -12756
rect 5158 -12808 5172 -12756
rect 5092 -12822 5172 -12808
<< via2 >>
rect 240 2370 296 2372
rect 240 2318 242 2370
rect 242 2318 294 2370
rect 294 2318 296 2370
rect 240 2316 296 2318
rect 582 2227 638 2229
rect 582 2175 584 2227
rect 584 2175 636 2227
rect 636 2175 638 2227
rect 582 2173 638 2175
rect 468 1696 524 1698
rect 468 1644 470 1696
rect 470 1644 522 1696
rect 522 1644 524 1696
rect 468 1642 524 1644
rect 354 1536 410 1538
rect 354 1484 356 1536
rect 356 1484 408 1536
rect 408 1484 410 1536
rect 354 1482 410 1484
rect 3000 2370 3056 2372
rect 3000 2318 3002 2370
rect 3002 2318 3054 2370
rect 3054 2318 3056 2370
rect 3000 2316 3056 2318
rect 3280 2230 3336 2232
rect 3280 2178 3282 2230
rect 3282 2178 3334 2230
rect 3334 2178 3336 2230
rect 3280 2176 3336 2178
rect 3347 1696 3403 1698
rect 3347 1644 3349 1696
rect 3349 1644 3401 1696
rect 3401 1644 3403 1696
rect 3347 1642 3403 1644
rect 3347 1536 3403 1538
rect 3347 1484 3349 1536
rect 3349 1484 3401 1536
rect 3401 1484 3403 1536
rect 3347 1482 3403 1484
rect 696 -460 752 -458
rect 696 -512 698 -460
rect 698 -512 750 -460
rect 750 -512 752 -460
rect 696 -514 752 -512
rect 810 -1161 866 -1159
rect 810 -1213 812 -1161
rect 812 -1213 864 -1161
rect 864 -1213 866 -1161
rect 810 -1215 866 -1213
rect 580 -1857 636 -1855
rect 580 -1909 582 -1857
rect 582 -1909 634 -1857
rect 634 -1909 636 -1857
rect 580 -1911 636 -1909
rect 468 -2564 524 -2562
rect 468 -2616 470 -2564
rect 470 -2616 522 -2564
rect 522 -2616 524 -2564
rect 468 -2618 524 -2616
rect 3872 -460 3928 -458
rect 3872 -512 3874 -460
rect 3874 -512 3926 -460
rect 3926 -512 3928 -460
rect 3872 -514 3928 -512
rect 3326 -1161 3382 -1159
rect 3326 -1213 3328 -1161
rect 3328 -1213 3380 -1161
rect 3380 -1213 3382 -1161
rect 3326 -1215 3382 -1213
rect 3326 -1856 3382 -1854
rect 3326 -1908 3328 -1856
rect 3328 -1908 3380 -1856
rect 3380 -1908 3382 -1856
rect 3326 -1910 3382 -1908
rect 3872 -2564 3928 -2562
rect 3872 -2616 3874 -2564
rect 3874 -2616 3926 -2564
rect 3926 -2616 3928 -2564
rect 3872 -2618 3928 -2616
rect 582 -6183 638 -6181
rect 582 -6235 584 -6183
rect 584 -6235 636 -6183
rect 636 -6235 638 -6183
rect 582 -6237 638 -6235
rect 468 -6914 524 -6912
rect 468 -6966 470 -6914
rect 470 -6966 522 -6914
rect 522 -6966 524 -6914
rect 468 -6968 524 -6966
rect 3932 -6183 3988 -6181
rect 3932 -6235 3934 -6183
rect 3934 -6235 3986 -6183
rect 3986 -6235 3988 -6183
rect 3932 -6237 3988 -6235
rect 3366 -6914 3422 -6912
rect 3366 -6966 3368 -6914
rect 3368 -6966 3420 -6914
rect 3420 -6966 3422 -6914
rect 3366 -6968 3422 -6966
rect 240 -7552 296 -7550
rect 240 -7604 242 -7552
rect 242 -7604 294 -7552
rect 294 -7604 296 -7552
rect 240 -7606 296 -7604
rect 354 -8287 410 -8285
rect 354 -8339 356 -8287
rect 356 -8339 408 -8287
rect 408 -8339 410 -8287
rect 354 -8341 410 -8339
rect 3366 -7552 3422 -7550
rect 3366 -7604 3368 -7552
rect 3368 -7604 3420 -7552
rect 3420 -7604 3422 -7552
rect 3366 -7606 3422 -7604
rect 3932 -8287 3988 -8285
rect 3932 -8339 3934 -8287
rect 3934 -8339 3986 -8287
rect 3986 -8339 3988 -8287
rect 3932 -8341 3988 -8339
rect 810 -9002 866 -9000
rect 810 -9054 812 -9002
rect 812 -9054 864 -9002
rect 864 -9054 866 -9002
rect 810 -9056 866 -9054
rect 696 -9702 752 -9700
rect 696 -9754 698 -9702
rect 698 -9754 750 -9702
rect 750 -9754 752 -9702
rect 696 -9756 752 -9754
rect 354 -10398 410 -10396
rect 354 -10450 356 -10398
rect 356 -10450 408 -10398
rect 408 -10450 410 -10398
rect 354 -10452 410 -10450
rect 240 -11105 296 -11103
rect 240 -11157 242 -11105
rect 242 -11157 294 -11105
rect 294 -11157 296 -11105
rect 240 -11159 296 -11157
rect 3872 -9001 3928 -8999
rect 3872 -9053 3874 -9001
rect 3874 -9053 3926 -9001
rect 3926 -9053 3928 -9001
rect 3872 -9055 3928 -9053
rect 3326 -9702 3382 -9700
rect 3326 -9754 3328 -9702
rect 3328 -9754 3380 -9702
rect 3380 -9754 3382 -9702
rect 3326 -9756 3382 -9754
rect 3326 -10397 3382 -10395
rect 3326 -10449 3328 -10397
rect 3328 -10449 3380 -10397
rect 3380 -10449 3382 -10397
rect 3326 -10451 3382 -10449
rect 3872 -11105 3928 -11103
rect 3872 -11157 3874 -11105
rect 3874 -11157 3926 -11105
rect 3926 -11157 3928 -11105
rect 3872 -11159 3928 -11157
<< metal3 >>
rect 218 2373 318 2393
rect 2978 2373 3078 2393
rect 218 2372 3078 2373
rect 218 2316 240 2372
rect 296 2316 3000 2372
rect 3056 2316 3078 2372
rect 218 2313 3078 2316
rect 218 2293 318 2313
rect 2978 2293 3078 2313
rect 560 2233 660 2250
rect 3258 2233 3358 2253
rect 560 2232 3358 2233
rect 560 2229 3280 2232
rect 560 2173 582 2229
rect 638 2176 3280 2229
rect 3336 2176 3358 2232
rect 638 2173 3358 2176
rect 560 2150 660 2173
rect 3258 2153 3358 2173
rect 446 1699 546 1719
rect 3325 1699 3425 1719
rect 446 1698 3425 1699
rect 446 1642 468 1698
rect 524 1642 3347 1698
rect 3403 1642 3425 1698
rect 446 1639 3425 1642
rect 446 1619 546 1639
rect 3325 1619 3425 1639
rect 332 1539 432 1559
rect 3325 1539 3425 1559
rect 332 1538 3425 1539
rect 332 1482 354 1538
rect 410 1482 3347 1538
rect 3403 1482 3425 1538
rect 332 1479 3425 1482
rect 332 1459 432 1479
rect 3325 1459 3425 1479
rect 674 -457 774 -437
rect 3850 -457 3950 -437
rect 674 -458 3950 -457
rect 674 -514 696 -458
rect 752 -514 3872 -458
rect 3928 -514 3950 -458
rect 674 -517 3950 -514
rect 674 -537 774 -517
rect 3850 -537 3950 -517
rect 788 -1158 888 -1138
rect 3304 -1158 3404 -1138
rect 788 -1159 3404 -1158
rect 788 -1215 810 -1159
rect 866 -1215 3326 -1159
rect 3382 -1215 3404 -1159
rect 788 -1218 3404 -1215
rect 788 -1238 888 -1218
rect 3304 -1238 3404 -1218
rect 558 -1852 658 -1834
rect 3304 -1852 3404 -1833
rect 558 -1854 3404 -1852
rect 558 -1855 3326 -1854
rect 558 -1911 580 -1855
rect 636 -1910 3326 -1855
rect 3382 -1910 3404 -1854
rect 636 -1911 3404 -1910
rect 558 -1912 3404 -1911
rect 558 -1934 658 -1912
rect 3304 -1933 3404 -1912
rect 446 -2561 546 -2541
rect 3850 -2561 3950 -2541
rect 446 -2562 3950 -2561
rect 446 -2618 468 -2562
rect 524 -2618 3872 -2562
rect 3928 -2618 3950 -2562
rect 446 -2621 3950 -2618
rect 446 -2641 546 -2621
rect 3850 -2641 3950 -2621
rect 560 -6180 660 -6158
rect 3910 -6180 4010 -6158
rect 560 -6181 4010 -6180
rect 560 -6237 582 -6181
rect 638 -6237 3932 -6181
rect 3988 -6237 4010 -6181
rect 560 -6240 4010 -6237
rect 560 -6258 660 -6240
rect 3910 -6258 4010 -6240
rect 446 -6910 546 -6889
rect 3344 -6910 3444 -6889
rect 446 -6912 3444 -6910
rect 446 -6968 468 -6912
rect 524 -6968 3366 -6912
rect 3422 -6968 3444 -6912
rect 446 -6970 3444 -6968
rect 446 -6989 546 -6970
rect 3344 -6989 3444 -6970
rect 218 -7548 318 -7527
rect 3344 -7548 3444 -7527
rect 218 -7550 3444 -7548
rect 218 -7606 240 -7550
rect 296 -7606 3366 -7550
rect 3422 -7606 3444 -7550
rect 218 -7608 3444 -7606
rect 218 -7627 318 -7608
rect 3344 -7627 3444 -7608
rect 332 -8282 432 -8262
rect 3910 -8282 4010 -8262
rect 332 -8285 4010 -8282
rect 332 -8341 354 -8285
rect 410 -8341 3932 -8285
rect 3988 -8341 4010 -8285
rect 332 -8342 4010 -8341
rect 332 -8362 432 -8342
rect 3910 -8362 4010 -8342
rect 788 -8998 888 -8979
rect 3850 -8998 3950 -8978
rect 788 -8999 3950 -8998
rect 788 -9000 3872 -8999
rect 788 -9056 810 -9000
rect 866 -9055 3872 -9000
rect 3928 -9055 3950 -8999
rect 866 -9056 3950 -9055
rect 788 -9058 3950 -9056
rect 788 -9079 888 -9058
rect 3850 -9078 3950 -9058
rect 674 -9699 774 -9679
rect 3304 -9699 3404 -9679
rect 674 -9700 3404 -9699
rect 674 -9756 696 -9700
rect 752 -9756 3326 -9700
rect 3382 -9756 3404 -9700
rect 674 -9759 3404 -9756
rect 674 -9779 774 -9759
rect 3304 -9779 3404 -9759
rect 332 -10393 432 -10375
rect 3304 -10393 3404 -10374
rect 332 -10395 3404 -10393
rect 332 -10396 3326 -10395
rect 332 -10452 354 -10396
rect 410 -10451 3326 -10396
rect 3382 -10451 3404 -10395
rect 410 -10452 3404 -10451
rect 332 -10453 3404 -10452
rect 332 -10475 432 -10453
rect 3304 -10474 3404 -10453
rect 218 -11102 318 -11082
rect 3850 -11102 3950 -11082
rect 218 -11103 3950 -11102
rect 218 -11159 240 -11103
rect 296 -11159 3872 -11103
rect 3928 -11159 3950 -11103
rect 218 -11162 3950 -11159
rect 218 -11182 318 -11162
rect 3850 -11182 3950 -11162
<< labels >>
flabel metal1 s 930 2283 974 2329 2 FreeSans 2000 0 0 0 GND
port 1 nsew
flabel metal1 s 10 2278 71 2338 2 FreeSans 2500 0 0 0 x0
port 2 nsew
flabel metal1 s 123 2217 184 2277 2 FreeSans 2500 0 0 0 x0_bar
port 3 nsew
flabel metal1 s 238 2278 299 2338 2 FreeSans 2500 0 0 0 x1
port 4 nsew
flabel metal1 s 352 2217 413 2277 2 FreeSans 2500 0 0 0 x1_bar
port 5 nsew
flabel metal1 s 467 2282 528 2342 2 FreeSans 2500 0 0 0 x2
port 6 nsew
flabel metal1 s 579 2218 640 2278 2 FreeSans 2500 0 0 0 x2_bar
port 7 nsew
flabel metal1 s 694 2279 755 2339 2 FreeSans 2500 0 0 0 x3
port 8 nsew
flabel metal1 s 808 2218 869 2278 2 FreeSans 2500 0 0 0 x3_bar
port 9 nsew
flabel metal2 s 1158 2397 1181 2421 2 FreeSans 2000 0 0 0 Dis1
port 10 nsew
flabel metal2 s 1038 2391 1069 2422 2 FreeSans 2000 0 0 0 CLK1
port 11 nsew
flabel metal2 s 5853 2452 5887 2486 2 FreeSans 2000 0 0 0 CLK2
port 12 nsew
flabel metal2 s 5770 2424 5795 2448 2 FreeSans 2000 0 0 0 Dis2
port 13 nsew
flabel metal2 s 5486 2441 5511 2466 2 FreeSans 2000 0 0 0 CLK3
port 14 nsew
flabel metal2 s 5954 2442 5973 2463 2 FreeSans 2000 0 0 0 Dis3
port 15 nsew
flabel metal2 s 7458 711 7477 730 2 FreeSans 2000 0 0 0 s0
port 16 nsew
flabel metal2 s 7459 590 7480 609 2 FreeSans 2000 0 0 0 s0_bar
port 17 nsew
flabel metal2 s 7227 -3705 7248 -3685 2 FreeSans 2000 0 0 0 s1_bar
port 18 nsew
flabel metal2 s 7229 -3811 7250 -3790 2 FreeSans 2000 0 0 0 s1
port 19 nsew
flabel metal2 s 7494 -4989 7514 -4969 2 FreeSans 2000 0 0 0 s2
port 20 nsew
flabel metal2 s 7499 -5116 7521 -5095 2 FreeSans 2000 0 0 0 s2_bar
port 21 nsew
flabel metal2 s 7231 -12247 7251 -12228 2 FreeSans 2000 0 0 0 s3_bar
port 22 nsew
flabel metal2 s 7232 -12353 7253 -12332 2 FreeSans 2000 0 0 0 s3
port 23 nsew
flabel metal1 930 -10103 974 -10057 2 FreeSans 2000 0 0 0 EESPFAL_s3_0/GND
flabel metal1 10 -9084 71 -9024 2 FreeSans 2500 0 0 0 EESPFAL_s3_0/x0
flabel metal1 123 -9145 184 -9085 2 FreeSans 2500 0 0 0 EESPFAL_s3_0/x0_bar
flabel metal1 238 -9084 299 -9024 2 FreeSans 2500 0 0 0 EESPFAL_s3_0/x1
flabel metal1 352 -9145 413 -9085 2 FreeSans 2500 0 0 0 EESPFAL_s3_0/x1_bar
flabel metal1 467 -9080 528 -9020 2 FreeSans 2500 0 0 0 EESPFAL_s3_0/x2
flabel metal1 579 -9144 640 -9084 2 FreeSans 2500 0 0 0 EESPFAL_s3_0/x2_bar
flabel metal1 694 -9083 755 -9023 2 FreeSans 2500 0 0 0 EESPFAL_s3_0/x3
flabel metal1 808 -9144 869 -9084 2 FreeSans 2500 0 0 0 EESPFAL_s3_0/x3_bar
flabel metal2 7260 -12247 7280 -12227 2 FreeSans 2000 0 0 0 EESPFAL_s3_0/s3_bar
flabel metal2 7260 -12353 7280 -12332 2 FreeSans 2000 0 0 0 EESPFAL_s3_0/s3
flabel metal2 1080 -8901 1111 -8870 2 FreeSans 2000 0 0 0 EESPFAL_s3_0/CLK1
flabel metal2 1200 -8895 1223 -8871 2 FreeSans 2000 0 0 0 EESPFAL_s3_0/Dis1
flabel metal2 5167 -8888 5186 -8867 2 FreeSans 2000 0 0 0 EESPFAL_s3_0/Dis3
flabel metal2 5278 -8891 5303 -8866 2 FreeSans 2000 0 0 0 EESPFAL_s3_0/CLK3
flabel metal2 5426 -8889 5451 -8865 2 FreeSans 2000 0 0 0 EESPFAL_s3_0/Dis2
flabel metal2 7014 -8899 7048 -8865 2 FreeSans 2000 0 0 0 EESPFAL_s3_0/CLK2
rlabel metal1 2191 -12240 2231 -12200 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/OUT_bar
rlabel metal1 2141 -12920 2181 -12880 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/GND!
rlabel metal1 2141 -11740 2181 -11700 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/CLK
rlabel locali 2091 -12365 2131 -12325 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/OUT
rlabel locali 1181 -11850 1201 -11830 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A
rlabel locali 1181 -12160 1201 -12140 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A_bar
rlabel locali 1181 -11970 1201 -11950 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B
rlabel locali 1181 -12240 1201 -12220 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B_bar
rlabel locali 1181 -12080 1201 -12060 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C
rlabel locali 1181 -12340 1201 -12320 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C_bar
rlabel locali 1941 -12800 1981 -12760 4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/Dis
rlabel metal1 4241 -12240 4281 -12200 4 EESPFAL_s3_0/EESPFAL_INV4_0/OUT
rlabel metal1 4191 -12920 4231 -12880 4 EESPFAL_s3_0/EESPFAL_INV4_0/GND!
rlabel metal1 4191 -11740 4231 -11700 4 EESPFAL_s3_0/EESPFAL_INV4_0/CLK
rlabel locali 4141 -12365 4181 -12325 4 EESPFAL_s3_0/EESPFAL_INV4_0/OUT_bar
rlabel locali 4771 -12120 4811 -12080 4 EESPFAL_s3_0/EESPFAL_INV4_0/A
rlabel locali 3611 -12360 3651 -12320 4 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar
rlabel locali 3991 -12800 4031 -12760 4 EESPFAL_s3_0/EESPFAL_INV4_0/Dis
rlabel metal1 6181 -12241 6221 -12201 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/OUT_bar
rlabel metal1 6231 -12921 6271 -12881 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/GND!
rlabel metal1 6231 -11741 6271 -11701 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/CLK
rlabel locali 6281 -12366 6321 -12326 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/OUT
rlabel locali 7211 -11861 7231 -11841 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/A
rlabel locali 7211 -12161 7231 -12141 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/A_bar
rlabel locali 7211 -11971 7231 -11951 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/B
rlabel locali 7211 -12281 7231 -12261 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/B_bar
rlabel locali 7211 -12071 7231 -12051 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C
rlabel locali 7211 -12381 7231 -12361 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar
rlabel locali 6431 -12801 6471 -12761 6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/Dis
rlabel metal1 2190 -10780 2230 -10740 2 EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT_bar
rlabel metal1 2140 -10100 2180 -10060 2 EESPFAL_s3_0/EESPFAL_XOR_v3_1/GND!
rlabel metal1 2140 -11280 2180 -11240 2 EESPFAL_s3_0/EESPFAL_XOR_v3_1/CLK
rlabel locali 2090 -10655 2130 -10615 2 EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT
rlabel locali 1030 -11140 1050 -11120 2 EESPFAL_s3_0/EESPFAL_XOR_v3_1/A
rlabel locali 1030 -11040 1050 -11020 2 EESPFAL_s3_0/EESPFAL_XOR_v3_1/A_bar
rlabel locali 1030 -10940 1050 -10920 2 EESPFAL_s3_0/EESPFAL_XOR_v3_1/B
rlabel locali 1030 -10840 1050 -10820 2 EESPFAL_s3_0/EESPFAL_XOR_v3_1/B_bar
rlabel locali 1940 -10220 1980 -10180 2 EESPFAL_s3_0/EESPFAL_XOR_v3_1/Dis
rlabel metal1 4380 -10780 4420 -10740 2 EESPFAL_s3_0/EESPFAL_INV4_1/OUT
rlabel metal1 4330 -10100 4370 -10060 2 EESPFAL_s3_0/EESPFAL_INV4_1/GND!
rlabel metal1 4330 -11280 4370 -11240 2 EESPFAL_s3_0/EESPFAL_INV4_1/CLK
rlabel locali 4280 -10655 4320 -10615 2 EESPFAL_s3_0/EESPFAL_INV4_1/OUT_bar
rlabel locali 4910 -10900 4950 -10860 2 EESPFAL_s3_0/EESPFAL_INV4_1/A
rlabel locali 3750 -10660 3790 -10620 2 EESPFAL_s3_0/EESPFAL_INV4_1/A_bar
rlabel locali 4130 -10220 4170 -10180 2 EESPFAL_s3_0/EESPFAL_INV4_1/Dis
rlabel metal1 6260 -10780 6300 -10740 2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar
rlabel metal1 6210 -10100 6250 -10060 2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/GND!
rlabel metal1 6210 -11280 6250 -11240 2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/CLK
rlabel locali 6160 -10655 6200 -10615 2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT
rlabel locali 5400 -11040 5420 -11020 2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A
rlabel locali 5400 -10820 5420 -10800 2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar
rlabel locali 5400 -10920 5420 -10900 2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B
rlabel locali 5400 -10720 5420 -10700 2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar
rlabel locali 6010 -10220 6050 -10180 2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/Dis
rlabel metal1 2190 -9420 2230 -9380 4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT_bar
rlabel metal1 2140 -10100 2180 -10060 4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/GND!
rlabel metal1 2140 -8920 2180 -8880 4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/CLK
rlabel locali 2090 -9545 2130 -9505 4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT
rlabel locali 1030 -9040 1050 -9020 4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/A
rlabel locali 1030 -9140 1050 -9120 4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/A_bar
rlabel locali 1030 -9240 1050 -9220 4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/B
rlabel locali 1030 -9340 1050 -9320 4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/B_bar
rlabel locali 1940 -9980 1980 -9940 4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/Dis
rlabel metal1 4380 -9420 4420 -9380 4 EESPFAL_s3_0/EESPFAL_INV4_2/OUT
rlabel metal1 4330 -10100 4370 -10060 4 EESPFAL_s3_0/EESPFAL_INV4_2/GND!
rlabel metal1 4330 -8920 4370 -8880 4 EESPFAL_s3_0/EESPFAL_INV4_2/CLK
rlabel locali 4280 -9545 4320 -9505 4 EESPFAL_s3_0/EESPFAL_INV4_2/OUT_bar
rlabel locali 4910 -9300 4950 -9260 4 EESPFAL_s3_0/EESPFAL_INV4_2/A
rlabel locali 3750 -9540 3790 -9500 4 EESPFAL_s3_0/EESPFAL_INV4_2/A_bar
rlabel locali 4130 -9980 4170 -9940 4 EESPFAL_s3_0/EESPFAL_INV4_2/Dis
rlabel metal1 6260 -9420 6300 -9380 4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar
rlabel metal1 6210 -10100 6250 -10060 4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/GND!
rlabel metal1 6210 -8920 6250 -8880 4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/CLK
rlabel locali 6160 -9545 6200 -9505 4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT
rlabel locali 5400 -9140 5420 -9120 4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A
rlabel locali 5400 -9360 5420 -9340 4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar
rlabel locali 5400 -9260 5420 -9240 4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B
rlabel locali 5400 -9460 5420 -9440 4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar
rlabel locali 6010 -9980 6050 -9940 4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/Dis
flabel metal1 935 -7277 969 -7243 4 FreeSans 2000 0 0 0 EESPFAL_s2_0/GND
flabel metal1 10 -8316 71 -8256 4 FreeSans 3126 0 0 0 EESPFAL_s2_0/x0
flabel metal1 123 -8255 184 -8195 4 FreeSans 3126 0 0 0 EESPFAL_s2_0/x0_bar
flabel metal1 238 -8316 299 -8256 4 FreeSans 3126 0 0 0 EESPFAL_s2_0/x1
flabel metal1 352 -8255 413 -8195 4 FreeSans 3126 0 0 0 EESPFAL_s2_0/x1_bar
flabel metal1 466 -8317 527 -8257 4 FreeSans 3126 0 0 0 EESPFAL_s2_0/x2
flabel metal1 579 -8256 640 -8196 4 FreeSans 3126 0 0 0 EESPFAL_s2_0/x2_bar
flabel metal1 694 -8317 755 -8257 4 FreeSans 3126 0 0 0 EESPFAL_s2_0/x3
flabel metal1 808 -8256 869 -8196 4 FreeSans 3126 0 0 0 EESPFAL_s2_0/x3_bar
flabel metal2 7520 -5115 7540 -5095 4 FreeSans 2000 0 0 0 EESPFAL_s2_0/s2_bar
flabel metal2 7520 -4989 7540 -4969 4 FreeSans 2000 0 0 0 EESPFAL_s2_0/s2
flabel metal2 1151 -8475 1171 -8455 4 FreeSans 2000 0 0 0 EESPFAL_s2_0/CLK1
flabel metal2 1522 -8472 1542 -8452 4 FreeSans 2000 0 0 0 EESPFAL_s2_0/Dis1
flabel metal2 5342 -8474 5362 -8454 4 FreeSans 2000 0 0 0 EESPFAL_s2_0/Dis3
flabel metal2 5488 -8474 5508 -8454 4 FreeSans 2000 0 0 0 EESPFAL_s2_0/Dis2
flabel metal2 5576 -8474 5596 -8454 4 FreeSans 2000 0 0 0 EESPFAL_s2_0/CLK3
flabel metal2 5720 -8474 5740 -8454 4 FreeSans 2000 0 0 0 EESPFAL_s2_0/CLK2
rlabel metal1 2230 -6600 2270 -6560 4 EESPFAL_s2_0/EESPFAL_XOR_v3_1/OUT_bar
rlabel metal1 2180 -7280 2220 -7240 4 EESPFAL_s2_0/EESPFAL_XOR_v3_1/GND!
rlabel metal1 2180 -6100 2220 -6060 4 EESPFAL_s2_0/EESPFAL_XOR_v3_1/CLK
rlabel locali 2130 -6725 2170 -6685 4 EESPFAL_s2_0/EESPFAL_XOR_v3_1/OUT
rlabel locali 1070 -6220 1090 -6200 4 EESPFAL_s2_0/EESPFAL_XOR_v3_1/A
rlabel locali 1070 -6320 1090 -6300 4 EESPFAL_s2_0/EESPFAL_XOR_v3_1/A_bar
rlabel locali 1070 -6420 1090 -6400 4 EESPFAL_s2_0/EESPFAL_XOR_v3_1/B
rlabel locali 1070 -6520 1090 -6500 4 EESPFAL_s2_0/EESPFAL_XOR_v3_1/B_bar
rlabel locali 1980 -7160 2020 -7120 4 EESPFAL_s2_0/EESPFAL_XOR_v3_1/Dis
rlabel locali 2130 -5229 2170 -5189 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/OUT
rlabel locali 1070 -5819 1090 -5799 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/A
rlabel locali 1070 -5359 1090 -5339 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/A_bar
rlabel locali 1070 -5699 1090 -5679 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/B
rlabel locali 1070 -5259 1090 -5239 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/B_bar
rlabel locali 1070 -5579 1090 -5559 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/C
rlabel locali 1070 -5159 1090 -5139 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/C_bar
rlabel locali 1070 -5459 1090 -5439 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/D
rlabel locali 1070 -5059 1090 -5039 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/D_bar
rlabel locali 1980 -4579 2020 -4539 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/Dis
rlabel metal1 2230 -5369 2270 -5329 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/OUT_bar
rlabel metal1 2180 -4459 2220 -4419 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/GND!
rlabel metal1 2180 -5959 2220 -5919 2 EESPFAL_s2_0/EESPFAL_4in_NAND_0/CLK
rlabel metal1 4440 -6600 4480 -6560 4 EESPFAL_s2_0/EESPFAL_INV4_0/OUT
rlabel metal1 4390 -7280 4430 -7240 4 EESPFAL_s2_0/EESPFAL_INV4_0/GND!
rlabel metal1 4390 -6100 4430 -6060 4 EESPFAL_s2_0/EESPFAL_INV4_0/CLK
rlabel locali 4340 -6725 4380 -6685 4 EESPFAL_s2_0/EESPFAL_INV4_0/OUT_bar
rlabel locali 4970 -6480 5010 -6440 4 EESPFAL_s2_0/EESPFAL_INV4_0/A
rlabel locali 3810 -6720 3850 -6680 4 EESPFAL_s2_0/EESPFAL_INV4_0/A_bar
rlabel locali 4190 -7160 4230 -7120 4 EESPFAL_s2_0/EESPFAL_INV4_0/Dis
rlabel metal1 4441 -5140 4481 -5100 2 EESPFAL_s2_0/EESPFAL_INV4_2/OUT
rlabel metal1 4391 -4460 4431 -4420 2 EESPFAL_s2_0/EESPFAL_INV4_2/GND!
rlabel metal1 4391 -5640 4431 -5600 2 EESPFAL_s2_0/EESPFAL_INV4_2/CLK
rlabel locali 4341 -5015 4381 -4975 2 EESPFAL_s2_0/EESPFAL_INV4_2/OUT_bar
rlabel locali 4971 -5260 5011 -5220 2 EESPFAL_s2_0/EESPFAL_INV4_2/A
rlabel locali 3811 -5020 3851 -4980 2 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar
rlabel locali 4191 -4580 4231 -4540 2 EESPFAL_s2_0/EESPFAL_INV4_2/Dis
rlabel metal1 6319 -6600 6359 -6560 4 EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT_bar
rlabel metal1 6269 -7280 6309 -7240 4 EESPFAL_s2_0/EESPFAL_NAND_v3_0/GND!
rlabel metal1 6269 -6100 6309 -6060 4 EESPFAL_s2_0/EESPFAL_NAND_v3_0/CLK
rlabel locali 6219 -6725 6259 -6685 4 EESPFAL_s2_0/EESPFAL_NAND_v3_0/OUT
rlabel locali 5459 -6320 5479 -6300 4 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A
rlabel locali 5459 -6540 5479 -6520 4 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar
rlabel locali 5459 -6440 5479 -6420 4 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B
rlabel locali 5459 -6640 5479 -6620 4 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar
rlabel locali 6069 -7160 6109 -7120 4 EESPFAL_s2_0/EESPFAL_NAND_v3_0/Dis
rlabel metal1 6400 -5140 6440 -5100 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/OUT_bar
rlabel metal1 6450 -4460 6490 -4420 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/GND!
rlabel metal1 6450 -5640 6490 -5600 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/CLK
rlabel locali 6500 -5015 6540 -4975 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/OUT
rlabel locali 7430 -5500 7450 -5480 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/A
rlabel locali 7430 -5200 7450 -5180 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/A_bar
rlabel locali 7430 -5390 7450 -5370 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B
rlabel locali 7430 -5080 7450 -5060 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar
rlabel locali 7430 -5290 7450 -5270 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C
rlabel locali 7430 -4980 7450 -4960 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar
rlabel locali 6650 -4580 6690 -4540 8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/Dis
rlabel metal1 2230 -7960 2270 -7920 2 EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT_bar
rlabel metal1 2180 -7280 2220 -7240 2 EESPFAL_s2_0/EESPFAL_XOR_v3_0/GND!
rlabel metal1 2180 -8460 2220 -8420 2 EESPFAL_s2_0/EESPFAL_XOR_v3_0/CLK
rlabel locali 2130 -7835 2170 -7795 2 EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT
rlabel locali 1070 -8320 1090 -8300 2 EESPFAL_s2_0/EESPFAL_XOR_v3_0/A
rlabel locali 1070 -8220 1090 -8200 2 EESPFAL_s2_0/EESPFAL_XOR_v3_0/A_bar
rlabel locali 1070 -8120 1090 -8100 2 EESPFAL_s2_0/EESPFAL_XOR_v3_0/B
rlabel locali 1070 -8020 1090 -8000 2 EESPFAL_s2_0/EESPFAL_XOR_v3_0/B_bar
rlabel locali 1980 -7400 2020 -7360 2 EESPFAL_s2_0/EESPFAL_XOR_v3_0/Dis
rlabel metal1 4440 -7960 4480 -7920 2 EESPFAL_s2_0/EESPFAL_INV4_1/OUT
rlabel metal1 4390 -7280 4430 -7240 2 EESPFAL_s2_0/EESPFAL_INV4_1/GND!
rlabel metal1 4390 -8460 4430 -8420 2 EESPFAL_s2_0/EESPFAL_INV4_1/CLK
rlabel locali 4340 -7835 4380 -7795 2 EESPFAL_s2_0/EESPFAL_INV4_1/OUT_bar
rlabel locali 4970 -8080 5010 -8040 2 EESPFAL_s2_0/EESPFAL_INV4_1/A
rlabel locali 3810 -7840 3850 -7800 2 EESPFAL_s2_0/EESPFAL_INV4_1/A_bar
rlabel locali 4190 -7400 4230 -7360 2 EESPFAL_s2_0/EESPFAL_INV4_1/Dis
rlabel metal1 6319 -7960 6359 -7920 2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar
rlabel metal1 6269 -7280 6309 -7240 2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/GND!
rlabel metal1 6269 -8460 6309 -8420 2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/CLK
rlabel locali 6219 -7835 6259 -7795 2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT
rlabel locali 5459 -8220 5479 -8200 2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A
rlabel locali 5459 -8000 5479 -7980 2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar
rlabel locali 5459 -8100 5479 -8080 2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B
rlabel locali 5459 -7900 5479 -7880 2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar
rlabel locali 6069 -7400 6109 -7360 2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/Dis
flabel metal1 930 -1562 974 -1516 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/GND
flabel metal1 10 -543 71 -483 2 FreeSans 2500 0 0 0 EESPFAL_s1_0/x0
flabel metal1 123 -604 184 -544 2 FreeSans 2500 0 0 0 EESPFAL_s1_0/x0_bar
flabel metal1 238 -543 299 -483 2 FreeSans 2500 0 0 0 EESPFAL_s1_0/x1
flabel metal1 352 -604 413 -544 2 FreeSans 2500 0 0 0 EESPFAL_s1_0/x1_bar
flabel metal1 466 -542 527 -482 2 FreeSans 2500 0 0 0 EESPFAL_s1_0/x2
flabel metal1 579 -603 640 -543 2 FreeSans 2500 0 0 0 EESPFAL_s1_0/x2_bar
flabel metal1 694 -542 755 -482 2 FreeSans 2500 0 0 0 EESPFAL_s1_0/x3
flabel metal1 808 -603 869 -543 2 FreeSans 2500 0 0 0 EESPFAL_s1_0/x3_bar
flabel metal2 7260 -3706 7280 -3686 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/s1_bar
flabel metal2 7260 -3812 7280 -3791 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/s1
flabel metal2 7271 -3697 7271 -3697 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/s1_bar
flabel metal2 7270 -3802 7270 -3802 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/s1
flabel metal2 7271 -3697 7271 -3697 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/s1_bar
flabel metal2 7270 -3802 7270 -3802 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/s1
flabel metal2 7271 -3697 7271 -3697 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/s1_bar
flabel metal2 7270 -3802 7270 -3802 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/s1
flabel metal2 1080 -360 1111 -329 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/CLK1
flabel metal2 1200 -354 1223 -330 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/Dis1
flabel metal2 5167 -347 5186 -326 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/Dis3
flabel metal2 5278 -350 5303 -325 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/CLK3
flabel metal2 5406 -348 5431 -324 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/Dis2
flabel metal2 7014 -367 7048 -333 2 FreeSans 2000 0 0 0 EESPFAL_s1_0/CLK2
rlabel metal1 2191 -3699 2231 -3659 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/OUT_bar
rlabel metal1 2141 -4379 2181 -4339 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/GND!
rlabel metal1 2141 -3199 2181 -3159 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/CLK
rlabel locali 2091 -3824 2131 -3784 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/OUT
rlabel locali 1181 -3309 1201 -3289 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A
rlabel locali 1181 -3619 1201 -3599 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A_bar
rlabel locali 1181 -3429 1201 -3409 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B
rlabel locali 1181 -3699 1201 -3679 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B_bar
rlabel locali 1181 -3539 1201 -3519 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C
rlabel locali 1181 -3799 1201 -3779 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C_bar
rlabel locali 1941 -4259 1981 -4219 4 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/Dis
rlabel metal1 4241 -3699 4281 -3659 4 EESPFAL_s1_0/EESPFAL_INV4_0/OUT
rlabel metal1 4191 -4379 4231 -4339 4 EESPFAL_s1_0/EESPFAL_INV4_0/GND!
rlabel metal1 4191 -3199 4231 -3159 4 EESPFAL_s1_0/EESPFAL_INV4_0/CLK
rlabel locali 4141 -3824 4181 -3784 4 EESPFAL_s1_0/EESPFAL_INV4_0/OUT_bar
rlabel locali 4771 -3579 4811 -3539 4 EESPFAL_s1_0/EESPFAL_INV4_0/A
rlabel locali 3611 -3819 3651 -3779 4 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar
rlabel locali 3991 -4259 4031 -4219 4 EESPFAL_s1_0/EESPFAL_INV4_0/Dis
rlabel metal1 6181 -3700 6221 -3660 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/OUT_bar
rlabel metal1 6231 -4380 6271 -4340 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/GND!
rlabel metal1 6231 -3200 6271 -3160 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/CLK
rlabel locali 6281 -3825 6321 -3785 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/OUT
rlabel locali 7211 -3320 7231 -3300 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/A
rlabel locali 7211 -3620 7231 -3600 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/A_bar
rlabel locali 7211 -3430 7231 -3410 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/B
rlabel locali 7211 -3740 7231 -3720 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/B_bar
rlabel locali 7211 -3530 7231 -3510 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C
rlabel locali 7211 -3840 7231 -3820 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar
rlabel locali 6431 -4260 6471 -4220 6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/Dis
rlabel metal1 2190 -2239 2230 -2199 2 EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT_bar
rlabel metal1 2140 -1559 2180 -1519 2 EESPFAL_s1_0/EESPFAL_XOR_v3_1/GND!
rlabel metal1 2140 -2739 2180 -2699 2 EESPFAL_s1_0/EESPFAL_XOR_v3_1/CLK
rlabel locali 2090 -2114 2130 -2074 2 EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT
rlabel locali 1030 -2599 1050 -2579 2 EESPFAL_s1_0/EESPFAL_XOR_v3_1/A
rlabel locali 1030 -2499 1050 -2479 2 EESPFAL_s1_0/EESPFAL_XOR_v3_1/A_bar
rlabel locali 1030 -2399 1050 -2379 2 EESPFAL_s1_0/EESPFAL_XOR_v3_1/B
rlabel locali 1030 -2299 1050 -2279 2 EESPFAL_s1_0/EESPFAL_XOR_v3_1/B_bar
rlabel locali 1940 -1679 1980 -1639 2 EESPFAL_s1_0/EESPFAL_XOR_v3_1/Dis
rlabel metal1 4380 -2239 4420 -2199 2 EESPFAL_s1_0/EESPFAL_INV4_1/OUT
rlabel metal1 4330 -1559 4370 -1519 2 EESPFAL_s1_0/EESPFAL_INV4_1/GND!
rlabel metal1 4330 -2739 4370 -2699 2 EESPFAL_s1_0/EESPFAL_INV4_1/CLK
rlabel locali 4280 -2114 4320 -2074 2 EESPFAL_s1_0/EESPFAL_INV4_1/OUT_bar
rlabel locali 4910 -2359 4950 -2319 2 EESPFAL_s1_0/EESPFAL_INV4_1/A
rlabel locali 3750 -2119 3790 -2079 2 EESPFAL_s1_0/EESPFAL_INV4_1/A_bar
rlabel locali 4130 -1679 4170 -1639 2 EESPFAL_s1_0/EESPFAL_INV4_1/Dis
rlabel metal1 6260 -2239 6300 -2199 2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar
rlabel metal1 6210 -1559 6250 -1519 2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/GND!
rlabel metal1 6210 -2739 6250 -2699 2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/CLK
rlabel locali 6160 -2114 6200 -2074 2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT
rlabel locali 5400 -2499 5420 -2479 2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A
rlabel locali 5400 -2279 5420 -2259 2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar
rlabel locali 5400 -2379 5420 -2359 2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B
rlabel locali 5400 -2179 5420 -2159 2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar
rlabel locali 6010 -1679 6050 -1639 2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/Dis
rlabel metal1 2190 -879 2230 -839 4 EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT_bar
rlabel metal1 2140 -1559 2180 -1519 4 EESPFAL_s1_0/EESPFAL_XOR_v3_0/GND!
rlabel metal1 2140 -379 2180 -339 4 EESPFAL_s1_0/EESPFAL_XOR_v3_0/CLK
rlabel locali 2090 -1004 2130 -964 4 EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT
rlabel locali 1030 -499 1050 -479 4 EESPFAL_s1_0/EESPFAL_XOR_v3_0/A
rlabel locali 1030 -599 1050 -579 4 EESPFAL_s1_0/EESPFAL_XOR_v3_0/A_bar
rlabel locali 1030 -699 1050 -679 4 EESPFAL_s1_0/EESPFAL_XOR_v3_0/B
rlabel locali 1030 -799 1050 -779 4 EESPFAL_s1_0/EESPFAL_XOR_v3_0/B_bar
rlabel locali 1940 -1439 1980 -1399 4 EESPFAL_s1_0/EESPFAL_XOR_v3_0/Dis
rlabel metal1 4380 -879 4420 -839 4 EESPFAL_s1_0/EESPFAL_INV4_2/OUT
rlabel metal1 4330 -1559 4370 -1519 4 EESPFAL_s1_0/EESPFAL_INV4_2/GND!
rlabel metal1 4330 -379 4370 -339 4 EESPFAL_s1_0/EESPFAL_INV4_2/CLK
rlabel locali 4280 -1004 4320 -964 4 EESPFAL_s1_0/EESPFAL_INV4_2/OUT_bar
rlabel locali 4910 -759 4950 -719 4 EESPFAL_s1_0/EESPFAL_INV4_2/A
rlabel locali 3750 -999 3790 -959 4 EESPFAL_s1_0/EESPFAL_INV4_2/A_bar
rlabel locali 4130 -1439 4170 -1399 4 EESPFAL_s1_0/EESPFAL_INV4_2/Dis
rlabel metal1 6260 -879 6300 -839 4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar
rlabel metal1 6210 -1559 6250 -1519 4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/GND!
rlabel metal1 6210 -379 6250 -339 4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/CLK
rlabel locali 6160 -1004 6200 -964 4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT
rlabel locali 5400 -599 5420 -579 4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A
rlabel locali 5400 -819 5420 -799 4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar
rlabel locali 5400 -719 5420 -699 4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B
rlabel locali 5400 -919 5420 -899 4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar
rlabel locali 6010 -1439 6050 -1399 4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/Dis
flabel metal1 930 1258 975 1303 2 FreeSans 2000 0 0 0 EESPFAL_s0_0/GND
flabel metal1 10 2277 71 2337 2 FreeSans 2500 0 0 0 EESPFAL_s0_0/x0
flabel metal1 123 2216 184 2276 2 FreeSans 2500 0 0 0 EESPFAL_s0_0/x0_bar
flabel metal1 238 2277 299 2337 2 FreeSans 2500 0 0 0 EESPFAL_s0_0/x1
flabel metal1 352 2216 413 2276 2 FreeSans 2500 0 0 0 EESPFAL_s0_0/x1_bar
flabel metal1 466 2278 527 2338 2 FreeSans 2500 0 0 0 EESPFAL_s0_0/x2
flabel metal1 579 2217 640 2277 2 FreeSans 2500 0 0 0 EESPFAL_s0_0/x2_bar
flabel metal1 694 2278 755 2338 2 FreeSans 2500 0 0 0 EESPFAL_s0_0/x3
flabel metal1 808 2217 869 2277 2 FreeSans 2500 0 0 0 EESPFAL_s0_0/x3_bar
flabel metal2 7485 711 7500 726 2 FreeSans 2000 0 0 0 EESPFAL_s0_0/s0
flabel metal2 7485 591 7500 606 2 FreeSans 2000 0 0 0 EESPFAL_s0_0/s0_bar
flabel metal2 1038 2445 1078 2485 2 FreeSans 2000 0 0 0 EESPFAL_s0_0/CLK1
flabel metal2 1160 2461 1180 2481 2 FreeSans 2000 0 0 0 EESPFAL_s0_0/Dis1
flabel metal2 5770 2476 5785 2491 2 FreeSans 2000 0 0 0 EESPFAL_s0_0/Dis2
flabel metal2 5860 2476 5875 2491 2 FreeSans 2000 0 0 0 EESPFAL_s0_0/CLK2
flabel metal2 5955 2476 5970 2491 2 FreeSans 2000 0 0 0 EESPFAL_s0_0/Dis3
flabel metal2 5488 2473 5508 2493 2 FreeSans 2000 0 0 0 EESPFAL_s0_0/CLK3
rlabel metal1 2190 1941 2230 1981 4 EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT_bar
rlabel metal1 2140 1261 2180 1301 4 EESPFAL_s0_0/EESPFAL_XOR_v3_0/GND!
rlabel metal1 2140 2441 2180 2481 4 EESPFAL_s0_0/EESPFAL_XOR_v3_0/CLK
rlabel locali 2090 1816 2130 1856 4 EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT
rlabel locali 1030 2321 1050 2341 4 EESPFAL_s0_0/EESPFAL_XOR_v3_0/A
rlabel locali 1030 2221 1050 2241 4 EESPFAL_s0_0/EESPFAL_XOR_v3_0/A_bar
rlabel locali 1030 2121 1050 2141 4 EESPFAL_s0_0/EESPFAL_XOR_v3_0/B
rlabel locali 1030 2021 1050 2041 4 EESPFAL_s0_0/EESPFAL_XOR_v3_0/B_bar
rlabel locali 1940 1381 1980 1421 4 EESPFAL_s0_0/EESPFAL_XOR_v3_0/Dis
rlabel metal1 2190 581 2230 621 2 EESPFAL_s0_0/EESPFAL_NAND_v3_2/OUT_bar
rlabel metal1 2140 1261 2180 1301 2 EESPFAL_s0_0/EESPFAL_NAND_v3_2/GND!
rlabel metal1 2140 81 2180 121 2 EESPFAL_s0_0/EESPFAL_NAND_v3_2/CLK
rlabel locali 2090 706 2130 746 2 EESPFAL_s0_0/EESPFAL_NAND_v3_2/OUT
rlabel locali 1330 321 1350 341 2 EESPFAL_s0_0/EESPFAL_NAND_v3_2/A
rlabel locali 1330 541 1350 561 2 EESPFAL_s0_0/EESPFAL_NAND_v3_2/A_bar
rlabel locali 1330 441 1350 461 2 EESPFAL_s0_0/EESPFAL_NAND_v3_2/B
rlabel locali 1330 641 1350 661 2 EESPFAL_s0_0/EESPFAL_NAND_v3_2/B_bar
rlabel locali 1940 1141 1980 1181 2 EESPFAL_s0_0/EESPFAL_NAND_v3_2/Dis
rlabel locali 4410 1816 4450 1856 4 EESPFAL_s0_0/EESPFAL_NOR_v3_1/OUT
rlabel locali 3650 2191 3670 2211 4 EESPFAL_s0_0/EESPFAL_NOR_v3_1/A
rlabel locali 3650 1871 3670 1891 4 EESPFAL_s0_0/EESPFAL_NOR_v3_1/A_bar
rlabel locali 3650 2071 3670 2091 4 EESPFAL_s0_0/EESPFAL_NOR_v3_1/B
rlabel locali 3650 1971 3670 1991 4 EESPFAL_s0_0/EESPFAL_NOR_v3_1/B_bar
rlabel locali 4260 1381 4300 1421 4 EESPFAL_s0_0/EESPFAL_NOR_v3_1/Dis
rlabel metal1 4510 1941 4550 1981 4 EESPFAL_s0_0/EESPFAL_NOR_v3_1/OUT_bar
rlabel metal1 4460 1261 4500 1301 4 EESPFAL_s0_0/EESPFAL_NOR_v3_1/GND!
rlabel metal1 4460 2441 4500 2481 4 EESPFAL_s0_0/EESPFAL_NOR_v3_1/CLK
rlabel metal1 4510 581 4550 621 2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/OUT_bar
rlabel metal1 4460 1261 4500 1301 2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/GND!
rlabel metal1 4460 81 4500 121 2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/CLK
rlabel locali 4410 706 4450 746 2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/OUT
rlabel locali 3650 321 3670 341 2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/A
rlabel locali 3650 541 3670 561 2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/A_bar
rlabel locali 3650 441 3670 461 2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B
rlabel locali 3650 641 3670 661 2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar
rlabel locali 4260 1141 4300 1181 2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/Dis
rlabel locali 6530 706 6570 746 8 EESPFAL_s0_0/EESPFAL_NOR_v3_0/OUT
rlabel locali 7310 351 7330 371 8 EESPFAL_s0_0/EESPFAL_NOR_v3_0/A
rlabel locali 7310 671 7330 691 8 EESPFAL_s0_0/EESPFAL_NOR_v3_0/A_bar
rlabel locali 7310 471 7330 491 8 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B
rlabel locali 7310 571 7330 591 8 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar
rlabel locali 6680 1141 6720 1181 8 EESPFAL_s0_0/EESPFAL_NOR_v3_0/Dis
rlabel metal1 6430 581 6470 621 8 EESPFAL_s0_0/EESPFAL_NOR_v3_0/OUT_bar
rlabel metal1 6480 1261 6520 1301 8 EESPFAL_s0_0/EESPFAL_NOR_v3_0/GND!
rlabel metal1 6480 81 6520 121 8 EESPFAL_s0_0/EESPFAL_NOR_v3_0/CLK
rlabel metal1 6530 1941 6570 1981 4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar
rlabel metal1 6480 1261 6520 1301 4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/GND!
rlabel metal1 6480 2441 6520 2481 4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/CLK
rlabel locali 6430 1816 6470 1856 4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT
rlabel locali 5670 2221 5690 2241 4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A
rlabel locali 5670 2001 5690 2021 4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar
rlabel locali 5670 2101 5690 2121 4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B
rlabel locali 5670 1901 5690 1921 4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar
rlabel locali 6280 1381 6320 1421 4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/Dis
<< end >>
