magic
tech sky130A
magscale 1 2
timestamp 1670967196
<< locali >>
rect -34 600 34 657
rect -34 -657 34 -600
<< rlocali >>
rect -34 -600 34 600
<< properties >>
string gencell sky130_fd_pr__res_generic_l1
string library sky130
string parameters w 0.34 l 6 m 1 nx 1 wmin 0.17 lmin 0.17 rho 12.8 val 225.882 dummy 0 dw 0.0 term 0.0 snake 0 roverlap 0
<< end >>
