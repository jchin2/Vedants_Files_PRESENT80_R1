.subckt Power_Amp_LVS_1 Input VDD Ground
*.PININFO Input:I VDD:I Ground:B
XM1 VDD Input Ground Ground sky130_fd_pr__nfet_01v8_lvt L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20 
XC1 VDD Ground sky130_fd_pr__cap_mim_m3_1 W=12.05 L=12.05 MF=1 m=1
R1 Ground net1 sky130_fd_pr__res_generic_po W=1.6 L=1.66 m=1
XC2 VDD net1 sky130_fd_pr__cap_mim_m3_1 W=8.8 L=9 MF=1 m=1
.ends
** flattened .save nodes
.end
