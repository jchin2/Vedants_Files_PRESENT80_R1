magic
tech sky130A
magscale 1 2
timestamp 1670990700
<< xpolycontact >>
rect -35 98 35 530
rect -35 -530 35 -98
<< ppolyres >>
rect -35 -98 35 98
<< viali >>
rect -19 115 19 512
rect -19 -512 19 -115
<< metal1 >>
rect -25 512 25 524
rect -25 115 -19 512
rect 19 115 25 512
rect -25 103 25 115
rect -25 -115 25 -103
rect -25 -512 -19 -115
rect 19 -512 25 -115
rect -25 -524 25 -512
<< res0p35 >>
rect -37 -100 37 100
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 0.98 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 2.008k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 0 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
