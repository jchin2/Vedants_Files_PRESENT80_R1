* NGSPICE file created from CMOS_s2_flat.ext - technology: sky130A

.subckt CMOS_s2_flat GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar s2 VDD
X0 s2.t1 a_2442_n779# GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_2592_n1689# CMOS_AND_1/AND VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X2 VDD.t1 x0.t0 a_1735_499# VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X3 a_2592_n111# x2_bar.t0 GND.t9 GND.t0 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_2592_499# CMOS_AND_0/A a_2592_n111# GND.t30 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 CMOS_AND_1/AND a_1380_n1689# GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_1380_n1689# x1_bar.t0 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X7 a_2742_n1689# CMOS_AND_0/AND a_2592_n1689# VDD.t41 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X8 VDD.t28 x2.t0 a_177_499# VDD.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X9 CMOS_AND_1/A a_27_n111# VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X10 GND.t1 CMOS_AND_1/AND a_2442_n779# GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X11 a_2442_n779# CMOS_AND_0/AND GND.t36 GND.t30 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 VDD.t11 CMOS_AND_1/A a_1380_n1689# VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X13 GND.t25 x3_bar.t0 a_177_n111# GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X14 a_27_n111# x2.t1 a_n123_n111# GND.t22 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X15 a_n178_n1689# x1.t0 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=3.6e+12p pd=1.44e+07u as=0p ps=0u w=3e+06u l=150000u
X16 a_27_n111# x3.t0 a_n123_499# VDD.t32 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X17 CMOS_4in_AND_0/OUT.t0 a_n178_n1689# GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 GND.t18 CMOS_4in_AND_0/OUT.t2 a_2442_n779# GND.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_n178_n1689# x2.t2 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X20 CMOS_AND_0/AND a_2592_499# VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X21 a_1435_n111# x1.t1 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X22 a_1380_n779# x1_bar.t1 GND.t29 GND.t28 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X23 a_1380_n1689# CMOS_AND_1/A a_1380_n779# GND.t8 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X24 s2.t0 a_2442_n779# VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X25 a_1435_499# x0_bar.t0 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X26 a_n123_499# x2_bar.t1 VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X27 a_n28_n779# x0.t1 a_n178_n779# GND.t12 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X28 a_122_n779# x1.t2 a_n28_n779# GND.t23 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X29 VDD.t34 CMOS_AND_0/A a_2592_499# VDD.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X30 VDD.t13 x0.t2 a_n178_n1689# VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X31 CMOS_AND_1/AND a_1380_n1689# VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X32 a_1735_499# x1_bar.t2 CMOS_AND_0/A VDD.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X33 a_177_499# x3_bar.t1 a_27_n111# VDD.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X34 CMOS_AND_0/A x0.t3 a_1435_n111# GND.t14 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X35 a_1735_n111# x0_bar.t1 CMOS_AND_0/A GND.t19 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X36 CMOS_AND_0/AND a_2592_499# GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X37 a_2442_n779# CMOS_4in_AND_0/OUT.t3 a_2742_n1689# VDD.t18 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X38 a_n123_n111# x3.t1 GND.t27 GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X39 a_n178_n779# x2.t3 GND.t33 GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X40 CMOS_4in_AND_0/OUT.t1 a_n178_n1689# VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X41 a_177_n111# x2_bar.t2 a_27_n111# GND.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X42 VDD.t30 x3_bar.t2 a_n178_n1689# VDD.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X43 a_2592_499# x2_bar.t3 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X44 CMOS_AND_1/A a_27_n111# GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X45 GND.t16 x1_bar.t3 a_1735_n111# GND.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X46 CMOS_AND_0/A x1.t3 a_1435_499# VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X47 a_n178_n1689# x3_bar.t3 a_122_n779# GND.t31 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
R0 GND.n104 GND.t22 150.98
R1 GND.n80 GND.t14 150.98
R2 GND.n92 GND.t26 133.725
R3 GND.n160 GND.t20 133.725
R4 GND.n112 GND.t13 125.098
R5 GND.n72 GND.t19 125.098
R6 GND.n138 GND.t6 103.529
R7 GND.n92 GND.t32 103.529
R8 GND.n45 GND.t0 103.529
R9 GND.n160 GND.t28 103.529
R10 GND.n120 GND.t24 99.215
R11 GND.n63 GND.t15 99.215
R12 GND.n143 GND.t4 77.647
R13 GND.n101 GND.t12 77.647
R14 GND.n5 GND.t2 77.647
R15 GND.n36 GND.t30 77.647
R16 GND.n168 GND.t8 77.647
R17 GND.n108 GND.t23 51.764
R18 GND.n14 GND.t34 51.764
R19 GND.n28 GND.t17 51.764
R20 GND.n63 GND.t10 51.764
R21 GND.n85 GND 37.93
R22 GND.n91 GND.t27 30.21
R23 GND.n86 GND.t33 30.21
R24 GND.n137 GND.t7 30.21
R25 GND.n154 GND.t29 30.21
R26 GND.n67 GND.t11 30.21
R27 GND.n27 GND.t18 30.21
R28 GND.n9 GND.t3 30.21
R29 GND.n18 GND.t35 30.21
R30 GND.n53 GND.t9 30.21
R31 GND.n62 GND.t16 30.21
R32 GND.n159 GND.t21 30.21
R33 GND.n142 GND.t5 30.21
R34 GND.n124 GND.t25 30.21
R35 GND.n116 GND.t31 25.882
R36 GND.n0 GND.t36 24
R37 GND.n0 GND.t1 24
R38 GND.n38 GND.n35 11.52
R39 GND.n106 GND.n103 11.52
R40 GND.n3 GND.n2 9.154
R41 GND.n60 GND.n59 9.154
R42 GND.n65 GND.n64 9.154
R43 GND.n64 GND.n63 9.154
R44 GND.n70 GND.n69 9.154
R45 GND.n69 GND.n68 9.154
R46 GND.n74 GND.n73 9.154
R47 GND.n73 GND.n72 9.154
R48 GND.n78 GND.n77 9.154
R49 GND.n77 GND.n76 9.154
R50 GND.n82 GND.n81 9.154
R51 GND.n81 GND.n80 9.154
R52 GND.n170 GND.n169 9.154
R53 GND.n169 GND.n168 9.154
R54 GND.n166 GND.n165 9.154
R55 GND.n165 GND.n164 9.154
R56 GND.n162 GND.n161 9.154
R57 GND.n161 GND.n160 9.154
R58 GND.n157 GND.n156 9.154
R59 GND.n7 GND.n6 9.154
R60 GND.n6 GND.n5 9.154
R61 GND.n12 GND.n11 9.154
R62 GND.n11 GND.n10 9.154
R63 GND.n16 GND.n15 9.154
R64 GND.n15 GND.n14 9.154
R65 GND.n21 GND.n20 9.154
R66 GND.n20 GND.n19 9.154
R67 GND.n25 GND.n24 9.154
R68 GND.n24 GND.n23 9.154
R69 GND.n30 GND.n29 9.154
R70 GND.n29 GND.n28 9.154
R71 GND.n35 GND.n34 9.154
R72 GND.n34 GND.n33 9.154
R73 GND.n38 GND.n37 9.154
R74 GND.n37 GND.n36 9.154
R75 GND.n42 GND.n41 9.154
R76 GND.n41 GND.n40 9.154
R77 GND.n47 GND.n46 9.154
R78 GND.n46 GND.n45 9.154
R79 GND.n51 GND.n50 9.154
R80 GND.n149 GND.n148 9.154
R81 GND.n145 GND.n144 9.154
R82 GND.n144 GND.n143 9.154
R83 GND.n140 GND.n139 9.154
R84 GND.n139 GND.n138 9.154
R85 GND.n135 GND.n134 9.154
R86 GND.n134 GND.n133 9.154
R87 GND.n131 GND.n130 9.154
R88 GND.n130 GND.n129 9.154
R89 GND.n127 GND.n126 9.154
R90 GND.n126 GND.n125 9.154
R91 GND.n122 GND.n121 9.154
R92 GND.n121 GND.n120 9.154
R93 GND.n118 GND.n117 9.154
R94 GND.n117 GND.n116 9.154
R95 GND.n114 GND.n113 9.154
R96 GND.n113 GND.n112 9.154
R97 GND.n110 GND.n109 9.154
R98 GND.n109 GND.n108 9.154
R99 GND.n106 GND.n105 9.154
R100 GND.n105 GND.n104 9.154
R101 GND.n103 GND.n102 9.154
R102 GND.n102 GND.n101 9.154
R103 GND.n98 GND.n97 9.154
R104 GND.n97 GND.n96 9.154
R105 GND.n94 GND.n93 9.154
R106 GND.n93 GND.n92 9.154
R107 GND.n89 GND.n88 9.154
R108 GND.n2 GND.n1 8.108
R109 GND.n44 GND.n0 6.21
R110 GND.n86 GND.n85 4.706
R111 GND.n153 GND.n84 4.65
R112 GND.n61 GND.n60 4.65
R113 GND.n66 GND.n65 4.65
R114 GND.n71 GND.n70 4.65
R115 GND.n75 GND.n74 4.65
R116 GND.n79 GND.n78 4.65
R117 GND.n83 GND.n82 4.65
R118 GND.n171 GND.n170 4.65
R119 GND.n167 GND.n166 4.65
R120 GND.n163 GND.n162 4.65
R121 GND.n158 GND.n157 4.65
R122 GND.n57 GND.n56 4.65
R123 GND.n55 GND.n54 4.65
R124 GND.n8 GND.n7 4.65
R125 GND.n13 GND.n12 4.65
R126 GND.n17 GND.n16 4.65
R127 GND.n22 GND.n21 4.65
R128 GND.n26 GND.n25 4.65
R129 GND.n31 GND.n30 4.65
R130 GND.n35 GND.n32 4.65
R131 GND.n39 GND.n38 4.65
R132 GND.n43 GND.n42 4.65
R133 GND.n48 GND.n47 4.65
R134 GND.n52 GND.n51 4.65
R135 GND.n150 GND.n149 4.65
R136 GND.n146 GND.n145 4.65
R137 GND.n141 GND.n140 4.65
R138 GND.n136 GND.n135 4.65
R139 GND.n132 GND.n131 4.65
R140 GND.n128 GND.n127 4.65
R141 GND.n123 GND.n122 4.65
R142 GND.n119 GND.n118 4.65
R143 GND.n115 GND.n114 4.65
R144 GND.n111 GND.n110 4.65
R145 GND.n107 GND.n106 4.65
R146 GND.n103 GND.n100 4.65
R147 GND.n99 GND.n98 4.65
R148 GND.n95 GND.n94 4.65
R149 GND.n90 GND.n89 4.65
R150 GND.n152 GND.n151 4.65
R151 GND.n50 GND.n49 2.759
R152 GND.n4 GND.n3 2.562
R153 GND.n8 GND.n4 1.145
R154 GND.n57 GND.n55 0.525
R155 GND.n153 GND.n152 0.507
R156 GND.n17 GND.n13 0.09
R157 GND.n26 GND.n22 0.09
R158 GND.n32 GND.n31 0.09
R159 GND.n43 GND.n39 0.09
R160 GND.n52 GND.n48 0.09
R161 GND.n61 GND.n57 0.09
R162 GND.n75 GND.n71 0.09
R163 GND.n79 GND.n75 0.09
R164 GND.n83 GND.n79 0.09
R165 GND.n171 GND.n167 0.09
R166 GND.n167 GND.n163 0.09
R167 GND.n152 GND.n150 0.09
R168 GND.n150 GND.n146 0.09
R169 GND.n136 GND.n132 0.09
R170 GND.n132 GND.n128 0.09
R171 GND.n123 GND.n119 0.09
R172 GND.n119 GND.n115 0.09
R173 GND.n115 GND.n111 0.09
R174 GND.n111 GND.n107 0.09
R175 GND.n100 GND.n99 0.09
R176 GND.n99 GND.n95 0.09
R177 GND.n148 GND.n147 0.088
R178 GND.n18 GND.n17 0.078
R179 GND.n31 GND.n27 0.078
R180 GND.n67 GND.n66 0.078
R181 GND.n156 GND.n155 0.074
R182 GND.n88 GND.n87 0.074
R183 GND.n9 GND.n8 0.072
R184 GND.n146 GND.n142 0.071
R185 GND.n39 CMOS_AND_0/GND 0.065
R186 GND.n66 GND.n62 0.065
R187 CMOS_AND_1/GND GND.n171 0.065
R188 GND.n124 GND.n123 0.065
R189 GND.n100 GND 0.065
R190 GND.n48 GND.n44 0.063
R191 GND.n141 GND.n137 0.063
R192 GND.n55 GND.n53 0.056
R193 GND.n154 GND.n153 0.056
R194 GND.n163 GND.n159 0.055
R195 GND.n95 GND.n91 0.055
R196 GND.n59 GND.n58 0.047
R197 GND.n159 GND.n158 0.035
R198 GND.n91 GND.n90 0.035
R199 GND.n53 GND.n52 0.033
R200 GND.n158 GND.n154 0.033
R201 GND.n90 GND.n86 0.033
R202 GND.n44 GND.n43 0.026
R203 GND.n137 GND.n136 0.026
R204 GND.n32 CMOS_AND_0/GND 0.025
R205 GND.n62 GND.n61 0.025
R206 CMOS_AND_1/GND GND.n83 0.025
R207 GND.n128 GND.n124 0.025
R208 GND.n107 GND 0.025
R209 GND.n142 GND.n141 0.018
R210 GND.n13 GND.n9 0.017
R211 GND.n22 GND.n18 0.011
R212 GND.n27 GND.n26 0.011
R213 GND.n71 GND.n67 0.011
R214 s2.n2 s2.t0 120.552
R215 s2.n1 s2.t1 98.438
R216 s2 s2.n2 7.84
R217 s2 s2.n1 3.68
R218 s2.n1 s2.n0 3.084
R219 s2.n0 s2 0.374
R220 VDD.n72 VDD.t26 38.206
R221 VDD.n135 VDD.t32 36.141
R222 VDD.n311 VDD.t35 32.01
R223 VDD.n80 VDD.t21 32.01
R224 VDD.n127 VDD.t31 29.945
R225 VDD.n60 VDD.t23 29.945
R226 VDD.n34 VDD.t37 24.782
R227 VDD.n180 VDD.t2 24.782
R228 VDD.n227 VDD.t16 24.782
R229 VDD.n244 VDD.t8 24.782
R230 VDD.n292 VDD.t19 24.782
R231 VDD.n119 VDD.t27 23.75
R232 VDD.n52 VDD.t0 23.75
R233 VDD.n310 VDD.t36 22.029
R234 VDD.n118 VDD.t28 22.029
R235 VDD.n101 VDD.t7 22.029
R236 VDD.n84 VDD.t22 22.029
R237 VDD.n51 VDD.t1 22.029
R238 VDD.n42 VDD.t38 22.029
R239 VDD.n21 VDD.t34 22.029
R240 VDD.n8 VDD.t40 22.029
R241 VDD.n147 VDD.t5 22.029
R242 VDD.n188 VDD.t3 22.029
R243 VDD.n201 VDD.t15 22.029
R244 VDD.n214 VDD.t11 22.029
R245 VDD.n235 VDD.t17 22.029
R246 VDD.n248 VDD.t9 22.029
R247 VDD.n265 VDD.t30 22.029
R248 VDD.n300 VDD.t20 22.029
R249 VDD.n278 VDD.t25 19.7
R250 VDD.n278 VDD.t13 19.7
R251 VDD.n97 VDD.t6 18.586
R252 VDD.n26 VDD.t33 18.586
R253 VDD.n143 VDD.t4 18.586
R254 VDD.n172 VDD.t41 18.586
R255 VDD.n219 VDD.t10 18.586
R256 VDD.n284 VDD.t12 18.586
R257 VDD.n4 VDD.t39 12.391
R258 VDD.n164 VDD.t18 12.391
R259 VDD.n197 VDD.t14 12.391
R260 VDD.n274 VDD.t24 12.391
R261 VDD.n74 VDD.n71 11.52
R262 VDD.n28 VDD.n25 11.52
R263 VDD.n174 VDD.n171 11.52
R264 VDD.n221 VDD.n218 11.52
R265 VDD.n286 VDD.n283 11.52
R266 VDD.n141 VDD.n140 8.855
R267 VDD.n195 VDD.n194 8.855
R268 VDD.n242 VDD.n241 8.855
R269 VDD.n246 VDD.n245 8.855
R270 VDD.n245 VDD.n244 8.855
R271 VDD.n251 VDD.n250 8.855
R272 VDD.n250 VDD.n249 8.855
R273 VDD.n255 VDD.n254 8.855
R274 VDD.n254 VDD.n253 8.855
R275 VDD.n259 VDD.n258 8.855
R276 VDD.n258 VDD.n257 8.855
R277 VDD.n263 VDD.n262 8.855
R278 VDD.n262 VDD.n261 8.855
R279 VDD.n268 VDD.n267 8.855
R280 VDD.n267 VDD.n266 8.855
R281 VDD.n272 VDD.n271 8.855
R282 VDD.n271 VDD.n270 8.855
R283 VDD.n276 VDD.n275 8.855
R284 VDD.n275 VDD.n274 8.855
R285 VDD.n283 VDD.n282 8.855
R286 VDD.n282 VDD.n281 8.855
R287 VDD.n286 VDD.n285 8.855
R288 VDD.n285 VDD.n284 8.855
R289 VDD.n290 VDD.n289 8.855
R290 VDD.n289 VDD.n288 8.855
R291 VDD.n294 VDD.n293 8.855
R292 VDD.n293 VDD.n292 8.855
R293 VDD.n298 VDD.n297 8.855
R294 VDD.n199 VDD.n198 8.855
R295 VDD.n198 VDD.n197 8.855
R296 VDD.n204 VDD.n203 8.855
R297 VDD.n203 VDD.n202 8.855
R298 VDD.n208 VDD.n207 8.855
R299 VDD.n207 VDD.n206 8.855
R300 VDD.n212 VDD.n211 8.855
R301 VDD.n211 VDD.n210 8.855
R302 VDD.n218 VDD.n217 8.855
R303 VDD.n217 VDD.n216 8.855
R304 VDD.n221 VDD.n220 8.855
R305 VDD.n220 VDD.n219 8.855
R306 VDD.n225 VDD.n224 8.855
R307 VDD.n224 VDD.n223 8.855
R308 VDD.n229 VDD.n228 8.855
R309 VDD.n228 VDD.n227 8.855
R310 VDD.n233 VDD.n232 8.855
R311 VDD.n145 VDD.n144 8.855
R312 VDD.n144 VDD.n143 8.855
R313 VDD.n150 VDD.n149 8.855
R314 VDD.n149 VDD.n148 8.855
R315 VDD.n154 VDD.n153 8.855
R316 VDD.n153 VDD.n152 8.855
R317 VDD.n158 VDD.n157 8.855
R318 VDD.n157 VDD.n156 8.855
R319 VDD.n162 VDD.n161 8.855
R320 VDD.n161 VDD.n160 8.855
R321 VDD.n166 VDD.n165 8.855
R322 VDD.n165 VDD.n164 8.855
R323 VDD.n171 VDD.n170 8.855
R324 VDD.n170 VDD.n169 8.855
R325 VDD.n174 VDD.n173 8.855
R326 VDD.n173 VDD.n172 8.855
R327 VDD.n178 VDD.n177 8.855
R328 VDD.n177 VDD.n176 8.855
R329 VDD.n182 VDD.n181 8.855
R330 VDD.n181 VDD.n180 8.855
R331 VDD.n186 VDD.n185 8.855
R332 VDD.n2 VDD.n1 8.855
R333 VDD.n6 VDD.n5 8.855
R334 VDD.n5 VDD.n4 8.855
R335 VDD.n11 VDD.n10 8.855
R336 VDD.n10 VDD.n9 8.855
R337 VDD.n15 VDD.n14 8.855
R338 VDD.n14 VDD.n13 8.855
R339 VDD.n19 VDD.n18 8.855
R340 VDD.n18 VDD.n17 8.855
R341 VDD.n25 VDD.n24 8.855
R342 VDD.n24 VDD.n23 8.855
R343 VDD.n28 VDD.n27 8.855
R344 VDD.n27 VDD.n26 8.855
R345 VDD.n32 VDD.n31 8.855
R346 VDD.n31 VDD.n30 8.855
R347 VDD.n36 VDD.n35 8.855
R348 VDD.n35 VDD.n34 8.855
R349 VDD.n40 VDD.n39 8.855
R350 VDD.n49 VDD.n48 8.855
R351 VDD.n54 VDD.n53 8.855
R352 VDD.n53 VDD.n52 8.855
R353 VDD.n58 VDD.n57 8.855
R354 VDD.n57 VDD.n56 8.855
R355 VDD.n62 VDD.n61 8.855
R356 VDD.n61 VDD.n60 8.855
R357 VDD.n66 VDD.n65 8.855
R358 VDD.n65 VDD.n64 8.855
R359 VDD.n71 VDD.n70 8.855
R360 VDD.n70 VDD.n69 8.855
R361 VDD.n74 VDD.n73 8.855
R362 VDD.n73 VDD.n72 8.855
R363 VDD.n78 VDD.n77 8.855
R364 VDD.n77 VDD.n76 8.855
R365 VDD.n82 VDD.n81 8.855
R366 VDD.n81 VDD.n80 8.855
R367 VDD.n87 VDD.n86 8.855
R368 VDD.n95 VDD.n94 8.855
R369 VDD.n99 VDD.n98 8.855
R370 VDD.n98 VDD.n97 8.855
R371 VDD.n104 VDD.n103 8.855
R372 VDD.n103 VDD.n102 8.855
R373 VDD.n108 VDD.n107 8.855
R374 VDD.n107 VDD.n106 8.855
R375 VDD.n112 VDD.n111 8.855
R376 VDD.n111 VDD.n110 8.855
R377 VDD.n116 VDD.n115 8.855
R378 VDD.n115 VDD.n114 8.855
R379 VDD.n121 VDD.n120 8.855
R380 VDD.n120 VDD.n119 8.855
R381 VDD.n125 VDD.n124 8.855
R382 VDD.n124 VDD.n123 8.855
R383 VDD.n129 VDD.n128 8.855
R384 VDD.n128 VDD.n127 8.855
R385 VDD.n133 VDD.n132 8.855
R386 VDD.n132 VDD.n131 8.855
R387 VDD.n137 VDD.n136 8.855
R388 VDD.n136 VDD.n135 8.855
R389 VDD.n321 VDD.n320 8.855
R390 VDD.n320 VDD.n319 8.855
R391 VDD.n317 VDD.n316 8.855
R392 VDD.n316 VDD.n315 8.855
R393 VDD.n313 VDD.n312 8.855
R394 VDD.n312 VDD.n311 8.855
R395 VDD.n308 VDD.n307 8.855
R396 VDD.n266 VDD.t29 6.195
R397 VDD.n303 VDD.n302 4.91
R398 VDD.n302 VDD.n301 4.65
R399 VDD.n243 VDD.n242 4.65
R400 VDD.n247 VDD.n246 4.65
R401 VDD.n252 VDD.n251 4.65
R402 VDD.n256 VDD.n255 4.65
R403 VDD.n260 VDD.n259 4.65
R404 VDD.n264 VDD.n263 4.65
R405 VDD.n269 VDD.n268 4.65
R406 VDD.n273 VDD.n272 4.65
R407 VDD.n277 VDD.n276 4.65
R408 VDD.n283 VDD.n280 4.65
R409 VDD.n287 VDD.n286 4.65
R410 VDD.n291 VDD.n290 4.65
R411 VDD.n295 VDD.n294 4.65
R412 VDD.n299 VDD.n298 4.65
R413 VDD.n239 VDD.n238 4.65
R414 VDD.n237 VDD.n236 4.65
R415 VDD.n196 VDD.n195 4.65
R416 VDD.n200 VDD.n199 4.65
R417 VDD.n205 VDD.n204 4.65
R418 VDD.n209 VDD.n208 4.65
R419 VDD.n213 VDD.n212 4.65
R420 VDD.n218 VDD.n215 4.65
R421 VDD.n222 VDD.n221 4.65
R422 VDD.n226 VDD.n225 4.65
R423 VDD.n230 VDD.n229 4.65
R424 VDD.n234 VDD.n233 4.65
R425 VDD.n192 VDD.n191 4.65
R426 VDD.n190 VDD.n189 4.65
R427 VDD.n146 VDD.n145 4.65
R428 VDD.n151 VDD.n150 4.65
R429 VDD.n155 VDD.n154 4.65
R430 VDD.n159 VDD.n158 4.65
R431 VDD.n163 VDD.n162 4.65
R432 VDD.n167 VDD.n166 4.65
R433 VDD.n171 VDD.n168 4.65
R434 VDD.n175 VDD.n174 4.65
R435 VDD.n179 VDD.n178 4.65
R436 VDD.n183 VDD.n182 4.65
R437 VDD.n187 VDD.n186 4.65
R438 VDD.n7 VDD.n6 4.65
R439 VDD.n12 VDD.n11 4.65
R440 VDD.n16 VDD.n15 4.65
R441 VDD.n20 VDD.n19 4.65
R442 VDD.n25 VDD.n22 4.65
R443 VDD.n29 VDD.n28 4.65
R444 VDD.n33 VDD.n32 4.65
R445 VDD.n37 VDD.n36 4.65
R446 VDD.n41 VDD.n40 4.65
R447 VDD.n44 VDD.n43 4.65
R448 VDD.n46 VDD.n45 4.65
R449 VDD.n50 VDD.n49 4.65
R450 VDD.n55 VDD.n54 4.65
R451 VDD.n59 VDD.n58 4.65
R452 VDD.n63 VDD.n62 4.65
R453 VDD.n67 VDD.n66 4.65
R454 VDD.n71 VDD.n68 4.65
R455 VDD.n75 VDD.n74 4.65
R456 VDD.n79 VDD.n78 4.65
R457 VDD.n83 VDD.n82 4.65
R458 VDD.n88 VDD.n87 4.65
R459 VDD.n90 VDD.n89 4.65
R460 VDD.n92 VDD.n91 4.65
R461 VDD.n96 VDD.n95 4.65
R462 VDD.n100 VDD.n99 4.65
R463 VDD.n105 VDD.n104 4.65
R464 VDD.n109 VDD.n108 4.65
R465 VDD.n113 VDD.n112 4.65
R466 VDD.n117 VDD.n116 4.65
R467 VDD.n122 VDD.n121 4.65
R468 VDD.n126 VDD.n125 4.65
R469 VDD.n130 VDD.n129 4.65
R470 VDD.n134 VDD.n133 4.65
R471 VDD.n138 VDD.n137 4.65
R472 VDD.n322 VDD.n321 4.65
R473 VDD.n318 VDD.n317 4.65
R474 VDD.n314 VDD.n313 4.65
R475 VDD.n309 VDD.n308 4.65
R476 VDD.n305 VDD.n304 4.65
R477 VDD.n1 VDD.n0 4.288
R478 VDD.n48 VDD.n47 4.288
R479 VDD.n94 VDD.n93 4.288
R480 VDD.n140 VDD.n139 4.288
R481 VDD.n194 VDD.n193 4.288
R482 VDD.n241 VDD.n240 4.288
R483 VDD.n297 VDD.n296 4.288
R484 VDD.n232 VDD.n231 4.288
R485 VDD.n185 VDD.n184 4.288
R486 VDD.n39 VDD.n38 4.288
R487 VDD.n86 VDD.n85 4.288
R488 VDD.n307 VDD.n306 4.288
R489 VDD.n3 VDD.n2 2.562
R490 VDD.n142 VDD.n141 2.562
R491 VDD.n279 VDD.n278 2.329
R492 VDD.n7 VDD.n3 1.145
R493 VDD.n146 VDD.n142 1.145
R494 VDD.n239 VDD.n237 0.597
R495 VDD.n192 VDD.n190 0.525
R496 VDD.n46 VDD.n44 0.525
R497 VDD.n92 VDD.n90 0.507
R498 VDD.n305 VDD.n303 0.135
R499 VDD.n155 VDD.n151 0.09
R500 VDD.n159 VDD.n155 0.09
R501 VDD.n163 VDD.n159 0.09
R502 VDD.n167 VDD.n163 0.09
R503 VDD.n168 VDD.n167 0.09
R504 VDD.n179 VDD.n175 0.09
R505 VDD.n183 VDD.n179 0.09
R506 VDD.n187 VDD.n183 0.09
R507 VDD.n196 VDD.n192 0.09
R508 VDD.n200 VDD.n196 0.09
R509 VDD.n209 VDD.n205 0.09
R510 VDD.n213 VDD.n209 0.09
R511 VDD.n215 VDD.n213 0.09
R512 VDD.n226 VDD.n222 0.09
R513 VDD.n230 VDD.n226 0.09
R514 VDD.n234 VDD.n230 0.09
R515 VDD.n243 VDD.n239 0.09
R516 VDD.n247 VDD.n243 0.09
R517 VDD.n256 VDD.n252 0.09
R518 VDD.n260 VDD.n256 0.09
R519 VDD.n264 VDD.n260 0.09
R520 VDD.n273 VDD.n269 0.09
R521 VDD.n277 VDD.n273 0.09
R522 VDD.n280 VDD.n277 0.09
R523 VDD.n291 VDD.n287 0.09
R524 VDD.n295 VDD.n291 0.09
R525 VDD.n299 VDD.n295 0.09
R526 VDD.n16 VDD.n12 0.09
R527 VDD.n20 VDD.n16 0.09
R528 VDD.n22 VDD.n20 0.09
R529 VDD.n33 VDD.n29 0.09
R530 VDD.n37 VDD.n33 0.09
R531 VDD.n41 VDD.n37 0.09
R532 VDD.n50 VDD.n46 0.09
R533 VDD.n59 VDD.n55 0.09
R534 VDD.n63 VDD.n59 0.09
R535 VDD.n67 VDD.n63 0.09
R536 VDD.n68 VDD.n67 0.09
R537 VDD.n79 VDD.n75 0.09
R538 VDD.n83 VDD.n79 0.09
R539 VDD.n90 VDD.n88 0.09
R540 VDD.n96 VDD.n92 0.09
R541 VDD.n100 VDD.n96 0.09
R542 VDD.n109 VDD.n105 0.09
R543 VDD.n113 VDD.n109 0.09
R544 VDD.n117 VDD.n113 0.09
R545 VDD.n126 VDD.n122 0.09
R546 VDD.n130 VDD.n126 0.09
R547 VDD.n134 VDD.n130 0.09
R548 VDD.n138 VDD.n134 0.09
R549 VDD.n322 VDD.n318 0.09
R550 VDD.n318 VDD.n314 0.09
R551 VDD.n309 VDD.n305 0.09
R552 VDD.n269 VDD.n265 0.086
R553 VDD.n201 VDD.n200 0.078
R554 VDD.n8 VDD.n7 0.078
R555 VDD.n101 VDD.n100 0.071
R556 VDD.n147 VDD.n146 0.07
R557 VDD.n175 CMOS_3in_OR_0/VDD 0.065
R558 VDD.n222 CMOS_AND_1/VDD 0.065
R559 VDD.n287 VDD 0.065
R560 VDD.n29 CMOS_AND_0/VDD 0.065
R561 VDD.n55 VDD.n51 0.065
R562 VDD.n75 CMOS_XOR_0/VDD 0.065
R563 VDD.n122 VDD.n118 0.065
R564 CMOS_XNOR_0/VDD VDD.n322 0.065
R565 VDD.n248 VDD.n247 0.063
R566 VDD.n190 VDD.n188 0.056
R567 VDD.n237 VDD.n235 0.056
R568 VDD.n302 VDD.n300 0.056
R569 VDD.n44 VDD.n42 0.056
R570 VDD.n84 VDD.n83 0.055
R571 VDD.n314 VDD.n310 0.055
R572 VDD.n88 VDD.n84 0.035
R573 VDD.n310 VDD.n309 0.035
R574 VDD.n188 VDD.n187 0.033
R575 VDD.n235 VDD.n234 0.033
R576 VDD.n300 VDD.n299 0.033
R577 VDD.n42 VDD.n41 0.033
R578 VDD.n303 VDD 0.027
R579 VDD.n252 VDD.n248 0.026
R580 VDD.n168 CMOS_3in_OR_0/VDD 0.025
R581 VDD.n51 VDD.n50 0.025
R582 VDD.n68 CMOS_XOR_0/VDD 0.025
R583 VDD.n118 VDD.n117 0.025
R584 CMOS_XNOR_0/VDD VDD.n138 0.025
R585 VDD.n151 VDD.n147 0.02
R586 VDD.n280 VDD.n279 0.018
R587 VDD.n105 VDD.n101 0.018
R588 VDD.n215 VDD.n214 0.017
R589 VDD.n22 VDD.n21 0.017
R590 VDD.n205 VDD.n201 0.011
R591 VDD.n12 VDD.n8 0.011
R592 VDD.n214 CMOS_AND_1/VDD 0.007
R593 VDD.n21 CMOS_AND_0/VDD 0.007
R594 VDD.n279 VDD 0.006
R595 VDD.n265 VDD.n264 0.003
R596 x0.t0 x0.t3 924.95
R597 CMOS_XOR_0/B x0.t0 633.02
R598 x0.n0 x0.t1 570.366
R599 x0.n0 x0.t2 570.366
R600 x0.n1 x0 425.672
R601 x0 x0.n0 78.72
R602 CMOS_XOR_0/B x0.n1 45.032
R603 x0.n1 x0 0.156
R604 x2_bar.n0 x2_bar.t1 683.32
R605 x2_bar.n1 x2_bar.t0 579.86
R606 x2_bar.n1 x2_bar.t3 547.727
R607 x2_bar.n0 x2_bar.t2 528.72
R608 CMOS_XNOR_0/B_bar x2_bar.n3 198.92
R609 x2_bar.n3 x2_bar.n2 19.691
R610 x2_bar.n2 x2_bar.n1 8.764
R611 CMOS_XNOR_0/B_bar x2_bar.n0 3.68
R612 x2_bar.n2 x2_bar 2.72
R613 x2_bar.n3 x2_bar 1.205
R614 x1_bar.t3 x1_bar.t2 1345.61
R615 x1_bar.n0 x1_bar.t1 579.86
R616 x1_bar.n0 x1_bar.t0 547.727
R617 CMOS_XOR_0/A_bar x1_bar.t3 392.02
R618 CMOS_XOR_0/A_bar x1_bar.n2 44.912
R619 x1_bar.n2 x1_bar.n1 12.665
R620 x1_bar.n1 x1_bar.n0 8.764
R621 x1_bar.n1 x1_bar 2.72
R622 x1_bar.n2 x1_bar 2.663
R623 x2.t2 x2.t3 1221.07
R624 x2.t0 x2.t1 924.95
R625 x2 x2.t2 633.02
R626 CMOS_XNOR_0/B x2.t0 633.02
R627 CMOS_XNOR_0/B x2.n0 389.96
R628 x2.n0 x2 232.934
R629 x2.n0 x2 0.154
R630 x3_bar.t0 x3_bar.t1 1345.61
R631 x3_bar.n0 x3_bar.t2 811.366
R632 CMOS_XNOR_0/A_bar x3_bar.t0 392.02
R633 x3_bar.n0 x3_bar.t3 329.366
R634 CMOS_XNOR_0/A_bar x3_bar.n1 286.14
R635 x3_bar.n1 x3_bar 265.317
R636 x3_bar x3_bar.n0 78.72
R637 x3_bar.n1 x3_bar 2.112
R638 x1.t2 x1.t0 1221.07
R639 x1.n0 x1.t3 993.097
R640 x1.n2 x1.t2 389.3
R641 x1.n0 x1.t1 356.59
R642 x1.n2 x1.n1 183.871
R643 x1.n1 x1.n0 8.764
R644 x1.n1 CMOS_XOR_0/A 2.72
R645 x1 x1.n2 2.72
R646 x3.n0 x3.t0 993.097
R647 x3.n0 x3.t1 356.59
R648 x3 x3.n0 78.72
R649 CMOS_4in_AND_0/OUT.t3 CMOS_4in_AND_0/OUT.t2 1221.07
R650 CMOS_3in_OR_0/C CMOS_4in_AND_0/OUT.n0 739.238
R651 CMOS_3in_OR_0/C CMOS_4in_AND_0/OUT.t3 633.02
R652 CMOS_4in_AND_0/OUT CMOS_4in_AND_0/OUT.t0 114.438
R653 CMOS_4in_AND_0/OUT.n0 CMOS_4in_AND_0/OUT 95.237
R654 CMOS_4in_AND_0/OUT.n0 CMOS_4in_AND_0/OUT.t1 45.156
R655 x0_bar.n0 x0_bar.t0 616.084
R656 x0_bar.n0 x0_bar.t1 528.72
R657 x0_bar.n0 x0_bar 16.711
R658 x0_bar x0_bar.n0 3.68
C0 a_2742_n1689# s2 0.00fF
C1 s2 a_2592_n1689# 0.00fF
C2 CMOS_AND_1/AND a_2742_n1689# 0.00fF
C3 CMOS_4in_AND_0/OUT a_2592_n1689# 0.01fF
C4 a_2742_n1689# CMOS_4in_AND_0/OUT 0.01fF
C5 CMOS_AND_1/AND a_2592_n1689# 0.01fF
C6 CMOS_AND_1/AND s2 0.01fF
C7 a_1380_n1689# a_2592_n1689# 0.00fF
C8 a_1380_n1689# a_2742_n1689# 0.00fF
C9 CMOS_4in_AND_0/OUT s2 0.00fF
C10 a_1380_n779# CMOS_AND_1/AND 0.00fF
C11 a_1380_n779# CMOS_4in_AND_0/OUT 0.01fF
C12 a_1380_n1689# s2 0.00fF
C13 a_1380_n779# a_n178_n1689# 0.00fF
C14 a_122_n779# CMOS_4in_AND_0/OUT 0.00fF
C15 a_1380_n779# a_1380_n1689# 0.01fF
C16 a_122_n779# a_n178_n1689# 0.01fF
C17 a_122_n779# a_1380_n1689# 0.00fF
C18 CMOS_4in_AND_0/OUT a_n28_n779# 0.00fF
C19 a_n178_n1689# a_n28_n779# 0.01fF
C20 a_n178_n779# CMOS_4in_AND_0/OUT 0.00fF
C21 a_1380_n1689# a_n28_n779# 0.00fF
C22 a_n178_n779# a_n178_n1689# 0.00fF
C23 a_2742_n1689# CMOS_AND_0/AND 0.00fF
C24 CMOS_AND_1/AND CMOS_4in_AND_0/OUT 0.10fF
C25 CMOS_AND_1/AND a_n178_n1689# 0.00fF
C26 CMOS_AND_0/AND a_2592_n1689# 0.00fF
C27 CMOS_4in_AND_0/OUT a_n178_n1689# 0.05fF
C28 a_1380_n1689# CMOS_AND_1/AND 0.07fF
C29 CMOS_AND_0/AND s2 0.04fF
C30 a_1380_n1689# CMOS_4in_AND_0/OUT 0.10fF
C31 a_1380_n1689# a_n178_n1689# 0.01fF
C32 a_2742_n1689# a_2592_499# 0.00fF
C33 a_2592_499# a_2592_n1689# 0.00fF
C34 CMOS_AND_0/A a_2592_n1689# 0.00fF
C35 a_1380_n779# CMOS_AND_1/A 0.01fF
C36 a_1435_n111# a_1380_n1689# 0.00fF
C37 a_1735_n111# a_1380_n1689# 0.00fF
C38 s2 x1_bar 0.00fF
C39 a_1380_n779# x1_bar 0.01fF
C40 a_1380_n779# x1 0.00fF
C41 a_122_n779# x1_bar 0.01fF
C42 a_1380_n779# x0_bar 0.00fF
C43 CMOS_AND_1/AND CMOS_AND_0/AND 0.04fF
C44 a_122_n779# x1 0.00fF
C45 a_122_n779# x0_bar 0.00fF
C46 a_177_n111# a_n178_n1689# 0.00fF
C47 CMOS_AND_0/AND CMOS_4in_AND_0/OUT 0.06fF
C48 a_n28_n779# x1_bar 0.01fF
C49 CMOS_AND_1/A CMOS_AND_1/AND 0.00fF
C50 a_1735_499# a_1380_n1689# 0.00fF
C51 a_122_n779# a_27_n111# 0.00fF
C52 a_1380_n1689# CMOS_AND_0/AND 0.00fF
C53 s2 x2_bar 0.00fF
C54 CMOS_AND_1/A CMOS_4in_AND_0/OUT 0.02fF
C55 x1 a_n28_n779# 0.00fF
C56 a_n178_n779# x1_bar 0.01fF
C57 a_n28_n779# x0_bar 0.00fF
C58 a_n178_n1689# a_n123_n111# 0.00fF
C59 CMOS_AND_1/A a_n178_n1689# 0.00fF
C60 x1 a_n178_n779# 0.00fF
C61 VDD a_2592_n1689# 0.06fF
C62 CMOS_4in_AND_0/OUT a_2592_499# 0.00fF
C63 VDD a_2742_n1689# 0.06fF
C64 a_177_499# a_n178_n1689# 0.00fF
C65 a_n178_n779# x0_bar 0.00fF
C66 a_1380_n1689# CMOS_AND_1/A 0.05fF
C67 a_n28_n779# a_27_n111# 0.00fF
C68 a_1380_n1689# a_1435_499# 0.00fF
C69 a_1380_n779# x2_bar 0.01fF
C70 CMOS_AND_0/A CMOS_4in_AND_0/OUT 0.00fF
C71 CMOS_AND_1/AND CMOS_AND_0/A 0.02fF
C72 a_2592_n111# CMOS_AND_0/AND 0.01fF
C73 a_122_n779# x3_bar 0.00fF
C74 a_122_n779# x2_bar 0.01fF
C75 a_1435_n111# CMOS_AND_0/AND 0.00fF
C76 a_1735_n111# CMOS_AND_0/AND 0.00fF
C77 a_122_n779# x0 0.00fF
C78 VDD s2 0.37fF
C79 a_1380_n1689# CMOS_AND_0/A 0.01fF
C80 a_122_n779# x3 0.00fF
C81 CMOS_4in_AND_0/OUT x1_bar 0.08fF
C82 CMOS_AND_1/AND x1_bar 0.01fF
C83 a_n28_n779# x3_bar 0.00fF
C84 a_122_n779# x2 0.00fF
C85 a_1380_n779# VDD 0.00fF
C86 x1 CMOS_4in_AND_0/OUT 0.03fF
C87 a_2592_n111# a_2592_499# 0.01fF
C88 x0 a_n28_n779# 0.00fF
C89 a_1435_n111# CMOS_AND_1/A 0.00fF
C90 CMOS_4in_AND_0/OUT x0_bar 0.00fF
C91 a_1735_n111# CMOS_AND_1/A 0.00fF
C92 x2_bar a_n28_n779# 0.01fF
C93 a_n178_n779# x3_bar 0.00fF
C94 a_n178_n1689# x1_bar 0.14fF
C95 x3 a_n28_n779# 0.00fF
C96 a_1735_n111# a_2592_499# 0.00fF
C97 a_n178_n779# x0 0.00fF
C98 a_n178_n779# x2_bar 0.01fF
C99 VDD a_122_n779# 0.01fF
C100 a_1435_n111# a_2592_499# 0.00fF
C101 a_1380_n1689# x1_bar 0.07fF
C102 a_1380_n1689# x1 0.01fF
C103 x1 a_n178_n1689# 0.10fF
C104 a_n178_n779# x3 0.00fF
C105 x2 a_n28_n779# 0.00fF
C106 a_n178_n1689# x0_bar 0.01fF
C107 a_2592_n111# CMOS_AND_0/A 0.01fF
C108 CMOS_4in_AND_0/OUT a_27_n111# 0.01fF
C109 a_1380_n1689# x0_bar 0.00fF
C110 a_n178_n779# x2 0.00fF
C111 a_1735_n111# CMOS_AND_0/A 0.01fF
C112 a_n178_n1689# a_27_n111# 0.01fF
C113 a_1435_n111# CMOS_AND_0/A 0.01fF
C114 VDD a_n28_n779# 0.01fF
C115 VDD a_n178_n779# 0.01fF
C116 a_1735_499# CMOS_AND_0/AND 0.00fF
C117 a_2592_n111# x0_bar 0.00fF
C118 CMOS_AND_1/AND x0 0.00fF
C119 CMOS_4in_AND_0/OUT x3_bar 0.00fF
C120 a_1435_n111# x1_bar 0.00fF
C121 a_1735_n111# x1_bar 0.01fF
C122 a_1735_n111# x1 0.00fF
C123 a_2592_n111# x1 0.00fF
C124 CMOS_AND_1/AND x2_bar 0.03fF
C125 a_1435_n111# x0_bar 0.01fF
C126 CMOS_4in_AND_0/OUT x0 0.00fF
C127 a_1735_n111# x0_bar 0.00fF
C128 a_n178_n1689# x3_bar 0.14fF
C129 a_1435_n111# x1 0.00fF
C130 CMOS_4in_AND_0/OUT x2_bar 0.02fF
C131 CMOS_4in_AND_0/OUT x3 0.00fF
C132 x0 a_n178_n1689# 0.07fF
C133 CMOS_AND_1/A a_177_n111# 0.00fF
C134 a_1380_n1689# x3_bar 0.00fF
C135 x2_bar a_n178_n1689# 0.04fF
C136 a_1380_n1689# x0 0.02fF
C137 a_1735_499# CMOS_AND_1/A 0.00fF
C138 CMOS_AND_0/AND a_1435_499# 0.00fF
C139 CMOS_4in_AND_0/OUT x2 0.00fF
C140 a_1380_n1689# x2_bar 0.03fF
C141 CMOS_AND_1/A CMOS_AND_0/AND 0.01fF
C142 a_1435_n111# a_27_n111# 0.00fF
C143 x3 a_n178_n1689# 0.01fF
C144 CMOS_AND_0/AND a_2592_499# 0.08fF
C145 x2 a_n178_n1689# 0.03fF
C146 CMOS_AND_1/A a_n123_n111# 0.00fF
C147 a_1735_499# a_2592_499# 0.00fF
C148 VDD CMOS_AND_1/AND 0.53fF
C149 a_177_n111# CMOS_AND_0/A 0.00fF
C150 a_1380_n1689# x2 0.00fF
C151 VDD CMOS_4in_AND_0/OUT 2.11fF
C152 a_1735_499# CMOS_AND_0/A 0.03fF
C153 a_177_499# CMOS_AND_1/A 0.00fF
C154 CMOS_AND_1/A a_1435_499# 0.01fF
C155 VDD a_n178_n1689# 1.61fF
C156 CMOS_AND_0/A CMOS_AND_0/AND 0.04fF
C157 CMOS_AND_1/A a_n123_499# 0.00fF
C158 a_2592_n111# x2_bar 0.01fF
C159 VDD a_1380_n1689# 0.75fF
C160 a_1435_499# a_2592_499# 0.00fF
C161 a_1435_n111# x2_bar 0.01fF
C162 a_177_n111# x1_bar 0.01fF
C163 a_1735_n111# x2_bar 0.01fF
C164 a_1435_n111# x0 0.01fF
C165 a_1735_n111# x0 0.01fF
C166 a_177_n111# x1 0.00fF
C167 a_1735_499# x1_bar 0.01fF
C168 CMOS_AND_0/A a_1435_499# 0.02fF
C169 CMOS_AND_1/A CMOS_AND_0/A 0.05fF
C170 CMOS_AND_0/A a_2592_499# 0.09fF
C171 a_177_499# CMOS_AND_0/A 0.00fF
C172 CMOS_AND_0/AND x1_bar 0.00fF
C173 a_177_n111# x0_bar 0.01fF
C174 CMOS_AND_0/AND x0_bar 0.00fF
C175 VDD a_2592_n111# 0.01fF
C176 x1_bar a_n123_n111# 0.01fF
C177 x1 CMOS_AND_0/AND 0.00fF
C178 a_1735_499# x0_bar 0.00fF
C179 a_n123_n111# x0_bar 0.01fF
C180 a_1735_n111# VDD 0.01fF
C181 a_177_n111# a_27_n111# 0.01fF
C182 x1 a_n123_n111# 0.00fF
C183 VDD a_1435_n111# 0.01fF
C184 a_177_499# x1_bar 0.00fF
C185 a_1435_499# x1_bar 0.00fF
C186 CMOS_AND_1/A x1_bar 0.09fF
C187 a_1435_499# x0_bar 0.01fF
C188 a_n123_499# x1_bar 0.00fF
C189 a_2592_499# x1_bar 0.00fF
C190 CMOS_AND_1/A x0_bar 0.06fF
C191 a_177_499# x1 0.00fF
C192 CMOS_AND_1/A x1 0.08fF
C193 a_177_499# x0_bar 0.01fF
C194 x1 a_n123_499# 0.00fF
C195 x1 a_2592_499# 0.00fF
C196 a_n123_499# x0_bar 0.01fF
C197 a_27_n111# a_n123_n111# 0.01fF
C198 a_2592_499# x0_bar 0.00fF
C199 CMOS_AND_1/A a_27_n111# 0.08fF
C200 a_177_n111# x3_bar 0.01fF
C201 a_177_499# a_27_n111# 0.03fF
C202 a_1435_499# a_27_n111# 0.00fF
C203 CMOS_AND_0/A x1_bar 0.14fF
C204 a_177_n111# x0 0.00fF
C205 a_n123_499# a_27_n111# 0.02fF
C206 CMOS_AND_0/A x0_bar 0.15fF
C207 a_177_n111# x2_bar 0.01fF
C208 x1 CMOS_AND_0/A 0.09fF
C209 a_177_n111# x3 0.00fF
C210 CMOS_AND_0/AND x2_bar 0.06fF
C211 a_1735_499# x0 0.03fF
C212 CMOS_AND_0/AND x0 0.00fF
C213 a_1735_499# x2_bar 0.00fF
C214 a_177_n111# x2 0.01fF
C215 x0 a_n123_n111# 0.00fF
C216 a_n123_n111# x3_bar 0.01fF
C217 x2_bar a_n123_n111# 0.01fF
C218 CMOS_AND_0/A a_27_n111# 0.04fF
C219 CMOS_AND_1/A x3_bar 0.01fF
C220 x1_bar x0_bar 0.42fF
C221 x3 a_n123_n111# 0.00fF
C222 x1 x1_bar 3.46fF
C223 x1 x0_bar 2.98fF
C224 CMOS_AND_1/A x2_bar 0.04fF
C225 a_n123_499# x3_bar 0.01fF
C226 a_177_499# x0 0.01fF
C227 a_1435_499# x0 0.01fF
C228 VDD a_177_n111# 0.01fF
C229 x2 a_n123_n111# 0.01fF
C230 a_177_499# x3_bar 0.01fF
C231 CMOS_AND_1/A x0 0.03fF
C232 a_177_499# x2_bar 0.01fF
C233 a_1435_499# x2_bar 0.00fF
C234 VDD CMOS_AND_0/AND 0.49fF
C235 x0 a_n123_499# 0.01fF
C236 a_2592_499# x0 0.01fF
C237 a_177_499# x3 0.00fF
C238 x2_bar a_n123_499# 0.01fF
C239 CMOS_AND_1/A x3 0.00fF
C240 VDD a_1735_499# 0.06fF
C241 x2_bar a_2592_499# 0.05fF
C242 a_27_n111# x1_bar 0.05fF
C243 CMOS_AND_1/A x2 0.01fF
C244 a_177_499# x2 0.03fF
C245 VDD a_n123_n111# 0.01fF
C246 x3 a_n123_499# 0.00fF
C247 x1 a_27_n111# 0.05fF
C248 CMOS_AND_0/A x3_bar 0.00fF
C249 x2 a_n123_499# 0.02fF
C250 CMOS_AND_0/A x2_bar 0.24fF
C251 a_27_n111# x0_bar 0.22fF
C252 CMOS_AND_0/A x0 0.35fF
C253 VDD CMOS_AND_1/A 0.51fF
C254 CMOS_AND_0/A x3 0.00fF
C255 VDD a_177_499# 0.05fF
C256 VDD a_1435_499# 0.06fF
C257 CMOS_AND_0/A x2 0.00fF
C258 VDD a_n123_499# 0.05fF
C259 VDD a_2592_499# 0.78fF
C260 x1_bar x3_bar 0.14fF
C261 x1 x3_bar 0.21fF
C262 x2_bar x1_bar 4.09fF
C263 VDD CMOS_AND_0/A 1.03fF
C264 x0_bar x3_bar 0.11fF
C265 x0 x1_bar 0.19fF
C266 x1 x2_bar 0.08fF
C267 x0 x0_bar 3.24fF
C268 x3 x1_bar 0.11fF
C269 x1 x3 0.03fF
C270 x1 x0 0.30fF
C271 x2_bar x0_bar 0.11fF
C272 x2 x1_bar 2.48fF
C273 x3 x0_bar 0.07fF
C274 a_27_n111# x3_bar 0.14fF
C275 x1 x2 0.05fF
C276 x0 a_27_n111# 0.15fF
C277 x2_bar a_27_n111# 0.18fF
C278 x2 x0_bar 0.11fF
C279 VDD x1_bar 1.04fF
C280 VDD x1 0.30fF
C281 x3 a_27_n111# 0.05fF
C282 x2 a_27_n111# 0.34fF
C283 VDD x0_bar 0.55fF
C284 x0 x3_bar 0.35fF
C285 VDD a_27_n111# 1.04fF
C286 x2_bar x3_bar 0.20fF
C287 x3 x3_bar 3.01fF
C288 x2_bar x0 0.14fF
C289 x3 x2_bar 2.83fF
C290 x2 x3_bar 0.15fF
C291 x3 x0 0.08fF
C292 x2 x0 0.25fF
C293 x2 x2_bar 3.04fF
C294 VDD x3_bar 0.38fF
C295 x2 x3 0.17fF
C296 VDD x0 1.57fF
C297 VDD x2_bar 0.81fF
C298 VDD x3 0.11fF
C299 VDD x2 1.39fF
C300 a_2442_n779# a_2742_n1689# 0.02fF
C301 a_2442_n779# a_2592_n1689# 0.02fF
C302 a_2442_n779# s2 0.06fF
C303 a_2442_n779# a_1380_n779# 0.00fF
C304 a_2442_n779# CMOS_AND_1/AND 0.10fF
C305 a_2442_n779# CMOS_4in_AND_0/OUT 0.05fF
C306 a_2442_n779# a_1380_n1689# 0.01fF
C307 a_2442_n779# a_2592_n111# 0.00fF
C308 a_2442_n779# CMOS_AND_0/AND 0.12fF
C309 a_2442_n779# CMOS_AND_1/A 0.00fF
C310 a_2442_n779# a_2592_499# 0.01fF
C311 a_2442_n779# CMOS_AND_0/A 0.01fF
C312 a_2442_n779# x1_bar 0.00fF
C313 a_2442_n779# x2_bar 0.02fF
C314 a_2442_n779# VDD 0.54fF
C315 a_2742_n1689# GND 0.02fF
C316 a_2592_n1689# GND 0.02fF
C317 s2 GND 0.55fF
C318 a_1380_n779# GND 0.03fF
C319 a_122_n779# GND 0.03fF
C320 a_n28_n779# GND 0.03fF
C321 a_n178_n779# GND 0.03fF
C322 a_2442_n779# GND 0.94fF
C323 CMOS_4in_AND_0/OUT GND 0.81fF $ **FLOATING
C324 CMOS_AND_1/AND GND 0.58fF
C325 a_1380_n1689# GND 0.49fF
C326 a_n178_n1689# GND 0.51fF
C327 a_2592_n111# GND 0.02fF
C328 a_1735_n111# GND 0.03fF
C329 a_1435_n111# GND 0.02fF
C330 a_177_n111# GND 0.02fF
C331 a_n123_n111# GND 0.02fF
C332 CMOS_AND_0/AND GND 1.97fF
C333 a_1735_499# GND 0.01fF
C334 a_1435_499# GND 0.01fF
C335 CMOS_AND_1/A GND 1.09fF
C336 a_177_499# GND 0.01fF
C337 a_n123_499# GND 0.01fF
C338 a_2592_499# GND 0.54fF
C339 CMOS_AND_0/A GND 1.15fF
C340 x1_bar GND 2.98fF
C341 x1 GND 8.02fF
C342 x0_bar GND 4.91fF
C343 a_27_n111# GND 0.63fF
C344 x3_bar GND 5.48fF
C345 x3 GND 5.76fF
C346 x2_bar GND 2.34fF
C347 x0 GND 2.59fF
C348 x2 GND 1.75fF
C349 VDD GND 24.99fF
C350 x0_bar.t1 GND 0.19fF
C351 x0_bar.t0 GND 0.18fF
C352 x0_bar.n0 GND 1.79fF $ **FLOATING
C353 CMOS_4in_AND_0/OUT.t2 GND 0.10fF
C354 CMOS_4in_AND_0/OUT.t3 GND 0.12fF
C355 CMOS_4in_AND_0/OUT.t1 GND 0.31fF
C356 CMOS_4in_AND_0/OUT.t0 GND 0.29fF
C357 CMOS_4in_AND_0/OUT.n0 GND 0.69fF $ **FLOATING
C358 CMOS_3in_OR_0/C GND 0.41fF $ **FLOATING
C359 x3.t0 GND 0.29fF
C360 x3.t1 GND 0.11fF
C361 x3.n0 GND 0.33fF $ **FLOATING
C362 x1.t3 GND 0.29fF
C363 x1.t1 GND 0.12fF
C364 x1.n0 GND 0.33fF $ **FLOATING
C365 CMOS_XOR_0/A GND 0.04fF $ **FLOATING
C366 x1.n1 GND 1.58fF $ **FLOATING
C367 x1.t0 GND 0.33fF
C368 x1.t2 GND 0.27fF
C369 x1.n2 GND 0.41fF $ **FLOATING
C370 x3_bar.t1 GND 0.33fF
C371 x3_bar.t0 GND 0.29fF
C372 x3_bar.t3 GND 0.10fF
C373 x3_bar.t2 GND 0.24fF
C374 x3_bar.n0 GND 0.25fF $ **FLOATING
C375 x3_bar.n1 GND 4.10fF $ **FLOATING
C376 CMOS_XNOR_0/A_bar GND 0.48fF $ **FLOATING
C377 x2.t1 GND 0.54fF
C378 x2.t0 GND 0.36fF
C379 x2.t3 GND 0.16fF
C380 x2.t2 GND 0.19fF
C381 x2.n0 GND 3.36fF $ **FLOATING
C382 CMOS_XNOR_0/B GND 0.42fF $ **FLOATING
C383 x1_bar.t2 GND 0.33fF
C384 x1_bar.t3 GND 0.29fF
C385 x1_bar.t1 GND 0.14fF
C386 x1_bar.t0 GND 0.21fF
C387 x1_bar.n0 GND 0.29fF $ **FLOATING
C388 x1_bar.n1 GND 0.92fF $ **FLOATING
C389 x1_bar.n2 GND 6.04fF $ **FLOATING
C390 CMOS_XOR_0/A_bar GND 0.55fF $ **FLOATING
C391 x2_bar.t2 GND 0.24fF
C392 x2_bar.t1 GND 0.24fF
C393 x2_bar.n0 GND 0.65fF $ **FLOATING
C394 x2_bar.t3 GND 0.21fF
C395 x2_bar.t0 GND 0.14fF
C396 x2_bar.n1 GND 0.29fF $ **FLOATING
C397 x2_bar.n2 GND 1.75fF $ **FLOATING
C398 x2_bar.n3 GND 5.49fF $ **FLOATING
C399 CMOS_XNOR_0/B_bar GND 0.23fF $ **FLOATING
C400 x0.t3 GND 0.43fF
C401 x0.t0 GND 0.29fF
C402 x0.t1 GND 0.08fF
C403 x0.t2 GND 0.12fF
C404 x0.n0 GND 0.14fF $ **FLOATING
C405 x0.n1 GND 3.69fF $ **FLOATING
C406 CMOS_XOR_0/B GND 0.33fF $ **FLOATING
C407 VDD.t28 GND 0.07fF
C408 VDD.t7 GND 0.07fF
C409 VDD.t22 GND 0.07fF
C410 CMOS_XOR_0/VDD GND 0.01fF $ **FLOATING
C411 VDD.t1 GND 0.07fF
C412 VDD.t38 GND 0.07fF
C413 CMOS_AND_0/VDD GND 0.01fF $ **FLOATING
C414 VDD.t40 GND 0.07fF
C415 VDD.n0 GND 0.20fF $ **FLOATING
C416 VDD.n1 GND 0.02fF $ **FLOATING
C417 VDD.n2 GND 0.01fF $ **FLOATING
C418 VDD.n3 GND 0.15fF $ **FLOATING
C419 VDD.t39 GND 0.10fF
C420 VDD.n4 GND 0.10fF $ **FLOATING
C421 VDD.n5 GND 0.02fF $ **FLOATING
C422 VDD.n6 GND 0.01fF $ **FLOATING
C423 VDD.n7 GND 0.05fF $ **FLOATING
C424 VDD.n8 GND 0.37fF $ **FLOATING
C425 VDD.n9 GND 0.17fF $ **FLOATING
C426 VDD.n10 GND 0.02fF $ **FLOATING
C427 VDD.n11 GND 0.01fF $ **FLOATING
C428 VDD.n12 GND 0.01fF $ **FLOATING
C429 VDD.n13 GND 0.17fF $ **FLOATING
C430 VDD.n14 GND 0.02fF $ **FLOATING
C431 VDD.n15 GND 0.01fF $ **FLOATING
C432 VDD.n16 GND 0.02fF $ **FLOATING
C433 VDD.n17 GND 0.17fF $ **FLOATING
C434 VDD.n18 GND 0.02fF $ **FLOATING
C435 VDD.n19 GND 0.01fF $ **FLOATING
C436 VDD.n20 GND 0.02fF $ **FLOATING
C437 VDD.t34 GND 0.07fF
C438 VDD.n21 GND 0.37fF $ **FLOATING
C439 VDD.n22 GND 0.01fF $ **FLOATING
C440 VDD.n23 GND 0.17fF $ **FLOATING
C441 VDD.n24 GND 0.02fF $ **FLOATING
C442 VDD.n25 GND 0.01fF $ **FLOATING
C443 VDD.t33 GND 0.09fF
C444 VDD.n26 GND 0.11fF $ **FLOATING
C445 VDD.n27 GND 0.02fF $ **FLOATING
C446 VDD.n28 GND 0.01fF $ **FLOATING
C447 VDD.n29 GND 0.02fF $ **FLOATING
C448 VDD.n30 GND 0.15fF $ **FLOATING
C449 VDD.n31 GND 0.02fF $ **FLOATING
C450 VDD.n32 GND 0.01fF $ **FLOATING
C451 VDD.n33 GND 0.02fF $ **FLOATING
C452 VDD.t37 GND 0.10fF
C453 VDD.n34 GND 0.11fF $ **FLOATING
C454 VDD.n35 GND 0.02fF $ **FLOATING
C455 VDD.n36 GND 0.01fF $ **FLOATING
C456 VDD.n37 GND 0.02fF $ **FLOATING
C457 VDD.n38 GND 0.19fF $ **FLOATING
C458 VDD.n39 GND 0.02fF $ **FLOATING
C459 VDD.n40 GND 0.01fF $ **FLOATING
C460 VDD.n41 GND 0.01fF $ **FLOATING
C461 VDD.n42 GND 0.37fF $ **FLOATING
C462 VDD.n43 GND 0.18fF $ **FLOATING
C463 VDD.n44 GND 0.06fF $ **FLOATING
C464 VDD.n45 GND 0.14fF $ **FLOATING
C465 VDD.n46 GND 0.06fF $ **FLOATING
C466 VDD.n47 GND 0.21fF $ **FLOATING
C467 VDD.n48 GND 0.02fF $ **FLOATING
C468 VDD.n49 GND 0.01fF $ **FLOATING
C469 VDD.n50 GND 0.01fF $ **FLOATING
C470 VDD.n51 GND 0.37fF $ **FLOATING
C471 VDD.t0 GND 0.09fF
C472 VDD.n52 GND 0.12fF $ **FLOATING
C473 VDD.n53 GND 0.02fF $ **FLOATING
C474 VDD.n54 GND 0.01fF $ **FLOATING
C475 VDD.n55 GND 0.02fF $ **FLOATING
C476 VDD.n56 GND 0.14fF $ **FLOATING
C477 VDD.n57 GND 0.02fF $ **FLOATING
C478 VDD.n58 GND 0.01fF $ **FLOATING
C479 VDD.n59 GND 0.02fF $ **FLOATING
C480 VDD.t23 GND 0.09fF
C481 VDD.n60 GND 0.12fF $ **FLOATING
C482 VDD.n61 GND 0.02fF $ **FLOATING
C483 VDD.n62 GND 0.01fF $ **FLOATING
C484 VDD.n63 GND 0.02fF $ **FLOATING
C485 VDD.n64 GND 0.14fF $ **FLOATING
C486 VDD.n65 GND 0.02fF $ **FLOATING
C487 VDD.n66 GND 0.01fF $ **FLOATING
C488 VDD.n67 GND 0.02fF $ **FLOATING
C489 VDD.n68 GND 0.01fF $ **FLOATING
C490 VDD.n69 GND 0.13fF $ **FLOATING
C491 VDD.n70 GND 0.02fF $ **FLOATING
C492 VDD.n71 GND 0.01fF $ **FLOATING
C493 VDD.t26 GND 0.09fF
C494 VDD.n72 GND 0.13fF $ **FLOATING
C495 VDD.n73 GND 0.02fF $ **FLOATING
C496 VDD.n74 GND 0.01fF $ **FLOATING
C497 VDD.n75 GND 0.02fF $ **FLOATING
C498 VDD.n76 GND 0.13fF $ **FLOATING
C499 VDD.n77 GND 0.02fF $ **FLOATING
C500 VDD.n78 GND 0.01fF $ **FLOATING
C501 VDD.n79 GND 0.02fF $ **FLOATING
C502 VDD.t21 GND 0.09fF
C503 VDD.n80 GND 0.13fF $ **FLOATING
C504 VDD.n81 GND 0.02fF $ **FLOATING
C505 VDD.n82 GND 0.01fF $ **FLOATING
C506 VDD.n83 GND 0.02fF $ **FLOATING
C507 VDD.n84 GND 0.37fF $ **FLOATING
C508 VDD.n85 GND 0.19fF $ **FLOATING
C509 VDD.n86 GND 0.02fF $ **FLOATING
C510 VDD.n87 GND 0.01fF $ **FLOATING
C511 VDD.n88 GND 0.01fF $ **FLOATING
C512 VDD.n89 GND 0.11fF $ **FLOATING
C513 VDD.n90 GND 0.06fF $ **FLOATING
C514 VDD.n91 GND 0.17fF $ **FLOATING
C515 VDD.n92 GND 0.06fF $ **FLOATING
C516 VDD.n93 GND 0.19fF $ **FLOATING
C517 VDD.n94 GND 0.02fF $ **FLOATING
C518 VDD.n95 GND 0.01fF $ **FLOATING
C519 VDD.n96 GND 0.02fF $ **FLOATING
C520 VDD.t6 GND 0.10fF
C521 VDD.n97 GND 0.11fF $ **FLOATING
C522 VDD.n98 GND 0.02fF $ **FLOATING
C523 VDD.n99 GND 0.01fF $ **FLOATING
C524 VDD.n100 GND 0.02fF $ **FLOATING
C525 VDD.n101 GND 0.37fF $ **FLOATING
C526 VDD.n102 GND 0.17fF $ **FLOATING
C527 VDD.n103 GND 0.02fF $ **FLOATING
C528 VDD.n104 GND 0.01fF $ **FLOATING
C529 VDD.n105 GND 0.01fF $ **FLOATING
C530 VDD.n106 GND 0.17fF $ **FLOATING
C531 VDD.n107 GND 0.02fF $ **FLOATING
C532 VDD.n108 GND 0.01fF $ **FLOATING
C533 VDD.n109 GND 0.02fF $ **FLOATING
C534 VDD.n110 GND 0.17fF $ **FLOATING
C535 VDD.n111 GND 0.02fF $ **FLOATING
C536 VDD.n112 GND 0.01fF $ **FLOATING
C537 VDD.n113 GND 0.02fF $ **FLOATING
C538 VDD.n114 GND 0.17fF $ **FLOATING
C539 VDD.n115 GND 0.02fF $ **FLOATING
C540 VDD.n116 GND 0.01fF $ **FLOATING
C541 VDD.n117 GND 0.01fF $ **FLOATING
C542 VDD.n118 GND 0.37fF $ **FLOATING
C543 VDD.t27 GND 0.09fF
C544 VDD.n119 GND 0.11fF $ **FLOATING
C545 VDD.n120 GND 0.02fF $ **FLOATING
C546 VDD.n121 GND 0.01fF $ **FLOATING
C547 VDD.n122 GND 0.02fF $ **FLOATING
C548 VDD.n123 GND 0.14fF $ **FLOATING
C549 VDD.n124 GND 0.02fF $ **FLOATING
C550 VDD.n125 GND 0.01fF $ **FLOATING
C551 VDD.n126 GND 0.02fF $ **FLOATING
C552 VDD.t31 GND 0.09fF
C553 VDD.n127 GND 0.12fF $ **FLOATING
C554 VDD.n128 GND 0.02fF $ **FLOATING
C555 VDD.n129 GND 0.01fF $ **FLOATING
C556 VDD.n130 GND 0.02fF $ **FLOATING
C557 VDD.n131 GND 0.14fF $ **FLOATING
C558 VDD.n132 GND 0.02fF $ **FLOATING
C559 VDD.n133 GND 0.01fF $ **FLOATING
C560 VDD.n134 GND 0.02fF $ **FLOATING
C561 VDD.t32 GND 0.09fF
C562 VDD.n135 GND 0.13fF $ **FLOATING
C563 VDD.n136 GND 0.02fF $ **FLOATING
C564 VDD.n137 GND 0.01fF $ **FLOATING
C565 VDD.n138 GND 0.01fF $ **FLOATING
C566 VDD.t36 GND 0.07fF
C567 VDD.t20 GND 0.07fF
C568 VDD.t30 GND 0.07fF
C569 VDD.t9 GND 0.07fF
C570 VDD.t17 GND 0.07fF
C571 CMOS_AND_1/VDD GND 0.01fF $ **FLOATING
C572 VDD.t15 GND 0.07fF
C573 VDD.t3 GND 0.07fF
C574 CMOS_3in_OR_0/VDD GND 0.01fF $ **FLOATING
C575 VDD.t5 GND 0.07fF
C576 VDD.n139 GND 0.20fF $ **FLOATING
C577 VDD.n140 GND 0.02fF $ **FLOATING
C578 VDD.n141 GND 0.01fF $ **FLOATING
C579 VDD.n142 GND 0.16fF $ **FLOATING
C580 VDD.t4 GND 0.10fF
C581 VDD.n143 GND 0.11fF $ **FLOATING
C582 VDD.n144 GND 0.02fF $ **FLOATING
C583 VDD.n145 GND 0.01fF $ **FLOATING
C584 VDD.n146 GND 0.05fF $ **FLOATING
C585 VDD.n147 GND 0.37fF $ **FLOATING
C586 VDD.n148 GND 0.17fF $ **FLOATING
C587 VDD.n149 GND 0.02fF $ **FLOATING
C588 VDD.n150 GND 0.01fF $ **FLOATING
C589 VDD.n151 GND 0.01fF $ **FLOATING
C590 VDD.n152 GND 0.17fF $ **FLOATING
C591 VDD.n153 GND 0.02fF $ **FLOATING
C592 VDD.n154 GND 0.01fF $ **FLOATING
C593 VDD.n155 GND 0.02fF $ **FLOATING
C594 VDD.n156 GND 0.17fF $ **FLOATING
C595 VDD.n157 GND 0.02fF $ **FLOATING
C596 VDD.n158 GND 0.01fF $ **FLOATING
C597 VDD.n159 GND 0.02fF $ **FLOATING
C598 VDD.n160 GND 0.17fF $ **FLOATING
C599 VDD.n161 GND 0.02fF $ **FLOATING
C600 VDD.n162 GND 0.01fF $ **FLOATING
C601 VDD.n163 GND 0.02fF $ **FLOATING
C602 VDD.t18 GND 0.09fF
C603 VDD.n164 GND 0.10fF $ **FLOATING
C604 VDD.n165 GND 0.02fF $ **FLOATING
C605 VDD.n166 GND 0.01fF $ **FLOATING
C606 VDD.n167 GND 0.02fF $ **FLOATING
C607 VDD.n168 GND 0.01fF $ **FLOATING
C608 VDD.n169 GND 0.16fF $ **FLOATING
C609 VDD.n170 GND 0.02fF $ **FLOATING
C610 VDD.n171 GND 0.01fF $ **FLOATING
C611 VDD.t41 GND 0.09fF
C612 VDD.n172 GND 0.11fF $ **FLOATING
C613 VDD.n173 GND 0.02fF $ **FLOATING
C614 VDD.n174 GND 0.01fF $ **FLOATING
C615 VDD.n175 GND 0.02fF $ **FLOATING
C616 VDD.n176 GND 0.15fF $ **FLOATING
C617 VDD.n177 GND 0.02fF $ **FLOATING
C618 VDD.n178 GND 0.01fF $ **FLOATING
C619 VDD.n179 GND 0.02fF $ **FLOATING
C620 VDD.t2 GND 0.10fF
C621 VDD.n180 GND 0.11fF $ **FLOATING
C622 VDD.n181 GND 0.02fF $ **FLOATING
C623 VDD.n182 GND 0.01fF $ **FLOATING
C624 VDD.n183 GND 0.02fF $ **FLOATING
C625 VDD.n184 GND 0.19fF $ **FLOATING
C626 VDD.n185 GND 0.02fF $ **FLOATING
C627 VDD.n186 GND 0.01fF $ **FLOATING
C628 VDD.n187 GND 0.01fF $ **FLOATING
C629 VDD.n188 GND 0.37fF $ **FLOATING
C630 VDD.n189 GND 0.18fF $ **FLOATING
C631 VDD.n190 GND 0.06fF $ **FLOATING
C632 VDD.n191 GND 0.16fF $ **FLOATING
C633 VDD.n192 GND 0.06fF $ **FLOATING
C634 VDD.n193 GND 0.19fF $ **FLOATING
C635 VDD.n194 GND 0.02fF $ **FLOATING
C636 VDD.n195 GND 0.01fF $ **FLOATING
C637 VDD.n196 GND 0.02fF $ **FLOATING
C638 VDD.t14 GND 0.10fF
C639 VDD.n197 GND 0.10fF $ **FLOATING
C640 VDD.n198 GND 0.02fF $ **FLOATING
C641 VDD.n199 GND 0.01fF $ **FLOATING
C642 VDD.n200 GND 0.02fF $ **FLOATING
C643 VDD.n201 GND 0.37fF $ **FLOATING
C644 VDD.n202 GND 0.17fF $ **FLOATING
C645 VDD.n203 GND 0.02fF $ **FLOATING
C646 VDD.n204 GND 0.01fF $ **FLOATING
C647 VDD.n205 GND 0.01fF $ **FLOATING
C648 VDD.n206 GND 0.17fF $ **FLOATING
C649 VDD.n207 GND 0.02fF $ **FLOATING
C650 VDD.n208 GND 0.01fF $ **FLOATING
C651 VDD.n209 GND 0.02fF $ **FLOATING
C652 VDD.n210 GND 0.17fF $ **FLOATING
C653 VDD.n211 GND 0.02fF $ **FLOATING
C654 VDD.n212 GND 0.01fF $ **FLOATING
C655 VDD.n213 GND 0.02fF $ **FLOATING
C656 VDD.t11 GND 0.07fF
C657 VDD.n214 GND 0.37fF $ **FLOATING
C658 VDD.n215 GND 0.01fF $ **FLOATING
C659 VDD.n216 GND 0.17fF $ **FLOATING
C660 VDD.n217 GND 0.02fF $ **FLOATING
C661 VDD.n218 GND 0.01fF $ **FLOATING
C662 VDD.t10 GND 0.09fF
C663 VDD.n219 GND 0.11fF $ **FLOATING
C664 VDD.n220 GND 0.02fF $ **FLOATING
C665 VDD.n221 GND 0.01fF $ **FLOATING
C666 VDD.n222 GND 0.02fF $ **FLOATING
C667 VDD.n223 GND 0.15fF $ **FLOATING
C668 VDD.n224 GND 0.02fF $ **FLOATING
C669 VDD.n225 GND 0.01fF $ **FLOATING
C670 VDD.n226 GND 0.02fF $ **FLOATING
C671 VDD.t16 GND 0.10fF
C672 VDD.n227 GND 0.11fF $ **FLOATING
C673 VDD.n228 GND 0.02fF $ **FLOATING
C674 VDD.n229 GND 0.01fF $ **FLOATING
C675 VDD.n230 GND 0.02fF $ **FLOATING
C676 VDD.n231 GND 0.19fF $ **FLOATING
C677 VDD.n232 GND 0.02fF $ **FLOATING
C678 VDD.n233 GND 0.01fF $ **FLOATING
C679 VDD.n234 GND 0.01fF $ **FLOATING
C680 VDD.n235 GND 0.37fF $ **FLOATING
C681 VDD.n236 GND 0.18fF $ **FLOATING
C682 VDD.n237 GND 0.07fF $ **FLOATING
C683 VDD.n238 GND 0.18fF $ **FLOATING
C684 VDD.n239 GND 0.07fF $ **FLOATING
C685 VDD.n240 GND 0.19fF $ **FLOATING
C686 VDD.n241 GND 0.02fF $ **FLOATING
C687 VDD.n242 GND 0.01fF $ **FLOATING
C688 VDD.n243 GND 0.02fF $ **FLOATING
C689 VDD.t8 GND 0.10fF
C690 VDD.n244 GND 0.11fF $ **FLOATING
C691 VDD.n245 GND 0.02fF $ **FLOATING
C692 VDD.n246 GND 0.01fF $ **FLOATING
C693 VDD.n247 GND 0.02fF $ **FLOATING
C694 VDD.n248 GND 0.37fF $ **FLOATING
C695 VDD.n249 GND 0.17fF $ **FLOATING
C696 VDD.n250 GND 0.02fF $ **FLOATING
C697 VDD.n251 GND 0.01fF $ **FLOATING
C698 VDD.n252 GND 0.01fF $ **FLOATING
C699 VDD.n253 GND 0.17fF $ **FLOATING
C700 VDD.n254 GND 0.02fF $ **FLOATING
C701 VDD.n255 GND 0.01fF $ **FLOATING
C702 VDD.n256 GND 0.02fF $ **FLOATING
C703 VDD.n257 GND 0.17fF $ **FLOATING
C704 VDD.n258 GND 0.02fF $ **FLOATING
C705 VDD.n259 GND 0.01fF $ **FLOATING
C706 VDD.n260 GND 0.02fF $ **FLOATING
C707 VDD.n261 GND 0.17fF $ **FLOATING
C708 VDD.n262 GND 0.02fF $ **FLOATING
C709 VDD.n263 GND 0.01fF $ **FLOATING
C710 VDD.n264 GND 0.01fF $ **FLOATING
C711 VDD.n265 GND 0.37fF $ **FLOATING
C712 VDD.t29 GND 0.09fF
C713 VDD.n266 GND 0.09fF $ **FLOATING
C714 VDD.n267 GND 0.02fF $ **FLOATING
C715 VDD.n268 GND 0.01fF $ **FLOATING
C716 VDD.n269 GND 0.02fF $ **FLOATING
C717 VDD.n270 GND 0.16fF $ **FLOATING
C718 VDD.n271 GND 0.02fF $ **FLOATING
C719 VDD.n272 GND 0.01fF $ **FLOATING
C720 VDD.n273 GND 0.02fF $ **FLOATING
C721 VDD.t24 GND 0.09fF
C722 VDD.n274 GND 0.10fF $ **FLOATING
C723 VDD.n275 GND 0.02fF $ **FLOATING
C724 VDD.n276 GND 0.01fF $ **FLOATING
C725 VDD.n277 GND 0.02fF $ **FLOATING
C726 VDD.t25 GND 0.05fF
C727 VDD.t13 GND 0.05fF
C728 VDD.n278 GND 0.19fF $ **FLOATING
C729 VDD.n279 GND 0.15fF $ **FLOATING
C730 VDD.n280 GND 0.01fF $ **FLOATING
C731 VDD.n281 GND 0.16fF $ **FLOATING
C732 VDD.n282 GND 0.02fF $ **FLOATING
C733 VDD.n283 GND 0.01fF $ **FLOATING
C734 VDD.t12 GND 0.09fF
C735 VDD.n284 GND 0.11fF $ **FLOATING
C736 VDD.n285 GND 0.02fF $ **FLOATING
C737 VDD.n286 GND 0.01fF $ **FLOATING
C738 VDD.n287 GND 0.02fF $ **FLOATING
C739 VDD.n288 GND 0.15fF $ **FLOATING
C740 VDD.n289 GND 0.02fF $ **FLOATING
C741 VDD.n290 GND 0.01fF $ **FLOATING
C742 VDD.n291 GND 0.02fF $ **FLOATING
C743 VDD.t19 GND 0.10fF
C744 VDD.n292 GND 0.11fF $ **FLOATING
C745 VDD.n293 GND 0.02fF $ **FLOATING
C746 VDD.n294 GND 0.01fF $ **FLOATING
C747 VDD.n295 GND 0.02fF $ **FLOATING
C748 VDD.n296 GND 0.19fF $ **FLOATING
C749 VDD.n297 GND 0.02fF $ **FLOATING
C750 VDD.n298 GND 0.01fF $ **FLOATING
C751 VDD.n299 GND 0.01fF $ **FLOATING
C752 VDD.n300 GND 0.37fF $ **FLOATING
C753 VDD.n301 GND 0.18fF $ **FLOATING
C754 VDD.n302 GND 0.35fF $ **FLOATING
C755 VDD.n303 GND 0.34fF $ **FLOATING
C756 VDD.n304 GND 0.11fF $ **FLOATING
C757 VDD.n305 GND 0.02fF $ **FLOATING
C758 VDD.n306 GND 0.19fF $ **FLOATING
C759 VDD.n307 GND 0.02fF $ **FLOATING
C760 VDD.n308 GND 0.01fF $ **FLOATING
C761 VDD.n309 GND 0.01fF $ **FLOATING
C762 VDD.n310 GND 0.37fF $ **FLOATING
C763 VDD.t35 GND 0.09fF
C764 VDD.n311 GND 0.13fF $ **FLOATING
C765 VDD.n312 GND 0.02fF $ **FLOATING
C766 VDD.n313 GND 0.01fF $ **FLOATING
C767 VDD.n314 GND 0.02fF $ **FLOATING
C768 VDD.n315 GND 0.13fF $ **FLOATING
C769 VDD.n316 GND 0.02fF $ **FLOATING
C770 VDD.n317 GND 0.01fF $ **FLOATING
C771 VDD.n318 GND 0.02fF $ **FLOATING
C772 VDD.n319 GND 0.13fF $ **FLOATING
C773 VDD.n320 GND 0.02fF $ **FLOATING
C774 VDD.n321 GND 0.01fF $ **FLOATING
C775 VDD.n322 GND 0.02fF $ **FLOATING
C776 CMOS_XNOR_0/VDD GND 0.01fF $ **FLOATING
.ends

