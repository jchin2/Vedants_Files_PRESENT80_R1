magic
tech sky130A
timestamp 1670967604
<< metal4 >>
rect -2530 14810 15070 14910
rect -2530 -2290 -2430 14810
rect -2230 14510 14770 14610
rect -2230 -1990 -2130 14510
rect -1930 14210 14470 14310
rect -1930 -1690 -1830 14210
rect -1630 13910 14170 14010
rect -1630 -1390 -1530 13910
rect -1330 13610 13870 13710
rect -1330 -1090 -1230 13610
rect -1030 13310 13570 13410
rect -1030 -790 -930 13310
rect -730 13010 13270 13110
rect -730 -490 -630 13010
rect -430 12710 12970 12810
rect -430 -190 -330 12710
rect -130 12410 12670 12510
rect -130 110 -30 12410
rect -130 10 6170 110
rect 12570 -190 12670 12410
rect -430 -290 12670 -190
rect 12870 -490 12970 12710
rect -730 -590 12970 -490
rect 13170 -790 13270 13010
rect -1030 -890 13270 -790
rect 13470 -1090 13570 13310
rect -1330 -1190 13570 -1090
rect 13770 -1390 13870 13610
rect -1630 -1490 13870 -1390
rect 14070 -1690 14170 13910
rect -1930 -1790 14170 -1690
rect 14370 -1990 14470 14210
rect -2230 -2090 14470 -1990
rect 14670 -2290 14770 14510
rect -2530 -2390 14770 -2290
rect 14970 -2590 15070 14810
rect 6170 -2690 15070 -2590
<< properties >>
string path 144.700 -23.400 146.700 -23.400 
<< end >>
