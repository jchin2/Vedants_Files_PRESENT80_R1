magic
tech sky130A
magscale 1 2
timestamp 1677167050
<< locali >>
rect -1031 1258 -951 1281
rect -1031 1224 -1008 1258
rect -974 1224 -951 1258
rect -1031 1189 -951 1224
rect 1660 1189 1740 1205
rect -1031 1186 247 1189
rect -1031 1152 -1008 1186
rect -974 1152 247 1186
rect -1031 1149 247 1152
rect 1660 1182 1805 1189
rect -1031 1114 -951 1149
rect 1660 1148 1683 1182
rect 1717 1149 1805 1182
rect 1717 1148 1740 1149
rect 1660 1125 1740 1148
rect -1031 1080 -1008 1114
rect -974 1080 -951 1114
rect -1031 1057 -951 1080
rect -917 524 -837 547
rect -917 490 -894 524
rect -860 490 -837 524
rect -917 455 -837 490
rect -917 452 -233 455
rect -917 418 -894 452
rect -860 418 -233 452
rect -917 415 -233 418
rect -917 380 -837 415
rect 3212 408 3319 431
rect -917 346 -894 380
rect -860 346 -837 380
rect 2056 360 2136 383
rect -917 323 -837 346
rect -803 333 -723 356
rect -803 299 -780 333
rect -746 299 -723 333
rect 2056 326 2079 360
rect 2113 326 2136 360
rect 2056 303 2136 326
rect 3212 374 3262 408
rect 3296 374 3319 408
rect 3212 336 3319 374
rect -803 264 -723 299
rect -803 261 -203 264
rect -803 227 -780 261
rect -746 227 -203 261
rect -803 224 -203 227
rect -803 189 -723 224
rect -803 155 -780 189
rect -746 155 -723 189
rect -803 132 -723 155
rect -689 -92 -609 -69
rect 828 -91 958 -51
rect -689 -126 -666 -92
rect -632 -109 -609 -92
rect -632 -126 -421 -109
rect -689 -149 -421 -126
rect -689 -164 -609 -149
rect -689 -198 -666 -164
rect -632 -198 -609 -164
rect -461 -161 -421 -149
rect -689 -236 -609 -198
rect -689 -270 -666 -236
rect -632 -270 -609 -236
rect -689 -293 -609 -270
rect -575 -206 -495 -183
rect -461 -201 247 -161
rect -575 -240 -552 -206
rect -518 -240 -495 -206
rect -575 -255 -495 -240
rect -575 -278 -353 -255
rect -575 -312 -552 -278
rect -518 -312 -353 -278
rect -575 -335 -353 -312
rect -1259 -372 -1179 -349
rect -1259 -406 -1236 -372
rect -1202 -406 -1179 -372
rect -1259 -441 -1179 -406
rect -575 -350 -495 -335
rect -575 -384 -552 -350
rect -518 -384 -495 -350
rect -575 -407 -495 -384
rect 556 -391 636 -373
rect -461 -431 42 -391
rect 122 -396 636 -391
rect 122 -430 579 -396
rect 613 -430 636 -396
rect 918 -389 958 -91
rect 1660 -160 1740 -137
rect 1660 -194 1683 -160
rect 1717 -161 1740 -160
rect 2077 -161 2117 303
rect 3212 302 3262 336
rect 3296 302 3319 336
rect 3212 279 3319 302
rect 1717 -194 1805 -161
rect 1660 -201 1805 -194
rect 2077 -201 2662 -161
rect 1660 -217 1740 -201
rect 918 -429 1450 -389
rect 3239 -393 3319 -373
rect 2742 -396 3319 -393
rect 122 -431 636 -430
rect -461 -441 -421 -431
rect -1259 -444 -421 -441
rect -1259 -478 -1236 -444
rect -1202 -478 -421 -444
rect 556 -453 636 -431
rect 2742 -430 3262 -396
rect 3296 -430 3319 -396
rect 2742 -433 3319 -430
rect 3239 -453 3319 -433
rect -1259 -481 -421 -478
rect -1259 -516 -1179 -481
rect -1259 -550 -1236 -516
rect -1202 -550 -1179 -516
rect -1259 -573 -1179 -550
rect -689 -754 -609 -731
rect -689 -788 -666 -754
rect -632 -788 -609 -754
rect -689 -826 -609 -788
rect -689 -860 -666 -826
rect -632 -839 -609 -826
rect -632 -860 192 -839
rect -689 -879 192 -860
rect -1487 -920 -1407 -897
rect -1487 -954 -1464 -920
rect -1430 -954 -1407 -920
rect -1487 -989 -1407 -954
rect -689 -898 -609 -879
rect -689 -932 -666 -898
rect -632 -932 -609 -898
rect -689 -955 -609 -932
rect 3303 -883 3383 -860
rect 3303 -917 3326 -883
rect 3360 -917 3383 -883
rect 3303 -955 3383 -917
rect 3303 -989 3326 -955
rect 3360 -989 3383 -955
rect -1487 -992 -108 -989
rect -1487 -1026 -1464 -992
rect -1430 -1026 -108 -992
rect -1487 -1029 -108 -1026
rect -1487 -1064 -1407 -1029
rect 2000 -1029 2512 -989
rect 3303 -1012 3383 -989
rect -1487 -1098 -1464 -1064
rect -1430 -1098 -1407 -1064
rect -1487 -1121 -1407 -1098
rect -1031 -1670 -951 -1647
rect -1031 -1704 -1008 -1670
rect -974 -1704 -951 -1670
rect -1031 -1739 -951 -1704
rect 702 -1739 742 -1669
rect -1031 -1742 -258 -1739
rect -1031 -1776 -1008 -1742
rect -974 -1776 -258 -1742
rect -1031 -1779 -258 -1776
rect 702 -1779 2832 -1739
rect -1031 -1814 -951 -1779
rect -1031 -1848 -1008 -1814
rect -974 -1848 -951 -1814
rect -1031 -1871 -951 -1848
<< viali >>
rect -1008 1224 -974 1258
rect -1008 1152 -974 1186
rect 1683 1148 1717 1182
rect -1008 1080 -974 1114
rect -894 490 -860 524
rect -894 418 -860 452
rect 1348 418 1382 452
rect 2505 412 2539 446
rect -894 346 -860 380
rect -780 299 -746 333
rect 2079 326 2113 360
rect 3262 374 3296 408
rect -780 227 -746 261
rect 1378 227 1412 261
rect -780 155 -746 189
rect -666 -126 -632 -92
rect -666 -198 -632 -164
rect -666 -270 -632 -236
rect -552 -240 -518 -206
rect -552 -312 -518 -278
rect -1236 -406 -1202 -372
rect -552 -384 -518 -350
rect 579 -430 613 -396
rect 1683 -194 1717 -160
rect 3262 302 3296 336
rect -1236 -478 -1202 -444
rect 3262 -430 3296 -396
rect -1236 -550 -1202 -516
rect -666 -788 -632 -754
rect -666 -860 -632 -826
rect -1464 -954 -1430 -920
rect -666 -932 -632 -898
rect 3326 -917 3360 -883
rect 3326 -989 3360 -955
rect -1464 -1026 -1430 -992
rect 1293 -1036 1327 -1002
rect -1464 -1098 -1430 -1064
rect -1008 -1704 -974 -1670
rect -1008 -1776 -974 -1742
rect -1008 -1848 -974 -1814
<< metal1 >>
rect -1487 1259 -1407 1333
rect -1487 1207 -1473 1259
rect -1421 1207 -1407 1259
rect -1487 1191 -1407 1207
rect -1487 1139 -1473 1191
rect -1421 1139 -1407 1191
rect -1487 1123 -1407 1139
rect -1487 1071 -1473 1123
rect -1421 1071 -1407 1123
rect -1487 -920 -1407 1071
rect -1487 -954 -1464 -920
rect -1430 -954 -1407 -920
rect -1487 -992 -1407 -954
rect -1487 -1026 -1464 -992
rect -1430 -1026 -1407 -992
rect -1487 -1064 -1407 -1026
rect -1487 -1098 -1464 -1064
rect -1430 -1098 -1407 -1064
rect -1487 -1924 -1407 -1098
rect -1373 -1924 -1293 1333
rect -1259 -372 -1179 1333
rect -1259 -406 -1236 -372
rect -1202 -406 -1179 -372
rect -1259 -444 -1179 -406
rect -1259 -478 -1236 -444
rect -1202 -478 -1179 -444
rect -1259 -516 -1179 -478
rect -1259 -550 -1236 -516
rect -1202 -550 -1179 -516
rect -1259 -1924 -1179 -550
rect -1145 -407 -1065 1333
rect -1145 -459 -1131 -407
rect -1079 -459 -1065 -407
rect -1145 -475 -1065 -459
rect -1145 -527 -1131 -475
rect -1079 -527 -1065 -475
rect -1145 -543 -1065 -527
rect -1145 -595 -1131 -543
rect -1079 -595 -1065 -543
rect -1145 -926 -1065 -595
rect -1145 -978 -1131 -926
rect -1079 -978 -1065 -926
rect -1145 -994 -1065 -978
rect -1145 -1046 -1131 -994
rect -1079 -1046 -1065 -994
rect -1145 -1062 -1065 -1046
rect -1145 -1114 -1131 -1062
rect -1079 -1114 -1065 -1062
rect -1145 -1924 -1065 -1114
rect -1031 1258 -951 1333
rect -1031 1224 -1008 1258
rect -974 1224 -951 1258
rect -1031 1186 -951 1224
rect -1031 1152 -1008 1186
rect -974 1152 -951 1186
rect -1031 1114 -951 1152
rect -1031 1080 -1008 1114
rect -974 1080 -951 1114
rect -1031 -563 -951 1080
rect -1031 -615 -1017 -563
rect -965 -615 -951 -563
rect -1031 -631 -951 -615
rect -1031 -683 -1017 -631
rect -965 -683 -951 -631
rect -1031 -699 -951 -683
rect -1031 -751 -1017 -699
rect -965 -751 -951 -699
rect -1031 -1670 -951 -751
rect -1031 -1704 -1008 -1670
rect -974 -1704 -951 -1670
rect -1031 -1742 -951 -1704
rect -1031 -1776 -1008 -1742
rect -974 -1776 -951 -1742
rect -1031 -1814 -951 -1776
rect -1031 -1848 -1008 -1814
rect -974 -1848 -951 -1814
rect -1031 -1923 -951 -1848
rect -917 524 -837 1333
rect -917 490 -894 524
rect -860 490 -837 524
rect -917 452 -837 490
rect -917 418 -894 452
rect -860 418 -837 452
rect -917 380 -837 418
rect -917 346 -894 380
rect -860 346 -837 380
rect -917 -87 -837 346
rect -917 -139 -903 -87
rect -851 -139 -837 -87
rect -917 -155 -837 -139
rect -917 -207 -903 -155
rect -851 -207 -837 -155
rect -917 -223 -837 -207
rect -917 -275 -903 -223
rect -851 -275 -837 -223
rect -917 -1924 -837 -275
rect -803 333 -723 1333
rect -803 299 -780 333
rect -746 299 -723 333
rect -803 261 -723 299
rect -803 227 -780 261
rect -746 227 -723 261
rect -803 189 -723 227
rect -803 155 -780 189
rect -746 155 -723 189
rect -803 -1923 -723 155
rect -689 -92 -609 1333
rect -689 -126 -666 -92
rect -632 -126 -609 -92
rect -689 -164 -609 -126
rect -689 -198 -666 -164
rect -632 -198 -609 -164
rect -689 -236 -609 -198
rect -689 -270 -666 -236
rect -632 -270 -609 -236
rect -689 -754 -609 -270
rect -689 -788 -666 -754
rect -632 -788 -609 -754
rect -689 -826 -609 -788
rect -689 -860 -666 -826
rect -632 -860 -609 -826
rect -689 -898 -609 -860
rect -689 -932 -666 -898
rect -632 -932 -609 -898
rect -689 -1923 -609 -932
rect -575 -206 -495 1333
rect -575 -240 -552 -206
rect -518 -240 -495 -206
rect -575 -278 -495 -240
rect -575 -312 -552 -278
rect -518 -312 -495 -278
rect -575 -350 -495 -312
rect -575 -384 -552 -350
rect -518 -384 -495 -350
rect -575 -1923 -495 -384
rect -461 1233 -353 1333
rect 873 1233 1205 1333
rect 2121 1233 2417 1333
rect -461 -1823 -381 1233
rect 1660 1191 1740 1205
rect 1660 1139 1674 1191
rect 1726 1139 1740 1191
rect 1660 1125 1740 1139
rect 1325 461 1405 475
rect 1325 409 1339 461
rect 1391 409 1405 461
rect 1325 395 1405 409
rect 2482 455 2562 469
rect 2482 403 2496 455
rect 2548 403 2562 455
rect 2482 389 2562 403
rect 3239 417 3319 431
rect 2056 369 2136 383
rect 2056 317 2070 369
rect 2122 317 2136 369
rect 2056 303 2136 317
rect 3239 365 3253 417
rect 3305 365 3319 417
rect 3239 345 3319 365
rect 3239 293 3253 345
rect 3305 293 3319 345
rect 1355 270 1435 284
rect 3239 279 3319 293
rect 1355 218 1369 270
rect 1421 218 1435 270
rect 1355 204 1435 218
rect 1660 -151 1740 -137
rect 1660 -203 1674 -151
rect 1726 -203 1740 -151
rect 1660 -217 1740 -203
rect 884 -345 1205 -245
rect 2085 -345 2417 -245
rect 556 -387 636 -373
rect 556 -439 570 -387
rect 622 -439 636 -387
rect 556 -453 636 -439
rect 3239 -387 3319 -373
rect 3239 -439 3253 -387
rect 3305 -439 3319 -387
rect 3239 -453 3319 -439
rect 3303 -874 3383 -860
rect 3303 -926 3317 -874
rect 3369 -926 3383 -874
rect 3303 -946 3383 -926
rect 1270 -993 1350 -979
rect 1270 -1045 1284 -993
rect 1336 -1045 1350 -993
rect 3303 -998 3317 -946
rect 3369 -998 3383 -946
rect 3303 -1012 3383 -998
rect 1270 -1059 1350 -1045
rect -461 -1923 -353 -1823
rect 657 -1923 1169 -1823
rect 2085 -1923 2417 -1823
<< via1 >>
rect -1473 1207 -1421 1259
rect -1473 1139 -1421 1191
rect -1473 1071 -1421 1123
rect -1131 -459 -1079 -407
rect -1131 -527 -1079 -475
rect -1131 -595 -1079 -543
rect -1131 -978 -1079 -926
rect -1131 -1046 -1079 -994
rect -1131 -1114 -1079 -1062
rect -1017 -615 -965 -563
rect -1017 -683 -965 -631
rect -1017 -751 -965 -699
rect -903 -139 -851 -87
rect -903 -207 -851 -155
rect -903 -275 -851 -223
rect 1674 1182 1726 1191
rect 1674 1148 1683 1182
rect 1683 1148 1717 1182
rect 1717 1148 1726 1182
rect 1674 1139 1726 1148
rect 1339 452 1391 461
rect 1339 418 1348 452
rect 1348 418 1382 452
rect 1382 418 1391 452
rect 1339 409 1391 418
rect 2496 446 2548 455
rect 2496 412 2505 446
rect 2505 412 2539 446
rect 2539 412 2548 446
rect 2496 403 2548 412
rect 2070 360 2122 369
rect 2070 326 2079 360
rect 2079 326 2113 360
rect 2113 326 2122 360
rect 2070 317 2122 326
rect 3253 408 3305 417
rect 3253 374 3262 408
rect 3262 374 3296 408
rect 3296 374 3305 408
rect 3253 365 3305 374
rect 3253 336 3305 345
rect 3253 302 3262 336
rect 3262 302 3296 336
rect 3296 302 3305 336
rect 3253 293 3305 302
rect 1369 261 1421 270
rect 1369 227 1378 261
rect 1378 227 1412 261
rect 1412 227 1421 261
rect 1369 218 1421 227
rect 1674 -160 1726 -151
rect 1674 -194 1683 -160
rect 1683 -194 1717 -160
rect 1717 -194 1726 -160
rect 1674 -203 1726 -194
rect 570 -396 622 -387
rect 570 -430 579 -396
rect 579 -430 613 -396
rect 613 -430 622 -396
rect 570 -439 622 -430
rect 3253 -396 3305 -387
rect 3253 -430 3262 -396
rect 3262 -430 3296 -396
rect 3296 -430 3305 -396
rect 3253 -439 3305 -430
rect 3317 -883 3369 -874
rect 3317 -917 3326 -883
rect 3326 -917 3360 -883
rect 3360 -917 3369 -883
rect 3317 -926 3369 -917
rect 1284 -1002 1336 -993
rect 1284 -1036 1293 -1002
rect 1293 -1036 1327 -1002
rect 1327 -1036 1336 -1002
rect 1284 -1045 1336 -1036
rect 3317 -955 3369 -946
rect 3317 -989 3326 -955
rect 3326 -989 3360 -955
rect 3360 -989 3369 -955
rect 3317 -998 3369 -989
<< metal2 >>
rect -1487 1259 -1407 1273
rect -1487 1207 -1473 1259
rect -1421 1207 -1407 1259
rect -1487 1191 -1407 1207
rect -1487 1139 -1473 1191
rect -1421 1185 -1407 1191
rect 1660 1191 1740 1205
rect 1660 1185 1674 1191
rect -1421 1145 1674 1185
rect -1421 1139 -1407 1145
rect -1487 1123 -1407 1139
rect 1660 1139 1674 1145
rect 1726 1139 1740 1191
rect 1660 1125 1740 1139
rect -1487 1071 -1473 1123
rect -1421 1071 -1407 1123
rect -1487 1057 -1407 1071
rect 1325 461 1405 475
rect 1325 455 1339 461
rect 980 415 1339 455
rect -917 -87 -837 -73
rect -917 -139 -903 -87
rect -851 -139 -837 -87
rect -917 -155 -837 -139
rect -917 -207 -903 -155
rect -851 -161 -837 -155
rect 980 -161 1020 415
rect 1325 409 1339 415
rect 1391 409 1405 461
rect 2482 455 2562 469
rect 2482 449 2496 455
rect 1325 395 1405 409
rect 2164 409 2496 449
rect 2056 369 2136 383
rect 2056 317 2070 369
rect 2122 317 2136 369
rect 2056 303 2136 317
rect 1355 270 1435 284
rect 1355 218 1369 270
rect 1421 218 1435 270
rect 1355 204 1435 218
rect -851 -201 1020 -161
rect -851 -207 -837 -201
rect -917 -223 -837 -207
rect -917 -275 -903 -223
rect -851 -275 -837 -223
rect -917 -289 -837 -275
rect 556 -387 636 -373
rect -1145 -407 -1065 -393
rect -1145 -459 -1131 -407
rect -1079 -459 -1065 -407
rect 556 -439 570 -387
rect 622 -393 636 -387
rect 1375 -393 1415 204
rect 1660 -151 1740 -137
rect 1660 -203 1674 -151
rect 1726 -203 1740 -151
rect 1660 -217 1740 -203
rect 622 -433 1415 -393
rect 622 -439 636 -433
rect 556 -453 636 -439
rect -1145 -475 -1065 -459
rect -1145 -527 -1131 -475
rect -1079 -481 -1065 -475
rect 1680 -481 1720 -217
rect -1079 -521 1720 -481
rect -1079 -527 -1065 -521
rect -1145 -543 -1065 -527
rect -1145 -595 -1131 -543
rect -1079 -595 -1065 -543
rect 2164 -549 2204 409
rect 2482 403 2496 409
rect 2548 403 2562 455
rect 2482 389 2562 403
rect 3239 417 3319 431
rect 3239 365 3253 417
rect 3305 365 3319 417
rect 3239 345 3319 365
rect 3239 293 3253 345
rect 3305 293 3319 345
rect 3239 279 3319 293
rect 3259 -373 3299 279
rect 3239 -387 3319 -373
rect 3239 -439 3253 -387
rect 3305 -439 3319 -387
rect 3239 -453 3319 -439
rect -1145 -609 -1065 -595
rect -1031 -563 2204 -549
rect -1031 -615 -1017 -563
rect -965 -589 2204 -563
rect -965 -615 -951 -589
rect -1031 -631 -951 -615
rect -1031 -683 -1017 -631
rect -965 -683 -951 -631
rect -1031 -699 -951 -683
rect -1031 -751 -1017 -699
rect -965 -751 -951 -699
rect -1031 -765 -951 -751
rect 3303 -874 3383 -860
rect -1145 -926 -1065 -912
rect -1145 -978 -1131 -926
rect -1079 -978 -1065 -926
rect -1145 -994 -1065 -978
rect 3303 -926 3317 -874
rect 3369 -916 3383 -874
rect 3369 -926 3428 -916
rect 3303 -946 3428 -926
rect -1145 -1046 -1131 -994
rect -1079 -1000 -1065 -994
rect 1270 -993 1350 -979
rect 1270 -1000 1284 -993
rect -1079 -1040 1284 -1000
rect -1079 -1046 -1065 -1040
rect -1145 -1062 -1065 -1046
rect 1270 -1045 1284 -1040
rect 1336 -1045 1350 -993
rect 3303 -998 3317 -946
rect 3369 -956 3428 -946
rect 3369 -998 3383 -956
rect 3303 -1012 3383 -998
rect 1270 -1059 1350 -1045
rect -1145 -1114 -1131 -1062
rect -1079 -1114 -1065 -1062
rect -1145 -1128 -1065 -1114
use CMOS_3in_OR  CMOS_3in_OR_0
timestamp 1505767276
transform 1 0 2922 0 -1 -1089
box -541 -870 542 870
use CMOS_4in_AND  CMOS_4in_AND_0
timestamp 1505767276
transform 1 0 227 0 -1 -1089
box -616 -870 616 870
use CMOS_AND  CMOS_AND_0
timestamp 1505767276
transform 1 0 2857 0 1 499
box -476 -870 476 870
use CMOS_AND  CMOS_AND_1
timestamp 1505767276
transform 1 0 1645 0 -1 -1089
box -476 -870 476 870
use CMOS_XNOR  CMOS_XNOR_0
timestamp 1505767276
transform 1 0 260 0 1 499
box -649 -870 650 870
use CMOS_XOR  CMOS_XOR_0
timestamp 1505767276
transform 1 0 1645 0 1 499
box -476 -870 476 870
<< labels >>
flabel metal1 s -552 -312 -518 -278 2 FreeSans 3125 0 0 0 GND
port 1 nsew
flabel metal1 s -1477 1267 -1416 1327 2 FreeSans 3907 0 0 0 x0
port 2 nsew
flabel metal1 s -1364 1206 -1303 1266 2 FreeSans 3907 0 0 0 x0_bar
port 3 nsew
flabel metal1 s -1249 1267 -1188 1327 2 FreeSans 3907 0 0 0 x1
port 4 nsew
flabel metal1 s -1135 1206 -1074 1266 2 FreeSans 3907 0 0 0 x1_bar
port 5 nsew
flabel metal1 s -1021 1268 -960 1328 2 FreeSans 3907 0 0 0 x2
port 6 nsew
flabel metal1 s -908 1207 -847 1267 2 FreeSans 3907 0 0 0 x2_bar
port 7 nsew
flabel metal1 s -793 1268 -732 1328 2 FreeSans 3907 0 0 0 x3
port 8 nsew
flabel metal1 s -443 1267 -409 1301 2 FreeSans 3125 0 0 0 VDD
port 9 nsew
flabel metal1 s -678 1208 -617 1268 2 FreeSans 3907 0 0 0 x3_bar
port 10 nsew
flabel metal2 s 3326 -917 3360 -883 2 FreeSans 3125 0 0 0 s1
port 11 nsew
<< end >>
