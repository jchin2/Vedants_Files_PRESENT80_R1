* NGSPICE file created from EESPFAL_s0_flat.ext - technology: sky130A

.subckt EESPFAL_s0_flat GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar Dis1 Dis2 Dis3
+ s0 s0_bar CLK3 CLK2 CLK1
X0 EESPFAL_NAND_v3_0/OUT_bar Dis2.t0 GND.t43 GND.t12 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_6340_2870# EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/OUT GND.t34 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X2 CLK2.t17 EESPFAL_NOR_v3_0/B_bar EESPFAL_NOR_v3_0/B CLK2.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/B CLK1.t21 CLK1.t20 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 CLK1.t0 x2_bar.t0 EESPFAL_NAND_v3_0/B GND.t3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X5 EESPFAL_NAND_v3_0/A.t4 EESPFAL_NAND_v3_0/A_bar.t6 CLK1.t33 CLK1.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 CLK1.t8 EESPFAL_NAND_v3_0/A_bar.t7 EESPFAL_NAND_v3_0/A.t3 CLK1.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 GND.t33 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar GND.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X8 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar GND.t32 GND.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 EESPFAL_NAND_v3_0/B x1.t0 CLK1.t29 GND.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 EESPFAL_NAND_v3_1/B_bar Dis1.t0 GND.t46 GND.t10 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X11 CLK1.t25 x2.t0 a_2000_2190# GND.t47 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X12 GND.t23 Dis3.t0 s0_bar.t1 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 GND.t27 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar GND.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 CLK3.t10 EESPFAL_NAND_v3_0/OUT s0.t5 GND.t30 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 s0.t1 EESPFAL_NOR_v3_0/B CLK3.t1 GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 EESPFAL_NAND_v3_0/A_bar.t2 x3.t0 a_740_2870# GND.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X17 a_2000_2870# x3_bar.t0 EESPFAL_NAND_v3_0/A.t0 GND.t8 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X18 EESPFAL_NOR_v3_0/B_bar EESPFAL_NAND_v3_0/A.t6 CLK2.t10 GND.t4 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X19 CLK3.t5 s0.t6 s0_bar.t0 CLK3.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X20 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_NAND_v3_0/OUT CLK2.t21 CLK2.t20 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X21 EESPFAL_NAND_v3_1/B_bar EESPFAL_NAND_v3_1/B CLK1.t13 CLK1.t12 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X22 CLK1.t11 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar CLK1.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X23 CLK1.t19 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar CLK1.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X24 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar CLK1.t17 CLK1.t16 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X25 GND.t51 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar GND.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X26 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar GND.t2 GND.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X27 CLK2.t9 EESPFAL_NAND_v3_0/A.t7 a_6340_2870# GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X28 GND.t38 Dis1.t1 EESPFAL_NAND_v3_0/B GND.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X29 EESPFAL_NOR_v3_0/B_bar Dis2.t1 GND.t42 GND.t41 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X30 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X31 GND.t49 Dis1.t2 EESPFAL_NAND_v3_1/B GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X32 a_3060_2870# x1_bar.t0 CLK1.t9 GND.t5 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X33 EESPFAL_NOR_v3_0/B_bar EESPFAL_NOR_v3_0/B CLK2.t8 CLK2.t7 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X34 CLK2.t19 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar CLK2.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X35 CLK1.t22 x1.t1 EESPFAL_NAND_v3_1/B_bar GND.t45 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X36 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar CLK1.t4 CLK1.t3 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X37 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar CLK2.t3 CLK2.t2 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X38 GND.t40 Dis2.t2 EESPFAL_NAND_v3_0/OUT GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X39 CLK1.t2 EESPFAL_NAND_v3_1/B_bar EESPFAL_NAND_v3_1/B CLK1.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X40 CLK1.t15 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/B CLK1.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X41 EESPFAL_NAND_v3_0/A_bar.t0 Dis1.t3 GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X42 GND.t21 EESPFAL_NAND_v3_0/A.t8 EESPFAL_NAND_v3_0/A_bar.t1 GND.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X43 CLK1.t24 x0.t0 a_2000_2870# GND.t47 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X44 s0.t0 Dis3.t1 GND.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X45 a_6340_2190# EESPFAL_NOR_v3_0/B_bar s0_bar.t4 GND.t34 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X46 GND.t15 EESPFAL_NOR_v3_0/B EESPFAL_NOR_v3_0/B_bar GND.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X47 a_4320_2190# EESPFAL_NAND_v3_1/B EESPFAL_NOR_v3_0/B GND.t3 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X48 CLK2.t11 EESPFAL_NAND_v3_0/A_bar.t8 a_4320_2190# GND.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X49 CLK2.t13 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/OUT_bar GND.t30 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X50 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_NAND_v3_0/A_bar.t9 CLK2.t12 GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X51 EESPFAL_NOR_v3_0/B EESPFAL_NOR_v3_0/B_bar GND.t50 GND.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X52 EESPFAL_NAND_v3_0/B_bar x2.t1 a_3060_2870# GND.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X53 a_440_2870# x3_bar.t1 EESPFAL_NAND_v3_0/A_bar.t3 GND.t28 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X54 s0.t3 s0_bar.t5 CLK3.t9 CLK3.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X55 EESPFAL_NAND_v3_1/B_bar x2_bar.t1 CLK1.t6 GND.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X56 a_2000_2190# x1_bar.t1 EESPFAL_NAND_v3_1/B GND.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X57 CLK2.t6 EESPFAL_NOR_v3_0/B EESPFAL_NOR_v3_0/B_bar CLK2.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X58 EESPFAL_NOR_v3_0/B EESPFAL_NOR_v3_0/B_bar CLK2.t15 CLK2.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X59 EESPFAL_NAND_v3_0/A_bar.t5 EESPFAL_NAND_v3_0/A.t9 CLK1.t31 CLK1.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X60 CLK1.t28 EESPFAL_NAND_v3_0/A.t10 EESPFAL_NAND_v3_0/A_bar.t4 CLK1.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X61 CLK2.t1 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_NAND_v3_0/OUT CLK2.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X62 EESPFAL_NAND_v3_0/B_bar Dis1.t4 GND.t44 GND.t41 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X63 EESPFAL_NAND_v3_0/A.t2 EESPFAL_NAND_v3_0/A_bar.t10 GND.t24 GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X64 a_2300_2870# x0_bar.t0 CLK1.t26 GND.t48 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X65 GND.t18 s0_bar.t6 s0.t2 GND.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X66 CLK3.t0 EESPFAL_NAND_v3_0/OUT_bar a_6340_2190# GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X67 GND.t36 Dis1.t5 EESPFAL_NAND_v3_0/A.t5 GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X68 EESPFAL_NAND_v3_0/A.t1 x3.t1 a_2300_2870# GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X69 s0_bar.t3 s0.t7 GND.t26 GND.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X70 GND.t39 Dis2.t3 EESPFAL_NOR_v3_0/B GND.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X71 CLK1.t5 x0_bar.t1 a_440_2870# GND.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X72 a_740_2870# x0.t1 CLK1.t23 GND.t45 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X73 CLK2.t4 EESPFAL_NAND_v3_1/B_bar EESPFAL_NOR_v3_0/B_bar GND.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X74 CLK3.t7 s0_bar.t7 s0.t4 CLK3.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X75 s0_bar.t2 s0.t8 CLK3.t3 CLK3.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
R0 Dis2.n0 Dis2.t2 504.5
R1 Dis2.n3 Dis2.n2 403.84
R2 Dis2.n2 Dis2.t3 389.3
R3 Dis2.n1 Dis2.t1 389.3
R4 Dis2.n0 Dis2.t0 389.3
R5 Dis2 Dis2.n3 149.76
R6 Dis2.n2 Dis2.n1 115.2
R7 Dis2.n3 Dis2 7.383
R8 Dis2.n1 EESPFAL_NAND_v3_1/Dis 3.2
R9 Dis2 Dis2.n0 3.2
R10 GND.n224 GND.t28 269.289
R11 GND.n168 GND.t29 269.289
R12 GND.n230 GND.t9 133.857
R13 GND.n175 GND.t48 133.857
R14 GND.n6 GND.t0 70.155
R15 GND.n80 GND.t30 70.155
R16 GND.n88 GND.t25 70.155
R17 GND.n162 GND.t5 70.155
R18 GND.n183 GND.t47 63.953
R19 GND.n208 GND.t35 63.953
R20 GND.n263 GND.t10 63.953
R21 GND.n238 GND.t45 63.953
R22 GND.n31 GND.t22 63.953
R23 GND.n55 GND.t12 63.953
R24 GND.n113 GND.t37 63.953
R25 GND.n137 GND.t41 63.953
R26 GND.n225 GND 31.565
R27 GND.n30 GND.t40 29.103
R28 GND.n59 GND.t43 29.103
R29 GND.n112 GND.t38 29.103
R30 GND.n141 GND.t44 29.103
R31 GND.n207 GND.t36 29.103
R32 GND.n262 GND.t11 29.103
R33 GND.n30 GND.t23 29.102
R34 GND.n59 GND.t13 29.102
R35 GND.n112 GND.t39 29.102
R36 GND.n141 GND.t42 29.102
R37 GND.n207 GND.t49 29.102
R38 GND.n262 GND.t46 29.102
R39 GND.n1 GND.t7 24
R40 GND.n1 GND.t27 24
R41 GND.n0 GND.t24 24
R42 GND.n0 GND.t21 24
R43 GND.n5 GND.t26 24
R44 GND.n5 GND.t18 24
R45 GND.n4 GND.t2 24
R46 GND.n4 GND.t51 24
R47 GND.n3 GND.t50 24
R48 GND.n3 GND.t15 24
R49 GND.n2 GND.t32 24
R50 GND.n2 GND.t33 24
R51 GND.n191 GND.t8 21.317
R52 GND.n216 GND.t6 21.317
R53 GND.n271 GND.t20 21.317
R54 GND.n246 GND.t19 21.317
R55 GND.n14 GND.t34 21.317
R56 GND.n39 GND.t1 21.317
R57 GND.n47 GND.t17 21.317
R58 GND.n72 GND.t16 21.317
R59 GND.n96 GND.t3 21.317
R60 GND.n121 GND.t31 21.317
R61 GND.n129 GND.t14 21.317
R62 GND.n154 GND.t4 21.317
R63 GND.n49 GND.n46 12.8
R64 GND.n131 GND.n128 12.8
R65 GND.n8 GND.n7 9.154
R66 GND.n90 GND.n89 9.154
R67 GND.n94 GND.n93 9.154
R68 GND.n93 GND.n92 9.154
R69 GND.n98 GND.n97 9.154
R70 GND.n97 GND.n96 9.154
R71 GND.n102 GND.n101 9.154
R72 GND.n101 GND.n100 9.154
R73 GND.n106 GND.n105 9.154
R74 GND.n105 GND.n104 9.154
R75 GND.n110 GND.n109 9.154
R76 GND.n109 GND.n108 9.154
R77 GND.n115 GND.n114 9.154
R78 GND.n114 GND.n113 9.154
R79 GND.n119 GND.n118 9.154
R80 GND.n118 GND.n117 9.154
R81 GND.n123 GND.n122 9.154
R82 GND.n122 GND.n121 9.154
R83 GND.n128 GND.n127 9.154
R84 GND.n127 GND.n126 9.154
R85 GND.n131 GND.n130 9.154
R86 GND.n130 GND.n129 9.154
R87 GND.n135 GND.n134 9.154
R88 GND.n134 GND.n133 9.154
R89 GND.n139 GND.n138 9.154
R90 GND.n138 GND.n137 9.154
R91 GND.n144 GND.n143 9.154
R92 GND.n143 GND.n142 9.154
R93 GND.n148 GND.n147 9.154
R94 GND.n147 GND.n146 9.154
R95 GND.n152 GND.n151 9.154
R96 GND.n151 GND.n150 9.154
R97 GND.n156 GND.n155 9.154
R98 GND.n155 GND.n154 9.154
R99 GND.n160 GND.n159 9.154
R100 GND.n159 GND.n158 9.154
R101 GND.n164 GND.n163 9.154
R102 GND.n12 GND.n11 9.154
R103 GND.n11 GND.n10 9.154
R104 GND.n16 GND.n15 9.154
R105 GND.n15 GND.n14 9.154
R106 GND.n20 GND.n19 9.154
R107 GND.n19 GND.n18 9.154
R108 GND.n24 GND.n23 9.154
R109 GND.n23 GND.n22 9.154
R110 GND.n28 GND.n27 9.154
R111 GND.n27 GND.n26 9.154
R112 GND.n33 GND.n32 9.154
R113 GND.n32 GND.n31 9.154
R114 GND.n37 GND.n36 9.154
R115 GND.n36 GND.n35 9.154
R116 GND.n41 GND.n40 9.154
R117 GND.n40 GND.n39 9.154
R118 GND.n46 GND.n45 9.154
R119 GND.n45 GND.n44 9.154
R120 GND.n49 GND.n48 9.154
R121 GND.n48 GND.n47 9.154
R122 GND.n53 GND.n52 9.154
R123 GND.n52 GND.n51 9.154
R124 GND.n57 GND.n56 9.154
R125 GND.n56 GND.n55 9.154
R126 GND.n62 GND.n61 9.154
R127 GND.n61 GND.n60 9.154
R128 GND.n66 GND.n65 9.154
R129 GND.n65 GND.n64 9.154
R130 GND.n70 GND.n69 9.154
R131 GND.n69 GND.n68 9.154
R132 GND.n74 GND.n73 9.154
R133 GND.n73 GND.n72 9.154
R134 GND.n78 GND.n77 9.154
R135 GND.n77 GND.n76 9.154
R136 GND.n82 GND.n81 9.154
R137 GND.n173 GND.n172 9.154
R138 GND.n172 GND.n171 9.154
R139 GND.n177 GND.n176 9.154
R140 GND.n176 GND.n175 9.154
R141 GND.n181 GND.n180 9.154
R142 GND.n180 GND.n179 9.154
R143 GND.n185 GND.n184 9.154
R144 GND.n184 GND.n183 9.154
R145 GND.n189 GND.n188 9.154
R146 GND.n188 GND.n187 9.154
R147 GND.n193 GND.n192 9.154
R148 GND.n192 GND.n191 9.154
R149 GND.n197 GND.n196 9.154
R150 GND.n196 GND.n195 9.154
R151 GND.n201 GND.n200 9.154
R152 GND.n200 GND.n199 9.154
R153 GND.n205 GND.n204 9.154
R154 GND.n204 GND.n203 9.154
R155 GND.n210 GND.n209 9.154
R156 GND.n209 GND.n208 9.154
R157 GND.n214 GND.n213 9.154
R158 GND.n213 GND.n212 9.154
R159 GND.n218 GND.n217 9.154
R160 GND.n217 GND.n216 9.154
R161 GND.n222 GND.n221 9.154
R162 GND.n221 GND.n220 9.154
R163 GND.n273 GND.n272 9.154
R164 GND.n272 GND.n271 9.154
R165 GND.n269 GND.n268 9.154
R166 GND.n268 GND.n267 9.154
R167 GND.n265 GND.n264 9.154
R168 GND.n264 GND.n263 9.154
R169 GND.n260 GND.n259 9.154
R170 GND.n259 GND.n258 9.154
R171 GND.n256 GND.n255 9.154
R172 GND.n255 GND.n254 9.154
R173 GND.n252 GND.n251 9.154
R174 GND.n251 GND.n250 9.154
R175 GND.n248 GND.n247 9.154
R176 GND.n247 GND.n246 9.154
R177 GND.n244 GND.n243 9.154
R178 GND.n243 GND.n242 9.154
R179 GND.n240 GND.n239 9.154
R180 GND.n239 GND.n238 9.154
R181 GND.n236 GND.n235 9.154
R182 GND.n235 GND.n234 9.154
R183 GND.n232 GND.n231 9.154
R184 GND.n231 GND.n230 9.154
R185 GND.n228 GND.n227 9.154
R186 GND.n227 GND.n226 9.154
R187 GND.n225 GND.n224 9.154
R188 GND.n169 GND.n168 9.154
R189 GND.n223 GND.n1 5.103
R190 GND.n223 GND.n0 5.103
R191 GND.n43 GND.n5 5.103
R192 GND.n43 GND.n4 5.103
R193 GND.n125 GND.n3 5.103
R194 GND.n125 GND.n2 5.103
R195 GND.n167 GND.n166 4.65
R196 GND.n91 GND.n90 4.65
R197 GND.n95 GND.n94 4.65
R198 GND.n99 GND.n98 4.65
R199 GND.n103 GND.n102 4.65
R200 GND.n107 GND.n106 4.65
R201 GND.n111 GND.n110 4.65
R202 GND.n116 GND.n115 4.65
R203 GND.n120 GND.n119 4.65
R204 GND.n124 GND.n123 4.65
R205 GND.n128 GND.n125 4.65
R206 GND.n132 GND.n131 4.65
R207 GND.n136 GND.n135 4.65
R208 GND.n140 GND.n139 4.65
R209 GND.n145 GND.n144 4.65
R210 GND.n149 GND.n148 4.65
R211 GND.n153 GND.n152 4.65
R212 GND.n157 GND.n156 4.65
R213 GND.n161 GND.n160 4.65
R214 GND.n165 GND.n164 4.65
R215 GND.n87 GND.n86 4.65
R216 GND.n85 GND.n84 4.65
R217 GND.n13 GND.n12 4.65
R218 GND.n17 GND.n16 4.65
R219 GND.n21 GND.n20 4.65
R220 GND.n25 GND.n24 4.65
R221 GND.n29 GND.n28 4.65
R222 GND.n34 GND.n33 4.65
R223 GND.n38 GND.n37 4.65
R224 GND.n42 GND.n41 4.65
R225 GND.n46 GND.n43 4.65
R226 GND.n50 GND.n49 4.65
R227 GND.n54 GND.n53 4.65
R228 GND.n58 GND.n57 4.65
R229 GND.n63 GND.n62 4.65
R230 GND.n67 GND.n66 4.65
R231 GND.n71 GND.n70 4.65
R232 GND.n75 GND.n74 4.65
R233 GND.n79 GND.n78 4.65
R234 GND.n83 GND.n82 4.65
R235 GND.n174 GND.n173 4.65
R236 GND.n178 GND.n177 4.65
R237 GND.n182 GND.n181 4.65
R238 GND.n186 GND.n185 4.65
R239 GND.n190 GND.n189 4.65
R240 GND.n194 GND.n193 4.65
R241 GND.n198 GND.n197 4.65
R242 GND.n202 GND.n201 4.65
R243 GND.n206 GND.n205 4.65
R244 GND.n211 GND.n210 4.65
R245 GND.n215 GND.n214 4.65
R246 GND.n219 GND.n218 4.65
R247 GND.n223 GND.n222 4.65
R248 GND.n274 GND.n273 4.65
R249 GND.n270 GND.n269 4.65
R250 GND.n266 GND.n265 4.65
R251 GND.n261 GND.n260 4.65
R252 GND.n257 GND.n256 4.65
R253 GND.n253 GND.n252 4.65
R254 GND.n249 GND.n248 4.65
R255 GND.n245 GND.n244 4.65
R256 GND.n241 GND.n240 4.65
R257 GND.n237 GND.n236 4.65
R258 GND.n233 GND.n232 4.65
R259 GND.n170 GND.n169 4.65
R260 GND.n7 GND.n6 2.791
R261 GND.n89 GND.n88 2.791
R262 GND.n163 GND.n162 2.791
R263 GND.n81 GND.n80 2.791
R264 GND.n229 GND.n225 2.739
R265 GND.n9 GND.n8 2.682
R266 GND.n229 GND.n228 2.682
R267 GND.n13 GND.n9 1.095
R268 GND.n233 GND.n229 1.095
R269 GND.n170 GND.n167 0.6
R270 GND.n87 GND.n85 0.525
R271 GND.n17 GND.n13 0.1
R272 GND.n21 GND.n17 0.1
R273 GND.n25 GND.n21 0.1
R274 GND.n29 GND.n25 0.1
R275 GND.n38 GND.n34 0.1
R276 GND.n42 GND.n38 0.1
R277 GND.n43 GND.n42 0.1
R278 GND.n54 GND.n50 0.1
R279 GND.n58 GND.n54 0.1
R280 GND.n67 GND.n63 0.1
R281 GND.n71 GND.n67 0.1
R282 GND.n75 GND.n71 0.1
R283 GND.n79 GND.n75 0.1
R284 GND.n83 GND.n79 0.1
R285 GND.n85 GND.n83 0.1
R286 GND.n91 GND.n87 0.1
R287 GND.n95 GND.n91 0.1
R288 GND.n99 GND.n95 0.1
R289 GND.n103 GND.n99 0.1
R290 GND.n107 GND.n103 0.1
R291 GND.n111 GND.n107 0.1
R292 GND.n120 GND.n116 0.1
R293 GND.n124 GND.n120 0.1
R294 GND.n125 GND.n124 0.1
R295 GND.n136 GND.n132 0.1
R296 GND.n140 GND.n136 0.1
R297 GND.n149 GND.n145 0.1
R298 GND.n153 GND.n149 0.1
R299 GND.n157 GND.n153 0.1
R300 GND.n161 GND.n157 0.1
R301 GND.n165 GND.n161 0.1
R302 GND.n167 GND.n165 0.1
R303 GND.n174 GND.n170 0.1
R304 GND.n178 GND.n174 0.1
R305 GND.n182 GND.n178 0.1
R306 GND.n186 GND.n182 0.1
R307 GND.n190 GND.n186 0.1
R308 GND.n194 GND.n190 0.1
R309 GND.n198 GND.n194 0.1
R310 GND.n202 GND.n198 0.1
R311 GND.n206 GND.n202 0.1
R312 GND.n215 GND.n211 0.1
R313 GND.n219 GND.n215 0.1
R314 GND.n223 GND.n219 0.1
R315 GND.n274 GND.n270 0.1
R316 GND.n270 GND.n266 0.1
R317 GND.n261 GND.n257 0.1
R318 GND.n257 GND.n253 0.1
R319 GND.n253 GND.n249 0.1
R320 GND.n249 GND.n245 0.1
R321 GND.n245 GND.n241 0.1
R322 GND.n241 GND.n237 0.1
R323 GND.n237 GND.n233 0.1
R324 GND.n34 GND.n30 0.075
R325 GND.n50 GND 0.075
R326 GND.n59 GND.n58 0.075
R327 GND.n116 GND.n112 0.075
R328 GND.n132 EESPFAL_NAND_v3_1/GND 0.075
R329 GND.n141 GND.n140 0.075
R330 GND.n211 GND.n207 0.075
R331 EESPFAL_NAND_v3_2/GND GND.n274 0.075
R332 GND.n266 GND.n262 0.075
R333 GND.n30 GND.n29 0.025
R334 GND.n43 GND 0.025
R335 GND.n63 GND.n59 0.025
R336 GND.n112 GND.n111 0.025
R337 GND.n125 EESPFAL_NAND_v3_1/GND 0.025
R338 GND.n145 GND.n141 0.025
R339 GND.n207 GND.n206 0.025
R340 EESPFAL_NAND_v3_2/GND GND.n223 0.025
R341 GND.n262 GND.n261 0.025
R342 CLK2.n103 CLK2.t17 44.338
R343 CLK2.n74 CLK2.t8 44.338
R344 CLK2.n171 CLK2.t21 44.337
R345 CLK2.n27 CLK2.t1 44.337
R346 CLK2.n47 CLK2.t15 39.4
R347 CLK2.n47 CLK2.t6 39.4
R348 CLK2.n0 CLK2.t3 39.4
R349 CLK2.n0 CLK2.t19 39.4
R350 CLK2.n2 CLK2.t9 30.775
R351 CLK2.n99 CLK2.t16 24.568
R352 CLK2.n75 CLK2.t7 24.568
R353 CLK2.n28 CLK2.t0 24.568
R354 CLK2.n172 CLK2.t20 24.568
R355 CLK2.n133 CLK2.t11 24
R356 CLK2.n48 CLK2.t10 24
R357 CLK2.n48 CLK2.t4 24
R358 CLK2.n137 CLK2.t12 24
R359 CLK2.n137 CLK2.t13 24
R360 CLK2.n89 CLK2.n86 12.8
R361 CLK2.n126 CLK2.n125 8.855
R362 CLK2.n122 CLK2.n121 8.855
R363 CLK2.n121 CLK2.n120 8.855
R364 CLK2.n118 CLK2.n117 8.855
R365 CLK2.n117 CLK2.n116 8.855
R366 CLK2.n114 CLK2.n113 8.855
R367 CLK2.n113 CLK2.n112 8.855
R368 CLK2.n110 CLK2.n109 8.855
R369 CLK2.n109 CLK2.n108 8.855
R370 CLK2.n106 CLK2.n105 8.855
R371 CLK2.n105 CLK2.n104 8.855
R372 CLK2.n101 CLK2.n100 8.855
R373 CLK2.n100 CLK2.n99 8.855
R374 CLK2.n97 CLK2.n96 8.855
R375 CLK2.n96 CLK2.n95 8.855
R376 CLK2.n93 CLK2.n92 8.855
R377 CLK2.n92 CLK2.n91 8.855
R378 CLK2.n89 CLK2.n88 8.855
R379 CLK2.n88 CLK2.n87 8.855
R380 CLK2.n86 CLK2.n85 8.855
R381 CLK2.n85 CLK2.n84 8.855
R382 CLK2.n81 CLK2.n80 8.855
R383 CLK2.n80 CLK2.n79 8.855
R384 CLK2.n77 CLK2.n76 8.855
R385 CLK2.n76 CLK2.n75 8.855
R386 CLK2.n72 CLK2.n71 8.855
R387 CLK2.n71 CLK2.n70 8.855
R388 CLK2.n68 CLK2.n67 8.855
R389 CLK2.n67 CLK2.n66 8.855
R390 CLK2.n64 CLK2.n63 8.855
R391 CLK2.n63 CLK2.n62 8.855
R392 CLK2.n60 CLK2.n59 8.855
R393 CLK2.n59 CLK2.n58 8.855
R394 CLK2.n55 CLK2.n54 8.855
R395 CLK2.n54 CLK2.n53 8.855
R396 CLK2.n51 CLK2.n50 8.855
R397 CLK2.n5 CLK2.n4 8.855
R398 CLK2.n9 CLK2.n8 8.855
R399 CLK2.n8 CLK2.n7 8.855
R400 CLK2.n13 CLK2.n12 8.855
R401 CLK2.n12 CLK2.n11 8.855
R402 CLK2.n17 CLK2.n16 8.855
R403 CLK2.n16 CLK2.n15 8.855
R404 CLK2.n21 CLK2.n20 8.855
R405 CLK2.n20 CLK2.n19 8.855
R406 CLK2.n25 CLK2.n24 8.855
R407 CLK2.n24 CLK2.n23 8.855
R408 CLK2.n30 CLK2.n29 8.855
R409 CLK2.n29 CLK2.n28 8.855
R410 CLK2.n34 CLK2.n33 8.855
R411 CLK2.n33 CLK2.n32 8.855
R412 CLK2.n38 CLK2.n37 8.855
R413 CLK2.n37 CLK2.n36 8.855
R414 CLK2.n42 CLK2.n41 8.855
R415 CLK2.n41 CLK2.n40 8.855
R416 CLK2.n182 CLK2.n181 8.855
R417 CLK2.n181 CLK2.n180 8.855
R418 CLK2.n178 CLK2.n177 8.855
R419 CLK2.n177 CLK2.n176 8.855
R420 CLK2.n174 CLK2.n173 8.855
R421 CLK2.n173 CLK2.n172 8.855
R422 CLK2.n169 CLK2.n168 8.855
R423 CLK2.n168 CLK2.n167 8.855
R424 CLK2.n165 CLK2.n164 8.855
R425 CLK2.n164 CLK2.n163 8.855
R426 CLK2.n161 CLK2.n160 8.855
R427 CLK2.n160 CLK2.n159 8.855
R428 CLK2.n157 CLK2.n156 8.855
R429 CLK2.n156 CLK2.n155 8.855
R430 CLK2.n151 CLK2.n149 8.855
R431 CLK2.n149 CLK2.n148 8.855
R432 CLK2.n145 CLK2.n144 8.855
R433 CLK2.n135 CLK2.n134 8.365
R434 CLK2.n91 CLK2.t14 8.189
R435 CLK2.n84 CLK2.t5 8.189
R436 CLK2.n36 CLK2.t2 8.189
R437 CLK2.n180 CLK2.t18 8.189
R438 CLK2.n136 CLK2.n135 7.422
R439 CLK2.n57 CLK2.n48 6.776
R440 CLK2.n90 CLK2.n47 4.938
R441 CLK2.n43 CLK2.n0 4.938
R442 CLK2.n128 CLK2.n46 4.675
R443 CLK2.n2 CLK2.n1 4.675
R444 CLK2.n127 CLK2.n126 4.65
R445 CLK2.n123 CLK2.n122 4.65
R446 CLK2.n119 CLK2.n118 4.65
R447 CLK2.n115 CLK2.n114 4.65
R448 CLK2.n111 CLK2.n110 4.65
R449 CLK2.n107 CLK2.n106 4.65
R450 CLK2.n102 CLK2.n101 4.65
R451 CLK2.n98 CLK2.n97 4.65
R452 CLK2.n94 CLK2.n93 4.65
R453 CLK2.n90 CLK2.n89 4.65
R454 CLK2.n86 CLK2.n83 4.65
R455 CLK2.n82 CLK2.n81 4.65
R456 CLK2.n78 CLK2.n77 4.65
R457 CLK2.n73 CLK2.n72 4.65
R458 CLK2.n69 CLK2.n68 4.65
R459 CLK2.n65 CLK2.n64 4.65
R460 CLK2.n61 CLK2.n60 4.65
R461 CLK2.n56 CLK2.n55 4.65
R462 CLK2.n132 CLK2.n131 4.65
R463 CLK2.n130 CLK2.n129 4.65
R464 CLK2.n141 CLK2.n45 4.65
R465 CLK2.n140 CLK2.n139 4.65
R466 CLK2.n6 CLK2.n5 4.65
R467 CLK2.n10 CLK2.n9 4.65
R468 CLK2.n14 CLK2.n13 4.65
R469 CLK2.n18 CLK2.n17 4.65
R470 CLK2.n22 CLK2.n21 4.65
R471 CLK2.n26 CLK2.n25 4.65
R472 CLK2.n31 CLK2.n30 4.65
R473 CLK2.n35 CLK2.n34 4.65
R474 CLK2.n39 CLK2.n38 4.65
R475 CLK2.n43 CLK2.n42 4.65
R476 CLK2.n183 CLK2.n182 4.65
R477 CLK2.n179 CLK2.n178 4.65
R478 CLK2.n175 CLK2.n174 4.65
R479 CLK2.n170 CLK2.n169 4.65
R480 CLK2.n166 CLK2.n165 4.65
R481 CLK2.n162 CLK2.n161 4.65
R482 CLK2.n158 CLK2.n157 4.65
R483 CLK2.n139 CLK2.n138 3.715
R484 CLK2.n152 CLK2.n151 3.033
R485 CLK2.n151 CLK2.n150 2.72
R486 CLK2.n52 CLK2.n51 2.682
R487 CLK2.n146 CLK2.n145 2.682
R488 CLK2.n134 CLK2.n133 2.57
R489 CLK2.n138 CLK2.n137 2.57
R490 CLK2.n153 CLK2.n142 2.251
R491 CLK2.n154 CLK2.n44 2.246
R492 CLK2.n130 CLK2.n128 2.203
R493 CLK2.n153 CLK2.n141 2.203
R494 CLK2.n4 CLK2.n3 1.655
R495 CLK2.n125 CLK2.n124 1.655
R496 CLK2.n50 CLK2.n49 1.655
R497 CLK2.n144 CLK2.n143 1.655
R498 CLK2.n56 CLK2.n52 1.095
R499 CLK2.n147 CLK2.n146 1.073
R500 CLK2.n142 CLK2 0.279
R501 CLK2.n132 CLK2.n130 0.125
R502 CLK2.n141 CLK2.n140 0.125
R503 CLK2.n140 CLK2.n136 0.125
R504 CLK2.n127 CLK2.n123 0.1
R505 CLK2.n123 CLK2.n119 0.1
R506 CLK2.n119 CLK2.n115 0.1
R507 CLK2.n115 CLK2.n111 0.1
R508 CLK2.n111 CLK2.n107 0.1
R509 CLK2.n102 CLK2.n98 0.1
R510 CLK2.n98 CLK2.n94 0.1
R511 CLK2.n94 CLK2.n90 0.1
R512 CLK2.n83 CLK2.n82 0.1
R513 CLK2.n82 CLK2.n78 0.1
R514 CLK2.n73 CLK2.n69 0.1
R515 CLK2.n69 CLK2.n65 0.1
R516 CLK2.n65 CLK2.n61 0.1
R517 CLK2.n10 CLK2.n6 0.1
R518 CLK2.n14 CLK2.n10 0.1
R519 CLK2.n18 CLK2.n14 0.1
R520 CLK2.n22 CLK2.n18 0.1
R521 CLK2.n26 CLK2.n22 0.1
R522 CLK2.n35 CLK2.n31 0.1
R523 CLK2.n39 CLK2.n35 0.1
R524 CLK2.n43 CLK2.n39 0.1
R525 CLK2.n183 CLK2.n179 0.1
R526 CLK2.n179 CLK2.n175 0.1
R527 CLK2.n170 CLK2.n166 0.1
R528 CLK2.n166 CLK2.n162 0.1
R529 CLK2.n162 CLK2.n158 0.1
R530 CLK2.n61 CLK2.n57 0.087
R531 CLK2.n158 CLK2.n154 0.077
R532 CLK2.n128 CLK2.n127 0.075
R533 CLK2.n103 CLK2.n102 0.075
R534 CLK2.n83 EESPFAL_NAND_v3_1/CLK 0.075
R535 CLK2.n78 CLK2.n74 0.075
R536 CLK2.n6 CLK2.n2 0.075
R537 CLK2.n31 CLK2.n27 0.075
R538 CLK2 CLK2.n183 0.075
R539 CLK2.n175 CLK2.n171 0.075
R540 CLK2.n135 CLK2.n132 0.062
R541 CLK2.n107 CLK2.n103 0.025
R542 CLK2.n90 EESPFAL_NAND_v3_1/CLK 0.025
R543 CLK2.n74 CLK2.n73 0.025
R544 CLK2.n27 CLK2.n26 0.025
R545 CLK2 CLK2.n43 0.025
R546 CLK2.n171 CLK2.n170 0.025
R547 CLK2.n152 CLK2.n147 0.021
R548 CLK2.n57 CLK2.n56 0.012
R549 CLK2.n153 CLK2.n152 0.012
R550 CLK2.n154 CLK2.n153 0.01
R551 CLK1.n27 CLK1.t2 44.338
R552 CLK1.n268 CLK1.t13 44.338
R553 CLK1.n200 CLK1.t31 44.337
R554 CLK1.n173 CLK1.t8 44.337
R555 CLK1.n106 CLK1.t21 44.337
R556 CLK1.n79 CLK1.t15 44.337
R557 CLK1.n48 CLK1.t33 39.4
R558 CLK1.n48 CLK1.t28 39.4
R559 CLK1.n52 CLK1.t17 39.4
R560 CLK1.n52 CLK1.t19 39.4
R561 CLK1.n0 CLK1.t4 39.4
R562 CLK1.n0 CLK1.t11 39.4
R563 CLK1.n2 CLK1.t25 30.776
R564 CLK1.n131 CLK1.t9 30.775
R565 CLK1.n174 CLK1.t7 24.568
R566 CLK1.n196 CLK1.t30 24.568
R567 CLK1.n80 CLK1.t14 24.568
R568 CLK1.n102 CLK1.t20 24.568
R569 CLK1.n28 CLK1.t1 24.568
R570 CLK1.n269 CLK1.t12 24.568
R571 CLK1.n45 CLK1.t23 24
R572 CLK1.n45 CLK1.t5 24
R573 CLK1.n49 CLK1.t26 24
R574 CLK1.n49 CLK1.t24 24
R575 CLK1.n53 CLK1.t29 24
R576 CLK1.n53 CLK1.t0 24
R577 CLK1.n44 CLK1.t6 24
R578 CLK1.n44 CLK1.t22 24
R579 CLK1.n190 CLK1.n187 12.8
R580 CLK1.n96 CLK1.n93 12.8
R581 CLK1.n56 CLK1.n55 8.855
R582 CLK1.n60 CLK1.n59 8.855
R583 CLK1.n59 CLK1.n58 8.855
R584 CLK1.n65 CLK1.n64 8.855
R585 CLK1.n64 CLK1.n63 8.855
R586 CLK1.n69 CLK1.n68 8.855
R587 CLK1.n68 CLK1.n67 8.855
R588 CLK1.n73 CLK1.n72 8.855
R589 CLK1.n72 CLK1.n71 8.855
R590 CLK1.n77 CLK1.n76 8.855
R591 CLK1.n76 CLK1.n75 8.855
R592 CLK1.n82 CLK1.n81 8.855
R593 CLK1.n81 CLK1.n80 8.855
R594 CLK1.n86 CLK1.n85 8.855
R595 CLK1.n85 CLK1.n84 8.855
R596 CLK1.n90 CLK1.n89 8.855
R597 CLK1.n89 CLK1.n88 8.855
R598 CLK1.n93 CLK1.n51 8.855
R599 CLK1.n51 CLK1.n50 8.855
R600 CLK1.n96 CLK1.n95 8.855
R601 CLK1.n95 CLK1.n94 8.855
R602 CLK1.n100 CLK1.n99 8.855
R603 CLK1.n99 CLK1.n98 8.855
R604 CLK1.n104 CLK1.n103 8.855
R605 CLK1.n103 CLK1.n102 8.855
R606 CLK1.n109 CLK1.n108 8.855
R607 CLK1.n108 CLK1.n107 8.855
R608 CLK1.n113 CLK1.n112 8.855
R609 CLK1.n112 CLK1.n111 8.855
R610 CLK1.n117 CLK1.n116 8.855
R611 CLK1.n116 CLK1.n115 8.855
R612 CLK1.n121 CLK1.n120 8.855
R613 CLK1.n120 CLK1.n119 8.855
R614 CLK1.n125 CLK1.n124 8.855
R615 CLK1.n124 CLK1.n123 8.855
R616 CLK1.n129 CLK1.n128 8.855
R617 CLK1.n138 CLK1.n137 8.855
R618 CLK1.n142 CLK1.n141 8.855
R619 CLK1.n141 CLK1.n140 8.855
R620 CLK1.n146 CLK1.n145 8.855
R621 CLK1.n145 CLK1.n144 8.855
R622 CLK1.n151 CLK1.n150 8.855
R623 CLK1.n150 CLK1.n149 8.855
R624 CLK1.n155 CLK1.n154 8.855
R625 CLK1.n154 CLK1.n153 8.855
R626 CLK1.n159 CLK1.n158 8.855
R627 CLK1.n158 CLK1.n157 8.855
R628 CLK1.n163 CLK1.n162 8.855
R629 CLK1.n162 CLK1.n161 8.855
R630 CLK1.n167 CLK1.n166 8.855
R631 CLK1.n166 CLK1.n165 8.855
R632 CLK1.n171 CLK1.n170 8.855
R633 CLK1.n170 CLK1.n169 8.855
R634 CLK1.n176 CLK1.n175 8.855
R635 CLK1.n175 CLK1.n174 8.855
R636 CLK1.n180 CLK1.n179 8.855
R637 CLK1.n179 CLK1.n178 8.855
R638 CLK1.n184 CLK1.n183 8.855
R639 CLK1.n183 CLK1.n182 8.855
R640 CLK1.n187 CLK1.n47 8.855
R641 CLK1.n47 CLK1.n46 8.855
R642 CLK1.n190 CLK1.n189 8.855
R643 CLK1.n189 CLK1.n188 8.855
R644 CLK1.n194 CLK1.n193 8.855
R645 CLK1.n193 CLK1.n192 8.855
R646 CLK1.n198 CLK1.n197 8.855
R647 CLK1.n197 CLK1.n196 8.855
R648 CLK1.n203 CLK1.n202 8.855
R649 CLK1.n202 CLK1.n201 8.855
R650 CLK1.n207 CLK1.n206 8.855
R651 CLK1.n206 CLK1.n205 8.855
R652 CLK1.n211 CLK1.n210 8.855
R653 CLK1.n210 CLK1.n209 8.855
R654 CLK1.n215 CLK1.n214 8.855
R655 CLK1.n214 CLK1.n213 8.855
R656 CLK1.n219 CLK1.n218 8.855
R657 CLK1.n218 CLK1.n217 8.855
R658 CLK1.n223 CLK1.n222 8.855
R659 CLK1.n222 CLK1.n221 8.855
R660 CLK1.n228 CLK1.n227 8.855
R661 CLK1.n227 CLK1.n226 8.855
R662 CLK1.n232 CLK1.n231 8.855
R663 CLK1.n231 CLK1.n230 8.855
R664 CLK1.n236 CLK1.n235 8.855
R665 CLK1.n5 CLK1.n4 8.855
R666 CLK1.n9 CLK1.n8 8.855
R667 CLK1.n8 CLK1.n7 8.855
R668 CLK1.n13 CLK1.n12 8.855
R669 CLK1.n12 CLK1.n11 8.855
R670 CLK1.n17 CLK1.n16 8.855
R671 CLK1.n16 CLK1.n15 8.855
R672 CLK1.n21 CLK1.n20 8.855
R673 CLK1.n20 CLK1.n19 8.855
R674 CLK1.n25 CLK1.n24 8.855
R675 CLK1.n24 CLK1.n23 8.855
R676 CLK1.n30 CLK1.n29 8.855
R677 CLK1.n29 CLK1.n28 8.855
R678 CLK1.n34 CLK1.n33 8.855
R679 CLK1.n33 CLK1.n32 8.855
R680 CLK1.n38 CLK1.n37 8.855
R681 CLK1.n37 CLK1.n36 8.855
R682 CLK1.n42 CLK1.n41 8.855
R683 CLK1.n41 CLK1.n40 8.855
R684 CLK1.n279 CLK1.n278 8.855
R685 CLK1.n278 CLK1.n277 8.855
R686 CLK1.n275 CLK1.n274 8.855
R687 CLK1.n274 CLK1.n273 8.855
R688 CLK1.n271 CLK1.n270 8.855
R689 CLK1.n270 CLK1.n269 8.855
R690 CLK1.n266 CLK1.n265 8.855
R691 CLK1.n265 CLK1.n264 8.855
R692 CLK1.n262 CLK1.n261 8.855
R693 CLK1.n261 CLK1.n260 8.855
R694 CLK1.n258 CLK1.n257 8.855
R695 CLK1.n257 CLK1.n256 8.855
R696 CLK1.n254 CLK1.n253 8.855
R697 CLK1.n253 CLK1.n252 8.855
R698 CLK1.n249 CLK1.n248 8.855
R699 CLK1.n248 CLK1.n247 8.855
R700 CLK1.n245 CLK1.n244 8.855
R701 CLK1.n182 CLK1.t32 8.189
R702 CLK1.n188 CLK1.t27 8.189
R703 CLK1.n88 CLK1.t16 8.189
R704 CLK1.n94 CLK1.t18 8.189
R705 CLK1.n36 CLK1.t3 8.189
R706 CLK1.n277 CLK1.t10 8.189
R707 CLK1.n225 CLK1.n45 6.776
R708 CLK1.n148 CLK1.n49 6.776
R709 CLK1.n62 CLK1.n53 6.776
R710 CLK1.n251 CLK1.n44 6.776
R711 CLK1.n242 CLK1.n240 6.312
R712 CLK1.n186 CLK1.n48 4.938
R713 CLK1.n92 CLK1.n52 4.938
R714 CLK1.n43 CLK1.n0 4.938
R715 CLK1.n2 CLK1.n1 4.675
R716 CLK1.n61 CLK1.n60 4.65
R717 CLK1.n66 CLK1.n65 4.65
R718 CLK1.n70 CLK1.n69 4.65
R719 CLK1.n74 CLK1.n73 4.65
R720 CLK1.n78 CLK1.n77 4.65
R721 CLK1.n83 CLK1.n82 4.65
R722 CLK1.n87 CLK1.n86 4.65
R723 CLK1.n91 CLK1.n90 4.65
R724 CLK1.n93 CLK1.n92 4.65
R725 CLK1.n97 CLK1.n96 4.65
R726 CLK1.n101 CLK1.n100 4.65
R727 CLK1.n105 CLK1.n104 4.65
R728 CLK1.n110 CLK1.n109 4.65
R729 CLK1.n114 CLK1.n113 4.65
R730 CLK1.n118 CLK1.n117 4.65
R731 CLK1.n122 CLK1.n121 4.65
R732 CLK1.n126 CLK1.n125 4.65
R733 CLK1.n130 CLK1.n129 4.65
R734 CLK1.n133 CLK1.n132 4.65
R735 CLK1.n135 CLK1.n134 4.65
R736 CLK1.n139 CLK1.n138 4.65
R737 CLK1.n143 CLK1.n142 4.65
R738 CLK1.n147 CLK1.n146 4.65
R739 CLK1.n152 CLK1.n151 4.65
R740 CLK1.n156 CLK1.n155 4.65
R741 CLK1.n160 CLK1.n159 4.65
R742 CLK1.n164 CLK1.n163 4.65
R743 CLK1.n168 CLK1.n167 4.65
R744 CLK1.n172 CLK1.n171 4.65
R745 CLK1.n177 CLK1.n176 4.65
R746 CLK1.n181 CLK1.n180 4.65
R747 CLK1.n185 CLK1.n184 4.65
R748 CLK1.n187 CLK1.n186 4.65
R749 CLK1.n191 CLK1.n190 4.65
R750 CLK1.n195 CLK1.n194 4.65
R751 CLK1.n199 CLK1.n198 4.65
R752 CLK1.n204 CLK1.n203 4.65
R753 CLK1.n208 CLK1.n207 4.65
R754 CLK1.n212 CLK1.n211 4.65
R755 CLK1.n216 CLK1.n215 4.65
R756 CLK1.n220 CLK1.n219 4.65
R757 CLK1.n224 CLK1.n223 4.65
R758 CLK1.n229 CLK1.n228 4.65
R759 CLK1.n233 CLK1.n232 4.65
R760 CLK1.n237 CLK1.n236 4.65
R761 CLK1.n239 CLK1.n238 4.65
R762 CLK1.n6 CLK1.n5 4.65
R763 CLK1.n10 CLK1.n9 4.65
R764 CLK1.n14 CLK1.n13 4.65
R765 CLK1.n18 CLK1.n17 4.65
R766 CLK1.n22 CLK1.n21 4.65
R767 CLK1.n26 CLK1.n25 4.65
R768 CLK1.n31 CLK1.n30 4.65
R769 CLK1.n35 CLK1.n34 4.65
R770 CLK1.n39 CLK1.n38 4.65
R771 CLK1.n43 CLK1.n42 4.65
R772 CLK1.n280 CLK1.n279 4.65
R773 CLK1.n276 CLK1.n275 4.65
R774 CLK1.n272 CLK1.n271 4.65
R775 CLK1.n267 CLK1.n266 4.65
R776 CLK1.n263 CLK1.n262 4.65
R777 CLK1.n259 CLK1.n258 4.65
R778 CLK1.n255 CLK1.n254 4.65
R779 CLK1.n250 CLK1.n249 4.65
R780 CLK1.n246 CLK1.n245 4.65
R781 CLK1.n242 CLK1.n241 4.65
R782 CLK1.n57 CLK1.n56 2.682
R783 CLK1.n240 CLK1.n239 2.325
R784 CLK1.n55 CLK1.n54 1.655
R785 CLK1.n137 CLK1.n136 1.655
R786 CLK1.n4 CLK1.n3 1.655
R787 CLK1.n128 CLK1.n127 1.655
R788 CLK1.n235 CLK1.n234 1.655
R789 CLK1.n244 CLK1.n243 1.655
R790 CLK1.n61 CLK1.n57 1.096
R791 CLK1.n135 CLK1.n133 0.6
R792 CLK1.n240 CLK1 0.131
R793 CLK1.n70 CLK1.n66 0.1
R794 CLK1.n74 CLK1.n70 0.1
R795 CLK1.n78 CLK1.n74 0.1
R796 CLK1.n87 CLK1.n83 0.1
R797 CLK1.n91 CLK1.n87 0.1
R798 CLK1.n92 CLK1.n91 0.1
R799 CLK1.n101 CLK1.n97 0.1
R800 CLK1.n105 CLK1.n101 0.1
R801 CLK1.n114 CLK1.n110 0.1
R802 CLK1.n118 CLK1.n114 0.1
R803 CLK1.n122 CLK1.n118 0.1
R804 CLK1.n126 CLK1.n122 0.1
R805 CLK1.n130 CLK1.n126 0.1
R806 CLK1.n139 CLK1.n135 0.1
R807 CLK1.n143 CLK1.n139 0.1
R808 CLK1.n147 CLK1.n143 0.1
R809 CLK1.n156 CLK1.n152 0.1
R810 CLK1.n160 CLK1.n156 0.1
R811 CLK1.n164 CLK1.n160 0.1
R812 CLK1.n168 CLK1.n164 0.1
R813 CLK1.n172 CLK1.n168 0.1
R814 CLK1.n181 CLK1.n177 0.1
R815 CLK1.n185 CLK1.n181 0.1
R816 CLK1.n186 CLK1.n185 0.1
R817 CLK1.n195 CLK1.n191 0.1
R818 CLK1.n199 CLK1.n195 0.1
R819 CLK1.n208 CLK1.n204 0.1
R820 CLK1.n212 CLK1.n208 0.1
R821 CLK1.n216 CLK1.n212 0.1
R822 CLK1.n220 CLK1.n216 0.1
R823 CLK1.n224 CLK1.n220 0.1
R824 CLK1.n233 CLK1.n229 0.1
R825 CLK1.n237 CLK1.n233 0.1
R826 CLK1.n239 CLK1.n237 0.1
R827 CLK1.n10 CLK1.n6 0.1
R828 CLK1.n14 CLK1.n10 0.1
R829 CLK1.n18 CLK1.n14 0.1
R830 CLK1.n22 CLK1.n18 0.1
R831 CLK1.n26 CLK1.n22 0.1
R832 CLK1.n35 CLK1.n31 0.1
R833 CLK1.n39 CLK1.n35 0.1
R834 CLK1.n43 CLK1.n39 0.1
R835 CLK1.n280 CLK1.n276 0.1
R836 CLK1.n276 CLK1.n272 0.1
R837 CLK1.n267 CLK1.n263 0.1
R838 CLK1.n263 CLK1.n259 0.1
R839 CLK1.n259 CLK1.n255 0.1
R840 CLK1.n250 CLK1.n246 0.1
R841 CLK1.n246 CLK1.n242 0.1
R842 CLK1.n66 CLK1.n62 0.087
R843 CLK1.n255 CLK1.n251 0.087
R844 CLK1.n83 CLK1.n79 0.075
R845 CLK1.n97 CLK1 0.075
R846 CLK1.n106 CLK1.n105 0.075
R847 CLK1.n131 CLK1.n130 0.075
R848 CLK1.n152 CLK1.n148 0.075
R849 CLK1.n177 CLK1.n173 0.075
R850 CLK1.n191 EESPFAL_XOR_v3_0/CLK 0.075
R851 CLK1.n200 CLK1.n199 0.075
R852 CLK1.n225 CLK1.n224 0.075
R853 CLK1.n6 CLK1.n2 0.075
R854 CLK1.n31 CLK1.n27 0.075
R855 EESPFAL_NAND_v3_2/CLK CLK1.n280 0.075
R856 CLK1.n272 CLK1.n268 0.075
R857 CLK1.n79 CLK1.n78 0.025
R858 CLK1.n92 CLK1 0.025
R859 CLK1.n110 CLK1.n106 0.025
R860 CLK1.n133 CLK1.n131 0.025
R861 CLK1.n148 CLK1.n147 0.025
R862 CLK1.n173 CLK1.n172 0.025
R863 CLK1.n186 EESPFAL_XOR_v3_0/CLK 0.025
R864 CLK1.n204 CLK1.n200 0.025
R865 CLK1.n229 CLK1.n225 0.025
R866 CLK1.n27 CLK1.n26 0.025
R867 EESPFAL_NAND_v3_2/CLK CLK1.n43 0.025
R868 CLK1.n268 CLK1.n267 0.025
R869 CLK1.n62 CLK1.n61 0.012
R870 CLK1.n251 CLK1.n250 0.012
R871 x2_bar x2_bar.t0 833.352
R872 EESPFAL_NAND_v3_2/A_bar x2_bar.t1 736.033
R873 EESPFAL_NAND_v3_2/A_bar x2_bar.n0 231.218
R874 x2_bar.n0 x2_bar 22.325
R875 x2_bar.n0 x2_bar 0.025
R876 EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_0/A_bar.t8 1074.82
R877 EESPFAL_NAND_v3_0/A_bar.t6 EESPFAL_NAND_v3_0/A_bar.t7 819.4
R878 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/A_bar.t9 736.033
R879 EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_NAND_v3_0/A_bar.t10 506.1
R880 EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_NAND_v3_0/A_bar.t6 313.3
R881 EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_NAND_v3_0/A_bar.t3 273.936
R882 EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_NAND_v3_1/A 180.175
R883 EESPFAL_XOR_v3_0/OUT_bar EESPFAL_NAND_v3_0/A_bar.n0 161.141
R884 EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_NAND_v3_0/A_bar.n1 128.334
R885 EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_NAND_v3_0/A_bar.n2 105.6
R886 EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_NAND_v3_0/A_bar.t2 81.937
R887 EESPFAL_NAND_v3_0/A_bar.n7 EESPFAL_NAND_v3_0/A_bar.n5 64
R888 EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_NAND_v3_0/A_bar.n3 57.939
R889 EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_NAND_v3_0/A_bar.n4 41.6
R890 EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_NAND_v3_0/A_bar.t4 39.4
R891 EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_NAND_v3_0/A_bar.t5 39.4
R892 EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_NAND_v3_0/A_bar 24.135
R893 EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_NAND_v3_0/A_bar.t1 24
R894 EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_NAND_v3_0/A_bar.t0 24
R895 EESPFAL_NAND_v3_0/A_bar.n7 EESPFAL_NAND_v3_0/A_bar.n6 8.764
R896 EESPFAL_XOR_v3_0/OUT_bar EESPFAL_NAND_v3_0/A_bar.n7 4.65
R897 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/A.t7 1074.82
R898 EESPFAL_NAND_v3_0/A.t10 EESPFAL_NAND_v3_0/A.t9 819.4
R899 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_0/A.t6 736.033
R900 EESPFAL_NAND_v3_0/A.n1 EESPFAL_NAND_v3_0/A.t10 514.133
R901 EESPFAL_NAND_v3_0/A.n1 EESPFAL_NAND_v3_0/A.t8 305.266
R902 EESPFAL_NAND_v3_0/A.n6 EESPFAL_NAND_v3_0/A.n5 192
R903 EESPFAL_NAND_v3_0/A.n4 EESPFAL_NAND_v3_0/A.n3 166.735
R904 EESPFAL_NAND_v3_0/A.n5 EESPFAL_NAND_v3_0/A.n4 105.6
R905 EESPFAL_NAND_v3_0/A.n5 EESPFAL_NAND_v3_0/A.t0 97.937
R906 EESPFAL_NAND_v3_0/A.n6 EESPFAL_NAND_v3_0/A.t1 97.937
R907 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/A.n7 76.565
R908 EESPFAL_NAND_v3_0/A.n2 EESPFAL_NAND_v3_0/A.n1 76
R909 EESPFAL_NAND_v3_0/A.n4 EESPFAL_NAND_v3_0/A.n0 73.937
R910 EESPFAL_NAND_v3_0/A.n4 EESPFAL_NAND_v3_0/A.n2 57.6
R911 EESPFAL_NAND_v3_0/A.n3 EESPFAL_NAND_v3_0/A.t3 39.4
R912 EESPFAL_NAND_v3_0/A.n3 EESPFAL_NAND_v3_0/A.t4 39.4
R913 EESPFAL_NAND_v3_0/A.n7 EESPFAL_NAND_v3_0/A.n6 25.6
R914 EESPFAL_NAND_v3_0/A.n0 EESPFAL_NAND_v3_0/A.t5 24
R915 EESPFAL_NAND_v3_0/A.n0 EESPFAL_NAND_v3_0/A.t2 24
R916 EESPFAL_NAND_v3_0/A.n7 EESPFAL_NAND_v3_1/A_bar 21.729
R917 EESPFAL_NAND_v3_0/A.n2 EESPFAL_XOR_v3_0/OUT 3.2
R918 x1 x1.t0 1026.78
R919 EESPFAL_NAND_v3_2/B_bar x1.t1 527.366
R920 EESPFAL_NAND_v3_2/B_bar x1 340.599
R921 Dis1.n2 Dis1 598.4
R922 Dis1.n1 Dis1.t1 504.5
R923 Dis1.n0 Dis1.t2 504.5
R924 Dis1.n3 Dis1.t3 389.3
R925 Dis1.n2 Dis1.t5 389.3
R926 Dis1.n1 Dis1.t4 389.3
R927 Dis1.n0 Dis1.t0 389.3
R928 EESPFAL_NAND_v3_2/Dis Dis1.n4 241.84
R929 Dis1.n4 EESPFAL_XOR_v3_0/Dis 240.897
R930 Dis1.n3 Dis1.n2 115.2
R931 Dis1.n4 Dis1 3.562
R932 Dis1 Dis1.n1 3.2
R933 EESPFAL_XOR_v3_0/Dis Dis1.n3 3.2
R934 EESPFAL_NAND_v3_2/Dis Dis1.n0 3.2
R935 EESPFAL_NAND_v3_2/A x2.t0 1074.82
R936 x2 x2.t1 687.833
R937 EESPFAL_NAND_v3_2/A x2.n0 267.222
R938 x2.n0 x2 22.914
R939 x2.n0 x2 0.95
R940 Dis3 Dis3.t0 392.5
R941 Dis3.n0 Dis3.t1 389.3
R942 Dis3 Dis3.n0 112
R943 Dis3.n0 Dis3 103.493
R944 s0_bar.t7 s0_bar.t5 819.4
R945 s0_bar.n4 s0_bar.t6 506.1
R946 s0_bar.n4 s0_bar.t7 313.3
R947 s0_bar.n1 s0_bar.t4 187.536
R948 s0_bar.n3 s0_bar.n2 128.334
R949 s0_bar.n1 s0_bar.n0 57.937
R950 s0_bar.n5 s0_bar.n3 57.6
R951 s0_bar.n3 s0_bar.n1 41.6
R952 s0_bar.n2 s0_bar.t0 39.4
R953 s0_bar.n2 s0_bar.t2 39.4
R954 s0_bar.n0 s0_bar.t1 24
R955 s0_bar.n0 s0_bar.t3 24
R956 s0_bar.n5 s0_bar.n4 8.764
R957 s0_bar s0_bar.n5 4.681
R958 s0.t8 s0.t6 819.4
R959 s0.n0 s0.t8 514.133
R960 s0.n0 s0.t7 305.266
R961 s0.n5 s0.n2 166.734
R962 s0.n5 s0.n4 99.2
R963 s0.n4 s0.n3 99.2
R964 s0.n4 s0.t1 97.937
R965 s0.n3 s0.t5 91.537
R966 s0 s0.n0 79.2
R967 s0.n5 s0.n1 73.937
R968 s0 s0.n5 54.4
R969 s0.n2 s0.t4 39.4
R970 s0.n2 s0.t3 39.4
R971 s0.n1 s0.t2 24
R972 s0.n1 s0.t0 24
R973 s0.n3 s0 12.491
R974 CLK3.n27 CLK3.t5 44.338
R975 CLK3.n72 CLK3.t9 44.338
R976 CLK3.n0 CLK3.t3 39.4
R977 CLK3.n0 CLK3.t7 39.4
R978 CLK3.n2 CLK3.t0 30.776
R979 CLK3.n28 CLK3.t4 24.568
R980 CLK3.n73 CLK3.t8 24.568
R981 CLK3.n44 CLK3.t1 24
R982 CLK3.n44 CLK3.t10 24
R983 CLK3.n46 CLK3 10.139
R984 CLK3.n5 CLK3.n4 8.855
R985 CLK3.n9 CLK3.n8 8.855
R986 CLK3.n8 CLK3.n7 8.855
R987 CLK3.n13 CLK3.n12 8.855
R988 CLK3.n12 CLK3.n11 8.855
R989 CLK3.n17 CLK3.n16 8.855
R990 CLK3.n16 CLK3.n15 8.855
R991 CLK3.n21 CLK3.n20 8.855
R992 CLK3.n20 CLK3.n19 8.855
R993 CLK3.n25 CLK3.n24 8.855
R994 CLK3.n24 CLK3.n23 8.855
R995 CLK3.n30 CLK3.n29 8.855
R996 CLK3.n29 CLK3.n28 8.855
R997 CLK3.n34 CLK3.n33 8.855
R998 CLK3.n33 CLK3.n32 8.855
R999 CLK3.n38 CLK3.n37 8.855
R1000 CLK3.n37 CLK3.n36 8.855
R1001 CLK3.n42 CLK3.n41 8.855
R1002 CLK3.n41 CLK3.n40 8.855
R1003 CLK3.n83 CLK3.n82 8.855
R1004 CLK3.n82 CLK3.n81 8.855
R1005 CLK3.n79 CLK3.n78 8.855
R1006 CLK3.n78 CLK3.n77 8.855
R1007 CLK3.n75 CLK3.n74 8.855
R1008 CLK3.n74 CLK3.n73 8.855
R1009 CLK3.n70 CLK3.n69 8.855
R1010 CLK3.n69 CLK3.n68 8.855
R1011 CLK3.n66 CLK3.n65 8.855
R1012 CLK3.n65 CLK3.n64 8.855
R1013 CLK3.n62 CLK3.n61 8.855
R1014 CLK3.n61 CLK3.n60 8.855
R1015 CLK3.n58 CLK3.n57 8.855
R1016 CLK3.n57 CLK3.n56 8.855
R1017 CLK3.n53 CLK3.n52 8.855
R1018 CLK3.n52 CLK3.n51 8.855
R1019 CLK3.n49 CLK3.n48 8.855
R1020 CLK3.n36 CLK3.t2 8.189
R1021 CLK3.n81 CLK3.t6 8.189
R1022 CLK3.n55 CLK3.n44 6.776
R1023 CLK3.n43 CLK3.n0 4.938
R1024 CLK3.n2 CLK3.n1 4.675
R1025 CLK3.n46 CLK3.n45 4.65
R1026 CLK3.n6 CLK3.n5 4.65
R1027 CLK3.n10 CLK3.n9 4.65
R1028 CLK3.n14 CLK3.n13 4.65
R1029 CLK3.n18 CLK3.n17 4.65
R1030 CLK3.n22 CLK3.n21 4.65
R1031 CLK3.n26 CLK3.n25 4.65
R1032 CLK3.n31 CLK3.n30 4.65
R1033 CLK3.n35 CLK3.n34 4.65
R1034 CLK3.n39 CLK3.n38 4.65
R1035 CLK3.n43 CLK3.n42 4.65
R1036 CLK3.n84 CLK3.n83 4.65
R1037 CLK3.n80 CLK3.n79 4.65
R1038 CLK3.n76 CLK3.n75 4.65
R1039 CLK3.n71 CLK3.n70 4.65
R1040 CLK3.n67 CLK3.n66 4.65
R1041 CLK3.n63 CLK3.n62 4.65
R1042 CLK3.n59 CLK3.n58 4.65
R1043 CLK3.n54 CLK3.n53 4.65
R1044 CLK3.n50 CLK3.n49 4.65
R1045 CLK3.n4 CLK3.n3 1.655
R1046 CLK3.n48 CLK3.n47 1.655
R1047 CLK3.n10 CLK3.n6 0.1
R1048 CLK3.n14 CLK3.n10 0.1
R1049 CLK3.n18 CLK3.n14 0.1
R1050 CLK3.n22 CLK3.n18 0.1
R1051 CLK3.n26 CLK3.n22 0.1
R1052 CLK3.n35 CLK3.n31 0.1
R1053 CLK3.n39 CLK3.n35 0.1
R1054 CLK3.n43 CLK3.n39 0.1
R1055 CLK3.n84 CLK3.n80 0.1
R1056 CLK3.n80 CLK3.n76 0.1
R1057 CLK3.n71 CLK3.n67 0.1
R1058 CLK3.n67 CLK3.n63 0.1
R1059 CLK3.n63 CLK3.n59 0.1
R1060 CLK3.n54 CLK3.n50 0.1
R1061 CLK3.n50 CLK3.n46 0.1
R1062 CLK3.n59 CLK3.n55 0.087
R1063 CLK3.n6 CLK3.n2 0.075
R1064 CLK3.n31 CLK3.n27 0.075
R1065 CLK3 CLK3.n84 0.075
R1066 CLK3.n76 CLK3.n72 0.075
R1067 CLK3.n27 CLK3.n26 0.025
R1068 CLK3 CLK3.n43 0.025
R1069 CLK3.n72 CLK3.n71 0.025
R1070 CLK3.n55 CLK3.n54 0.012
R1071 x3.n0 x3.t1 800.452
R1072 x3.n0 x3.t0 787.997
R1073 x3 x3.n0 169.6
R1074 x3_bar.n0 x3_bar.t0 810.772
R1075 x3_bar.n0 x3_bar.t1 694.566
R1076 x3_bar x3_bar.n0 25.6
R1077 EESPFAL_NAND_v3_2/B x1_bar.t1 881.55
R1078 x1_bar x1_bar.t0 479.166
R1079 EESPFAL_NAND_v3_2/B x1_bar.n0 303.264
R1080 x1_bar.n0 x1_bar 23.191
R1081 x1_bar.n0 x1_bar 1.103
R1082 x0.n0 x0.t1 1176.57
R1083 x0.n0 x0.t0 1149.49
R1084 x0 x0.n0 128
R1085 x0_bar.n0 x0_bar.t0 1069.04
R1086 x0_bar.n0 x0_bar.t1 1015.9
R1087 x0_bar x0_bar.n0 89.6
C0 x3 x0_bar 1.68fF
C1 x3 Dis1 0.04fF
C2 x0 x2 0.05fF
C3 a_740_2870# x0_bar 0.00fF
C4 EESPFAL_NAND_v3_0/A_bar s0_bar 0.01fF
C5 x3_bar EESPFAL_NAND_v3_1/B 0.03fF
C6 a_740_2870# Dis1 0.01fF
C7 x1_bar EESPFAL_NOR_v3_0/B 0.00fF
C8 s0 EESPFAL_NAND_v3_0/OUT 0.06fF
C9 EESPFAL_NAND_v3_0/A x1 0.94fF
C10 a_6340_2190# s0 0.00fF
C11 x3_bar EESPFAL_NAND_v3_0/B_bar 0.00fF
C12 x0 CLK1 1.16fF
C13 s0 EESPFAL_NOR_v3_0/B 0.07fF
C14 s0 CLK3 0.86fF
C15 x0_bar a_2000_2190# 0.00fF
C16 Dis1 a_2000_2190# 0.00fF
C17 a_2000_2870# EESPFAL_NAND_v3_0/A_bar 0.01fF
C18 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/B 1.05fF
C19 a_2300_2870# x0_bar 0.00fF
C20 a_2300_2870# Dis1 0.00fF
C21 x0 x1 0.23fF
C22 x0_bar EESPFAL_NAND_v3_1/B_bar 0.01fF
C23 Dis1 EESPFAL_NAND_v3_1/B_bar 0.25fF
C24 EESPFAL_NAND_v3_1/B_bar EESPFAL_NOR_v3_0/B 0.00fF
C25 x0 EESPFAL_NAND_v3_0/B 0.00fF
C26 x2 x0_bar 0.06fF
C27 Dis1 x2 0.07fF
C28 Dis2 EESPFAL_NAND_v3_0/OUT 0.10fF
C29 Dis2 Dis1 0.03fF
C30 CLK2 Dis3 0.32fF
C31 EESPFAL_NAND_v3_1/B x1_bar 0.14fF
C32 x3 EESPFAL_NAND_v3_1/B 0.00fF
C33 Dis3 a_6340_2870# 0.00fF
C34 x2 EESPFAL_NOR_v3_0/B 0.00fF
C35 x2 CLK3 0.00fF
C36 Dis2 EESPFAL_NOR_v3_0/B 0.19fF
C37 CLK1 EESPFAL_NAND_v3_0/OUT 0.00fF
C38 Dis2 CLK3 0.25fF
C39 CLK1 x0_bar 0.51fF
C40 s0 EESPFAL_NAND_v3_0/OUT_bar 0.10fF
C41 Dis1 CLK1 1.95fF
C42 EESPFAL_NAND_v3_0/B_bar x1_bar 0.02fF
C43 x3 EESPFAL_NAND_v3_0/B_bar 0.00fF
C44 s0 EESPFAL_NAND_v3_1/B 0.00fF
C45 s0 a_4320_2190# 0.00fF
C46 x3_bar x2_bar 0.07fF
C47 CLK1 EESPFAL_NOR_v3_0/B 0.02fF
C48 CLK1 CLK3 0.10fF
C49 EESPFAL_NAND_v3_0/OUT x1 0.00fF
C50 a_440_2870# x2_bar 0.00fF
C51 x0_bar x1 2.74fF
C52 s0 EESPFAL_NAND_v3_0/B_bar 0.01fF
C53 Dis1 x1 0.05fF
C54 EESPFAL_NAND_v3_1/B a_2000_2190# 0.01fF
C55 EESPFAL_NOR_v3_0/B_bar x1_bar 0.01fF
C56 CLK3 x1 0.01fF
C57 EESPFAL_NOR_v3_0/B x1 0.00fF
C58 EESPFAL_NAND_v3_0/A Dis3 0.13fF
C59 a_2300_2870# EESPFAL_NAND_v3_1/B 0.00fF
C60 CLK2 a_6340_2870# 0.01fF
C61 EESPFAL_NAND_v3_0/B x0_bar 0.00fF
C62 EESPFAL_NOR_v3_0/B_bar s0 0.68fF
C63 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/OUT 0.07fF
C64 Dis1 EESPFAL_NAND_v3_0/B 0.08fF
C65 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar 0.76fF
C66 a_2300_2870# EESPFAL_NAND_v3_0/B_bar 0.00fF
C67 EESPFAL_NAND_v3_0/B EESPFAL_NOR_v3_0/B 0.02fF
C68 EESPFAL_NAND_v3_0/B CLK3 0.05fF
C69 EESPFAL_NOR_v3_0/B_bar a_2000_2190# 0.00fF
C70 x3_bar a_2000_2870# 0.00fF
C71 Dis2 EESPFAL_NAND_v3_0/OUT_bar 0.24fF
C72 x2 EESPFAL_NAND_v3_1/B 0.05fF
C73 Dis2 EESPFAL_NAND_v3_1/B 0.02fF
C74 EESPFAL_NAND_v3_0/A CLK2 0.83fF
C75 Dis2 a_4320_2190# 0.00fF
C76 a_3060_2870# x1_bar 0.00fF
C77 x2 EESPFAL_NAND_v3_0/B_bar 0.03fF
C78 CLK1 EESPFAL_NAND_v3_0/OUT_bar 0.02fF
C79 EESPFAL_NOR_v3_0/B_bar EESPFAL_NAND_v3_1/B_bar 0.09fF
C80 EESPFAL_NAND_v3_0/A a_6340_2870# 0.01fF
C81 Dis2 EESPFAL_NAND_v3_0/B_bar 0.05fF
C82 CLK1 EESPFAL_NAND_v3_1/B 0.84fF
C83 x2_bar x1_bar 0.65fF
C84 CLK1 a_4320_2190# 0.00fF
C85 x3 x2_bar 1.72fF
C86 a_740_2870# x2_bar 0.00fF
C87 EESPFAL_NAND_v3_0/OUT_bar x1 0.01fF
C88 CLK1 EESPFAL_NAND_v3_0/B_bar 0.79fF
C89 x3_bar EESPFAL_NAND_v3_0/A_bar 0.34fF
C90 EESPFAL_NOR_v3_0/B_bar x2 0.01fF
C91 EESPFAL_NAND_v3_1/B x1 0.00fF
C92 a_440_2870# EESPFAL_NAND_v3_0/A_bar 0.01fF
C93 Dis2 EESPFAL_NOR_v3_0/B_bar 0.26fF
C94 a_4320_2190# x1 0.00fF
C95 EESPFAL_NAND_v3_0/B_bar x1 0.06fF
C96 x2_bar a_2000_2190# 0.00fF
C97 EESPFAL_NOR_v3_0/B_bar CLK1 0.06fF
C98 s0_bar s0 1.61fF
C99 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/OUT_bar 0.17fF
C100 Dis3 EESPFAL_NAND_v3_0/OUT 0.05fF
C101 Dis1 Dis3 0.00fF
C102 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_0/B 0.02fF
C103 EESPFAL_NAND_v3_0/B a_4320_2190# 0.00fF
C104 a_2300_2870# x2_bar 0.00fF
C105 a_2000_2870# x1_bar 0.01fF
C106 a_6340_2190# Dis3 0.00fF
C107 a_2000_2870# x3 0.00fF
C108 EESPFAL_NOR_v3_0/B_bar x1 0.00fF
C109 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar 0.74fF
C110 x2_bar EESPFAL_NAND_v3_1/B_bar 0.07fF
C111 Dis3 CLK3 0.18fF
C112 Dis3 EESPFAL_NOR_v3_0/B 0.03fF
C113 EESPFAL_NAND_v3_0/A x0 0.04fF
C114 x2 a_3060_2870# 0.01fF
C115 Dis2 a_3060_2870# 0.00fF
C116 x2_bar x2 2.88fF
C117 EESPFAL_NOR_v3_0/B_bar EESPFAL_NAND_v3_0/B 0.07fF
C118 Dis2 x2_bar 0.01fF
C119 CLK2 EESPFAL_NAND_v3_0/OUT 0.63fF
C120 Dis1 CLK2 0.06fF
C121 CLK1 a_3060_2870# 0.02fF
C122 EESPFAL_NAND_v3_0/A_bar x1_bar 0.13fF
C123 a_6340_2190# CLK2 0.00fF
C124 x3 EESPFAL_NAND_v3_0/A_bar 0.17fF
C125 a_6340_2870# EESPFAL_NAND_v3_0/OUT 0.01fF
C126 x2_bar CLK1 0.74fF
C127 CLK2 EESPFAL_NOR_v3_0/B 0.58fF
C128 CLK2 CLK3 0.54fF
C129 a_740_2870# EESPFAL_NAND_v3_0/A_bar 0.01fF
C130 Dis2 s0_bar 0.01fF
C131 a_2000_2870# EESPFAL_NAND_v3_1/B_bar 0.00fF
C132 a_3060_2870# x1 0.00fF
C133 a_6340_2870# CLK3 0.00fF
C134 EESPFAL_NAND_v3_0/A_bar s0 0.01fF
C135 a_6340_2870# EESPFAL_NOR_v3_0/B 0.00fF
C136 x2_bar x1 3.72fF
C137 EESPFAL_NAND_v3_0/A_bar a_2000_2190# 0.01fF
C138 Dis3 EESPFAL_NAND_v3_0/OUT_bar 0.12fF
C139 a_2000_2870# x2 0.01fF
C140 EESPFAL_NAND_v3_0/A x0_bar 0.03fF
C141 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/OUT 0.08fF
C142 EESPFAL_NAND_v3_0/B a_3060_2870# 0.00fF
C143 EESPFAL_NAND_v3_0/A Dis1 0.31fF
C144 a_2300_2870# EESPFAL_NAND_v3_0/A_bar 0.02fF
C145 EESPFAL_NAND_v3_0/A a_6340_2190# 0.00fF
C146 a_440_2870# x3_bar 0.00fF
C147 x2_bar EESPFAL_NAND_v3_0/B 0.05fF
C148 Dis3 EESPFAL_NAND_v3_0/B_bar 0.00fF
C149 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_1/B_bar 0.06fF
C150 EESPFAL_NAND_v3_0/A CLK3 0.04fF
C151 EESPFAL_NAND_v3_0/A EESPFAL_NOR_v3_0/B 0.03fF
C152 a_2000_2870# CLK1 0.02fF
C153 x0 x0_bar 4.47fF
C154 x0 Dis1 0.03fF
C155 s0_bar EESPFAL_NAND_v3_0/B 0.02fF
C156 CLK2 EESPFAL_NAND_v3_0/OUT_bar 1.22fF
C157 a_2000_2870# x1 0.00fF
C158 EESPFAL_NOR_v3_0/B_bar Dis3 0.07fF
C159 EESPFAL_NAND_v3_0/A_bar x2 0.20fF
C160 a_6340_2870# EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C161 Dis2 EESPFAL_NAND_v3_0/A_bar 0.05fF
C162 CLK2 EESPFAL_NAND_v3_1/B 0.37fF
C163 CLK2 a_4320_2190# 0.01fF
C164 CLK2 EESPFAL_NAND_v3_0/B_bar 0.06fF
C165 EESPFAL_NAND_v3_0/A_bar CLK1 1.34fF
C166 EESPFAL_NAND_v3_0/A_bar x1 0.10fF
C167 x3_bar x1_bar 0.12fF
C168 EESPFAL_NOR_v3_0/B_bar CLK2 1.24fF
C169 x3_bar x3 3.78fF
C170 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/OUT_bar 0.10fF
C171 a_440_2870# x1_bar 0.01fF
C172 a_440_2870# x3 0.00fF
C173 EESPFAL_NOR_v3_0/B_bar a_6340_2870# 0.01fF
C174 a_740_2870# x3_bar 0.00fF
C175 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/B 0.32fF
C176 EESPFAL_NAND_v3_0/A a_4320_2190# 0.00fF
C177 x2_bar Dis3 0.00fF
C178 Dis1 x0_bar 0.04fF
C179 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/B_bar 0.08fF
C180 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/B 0.38fF
C181 a_6340_2190# EESPFAL_NAND_v3_0/OUT 0.01fF
C182 x3_bar a_2000_2190# 0.00fF
C183 EESPFAL_NAND_v3_0/OUT CLK3 0.70fF
C184 EESPFAL_NAND_v3_0/OUT EESPFAL_NOR_v3_0/B 0.99fF
C185 Dis1 CLK3 0.00fF
C186 Dis1 EESPFAL_NOR_v3_0/B 0.01fF
C187 x0 EESPFAL_NAND_v3_1/B 0.00fF
C188 s0_bar Dis3 0.16fF
C189 a_6340_2190# CLK3 0.01fF
C190 a_6340_2190# EESPFAL_NOR_v3_0/B 0.00fF
C191 EESPFAL_NAND_v3_0/A EESPFAL_NOR_v3_0/B_bar 0.11fF
C192 CLK3 EESPFAL_NOR_v3_0/B 0.46fF
C193 x0 EESPFAL_NAND_v3_0/B_bar 0.00fF
C194 CLK2 a_3060_2870# 0.00fF
C195 x3_bar EESPFAL_NAND_v3_1/B_bar 0.05fF
C196 x2_bar CLK2 0.01fF
C197 x3_bar x2 0.08fF
C198 x3 x1_bar 0.07fF
C199 s0_bar CLK2 0.03fF
C200 a_440_2870# x2 0.01fF
C201 a_740_2870# x1_bar 0.01fF
C202 s0_bar a_6340_2870# 0.00fF
C203 a_740_2870# x3 0.01fF
C204 x3_bar CLK1 0.53fF
C205 EESPFAL_NAND_v3_0/A a_3060_2870# 0.01fF
C206 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar 0.72fF
C207 Dis1 EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C208 a_440_2870# CLK1 0.01fF
C209 a_6340_2190# EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C210 a_2000_2190# x1_bar 0.01fF
C211 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_0/OUT 0.00fF
C212 EESPFAL_NAND_v3_0/A x2_bar 0.18fF
C213 EESPFAL_NAND_v3_1/B x0_bar 0.01fF
C214 Dis1 EESPFAL_NAND_v3_1/B 0.11fF
C215 x3 a_2000_2190# 0.00fF
C216 EESPFAL_NAND_v3_0/A_bar Dis3 0.02fF
C217 x3_bar x1 0.05fF
C218 EESPFAL_NAND_v3_0/OUT_bar CLK3 0.34fF
C219 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_NOR_v3_0/B 0.01fF
C220 EESPFAL_NAND_v3_0/B_bar x0_bar 0.00fF
C221 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/OUT 0.01fF
C222 Dis1 EESPFAL_NAND_v3_0/B_bar 0.15fF
C223 a_2300_2870# x1_bar 0.01fF
C224 a_440_2870# x1 0.00fF
C225 EESPFAL_NAND_v3_1/B CLK3 0.02fF
C226 EESPFAL_NAND_v3_1/B EESPFAL_NOR_v3_0/B 0.08fF
C227 a_2300_2870# x3 0.00fF
C228 a_4320_2190# CLK3 0.01fF
C229 a_4320_2190# EESPFAL_NOR_v3_0/B 0.01fF
C230 EESPFAL_NAND_v3_0/A s0_bar 0.01fF
C231 x1_bar EESPFAL_NAND_v3_1/B_bar 0.21fF
C232 x3 EESPFAL_NAND_v3_1/B_bar 0.01fF
C233 EESPFAL_NAND_v3_0/B_bar EESPFAL_NOR_v3_0/B 0.01fF
C234 EESPFAL_NAND_v3_0/B_bar CLK3 0.02fF
C235 x0 x2_bar 0.03fF
C236 x3_bar EESPFAL_NAND_v3_0/B 0.00fF
C237 a_740_2870# EESPFAL_NAND_v3_1/B_bar 0.00fF
C238 EESPFAL_NOR_v3_0/B_bar Dis1 0.02fF
C239 EESPFAL_NOR_v3_0/B_bar EESPFAL_NAND_v3_0/OUT 0.08fF
C240 a_6340_2190# EESPFAL_NOR_v3_0/B_bar 0.02fF
C241 EESPFAL_NAND_v3_0/A_bar CLK2 0.85fF
C242 x2 x1_bar 5.54fF
C243 x3 x2 0.06fF
C244 a_2000_2870# EESPFAL_NAND_v3_0/A 0.01fF
C245 Dis2 x1_bar 0.00fF
C246 EESPFAL_NOR_v3_0/B_bar CLK3 0.37fF
C247 EESPFAL_NOR_v3_0/B_bar EESPFAL_NOR_v3_0/B 0.88fF
C248 a_2000_2190# EESPFAL_NAND_v3_1/B_bar 0.01fF
C249 a_740_2870# x2 0.01fF
C250 CLK1 x1_bar 1.07fF
C251 x3 CLK1 0.41fF
C252 Dis2 s0 0.02fF
C253 a_2300_2870# EESPFAL_NAND_v3_1/B_bar 0.00fF
C254 a_740_2870# CLK1 0.02fF
C255 x2 a_2000_2190# 0.01fF
C256 a_2000_2870# x0 0.00fF
C257 x1_bar x1 2.20fF
C258 x3 x1 0.07fF
C259 Dis1 a_3060_2870# 0.00fF
C260 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/A_bar 1.56fF
C261 a_2300_2870# x2 0.01fF
C262 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/OUT_bar 0.09fF
C263 a_740_2870# x1 0.00fF
C264 CLK1 a_2000_2190# 0.01fF
C265 x2_bar x0_bar 0.19fF
C266 x2_bar Dis1 0.07fF
C267 x2_bar EESPFAL_NAND_v3_0/OUT 0.00fF
C268 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_0/B_bar 0.02fF
C269 x2 EESPFAL_NAND_v3_1/B_bar 0.07fF
C270 a_3060_2870# CLK3 0.00fF
C271 EESPFAL_NAND_v3_0/B_bar a_4320_2190# 0.00fF
C272 Dis2 EESPFAL_NAND_v3_1/B_bar 0.00fF
C273 EESPFAL_NAND_v3_0/B x1_bar 0.01fF
C274 x3 EESPFAL_NAND_v3_0/B 0.00fF
C275 a_2300_2870# CLK1 0.01fF
C276 x2_bar EESPFAL_NOR_v3_0/B 0.01fF
C277 x2_bar CLK3 0.01fF
C278 a_2000_2190# x1 0.00fF
C279 s0_bar EESPFAL_NAND_v3_0/OUT 0.11fF
C280 EESPFAL_NOR_v3_0/B_bar EESPFAL_NAND_v3_0/OUT_bar 0.26fF
C281 EESPFAL_NAND_v3_0/A_bar x0 0.06fF
C282 CLK1 EESPFAL_NAND_v3_1/B_bar 1.16fF
C283 a_6340_2190# s0_bar 0.00fF
C284 s0 EESPFAL_NAND_v3_0/B 0.02fF
C285 EESPFAL_NOR_v3_0/B_bar EESPFAL_NAND_v3_1/B 0.14fF
C286 EESPFAL_NOR_v3_0/B_bar a_4320_2190# 0.00fF
C287 Dis2 x2 0.00fF
C288 a_2300_2870# x1 0.00fF
C289 s0_bar CLK3 0.86fF
C290 s0_bar EESPFAL_NOR_v3_0/B 0.85fF
C291 EESPFAL_NOR_v3_0/B_bar EESPFAL_NAND_v3_0/B_bar 0.02fF
C292 EESPFAL_NAND_v3_1/B_bar x1 0.09fF
C293 CLK1 x2 1.06fF
C294 Dis2 CLK1 0.08fF
C295 a_2000_2870# x0_bar 0.00fF
C296 a_2000_2870# Dis1 0.00fF
C297 a_2300_2870# EESPFAL_NAND_v3_0/B 0.00fF
C298 x2 x1 0.06fF
C299 Dis2 x1 0.01fF
C300 EESPFAL_NAND_v3_1/B a_3060_2870# 0.00fF
C301 x2_bar EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C302 CLK1 x1 1.72fF
C303 x2_bar EESPFAL_NAND_v3_1/B 0.02fF
C304 x2 EESPFAL_NAND_v3_0/B 0.02fF
C305 EESPFAL_NAND_v3_0/B_bar a_3060_2870# 0.00fF
C306 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/OUT 0.04fF
C307 EESPFAL_NAND_v3_0/A_bar x0_bar 0.07fF
C308 EESPFAL_NAND_v3_0/A_bar Dis1 0.36fF
C309 Dis2 EESPFAL_NAND_v3_0/B 0.05fF
C310 x2_bar EESPFAL_NAND_v3_0/B_bar 0.11fF
C311 s0_bar EESPFAL_NAND_v3_0/OUT_bar 0.05fF
C312 EESPFAL_NAND_v3_0/A_bar CLK3 0.12fF
C313 EESPFAL_NAND_v3_0/A_bar EESPFAL_NOR_v3_0/B 0.09fF
C314 CLK1 EESPFAL_NAND_v3_0/B 0.83fF
C315 s0_bar EESPFAL_NAND_v3_1/B 0.00fF
C316 x3_bar EESPFAL_NAND_v3_0/A 0.09fF
C317 s0_bar a_4320_2190# 0.00fF
C318 EESPFAL_NOR_v3_0/B_bar a_3060_2870# 0.00fF
C319 s0 Dis3 0.15fF
C320 a_440_2870# EESPFAL_NAND_v3_0/A 0.00fF
C321 s0_bar EESPFAL_NAND_v3_0/B_bar 0.00fF
C322 EESPFAL_NOR_v3_0/B_bar x2_bar 0.01fF
C323 EESPFAL_NAND_v3_0/B x1 0.05fF
C324 a_2000_2870# EESPFAL_NAND_v3_1/B 0.00fF
C325 x3_bar x0 0.08fF
C326 CLK2 x1_bar 0.01fF
C327 EESPFAL_NOR_v3_0/B_bar s0_bar 0.15fF
C328 a_440_2870# x0 0.00fF
C329 a_2000_2870# EESPFAL_NAND_v3_0/B_bar 0.00fF
C330 s0 CLK2 0.08fF
C331 s0 a_6340_2870# 0.00fF
C332 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/OUT_bar 0.06fF
C333 CLK2 a_2000_2190# 0.00fF
C334 x2_bar a_3060_2870# 0.00fF
C335 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_1/B 1.25fF
C336 Dis2 Dis3 0.35fF
C337 EESPFAL_NAND_v3_0/A_bar a_4320_2190# 0.01fF
C338 EESPFAL_NAND_v3_0/A x1_bar 0.14fF
C339 x3 EESPFAL_NAND_v3_0/A 0.07fF
C340 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/B_bar 0.35fF
C341 CLK1 Dis3 0.01fF
C342 CLK2 EESPFAL_NAND_v3_1/B_bar 0.03fF
C343 a_740_2870# EESPFAL_NAND_v3_0/A 0.00fF
C344 EESPFAL_NAND_v3_0/A s0 0.01fF
C345 x3_bar x0_bar 0.15fF
C346 x3_bar Dis1 0.11fF
C347 EESPFAL_NAND_v3_0/A_bar EESPFAL_NOR_v3_0/B_bar 0.13fF
C348 Dis3 x1 0.00fF
C349 a_440_2870# x0_bar 0.01fF
C350 x0 x1_bar 0.03fF
C351 a_440_2870# Dis1 0.02fF
C352 x3 x0 0.16fF
C353 x2 CLK2 0.02fF
C354 EESPFAL_NAND_v3_0/A a_2000_2190# 0.00fF
C355 Dis2 CLK2 0.70fF
C356 a_740_2870# x0 0.00fF
C357 Dis2 a_6340_2870# 0.00fF
C358 a_2300_2870# EESPFAL_NAND_v3_0/A 0.01fF
C359 a_2000_2870# x2_bar 0.00fF
C360 CLK1 CLK2 0.24fF
C361 Dis3 EESPFAL_NAND_v3_0/B 0.14fF
C362 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/B_bar 0.26fF
C363 x0 a_2000_2190# 0.00fF
C364 CLK2 x1 0.04fF
C365 EESPFAL_NAND_v3_0/A x2 0.23fF
C366 EESPFAL_NAND_v3_0/A_bar a_3060_2870# 0.00fF
C367 Dis2 EESPFAL_NAND_v3_0/A 0.05fF
C368 x0 EESPFAL_NAND_v3_1/B_bar 0.00fF
C369 EESPFAL_NAND_v3_0/A_bar x2_bar 0.61fF
C370 CLK2 EESPFAL_NAND_v3_0/B 0.44fF
C371 EESPFAL_NAND_v3_0/A CLK1 1.22fF
C372 x0_bar x1_bar 0.05fF
C373 Dis1 x1_bar 0.15fF
C374 a_6340_2190# GND 0.01fF
C375 a_4320_2190# GND 0.01fF
C376 a_2000_2190# GND 0.02fF
C377 s0 GND 0.92fF
C378 s0_bar GND 0.93fF
C379 EESPFAL_NOR_v3_0/B_bar GND 1.57fF
C380 EESPFAL_NOR_v3_0/B GND 1.11fF
C381 EESPFAL_NAND_v3_1/B_bar GND 1.36fF
C382 EESPFAL_NAND_v3_1/B GND 1.33fF
C383 Dis3 GND 1.69fF
C384 a_6340_2870# GND 0.02fF
C385 a_3060_2870# GND 0.02fF
C386 a_2300_2870# GND 0.01fF
C387 a_2000_2870# GND 0.01fF
C388 a_740_2870# GND 0.01fF
C389 a_440_2870# GND 0.01fF
C390 Dis2 GND 3.77fF
C391 x1_bar GND 2.62fF
C392 x2 GND 2.45fF
C393 x2_bar GND 2.49fF
C394 x1 GND 9.10fF
C395 Dis1 GND 5.66fF
C396 EESPFAL_NAND_v3_0/OUT_bar GND 1.73fF
C397 EESPFAL_NAND_v3_0/OUT GND 1.78fF
C398 EESPFAL_NAND_v3_0/B_bar GND 1.17fF
C399 EESPFAL_NAND_v3_0/B GND 1.33fF
C400 x3 GND 2.89fF
C401 x3_bar GND 3.22fF
C402 x0_bar GND 5.16fF
C403 EESPFAL_NAND_v3_0/A_bar GND 2.50fF $ **FLOATING
C404 EESPFAL_NAND_v3_0/A GND 3.08fF $ **FLOATING
C405 x0 GND 4.06fF
C406 CLK3 GND 3.77fF
C407 CLK2 GND 7.28fF
C408 CLK1 GND 11.53fF
C409 x0_bar.t0 GND 0.43fF
C410 x0_bar.t1 GND 0.24fF
C411 x0_bar.n0 GND 2.31fF $ **FLOATING
C412 x0.t0 GND 0.19fF
C413 x0.t1 GND 0.17fF
C414 x0.n0 GND 1.44fF $ **FLOATING
C415 x1_bar.t1 GND 0.30fF
C416 x1_bar.t0 GND 0.12fF
C417 x1_bar.n0 GND 4.66fF $ **FLOATING
C418 EESPFAL_NAND_v3_2/B GND 1.36fF $ **FLOATING
C419 x3_bar.t0 GND 0.34fF
C420 x3_bar.t1 GND 0.12fF
C421 x3_bar.n0 GND 1.13fF $ **FLOATING
C422 x3.t0 GND 0.11fF
C423 x3.t1 GND 0.12fF
C424 x3.n0 GND 1.36fF $ **FLOATING
C425 CLK3.t3 GND 0.02fF
C426 CLK3.t7 GND 0.02fF
C427 CLK3.n0 GND 0.06fF $ **FLOATING
C428 CLK3.t5 GND 0.03fF
C429 CLK3.t0 GND 0.04fF
C430 CLK3.n1 GND 0.07fF $ **FLOATING
C431 CLK3.n2 GND 0.20fF $ **FLOATING
C432 CLK3.n3 GND 0.04fF $ **FLOATING
C433 CLK3.n4 GND 0.02fF $ **FLOATING
C434 CLK3.n5 GND 0.01fF $ **FLOATING
C435 CLK3.n6 GND 0.01fF $ **FLOATING
C436 CLK3.n7 GND 0.03fF $ **FLOATING
C437 CLK3.n8 GND 0.02fF $ **FLOATING
C438 CLK3.n9 GND 0.01fF $ **FLOATING
C439 CLK3.n10 GND 0.02fF $ **FLOATING
C440 CLK3.n11 GND 0.03fF $ **FLOATING
C441 CLK3.n12 GND 0.02fF $ **FLOATING
C442 CLK3.n13 GND 0.01fF $ **FLOATING
C443 CLK3.n14 GND 0.02fF $ **FLOATING
C444 CLK3.n15 GND 0.03fF $ **FLOATING
C445 CLK3.n16 GND 0.02fF $ **FLOATING
C446 CLK3.n17 GND 0.01fF $ **FLOATING
C447 CLK3.n18 GND 0.02fF $ **FLOATING
C448 CLK3.n19 GND 0.07fF $ **FLOATING
C449 CLK3.n20 GND 0.02fF $ **FLOATING
C450 CLK3.n21 GND 0.01fF $ **FLOATING
C451 CLK3.n22 GND 0.02fF $ **FLOATING
C452 CLK3.n23 GND 0.10fF $ **FLOATING
C453 CLK3.n24 GND 0.02fF $ **FLOATING
C454 CLK3.n25 GND 0.01fF $ **FLOATING
C455 CLK3.n26 GND 0.01fF $ **FLOATING
C456 CLK3.n27 GND 0.16fF $ **FLOATING
C457 CLK3.t4 GND 0.05fF
C458 CLK3.n28 GND 0.06fF $ **FLOATING
C459 CLK3.n29 GND 0.02fF $ **FLOATING
C460 CLK3.n30 GND 0.01fF $ **FLOATING
C461 CLK3.n31 GND 0.01fF $ **FLOATING
C462 CLK3.n32 GND 0.09fF $ **FLOATING
C463 CLK3.n33 GND 0.02fF $ **FLOATING
C464 CLK3.n34 GND 0.01fF $ **FLOATING
C465 CLK3.n35 GND 0.02fF $ **FLOATING
C466 CLK3.t2 GND 0.05fF
C467 CLK3.n36 GND 0.05fF $ **FLOATING
C468 CLK3.n37 GND 0.02fF $ **FLOATING
C469 CLK3.n38 GND 0.01fF $ **FLOATING
C470 CLK3.n39 GND 0.02fF $ **FLOATING
C471 CLK3.n40 GND 0.09fF $ **FLOATING
C472 CLK3.n41 GND 0.02fF $ **FLOATING
C473 CLK3.n42 GND 0.01fF $ **FLOATING
C474 CLK3.n43 GND 0.10fF $ **FLOATING
C475 CLK3.t9 GND 0.03fF
C476 CLK3.t1 GND 0.02fF
C477 CLK3.t10 GND 0.02fF
C478 CLK3.n44 GND 0.09fF $ **FLOATING
C479 CLK3.n45 GND 0.07fF $ **FLOATING
C480 CLK3.n46 GND 0.14fF $ **FLOATING
C481 CLK3.n47 GND 0.04fF $ **FLOATING
C482 CLK3.n48 GND 0.02fF $ **FLOATING
C483 CLK3.n49 GND 0.01fF $ **FLOATING
C484 CLK3.n50 GND 0.02fF $ **FLOATING
C485 CLK3.n51 GND 0.03fF $ **FLOATING
C486 CLK3.n52 GND 0.02fF $ **FLOATING
C487 CLK3.n53 GND 0.01fF $ **FLOATING
C488 CLK3.n54 GND 0.01fF $ **FLOATING
C489 CLK3.n55 GND 0.10fF $ **FLOATING
C490 CLK3.n56 GND 0.03fF $ **FLOATING
C491 CLK3.n57 GND 0.02fF $ **FLOATING
C492 CLK3.n58 GND 0.01fF $ **FLOATING
C493 CLK3.n59 GND 0.02fF $ **FLOATING
C494 CLK3.n60 GND 0.03fF $ **FLOATING
C495 CLK3.n61 GND 0.02fF $ **FLOATING
C496 CLK3.n62 GND 0.01fF $ **FLOATING
C497 CLK3.n63 GND 0.02fF $ **FLOATING
C498 CLK3.n64 GND 0.07fF $ **FLOATING
C499 CLK3.n65 GND 0.02fF $ **FLOATING
C500 CLK3.n66 GND 0.01fF $ **FLOATING
C501 CLK3.n67 GND 0.02fF $ **FLOATING
C502 CLK3.n68 GND 0.10fF $ **FLOATING
C503 CLK3.n69 GND 0.02fF $ **FLOATING
C504 CLK3.n70 GND 0.01fF $ **FLOATING
C505 CLK3.n71 GND 0.01fF $ **FLOATING
C506 CLK3.n72 GND 0.16fF $ **FLOATING
C507 CLK3.t8 GND 0.05fF
C508 CLK3.n73 GND 0.06fF $ **FLOATING
C509 CLK3.n74 GND 0.02fF $ **FLOATING
C510 CLK3.n75 GND 0.01fF $ **FLOATING
C511 CLK3.n76 GND 0.01fF $ **FLOATING
C512 CLK3.n77 GND 0.09fF $ **FLOATING
C513 CLK3.n78 GND 0.02fF $ **FLOATING
C514 CLK3.n79 GND 0.01fF $ **FLOATING
C515 CLK3.n80 GND 0.02fF $ **FLOATING
C516 CLK3.t6 GND 0.05fF
C517 CLK3.n81 GND 0.05fF $ **FLOATING
C518 CLK3.n82 GND 0.02fF $ **FLOATING
C519 CLK3.n83 GND 0.01fF $ **FLOATING
C520 CLK3.n84 GND 0.01fF $ **FLOATING
C521 x2.t0 GND 0.33fF
C522 x2.t1 GND 0.17fF
C523 x2.n0 GND 5.02fF $ **FLOATING
C524 EESPFAL_NAND_v3_2/A GND 1.56fF $ **FLOATING
C525 Dis1.t2 GND 0.16fF
C526 Dis1.t0 GND 0.10fF
C527 Dis1.n0 GND 0.41fF $ **FLOATING
C528 Dis1.t1 GND 0.16fF
C529 Dis1.t4 GND 0.10fF
C530 Dis1.n1 GND 0.41fF $ **FLOATING
C531 Dis1.t5 GND 0.10fF
C532 Dis1.n2 GND 0.71fF $ **FLOATING
C533 Dis1.t3 GND 0.10fF
C534 Dis1.n3 GND 0.22fF $ **FLOATING
C535 EESPFAL_XOR_v3_0/Dis GND 0.22fF $ **FLOATING
C536 Dis1.n4 GND 1.13fF $ **FLOATING
C537 EESPFAL_NAND_v3_2/Dis GND 0.22fF $ **FLOATING
C538 x1.t1 GND 0.14fF
C539 x1.t0 GND 0.34fF
C540 EESPFAL_NAND_v3_2/B_bar GND 0.54fF $ **FLOATING
C541 EESPFAL_NAND_v3_0/A.t7 GND 0.08fF
C542 EESPFAL_NAND_v3_0/A.t6 GND 0.04fF
C543 EESPFAL_NAND_v3_1/A_bar GND 0.16fF $ **FLOATING
C544 EESPFAL_NAND_v3_0/A.t1 GND 0.12fF
C545 EESPFAL_NAND_v3_0/A.t0 GND 0.12fF
C546 EESPFAL_NAND_v3_0/A.t5 GND 0.03fF
C547 EESPFAL_NAND_v3_0/A.t2 GND 0.03fF
C548 EESPFAL_NAND_v3_0/A.n0 GND 0.10fF $ **FLOATING
C549 EESPFAL_NAND_v3_0/A.t9 GND 0.04fF
C550 EESPFAL_NAND_v3_0/A.t10 GND 0.04fF
C551 EESPFAL_NAND_v3_0/A.t8 GND 0.02fF
C552 EESPFAL_NAND_v3_0/A.n1 GND 0.04fF $ **FLOATING
C553 EESPFAL_XOR_v3_0/OUT GND 0.01fF $ **FLOATING
C554 EESPFAL_NAND_v3_0/A.n2 GND 0.02fF $ **FLOATING
C555 EESPFAL_NAND_v3_0/A.t3 GND 0.03fF
C556 EESPFAL_NAND_v3_0/A.t4 GND 0.03fF
C557 EESPFAL_NAND_v3_0/A.n3 GND 0.09fF $ **FLOATING
C558 EESPFAL_NAND_v3_0/A.n4 GND 0.13fF $ **FLOATING
C559 EESPFAL_NAND_v3_0/A.n5 GND 0.13fF $ **FLOATING
C560 EESPFAL_NAND_v3_0/A.n6 GND 0.11fF $ **FLOATING
C561 EESPFAL_NAND_v3_0/A.n7 GND 0.36fF $ **FLOATING
C562 EESPFAL_XOR_v3_0/OUT_bar GND 0.12fF $ **FLOATING
C563 EESPFAL_NAND_v3_0/A_bar.t9 GND 0.04fF
C564 EESPFAL_NAND_v3_0/A_bar.t8 GND 0.07fF
C565 EESPFAL_NAND_v3_1/A GND 0.34fF $ **FLOATING
C566 EESPFAL_NAND_v3_0/A_bar.n0 GND 0.63fF $ **FLOATING
C567 EESPFAL_NAND_v3_0/A_bar.t4 GND 0.03fF
C568 EESPFAL_NAND_v3_0/A_bar.t5 GND 0.03fF
C569 EESPFAL_NAND_v3_0/A_bar.n1 GND 0.07fF $ **FLOATING
C570 EESPFAL_NAND_v3_0/A_bar.t2 GND 0.11fF
C571 EESPFAL_NAND_v3_0/A_bar.t3 GND 0.18fF
C572 EESPFAL_NAND_v3_0/A_bar.n2 GND 0.16fF $ **FLOATING
C573 EESPFAL_NAND_v3_0/A_bar.t1 GND 0.03fF
C574 EESPFAL_NAND_v3_0/A_bar.t0 GND 0.03fF
C575 EESPFAL_NAND_v3_0/A_bar.n3 GND 0.08fF $ **FLOATING
C576 EESPFAL_NAND_v3_0/A_bar.n4 GND 0.07fF $ **FLOATING
C577 EESPFAL_NAND_v3_0/A_bar.n5 GND 0.08fF $ **FLOATING
C578 EESPFAL_NAND_v3_0/A_bar.t7 GND 0.04fF
C579 EESPFAL_NAND_v3_0/A_bar.t6 GND 0.03fF
C580 EESPFAL_NAND_v3_0/A_bar.t10 GND 0.03fF
C581 EESPFAL_NAND_v3_0/A_bar.n6 GND 0.04fF $ **FLOATING
C582 EESPFAL_NAND_v3_0/A_bar.n7 GND 0.01fF $ **FLOATING
C583 x2_bar.t1 GND 0.14fF
C584 x2_bar.t0 GND 0.27fF
C585 x2_bar.n0 GND 4.17fF $ **FLOATING
C586 EESPFAL_NAND_v3_2/A_bar GND 0.43fF $ **FLOATING
C587 CLK1.t4 GND 0.02fF
C588 CLK1.t11 GND 0.02fF
C589 CLK1.n0 GND 0.06fF $ **FLOATING
C590 CLK1.t2 GND 0.03fF
C591 CLK1.t25 GND 0.04fF
C592 CLK1.n1 GND 0.07fF $ **FLOATING
C593 CLK1.n2 GND 0.20fF $ **FLOATING
C594 CLK1.n3 GND 0.04fF $ **FLOATING
C595 CLK1.n4 GND 0.02fF $ **FLOATING
C596 CLK1.n5 GND 0.01fF $ **FLOATING
C597 CLK1.n6 GND 0.02fF $ **FLOATING
C598 CLK1.n7 GND 0.03fF $ **FLOATING
C599 CLK1.n8 GND 0.02fF $ **FLOATING
C600 CLK1.n9 GND 0.01fF $ **FLOATING
C601 CLK1.n10 GND 0.02fF $ **FLOATING
C602 CLK1.n11 GND 0.03fF $ **FLOATING
C603 CLK1.n12 GND 0.02fF $ **FLOATING
C604 CLK1.n13 GND 0.01fF $ **FLOATING
C605 CLK1.n14 GND 0.02fF $ **FLOATING
C606 CLK1.n15 GND 0.03fF $ **FLOATING
C607 CLK1.n16 GND 0.02fF $ **FLOATING
C608 CLK1.n17 GND 0.01fF $ **FLOATING
C609 CLK1.n18 GND 0.02fF $ **FLOATING
C610 CLK1.n19 GND 0.08fF $ **FLOATING
C611 CLK1.n20 GND 0.02fF $ **FLOATING
C612 CLK1.n21 GND 0.01fF $ **FLOATING
C613 CLK1.n22 GND 0.02fF $ **FLOATING
C614 CLK1.n23 GND 0.10fF $ **FLOATING
C615 CLK1.n24 GND 0.02fF $ **FLOATING
C616 CLK1.n25 GND 0.01fF $ **FLOATING
C617 CLK1.n26 GND 0.01fF $ **FLOATING
C618 CLK1.n27 GND 0.17fF $ **FLOATING
C619 CLK1.t1 GND 0.05fF
C620 CLK1.n28 GND 0.06fF $ **FLOATING
C621 CLK1.n29 GND 0.02fF $ **FLOATING
C622 CLK1.n30 GND 0.01fF $ **FLOATING
C623 CLK1.n31 GND 0.02fF $ **FLOATING
C624 CLK1.n32 GND 0.09fF $ **FLOATING
C625 CLK1.n33 GND 0.02fF $ **FLOATING
C626 CLK1.n34 GND 0.01fF $ **FLOATING
C627 CLK1.n35 GND 0.02fF $ **FLOATING
C628 CLK1.t3 GND 0.05fF
C629 CLK1.n36 GND 0.05fF $ **FLOATING
C630 CLK1.n37 GND 0.02fF $ **FLOATING
C631 CLK1.n38 GND 0.01fF $ **FLOATING
C632 CLK1.n39 GND 0.02fF $ **FLOATING
C633 CLK1.n40 GND 0.09fF $ **FLOATING
C634 CLK1.n41 GND 0.02fF $ **FLOATING
C635 CLK1.n42 GND 0.01fF $ **FLOATING
C636 CLK1.n43 GND 0.10fF $ **FLOATING
C637 CLK1.t13 GND 0.03fF
C638 CLK1.t6 GND 0.02fF
C639 CLK1.t22 GND 0.02fF
C640 CLK1.n44 GND 0.09fF $ **FLOATING
C641 CLK1.t23 GND 0.02fF
C642 CLK1.t5 GND 0.02fF
C643 CLK1.n45 GND 0.09fF $ **FLOATING
C644 CLK1.t31 GND 0.03fF
C645 EESPFAL_XOR_v3_0/CLK GND 0.01fF $ **FLOATING
C646 CLK1.n46 GND 0.09fF $ **FLOATING
C647 CLK1.n47 GND 0.02fF $ **FLOATING
C648 CLK1.t33 GND 0.02fF
C649 CLK1.t28 GND 0.02fF
C650 CLK1.n48 GND 0.06fF $ **FLOATING
C651 CLK1.t8 GND 0.03fF
C652 CLK1.t26 GND 0.02fF
C653 CLK1.t24 GND 0.02fF
C654 CLK1.n49 GND 0.09fF $ **FLOATING
C655 CLK1.t9 GND 0.04fF
C656 CLK1.t21 GND 0.03fF
C657 CLK1.n50 GND 0.09fF $ **FLOATING
C658 CLK1.n51 GND 0.02fF $ **FLOATING
C659 CLK1.t17 GND 0.02fF
C660 CLK1.t19 GND 0.02fF
C661 CLK1.n52 GND 0.06fF $ **FLOATING
C662 CLK1.t15 GND 0.03fF
C663 CLK1.t29 GND 0.02fF
C664 CLK1.t0 GND 0.02fF
C665 CLK1.n53 GND 0.09fF $ **FLOATING
C666 CLK1.n54 GND 0.04fF $ **FLOATING
C667 CLK1.n55 GND 0.02fF $ **FLOATING
C668 CLK1.n56 GND 0.01fF $ **FLOATING
C669 CLK1.n57 GND 0.07fF $ **FLOATING
C670 CLK1.n58 GND 0.03fF $ **FLOATING
C671 CLK1.n59 GND 0.02fF $ **FLOATING
C672 CLK1.n60 GND 0.01fF $ **FLOATING
C673 CLK1.n61 GND 0.04fF $ **FLOATING
C674 CLK1.n62 GND 0.11fF $ **FLOATING
C675 CLK1.n63 GND 0.03fF $ **FLOATING
C676 CLK1.n64 GND 0.02fF $ **FLOATING
C677 CLK1.n65 GND 0.01fF $ **FLOATING
C678 CLK1.n66 GND 0.02fF $ **FLOATING
C679 CLK1.n67 GND 0.03fF $ **FLOATING
C680 CLK1.n68 GND 0.02fF $ **FLOATING
C681 CLK1.n69 GND 0.01fF $ **FLOATING
C682 CLK1.n70 GND 0.02fF $ **FLOATING
C683 CLK1.n71 GND 0.08fF $ **FLOATING
C684 CLK1.n72 GND 0.02fF $ **FLOATING
C685 CLK1.n73 GND 0.01fF $ **FLOATING
C686 CLK1.n74 GND 0.02fF $ **FLOATING
C687 CLK1.n75 GND 0.10fF $ **FLOATING
C688 CLK1.n76 GND 0.02fF $ **FLOATING
C689 CLK1.n77 GND 0.01fF $ **FLOATING
C690 CLK1.n78 GND 0.01fF $ **FLOATING
C691 CLK1.n79 GND 0.17fF $ **FLOATING
C692 CLK1.t14 GND 0.05fF
C693 CLK1.n80 GND 0.06fF $ **FLOATING
C694 CLK1.n81 GND 0.02fF $ **FLOATING
C695 CLK1.n82 GND 0.01fF $ **FLOATING
C696 CLK1.n83 GND 0.02fF $ **FLOATING
C697 CLK1.n84 GND 0.09fF $ **FLOATING
C698 CLK1.n85 GND 0.02fF $ **FLOATING
C699 CLK1.n86 GND 0.01fF $ **FLOATING
C700 CLK1.n87 GND 0.02fF $ **FLOATING
C701 CLK1.t16 GND 0.05fF
C702 CLK1.n88 GND 0.05fF $ **FLOATING
C703 CLK1.n89 GND 0.02fF $ **FLOATING
C704 CLK1.n90 GND 0.01fF $ **FLOATING
C705 CLK1.n91 GND 0.02fF $ **FLOATING
C706 CLK1.n92 GND 0.10fF $ **FLOATING
C707 CLK1.n93 GND 0.01fF $ **FLOATING
C708 CLK1.t18 GND 0.05fF
C709 CLK1.n94 GND 0.05fF $ **FLOATING
C710 CLK1.n95 GND 0.02fF $ **FLOATING
C711 CLK1.n96 GND 0.01fF $ **FLOATING
C712 CLK1.n97 GND 0.02fF $ **FLOATING
C713 CLK1.n98 GND 0.09fF $ **FLOATING
C714 CLK1.n99 GND 0.02fF $ **FLOATING
C715 CLK1.n100 GND 0.01fF $ **FLOATING
C716 CLK1.n101 GND 0.02fF $ **FLOATING
C717 CLK1.t20 GND 0.05fF
C718 CLK1.n102 GND 0.06fF $ **FLOATING
C719 CLK1.n103 GND 0.02fF $ **FLOATING
C720 CLK1.n104 GND 0.01fF $ **FLOATING
C721 CLK1.n105 GND 0.02fF $ **FLOATING
C722 CLK1.n106 GND 0.17fF $ **FLOATING
C723 CLK1.n107 GND 0.10fF $ **FLOATING
C724 CLK1.n108 GND 0.02fF $ **FLOATING
C725 CLK1.n109 GND 0.01fF $ **FLOATING
C726 CLK1.n110 GND 0.01fF $ **FLOATING
C727 CLK1.n111 GND 0.08fF $ **FLOATING
C728 CLK1.n112 GND 0.02fF $ **FLOATING
C729 CLK1.n113 GND 0.01fF $ **FLOATING
C730 CLK1.n114 GND 0.02fF $ **FLOATING
C731 CLK1.n115 GND 0.03fF $ **FLOATING
C732 CLK1.n116 GND 0.02fF $ **FLOATING
C733 CLK1.n117 GND 0.01fF $ **FLOATING
C734 CLK1.n118 GND 0.02fF $ **FLOATING
C735 CLK1.n119 GND 0.03fF $ **FLOATING
C736 CLK1.n120 GND 0.02fF $ **FLOATING
C737 CLK1.n121 GND 0.01fF $ **FLOATING
C738 CLK1.n122 GND 0.02fF $ **FLOATING
C739 CLK1.n123 GND 0.03fF $ **FLOATING
C740 CLK1.n124 GND 0.02fF $ **FLOATING
C741 CLK1.n125 GND 0.01fF $ **FLOATING
C742 CLK1.n126 GND 0.02fF $ **FLOATING
C743 CLK1.n127 GND 0.04fF $ **FLOATING
C744 CLK1.n128 GND 0.02fF $ **FLOATING
C745 CLK1.n129 GND 0.01fF $ **FLOATING
C746 CLK1.n130 GND 0.02fF $ **FLOATING
C747 CLK1.n131 GND 0.19fF $ **FLOATING
C748 CLK1.n132 GND 0.07fF $ **FLOATING
C749 CLK1.n133 GND 0.05fF $ **FLOATING
C750 CLK1.n134 GND 0.12fF $ **FLOATING
C751 CLK1.n135 GND 0.06fF $ **FLOATING
C752 CLK1.n136 GND 0.04fF $ **FLOATING
C753 CLK1.n137 GND 0.02fF $ **FLOATING
C754 CLK1.n138 GND 0.01fF $ **FLOATING
C755 CLK1.n139 GND 0.02fF $ **FLOATING
C756 CLK1.n140 GND 0.03fF $ **FLOATING
C757 CLK1.n141 GND 0.02fF $ **FLOATING
C758 CLK1.n142 GND 0.01fF $ **FLOATING
C759 CLK1.n143 GND 0.02fF $ **FLOATING
C760 CLK1.n144 GND 0.03fF $ **FLOATING
C761 CLK1.n145 GND 0.02fF $ **FLOATING
C762 CLK1.n146 GND 0.01fF $ **FLOATING
C763 CLK1.n147 GND 0.01fF $ **FLOATING
C764 CLK1.n148 GND 0.11fF $ **FLOATING
C765 CLK1.n149 GND 0.03fF $ **FLOATING
C766 CLK1.n150 GND 0.02fF $ **FLOATING
C767 CLK1.n151 GND 0.01fF $ **FLOATING
C768 CLK1.n152 GND 0.02fF $ **FLOATING
C769 CLK1.n153 GND 0.03fF $ **FLOATING
C770 CLK1.n154 GND 0.02fF $ **FLOATING
C771 CLK1.n155 GND 0.01fF $ **FLOATING
C772 CLK1.n156 GND 0.02fF $ **FLOATING
C773 CLK1.n157 GND 0.03fF $ **FLOATING
C774 CLK1.n158 GND 0.02fF $ **FLOATING
C775 CLK1.n159 GND 0.01fF $ **FLOATING
C776 CLK1.n160 GND 0.02fF $ **FLOATING
C777 CLK1.n161 GND 0.03fF $ **FLOATING
C778 CLK1.n162 GND 0.02fF $ **FLOATING
C779 CLK1.n163 GND 0.01fF $ **FLOATING
C780 CLK1.n164 GND 0.02fF $ **FLOATING
C781 CLK1.n165 GND 0.08fF $ **FLOATING
C782 CLK1.n166 GND 0.02fF $ **FLOATING
C783 CLK1.n167 GND 0.01fF $ **FLOATING
C784 CLK1.n168 GND 0.02fF $ **FLOATING
C785 CLK1.n169 GND 0.10fF $ **FLOATING
C786 CLK1.n170 GND 0.02fF $ **FLOATING
C787 CLK1.n171 GND 0.01fF $ **FLOATING
C788 CLK1.n172 GND 0.01fF $ **FLOATING
C789 CLK1.n173 GND 0.17fF $ **FLOATING
C790 CLK1.t7 GND 0.05fF
C791 CLK1.n174 GND 0.06fF $ **FLOATING
C792 CLK1.n175 GND 0.02fF $ **FLOATING
C793 CLK1.n176 GND 0.01fF $ **FLOATING
C794 CLK1.n177 GND 0.02fF $ **FLOATING
C795 CLK1.n178 GND 0.09fF $ **FLOATING
C796 CLK1.n179 GND 0.02fF $ **FLOATING
C797 CLK1.n180 GND 0.01fF $ **FLOATING
C798 CLK1.n181 GND 0.02fF $ **FLOATING
C799 CLK1.t32 GND 0.05fF
C800 CLK1.n182 GND 0.05fF $ **FLOATING
C801 CLK1.n183 GND 0.02fF $ **FLOATING
C802 CLK1.n184 GND 0.01fF $ **FLOATING
C803 CLK1.n185 GND 0.02fF $ **FLOATING
C804 CLK1.n186 GND 0.10fF $ **FLOATING
C805 CLK1.n187 GND 0.01fF $ **FLOATING
C806 CLK1.t27 GND 0.05fF
C807 CLK1.n188 GND 0.05fF $ **FLOATING
C808 CLK1.n189 GND 0.02fF $ **FLOATING
C809 CLK1.n190 GND 0.01fF $ **FLOATING
C810 CLK1.n191 GND 0.02fF $ **FLOATING
C811 CLK1.n192 GND 0.09fF $ **FLOATING
C812 CLK1.n193 GND 0.02fF $ **FLOATING
C813 CLK1.n194 GND 0.01fF $ **FLOATING
C814 CLK1.n195 GND 0.02fF $ **FLOATING
C815 CLK1.t30 GND 0.05fF
C816 CLK1.n196 GND 0.06fF $ **FLOATING
C817 CLK1.n197 GND 0.02fF $ **FLOATING
C818 CLK1.n198 GND 0.01fF $ **FLOATING
C819 CLK1.n199 GND 0.02fF $ **FLOATING
C820 CLK1.n200 GND 0.17fF $ **FLOATING
C821 CLK1.n201 GND 0.10fF $ **FLOATING
C822 CLK1.n202 GND 0.02fF $ **FLOATING
C823 CLK1.n203 GND 0.01fF $ **FLOATING
C824 CLK1.n204 GND 0.01fF $ **FLOATING
C825 CLK1.n205 GND 0.08fF $ **FLOATING
C826 CLK1.n206 GND 0.02fF $ **FLOATING
C827 CLK1.n207 GND 0.01fF $ **FLOATING
C828 CLK1.n208 GND 0.02fF $ **FLOATING
C829 CLK1.n209 GND 0.03fF $ **FLOATING
C830 CLK1.n210 GND 0.02fF $ **FLOATING
C831 CLK1.n211 GND 0.01fF $ **FLOATING
C832 CLK1.n212 GND 0.02fF $ **FLOATING
C833 CLK1.n213 GND 0.03fF $ **FLOATING
C834 CLK1.n214 GND 0.02fF $ **FLOATING
C835 CLK1.n215 GND 0.01fF $ **FLOATING
C836 CLK1.n216 GND 0.02fF $ **FLOATING
C837 CLK1.n217 GND 0.03fF $ **FLOATING
C838 CLK1.n218 GND 0.02fF $ **FLOATING
C839 CLK1.n219 GND 0.01fF $ **FLOATING
C840 CLK1.n220 GND 0.02fF $ **FLOATING
C841 CLK1.n221 GND 0.03fF $ **FLOATING
C842 CLK1.n222 GND 0.02fF $ **FLOATING
C843 CLK1.n223 GND 0.01fF $ **FLOATING
C844 CLK1.n224 GND 0.02fF $ **FLOATING
C845 CLK1.n225 GND 0.11fF $ **FLOATING
C846 CLK1.n226 GND 0.03fF $ **FLOATING
C847 CLK1.n227 GND 0.02fF $ **FLOATING
C848 CLK1.n228 GND 0.01fF $ **FLOATING
C849 CLK1.n229 GND 0.01fF $ **FLOATING
C850 CLK1.n230 GND 0.03fF $ **FLOATING
C851 CLK1.n231 GND 0.02fF $ **FLOATING
C852 CLK1.n232 GND 0.01fF $ **FLOATING
C853 CLK1.n233 GND 0.02fF $ **FLOATING
C854 CLK1.n234 GND 0.04fF $ **FLOATING
C855 CLK1.n235 GND 0.02fF $ **FLOATING
C856 CLK1.n236 GND 0.01fF $ **FLOATING
C857 CLK1.n237 GND 0.02fF $ **FLOATING
C858 CLK1.n238 GND 0.12fF $ **FLOATING
C859 CLK1.n239 GND 0.03fF $ **FLOATING
C860 CLK1.n240 GND 0.30fF $ **FLOATING
C861 CLK1.n241 GND 0.07fF $ **FLOATING
C862 CLK1.n242 GND 0.20fF $ **FLOATING
C863 CLK1.n243 GND 0.04fF $ **FLOATING
C864 CLK1.n244 GND 0.02fF $ **FLOATING
C865 CLK1.n245 GND 0.01fF $ **FLOATING
C866 CLK1.n246 GND 0.02fF $ **FLOATING
C867 CLK1.n247 GND 0.03fF $ **FLOATING
C868 CLK1.n248 GND 0.02fF $ **FLOATING
C869 CLK1.n249 GND 0.01fF $ **FLOATING
C870 CLK1.n250 GND 0.01fF $ **FLOATING
C871 CLK1.n251 GND 0.11fF $ **FLOATING
C872 CLK1.n252 GND 0.03fF $ **FLOATING
C873 CLK1.n253 GND 0.02fF $ **FLOATING
C874 CLK1.n254 GND 0.01fF $ **FLOATING
C875 CLK1.n255 GND 0.02fF $ **FLOATING
C876 CLK1.n256 GND 0.03fF $ **FLOATING
C877 CLK1.n257 GND 0.02fF $ **FLOATING
C878 CLK1.n258 GND 0.01fF $ **FLOATING
C879 CLK1.n259 GND 0.02fF $ **FLOATING
C880 CLK1.n260 GND 0.08fF $ **FLOATING
C881 CLK1.n261 GND 0.02fF $ **FLOATING
C882 CLK1.n262 GND 0.01fF $ **FLOATING
C883 CLK1.n263 GND 0.02fF $ **FLOATING
C884 CLK1.n264 GND 0.10fF $ **FLOATING
C885 CLK1.n265 GND 0.02fF $ **FLOATING
C886 CLK1.n266 GND 0.01fF $ **FLOATING
C887 CLK1.n267 GND 0.01fF $ **FLOATING
C888 CLK1.n268 GND 0.17fF $ **FLOATING
C889 CLK1.t12 GND 0.05fF
C890 CLK1.n269 GND 0.06fF $ **FLOATING
C891 CLK1.n270 GND 0.02fF $ **FLOATING
C892 CLK1.n271 GND 0.01fF $ **FLOATING
C893 CLK1.n272 GND 0.02fF $ **FLOATING
C894 CLK1.n273 GND 0.09fF $ **FLOATING
C895 CLK1.n274 GND 0.02fF $ **FLOATING
C896 CLK1.n275 GND 0.01fF $ **FLOATING
C897 CLK1.n276 GND 0.02fF $ **FLOATING
C898 CLK1.t10 GND 0.05fF
C899 CLK1.n277 GND 0.05fF $ **FLOATING
C900 CLK1.n278 GND 0.02fF $ **FLOATING
C901 CLK1.n279 GND 0.01fF $ **FLOATING
C902 CLK1.n280 GND 0.02fF $ **FLOATING
C903 EESPFAL_NAND_v3_2/CLK GND 0.01fF $ **FLOATING
C904 CLK2.t3 GND 0.02fF
C905 CLK2.t19 GND 0.02fF
C906 CLK2.n0 GND 0.06fF $ **FLOATING
C907 CLK2.t1 GND 0.03fF
C908 CLK2.t9 GND 0.04fF
C909 CLK2.n1 GND 0.08fF $ **FLOATING
C910 CLK2.n2 GND 0.21fF $ **FLOATING
C911 CLK2.n3 GND 0.04fF $ **FLOATING
C912 CLK2.n4 GND 0.02fF $ **FLOATING
C913 CLK2.n5 GND 0.01fF $ **FLOATING
C914 CLK2.n6 GND 0.02fF $ **FLOATING
C915 CLK2.n7 GND 0.03fF $ **FLOATING
C916 CLK2.n8 GND 0.02fF $ **FLOATING
C917 CLK2.n9 GND 0.01fF $ **FLOATING
C918 CLK2.n10 GND 0.02fF $ **FLOATING
C919 CLK2.n11 GND 0.03fF $ **FLOATING
C920 CLK2.n12 GND 0.02fF $ **FLOATING
C921 CLK2.n13 GND 0.01fF $ **FLOATING
C922 CLK2.n14 GND 0.02fF $ **FLOATING
C923 CLK2.n15 GND 0.03fF $ **FLOATING
C924 CLK2.n16 GND 0.02fF $ **FLOATING
C925 CLK2.n17 GND 0.01fF $ **FLOATING
C926 CLK2.n18 GND 0.02fF $ **FLOATING
C927 CLK2.n19 GND 0.08fF $ **FLOATING
C928 CLK2.n20 GND 0.02fF $ **FLOATING
C929 CLK2.n21 GND 0.01fF $ **FLOATING
C930 CLK2.n22 GND 0.02fF $ **FLOATING
C931 CLK2.n23 GND 0.10fF $ **FLOATING
C932 CLK2.n24 GND 0.02fF $ **FLOATING
C933 CLK2.n25 GND 0.01fF $ **FLOATING
C934 CLK2.n26 GND 0.01fF $ **FLOATING
C935 CLK2.n27 GND 0.17fF $ **FLOATING
C936 CLK2.t0 GND 0.05fF
C937 CLK2.n28 GND 0.06fF $ **FLOATING
C938 CLK2.n29 GND 0.02fF $ **FLOATING
C939 CLK2.n30 GND 0.01fF $ **FLOATING
C940 CLK2.n31 GND 0.02fF $ **FLOATING
C941 CLK2.n32 GND 0.09fF $ **FLOATING
C942 CLK2.n33 GND 0.02fF $ **FLOATING
C943 CLK2.n34 GND 0.01fF $ **FLOATING
C944 CLK2.n35 GND 0.02fF $ **FLOATING
C945 CLK2.t2 GND 0.05fF
C946 CLK2.n36 GND 0.06fF $ **FLOATING
C947 CLK2.n37 GND 0.02fF $ **FLOATING
C948 CLK2.n38 GND 0.01fF $ **FLOATING
C949 CLK2.n39 GND 0.02fF $ **FLOATING
C950 CLK2.n40 GND 0.10fF $ **FLOATING
C951 CLK2.n41 GND 0.02fF $ **FLOATING
C952 CLK2.n42 GND 0.01fF $ **FLOATING
C953 CLK2.n43 GND 0.10fF $ **FLOATING
C954 CLK2.t21 GND 0.03fF
C955 CLK2.n44 GND 0.01fF $ **FLOATING
C956 CLK2.n45 GND 0.02fF $ **FLOATING
C957 CLK2.n46 GND 0.08fF $ **FLOATING
C958 CLK2.t17 GND 0.03fF
C959 CLK2.t15 GND 0.02fF
C960 CLK2.t6 GND 0.02fF
C961 CLK2.n47 GND 0.06fF $ **FLOATING
C962 EESPFAL_NAND_v3_1/CLK GND 0.01fF $ **FLOATING
C963 CLK2.t8 GND 0.03fF
C964 CLK2.t10 GND 0.02fF
C965 CLK2.t4 GND 0.02fF
C966 CLK2.n48 GND 0.09fF $ **FLOATING
C967 CLK2.n49 GND 0.04fF $ **FLOATING
C968 CLK2.n50 GND 0.02fF $ **FLOATING
C969 CLK2.n51 GND 0.01fF $ **FLOATING
C970 CLK2.n52 GND 0.08fF $ **FLOATING
C971 CLK2.n53 GND 0.03fF $ **FLOATING
C972 CLK2.n54 GND 0.02fF $ **FLOATING
C973 CLK2.n55 GND 0.01fF $ **FLOATING
C974 CLK2.n56 GND 0.04fF $ **FLOATING
C975 CLK2.n57 GND 0.11fF $ **FLOATING
C976 CLK2.n58 GND 0.03fF $ **FLOATING
C977 CLK2.n59 GND 0.02fF $ **FLOATING
C978 CLK2.n60 GND 0.01fF $ **FLOATING
C979 CLK2.n61 GND 0.02fF $ **FLOATING
C980 CLK2.n62 GND 0.03fF $ **FLOATING
C981 CLK2.n63 GND 0.02fF $ **FLOATING
C982 CLK2.n64 GND 0.01fF $ **FLOATING
C983 CLK2.n65 GND 0.02fF $ **FLOATING
C984 CLK2.n66 GND 0.08fF $ **FLOATING
C985 CLK2.n67 GND 0.02fF $ **FLOATING
C986 CLK2.n68 GND 0.01fF $ **FLOATING
C987 CLK2.n69 GND 0.02fF $ **FLOATING
C988 CLK2.n70 GND 0.10fF $ **FLOATING
C989 CLK2.n71 GND 0.02fF $ **FLOATING
C990 CLK2.n72 GND 0.01fF $ **FLOATING
C991 CLK2.n73 GND 0.01fF $ **FLOATING
C992 CLK2.n74 GND 0.17fF $ **FLOATING
C993 CLK2.t7 GND 0.05fF
C994 CLK2.n75 GND 0.06fF $ **FLOATING
C995 CLK2.n76 GND 0.02fF $ **FLOATING
C996 CLK2.n77 GND 0.01fF $ **FLOATING
C997 CLK2.n78 GND 0.02fF $ **FLOATING
C998 CLK2.n79 GND 0.09fF $ **FLOATING
C999 CLK2.n80 GND 0.02fF $ **FLOATING
C1000 CLK2.n81 GND 0.01fF $ **FLOATING
C1001 CLK2.n82 GND 0.02fF $ **FLOATING
C1002 CLK2.n83 GND 0.02fF $ **FLOATING
C1003 CLK2.t5 GND 0.05fF
C1004 CLK2.n84 GND 0.06fF $ **FLOATING
C1005 CLK2.n85 GND 0.02fF $ **FLOATING
C1006 CLK2.n86 GND 0.01fF $ **FLOATING
C1007 CLK2.n87 GND 0.10fF $ **FLOATING
C1008 CLK2.n88 GND 0.02fF $ **FLOATING
C1009 CLK2.n89 GND 0.01fF $ **FLOATING
C1010 CLK2.n90 GND 0.10fF $ **FLOATING
C1011 CLK2.t14 GND 0.05fF
C1012 CLK2.n91 GND 0.06fF $ **FLOATING
C1013 CLK2.n92 GND 0.02fF $ **FLOATING
C1014 CLK2.n93 GND 0.01fF $ **FLOATING
C1015 CLK2.n94 GND 0.02fF $ **FLOATING
C1016 CLK2.n95 GND 0.09fF $ **FLOATING
C1017 CLK2.n96 GND 0.02fF $ **FLOATING
C1018 CLK2.n97 GND 0.01fF $ **FLOATING
C1019 CLK2.n98 GND 0.02fF $ **FLOATING
C1020 CLK2.t16 GND 0.05fF
C1021 CLK2.n99 GND 0.06fF $ **FLOATING
C1022 CLK2.n100 GND 0.02fF $ **FLOATING
C1023 CLK2.n101 GND 0.01fF $ **FLOATING
C1024 CLK2.n102 GND 0.02fF $ **FLOATING
C1025 CLK2.n103 GND 0.17fF $ **FLOATING
C1026 CLK2.n104 GND 0.10fF $ **FLOATING
C1027 CLK2.n105 GND 0.02fF $ **FLOATING
C1028 CLK2.n106 GND 0.01fF $ **FLOATING
C1029 CLK2.n107 GND 0.01fF $ **FLOATING
C1030 CLK2.n108 GND 0.08fF $ **FLOATING
C1031 CLK2.n109 GND 0.02fF $ **FLOATING
C1032 CLK2.n110 GND 0.01fF $ **FLOATING
C1033 CLK2.n111 GND 0.02fF $ **FLOATING
C1034 CLK2.n112 GND 0.03fF $ **FLOATING
C1035 CLK2.n113 GND 0.02fF $ **FLOATING
C1036 CLK2.n114 GND 0.01fF $ **FLOATING
C1037 CLK2.n115 GND 0.02fF $ **FLOATING
C1038 CLK2.n116 GND 0.03fF $ **FLOATING
C1039 CLK2.n117 GND 0.02fF $ **FLOATING
C1040 CLK2.n118 GND 0.01fF $ **FLOATING
C1041 CLK2.n119 GND 0.02fF $ **FLOATING
C1042 CLK2.n120 GND 0.03fF $ **FLOATING
C1043 CLK2.n121 GND 0.02fF $ **FLOATING
C1044 CLK2.n122 GND 0.01fF $ **FLOATING
C1045 CLK2.n123 GND 0.02fF $ **FLOATING
C1046 CLK2.n124 GND 0.04fF $ **FLOATING
C1047 CLK2.n125 GND 0.02fF $ **FLOATING
C1048 CLK2.n126 GND 0.01fF $ **FLOATING
C1049 CLK2.n127 GND 0.02fF $ **FLOATING
C1050 CLK2.n128 GND 0.05fF $ **FLOATING
C1051 CLK2.n129 GND 0.02fF $ **FLOATING
C1052 CLK2.n130 GND 0.05fF $ **FLOATING
C1053 CLK2.n131 GND 0.01fF $ **FLOATING
C1054 CLK2.n132 GND 0.01fF $ **FLOATING
C1055 CLK2.t11 GND 0.02fF
C1056 CLK2.n133 GND 0.06fF $ **FLOATING
C1057 CLK2.n134 GND 0.01fF $ **FLOATING
C1058 CLK2.n135 GND 0.09fF $ **FLOATING
C1059 CLK2.n136 GND 0.09fF $ **FLOATING
C1060 CLK2.t12 GND 0.02fF
C1061 CLK2.t13 GND 0.02fF
C1062 CLK2.n137 GND 0.04fF $ **FLOATING
C1063 CLK2.n138 GND 0.01fF $ **FLOATING
C1064 CLK2.n139 GND 0.01fF $ **FLOATING
C1065 CLK2.n140 GND 0.01fF $ **FLOATING
C1066 CLK2.n141 GND 0.05fF $ **FLOATING
C1067 CLK2.n142 GND 0.01fF $ **FLOATING
C1068 CLK2.n143 GND 0.04fF $ **FLOATING
C1069 CLK2.n144 GND 0.02fF $ **FLOATING
C1070 CLK2.n145 GND 0.01fF $ **FLOATING
C1071 CLK2.n146 GND 0.08fF $ **FLOATING
C1072 CLK2.n147 GND 0.04fF $ **FLOATING
C1073 CLK2.n148 GND 0.03fF $ **FLOATING
C1074 CLK2.n149 GND 0.02fF $ **FLOATING
C1075 CLK2.n150 GND 0.01fF $ **FLOATING
C1076 CLK2.n151 GND 0.01fF $ **FLOATING
C1077 CLK2.n152 GND 0.00fF $ **FLOATING
C1078 CLK2.n153 GND 0.03fF $ **FLOATING
C1079 CLK2.n154 GND 0.01fF $ **FLOATING
C1080 CLK2.n155 GND 0.03fF $ **FLOATING
C1081 CLK2.n156 GND 0.02fF $ **FLOATING
C1082 CLK2.n157 GND 0.01fF $ **FLOATING
C1083 CLK2.n158 GND 0.02fF $ **FLOATING
C1084 CLK2.n159 GND 0.03fF $ **FLOATING
C1085 CLK2.n160 GND 0.02fF $ **FLOATING
C1086 CLK2.n161 GND 0.01fF $ **FLOATING
C1087 CLK2.n162 GND 0.02fF $ **FLOATING
C1088 CLK2.n163 GND 0.08fF $ **FLOATING
C1089 CLK2.n164 GND 0.02fF $ **FLOATING
C1090 CLK2.n165 GND 0.01fF $ **FLOATING
C1091 CLK2.n166 GND 0.02fF $ **FLOATING
C1092 CLK2.n167 GND 0.10fF $ **FLOATING
C1093 CLK2.n168 GND 0.02fF $ **FLOATING
C1094 CLK2.n169 GND 0.01fF $ **FLOATING
C1095 CLK2.n170 GND 0.01fF $ **FLOATING
C1096 CLK2.n171 GND 0.17fF $ **FLOATING
C1097 CLK2.t20 GND 0.05fF
C1098 CLK2.n172 GND 0.06fF $ **FLOATING
C1099 CLK2.n173 GND 0.02fF $ **FLOATING
C1100 CLK2.n174 GND 0.01fF $ **FLOATING
C1101 CLK2.n175 GND 0.02fF $ **FLOATING
C1102 CLK2.n176 GND 0.09fF $ **FLOATING
C1103 CLK2.n177 GND 0.02fF $ **FLOATING
C1104 CLK2.n178 GND 0.01fF $ **FLOATING
C1105 CLK2.n179 GND 0.02fF $ **FLOATING
C1106 CLK2.t18 GND 0.05fF
C1107 CLK2.n180 GND 0.06fF $ **FLOATING
C1108 CLK2.n181 GND 0.02fF $ **FLOATING
C1109 CLK2.n182 GND 0.01fF $ **FLOATING
C1110 CLK2.n183 GND 0.02fF $ **FLOATING
C1111 Dis2.t2 GND 0.18fF
C1112 Dis2.t0 GND 0.11fF
C1113 Dis2.n0 GND 0.45fF $ **FLOATING
C1114 Dis2.t3 GND 0.11fF
C1115 Dis2.t1 GND 0.11fF
C1116 EESPFAL_NAND_v3_1/Dis GND -0.30fF $ **FLOATING
C1117 Dis2.n1 GND 0.24fF $ **FLOATING
C1118 Dis2.n2 GND 0.61fF $ **FLOATING
C1119 Dis2.n3 GND 0.80fF $ **FLOATING
.ends

