* NGSPICE file created from EESPFAL_PRESENT80_R1.ext - technology: sky130A

.subckt EESPFAL_XOR_v3 OUT_bar GND OUT A A_bar B B_bar Dis CLK
X0 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X2 a_n840_410# A CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=7.5e+12p ps=3.22e+07u w=1.5e+06u l=150000u
X3 a_n1140_410# B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_420_410# B_bar OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X5 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X7 a_720_410# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar B a_n840_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 CLK A_bar a_n1140_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK A a_420_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 OUT B a_720_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_4in_XOR EESPFAL_XOR_v3_3/GND x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar
+ x2 x2_bar k2 k2_bar x3 x3_bar k3 k3_bar XOR0_bar XOR0 XOR1_bar XOR1 XOR2_bar XOR2
+ XOR3_bar XOR3 CLK Dis
XEESPFAL_XOR_v3_0 XOR0_bar EESPFAL_XOR_v3_3/GND XOR0 x0 x0_bar k0 k0_bar Dis CLK EESPFAL_XOR_v3
XEESPFAL_XOR_v3_1 XOR1_bar EESPFAL_XOR_v3_3/GND XOR1 x1 x1_bar k1 k1_bar Dis CLK EESPFAL_XOR_v3
XEESPFAL_XOR_v3_2 XOR2_bar EESPFAL_XOR_v3_3/GND XOR2 x2 x2_bar k2 k2_bar Dis CLK EESPFAL_XOR_v3
XEESPFAL_XOR_v3_3 XOR3_bar EESPFAL_XOR_v3_3/GND XOR3 x3 x3_bar k3 k3_bar Dis CLK EESPFAL_XOR_v3
.ends

.subckt EESPFAL_3in_NAND_v2 OUT_bar GND OUT A A_bar B B_bar C C_bar Dis CLK
X0 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u M=2
X1 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X2 a_n910_640# B a_n1060_640# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X4 CLK B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=7.7e+12p pd=3.36e+07u as=0p ps=0u w=1.5e+06u l=150000u
X5 CLK A a_n910_640# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n1060_640# C OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 OUT_bar A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 OUT_bar C_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_INV4 OUT GND OUT_bar A A_bar Dis CLK
X0 OUT A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=5.25e+12p ps=2.32e+07u w=1.5e+06u l=150000u
X1 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X2 GND Dis OUT_bar GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X3 GND OUT_bar OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X5 OUT_bar OUT GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 CLK A OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT Dis GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_3in_NOR_v2 OUT_bar GND OUT A A_bar B B_bar C C_bar Dis CLK
X0 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 OUT B CLK GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=7.7e+12p ps=3.36e+07u w=1.5e+06u l=150000u
X2 OUT_bar OUT CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X3 a_n1990_570# B_bar a_n2140_570# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X4 CLK A OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X6 CLK C OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n2140_570# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 OUT_bar C_bar a_n1990_570# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_NAND_v3 OUT_bar GND OUT A A_bar B B_bar Dis CLK
X0 CLK OUT_bar OUT CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X2 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X3 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X5 OUT_bar A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6e+12p ps=2.62e+07u w=1.5e+06u l=150000u
X6 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_501_n414# B OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 CLK A a_501_n414# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 CLK B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_s3 EESPFAL_INV4_2/GND x0 x1 x2 x2_bar x3 x3_bar s3_bar CLK1 s3 Dis1
+ Dis3 CLK3 Dis2 x0_bar CLK2 x1_bar EESPFAL_XOR_v3_0/OUT
XEESPFAL_3in_NAND_v2_0 EESPFAL_INV4_2/A_bar EESPFAL_INV4_2/GND EESPFAL_INV4_2/A x2_bar
+ x2 x0 x0_bar x3 x3_bar Dis1 CLK1 EESPFAL_3in_NAND_v2
XEESPFAL_INV4_0 EESPFAL_INV4_0/OUT EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/B x3_bar x3
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_INV4_1 EESPFAL_INV4_1/OUT EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/B x1 x1_bar
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_INV4_2 EESPFAL_INV4_2/OUT EESPFAL_INV4_2/GND EESPFAL_INV4_2/OUT_bar EESPFAL_INV4_2/A
+ EESPFAL_INV4_2/A_bar Dis2 CLK2 EESPFAL_INV4
XEESPFAL_XOR_v3_0 EESPFAL_NAND_v3_0/A EESPFAL_INV4_2/GND EESPFAL_XOR_v3_0/OUT x1 x1_bar
+ x0 x0_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_XOR_v3_1 EESPFAL_NAND_v3_1/A_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/A x2
+ x2_bar x3 x3_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_3in_NOR_v2_0 s3_bar EESPFAL_INV4_2/GND s3 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar
+ EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_2/OUT_bar EESPFAL_INV4_2/OUT
+ Dis3 CLK3 EESPFAL_3in_NOR_v2
XEESPFAL_NAND_v3_0 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/OUT
+ EESPFAL_NAND_v3_0/A EESPFAL_XOR_v3_0/OUT EESPFAL_NAND_v3_0/B EESPFAL_INV4_0/OUT
+ Dis2 CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_1 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/OUT
+ EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/B EESPFAL_INV4_1/OUT
+ Dis2 CLK2 EESPFAL_NAND_v3
.ends

.subckt EESPFAL_s1 EESPFAL_INV4_2/GND x0 x0_bar x1 x2 x2_bar x3 s1_bar s1 Dis1 Dis3
+ Dis2 x3_bar x1_bar CLK2 CLK1 CLK3
XEESPFAL_3in_NAND_v2_0 EESPFAL_INV4_2/A_bar EESPFAL_INV4_2/GND EESPFAL_INV4_2/A x3_bar
+ x3 x1 x1_bar x0_bar x0 Dis1 CLK1 EESPFAL_3in_NAND_v2
XEESPFAL_INV4_0 EESPFAL_INV4_0/OUT EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/B x3 x3_bar
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_INV4_1 EESPFAL_INV4_1/OUT EESPFAL_INV4_2/GND EESPFAL_INV4_1/OUT_bar x2 x2_bar
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_INV4_2 EESPFAL_INV4_2/OUT EESPFAL_INV4_2/GND EESPFAL_INV4_2/OUT_bar EESPFAL_INV4_2/A
+ EESPFAL_INV4_2/A_bar Dis2 CLK2 EESPFAL_INV4
XEESPFAL_XOR_v3_0 EESPFAL_NAND_v3_0/A EESPFAL_INV4_2/GND EESPFAL_XOR_v3_0/OUT x2 x2_bar
+ x0 x0_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_XOR_v3_1 EESPFAL_NAND_v3_1/A_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/A x1
+ x1_bar x3 x3_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_3in_NOR_v2_0 s1_bar EESPFAL_INV4_2/GND s1 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar
+ EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_2/OUT_bar EESPFAL_INV4_2/OUT
+ Dis3 CLK3 EESPFAL_3in_NOR_v2
XEESPFAL_NAND_v3_0 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/OUT
+ EESPFAL_NAND_v3_0/A EESPFAL_XOR_v3_0/OUT EESPFAL_NAND_v3_0/B EESPFAL_INV4_0/OUT
+ Dis2 CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_1 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/OUT
+ EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/A_bar EESPFAL_INV4_1/OUT EESPFAL_INV4_1/OUT_bar
+ Dis2 CLK2 EESPFAL_NAND_v3
.ends

.subckt EESPFAL_4in_NAND OUT_bar GND OUT A A_bar B B_bar C C_bar D D_bar Dis CLK
X0 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=3.6e+12p pd=1.68e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X1 CLK B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=8.5e+12p pd=3.68e+07u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n1040_180# B a_n1190_180# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 OUT_bar OUT CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u M=2
X4 CLK D_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n1340_180# D OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 OUT_bar A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar C_bar CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X11 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK A a_n1040_180# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_n1190_180# C a_n1340_180# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_s2 EESPFAL_INV4_2/GND x0 x1 x1_bar x2 x2_bar x3 x3_bar Dis1 Dis3 Dis2
+ CLK2 s2_bar s2 x0_bar CLK1 CLK3
XEESPFAL_4in_NAND_0 EESPFAL_INV4_1/A_bar EESPFAL_INV4_2/GND EESPFAL_INV4_1/A x3_bar
+ x3 x1 x1_bar x0 x0_bar x2 x2_bar Dis1 CLK1 EESPFAL_4in_NAND
XEESPFAL_INV4_0 EESPFAL_INV4_0/OUT EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/B x1_bar x1
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_INV4_1 EESPFAL_INV4_1/OUT EESPFAL_INV4_2/GND EESPFAL_INV4_1/OUT_bar EESPFAL_INV4_1/A
+ EESPFAL_INV4_1/A_bar Dis2 CLK2 EESPFAL_INV4
XEESPFAL_INV4_2 EESPFAL_INV4_2/OUT EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/B x2_bar x2
+ Dis1 CLK1 EESPFAL_INV4
XEESPFAL_XOR_v3_0 EESPFAL_NAND_v3_0/A EESPFAL_INV4_2/GND EESPFAL_XOR_v3_0/OUT x3 x3_bar
+ x2 x2_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_XOR_v3_1 EESPFAL_NAND_v3_1/A_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/A x1
+ x1_bar x0 x0_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_3in_NOR_v2_0 s2_bar EESPFAL_INV4_2/GND s2 EESPFAL_NAND_v3_0/OUT EESPFAL_NAND_v3_0/OUT_bar
+ EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_1/OUT_bar EESPFAL_INV4_1/OUT
+ Dis3 CLK3 EESPFAL_3in_NOR_v2
XEESPFAL_NAND_v3_0 EESPFAL_NAND_v3_0/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_0/OUT
+ EESPFAL_NAND_v3_0/A EESPFAL_XOR_v3_0/OUT EESPFAL_NAND_v3_0/B EESPFAL_INV4_0/OUT
+ Dis2 CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_1 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_INV4_2/GND EESPFAL_NAND_v3_1/OUT
+ EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/B EESPFAL_INV4_2/OUT
+ Dis2 CLK2 EESPFAL_NAND_v3
.ends

.subckt EESPFAL_NOR_v3 OUT_bar GND OUT A A_bar B B_bar Dis CLK
X0 a_n1820_550# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=6e+12p ps=2.62e+07u w=1.5e+06u l=150000u
X1 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X2 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u M=2
X3 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X4 OUT_bar B_bar a_n1820_550# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X6 OUT A CLK GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 CLK B OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt EESPFAL_s0 EESPFAL_XOR_v3_0/GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar Dis1
+ Dis2 CLK2 Dis3 s0 s0_bar CLK1 CLK3
XEESPFAL_XOR_v3_0 EESPFAL_NAND_v3_1/A EESPFAL_XOR_v3_0/GND EESPFAL_NAND_v3_0/A x0
+ x0_bar x3 x3_bar Dis1 CLK1 EESPFAL_XOR_v3
XEESPFAL_NOR_v3_0 s0_bar EESPFAL_XOR_v3_0/GND s0 EESPFAL_NOR_v3_0/A EESPFAL_NOR_v3_0/A_bar
+ EESPFAL_NOR_v3_0/B EESPFAL_NOR_v3_0/B_bar Dis3 CLK3 EESPFAL_NOR_v3
XEESPFAL_NOR_v3_1 EESPFAL_NAND_v3_0/B_bar EESPFAL_XOR_v3_0/GND EESPFAL_NAND_v3_0/B
+ x1 x1_bar x2_bar x2 Dis1 CLK1 EESPFAL_NOR_v3
XEESPFAL_NAND_v3_0 EESPFAL_NOR_v3_0/A_bar EESPFAL_XOR_v3_0/GND EESPFAL_NOR_v3_0/A
+ EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar
+ Dis2 CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_1 EESPFAL_NOR_v3_0/B_bar EESPFAL_XOR_v3_0/GND EESPFAL_NOR_v3_0/B
+ EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar
+ Dis2 CLK2 EESPFAL_NAND_v3
XEESPFAL_NAND_v3_2 EESPFAL_NAND_v3_1/B_bar EESPFAL_XOR_v3_0/GND EESPFAL_NAND_v3_1/B
+ x2 x2_bar x1_bar x1 Dis1 CLK1 EESPFAL_NAND_v3
.ends

.subckt EESPFAL_Sbox EESPFAL_s3_0/EESPFAL_INV4_2/GND x0 x1 x2_bar Dis1 CLK1 CLK2 Dis2
+ CLK3 Dis3 s0 s0_bar s1_bar s1 s2 s2_bar s3_bar s3 x3_bar x3 x2 EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT
+ x0_bar x1_bar
XEESPFAL_s3_0 EESPFAL_s3_0/EESPFAL_INV4_2/GND x0 x1 x2 x2_bar x3 x3_bar s3_bar CLK1
+ s3 Dis1 Dis3 CLK3 Dis2 x0_bar CLK2 x1_bar EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT EESPFAL_s3
XEESPFAL_s1_0 EESPFAL_s3_0/EESPFAL_INV4_2/GND x0 x0_bar x1 x2 x2_bar x3 s1_bar s1
+ Dis1 Dis3 Dis2 x3_bar x1_bar CLK2 CLK1 CLK3 EESPFAL_s1
XEESPFAL_s2_0 EESPFAL_s3_0/EESPFAL_INV4_2/GND x0 x1 x1_bar x2 x2_bar x3 x3_bar Dis1
+ Dis3 Dis2 CLK2 s2_bar s2 x0_bar CLK1 CLK3 EESPFAL_s2
XEESPFAL_s0_0 EESPFAL_s3_0/EESPFAL_INV4_2/GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar
+ Dis1 Dis2 CLK2 Dis3 s0 s0_bar CLK1 CLK3 EESPFAL_s0
.ends

.subckt EESPFAL_PRESENT80_R1 GND x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar x2 x2_bar
+ k2 k2_bar x3 x3_bar k3 k3_bar s0 s0_bar CLK0 Dis0 CLK1 Dis1 s2 s2_bar s3_bar s3
+ s1_bar s1 CLK3 Dis2 CLK2 Dis3
XEESPFAL_4in_XOR_0 GND x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar x2 x2_bar k2 k2_bar
+ x3 x3_bar k3 k3_bar EESPFAL_Sbox_0/x0_bar EESPFAL_Sbox_0/x0 EESPFAL_Sbox_0/x1_bar
+ EESPFAL_Sbox_0/x1 EESPFAL_Sbox_0/x2_bar EESPFAL_Sbox_0/x2 EESPFAL_Sbox_0/x3_bar
+ EESPFAL_Sbox_0/x3 CLK0 Dis0 EESPFAL_4in_XOR
XEESPFAL_Sbox_0 GND EESPFAL_Sbox_0/x0 EESPFAL_Sbox_0/x1 EESPFAL_Sbox_0/x2_bar Dis1
+ CLK1 CLK2 Dis2 CLK3 Dis3 s0 s0_bar s1_bar s1 s2 s2_bar s3_bar s3 EESPFAL_Sbox_0/x3_bar
+ EESPFAL_Sbox_0/x3 EESPFAL_Sbox_0/x2 EESPFAL_Sbox_0/EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT
+ EESPFAL_Sbox_0/x0_bar EESPFAL_Sbox_0/x1_bar EESPFAL_Sbox
.ends

