magic
tech sky130A
magscale 1 2
timestamp 1671080676
<< nwell >>
rect 4281 -4985 6583 -3725
<< pwell >>
rect 1892 -6449 4064 -5557
rect 4346 -6481 6518 -5479
rect 6800 -6449 8972 -5557
<< pmoslvt >>
rect 4613 -4850 4713 -3900
rect 4833 -4850 4933 -3900
rect 5053 -4850 5153 -3900
rect 5273 -4850 5373 -3900
rect 5493 -4850 5593 -3900
rect 5713 -4850 5813 -3900
rect 5933 -4850 6033 -3900
rect 6153 -4850 6253 -3900
<< nmoslvt >>
rect 2158 -6423 2258 -5583
rect 2378 -6423 2478 -5583
rect 2598 -6423 2698 -5583
rect 2818 -6423 2918 -5583
rect 3038 -6423 3138 -5583
rect 3258 -6423 3358 -5583
rect 3478 -6423 3578 -5583
rect 3698 -6423 3798 -5583
rect 4612 -6455 4712 -5505
rect 4832 -6455 4932 -5505
rect 5052 -6455 5152 -5505
rect 5272 -6455 5372 -5505
rect 5492 -6455 5592 -5505
rect 5712 -6455 5812 -5505
rect 5932 -6455 6032 -5505
rect 6152 -6455 6252 -5505
rect 7066 -6423 7166 -5583
rect 7286 -6423 7386 -5583
rect 7506 -6423 7606 -5583
rect 7726 -6423 7826 -5583
rect 7946 -6423 8046 -5583
rect 8166 -6423 8266 -5583
rect 8386 -6423 8486 -5583
rect 8606 -6423 8706 -5583
<< ndiff >>
rect 4492 -5555 4612 -5505
rect 2038 -5607 2158 -5583
rect 2038 -5641 2081 -5607
rect 2115 -5641 2158 -5607
rect 2038 -5675 2158 -5641
rect 2038 -5709 2081 -5675
rect 2115 -5709 2158 -5675
rect 2038 -5743 2158 -5709
rect 2038 -5777 2081 -5743
rect 2115 -5777 2158 -5743
rect 2038 -5811 2158 -5777
rect 2038 -5845 2081 -5811
rect 2115 -5845 2158 -5811
rect 2038 -5879 2158 -5845
rect 2038 -5913 2081 -5879
rect 2115 -5913 2158 -5879
rect 2038 -5947 2158 -5913
rect 2038 -5981 2081 -5947
rect 2115 -5981 2158 -5947
rect 2038 -6015 2158 -5981
rect 2038 -6049 2081 -6015
rect 2115 -6049 2158 -6015
rect 2038 -6083 2158 -6049
rect 2038 -6117 2081 -6083
rect 2115 -6117 2158 -6083
rect 2038 -6151 2158 -6117
rect 2038 -6185 2081 -6151
rect 2115 -6185 2158 -6151
rect 2038 -6219 2158 -6185
rect 2038 -6253 2081 -6219
rect 2115 -6253 2158 -6219
rect 2038 -6287 2158 -6253
rect 2038 -6321 2081 -6287
rect 2115 -6321 2158 -6287
rect 2038 -6355 2158 -6321
rect 2038 -6389 2081 -6355
rect 2115 -6389 2158 -6355
rect 2038 -6423 2158 -6389
rect 2258 -5607 2378 -5583
rect 2258 -5641 2301 -5607
rect 2335 -5641 2378 -5607
rect 2258 -5675 2378 -5641
rect 2258 -5709 2301 -5675
rect 2335 -5709 2378 -5675
rect 2258 -5743 2378 -5709
rect 2258 -5777 2301 -5743
rect 2335 -5777 2378 -5743
rect 2258 -5811 2378 -5777
rect 2258 -5845 2301 -5811
rect 2335 -5845 2378 -5811
rect 2258 -5879 2378 -5845
rect 2258 -5913 2301 -5879
rect 2335 -5913 2378 -5879
rect 2258 -5947 2378 -5913
rect 2258 -5981 2301 -5947
rect 2335 -5981 2378 -5947
rect 2258 -6015 2378 -5981
rect 2258 -6049 2301 -6015
rect 2335 -6049 2378 -6015
rect 2258 -6083 2378 -6049
rect 2258 -6117 2301 -6083
rect 2335 -6117 2378 -6083
rect 2258 -6151 2378 -6117
rect 2258 -6185 2301 -6151
rect 2335 -6185 2378 -6151
rect 2258 -6219 2378 -6185
rect 2258 -6253 2301 -6219
rect 2335 -6253 2378 -6219
rect 2258 -6287 2378 -6253
rect 2258 -6321 2301 -6287
rect 2335 -6321 2378 -6287
rect 2258 -6355 2378 -6321
rect 2258 -6389 2301 -6355
rect 2335 -6389 2378 -6355
rect 2258 -6423 2378 -6389
rect 2478 -5607 2598 -5583
rect 2478 -5641 2521 -5607
rect 2555 -5641 2598 -5607
rect 2478 -5675 2598 -5641
rect 2478 -5709 2521 -5675
rect 2555 -5709 2598 -5675
rect 2478 -5743 2598 -5709
rect 2478 -5777 2521 -5743
rect 2555 -5777 2598 -5743
rect 2478 -5811 2598 -5777
rect 2478 -5845 2521 -5811
rect 2555 -5845 2598 -5811
rect 2478 -5879 2598 -5845
rect 2478 -5913 2521 -5879
rect 2555 -5913 2598 -5879
rect 2478 -5947 2598 -5913
rect 2478 -5981 2521 -5947
rect 2555 -5981 2598 -5947
rect 2478 -6015 2598 -5981
rect 2478 -6049 2521 -6015
rect 2555 -6049 2598 -6015
rect 2478 -6083 2598 -6049
rect 2478 -6117 2521 -6083
rect 2555 -6117 2598 -6083
rect 2478 -6151 2598 -6117
rect 2478 -6185 2521 -6151
rect 2555 -6185 2598 -6151
rect 2478 -6219 2598 -6185
rect 2478 -6253 2521 -6219
rect 2555 -6253 2598 -6219
rect 2478 -6287 2598 -6253
rect 2478 -6321 2521 -6287
rect 2555 -6321 2598 -6287
rect 2478 -6355 2598 -6321
rect 2478 -6389 2521 -6355
rect 2555 -6389 2598 -6355
rect 2478 -6423 2598 -6389
rect 2698 -5607 2818 -5583
rect 2698 -5641 2741 -5607
rect 2775 -5641 2818 -5607
rect 2698 -5675 2818 -5641
rect 2698 -5709 2741 -5675
rect 2775 -5709 2818 -5675
rect 2698 -5743 2818 -5709
rect 2698 -5777 2741 -5743
rect 2775 -5777 2818 -5743
rect 2698 -5811 2818 -5777
rect 2698 -5845 2741 -5811
rect 2775 -5845 2818 -5811
rect 2698 -5879 2818 -5845
rect 2698 -5913 2741 -5879
rect 2775 -5913 2818 -5879
rect 2698 -5947 2818 -5913
rect 2698 -5981 2741 -5947
rect 2775 -5981 2818 -5947
rect 2698 -6015 2818 -5981
rect 2698 -6049 2741 -6015
rect 2775 -6049 2818 -6015
rect 2698 -6083 2818 -6049
rect 2698 -6117 2741 -6083
rect 2775 -6117 2818 -6083
rect 2698 -6151 2818 -6117
rect 2698 -6185 2741 -6151
rect 2775 -6185 2818 -6151
rect 2698 -6219 2818 -6185
rect 2698 -6253 2741 -6219
rect 2775 -6253 2818 -6219
rect 2698 -6287 2818 -6253
rect 2698 -6321 2741 -6287
rect 2775 -6321 2818 -6287
rect 2698 -6355 2818 -6321
rect 2698 -6389 2741 -6355
rect 2775 -6389 2818 -6355
rect 2698 -6423 2818 -6389
rect 2918 -5607 3038 -5583
rect 2918 -5641 2961 -5607
rect 2995 -5641 3038 -5607
rect 2918 -5675 3038 -5641
rect 2918 -5709 2961 -5675
rect 2995 -5709 3038 -5675
rect 2918 -5743 3038 -5709
rect 2918 -5777 2961 -5743
rect 2995 -5777 3038 -5743
rect 2918 -5811 3038 -5777
rect 2918 -5845 2961 -5811
rect 2995 -5845 3038 -5811
rect 2918 -5879 3038 -5845
rect 2918 -5913 2961 -5879
rect 2995 -5913 3038 -5879
rect 2918 -5947 3038 -5913
rect 2918 -5981 2961 -5947
rect 2995 -5981 3038 -5947
rect 2918 -6015 3038 -5981
rect 2918 -6049 2961 -6015
rect 2995 -6049 3038 -6015
rect 2918 -6083 3038 -6049
rect 2918 -6117 2961 -6083
rect 2995 -6117 3038 -6083
rect 2918 -6151 3038 -6117
rect 2918 -6185 2961 -6151
rect 2995 -6185 3038 -6151
rect 2918 -6219 3038 -6185
rect 2918 -6253 2961 -6219
rect 2995 -6253 3038 -6219
rect 2918 -6287 3038 -6253
rect 2918 -6321 2961 -6287
rect 2995 -6321 3038 -6287
rect 2918 -6355 3038 -6321
rect 2918 -6389 2961 -6355
rect 2995 -6389 3038 -6355
rect 2918 -6423 3038 -6389
rect 3138 -5607 3258 -5583
rect 3138 -5641 3181 -5607
rect 3215 -5641 3258 -5607
rect 3138 -5675 3258 -5641
rect 3138 -5709 3181 -5675
rect 3215 -5709 3258 -5675
rect 3138 -5743 3258 -5709
rect 3138 -5777 3181 -5743
rect 3215 -5777 3258 -5743
rect 3138 -5811 3258 -5777
rect 3138 -5845 3181 -5811
rect 3215 -5845 3258 -5811
rect 3138 -5879 3258 -5845
rect 3138 -5913 3181 -5879
rect 3215 -5913 3258 -5879
rect 3138 -5947 3258 -5913
rect 3138 -5981 3181 -5947
rect 3215 -5981 3258 -5947
rect 3138 -6015 3258 -5981
rect 3138 -6049 3181 -6015
rect 3215 -6049 3258 -6015
rect 3138 -6083 3258 -6049
rect 3138 -6117 3181 -6083
rect 3215 -6117 3258 -6083
rect 3138 -6151 3258 -6117
rect 3138 -6185 3181 -6151
rect 3215 -6185 3258 -6151
rect 3138 -6219 3258 -6185
rect 3138 -6253 3181 -6219
rect 3215 -6253 3258 -6219
rect 3138 -6287 3258 -6253
rect 3138 -6321 3181 -6287
rect 3215 -6321 3258 -6287
rect 3138 -6355 3258 -6321
rect 3138 -6389 3181 -6355
rect 3215 -6389 3258 -6355
rect 3138 -6423 3258 -6389
rect 3358 -5607 3478 -5583
rect 3358 -5641 3401 -5607
rect 3435 -5641 3478 -5607
rect 3358 -5675 3478 -5641
rect 3358 -5709 3401 -5675
rect 3435 -5709 3478 -5675
rect 3358 -5743 3478 -5709
rect 3358 -5777 3401 -5743
rect 3435 -5777 3478 -5743
rect 3358 -5811 3478 -5777
rect 3358 -5845 3401 -5811
rect 3435 -5845 3478 -5811
rect 3358 -5879 3478 -5845
rect 3358 -5913 3401 -5879
rect 3435 -5913 3478 -5879
rect 3358 -5947 3478 -5913
rect 3358 -5981 3401 -5947
rect 3435 -5981 3478 -5947
rect 3358 -6015 3478 -5981
rect 3358 -6049 3401 -6015
rect 3435 -6049 3478 -6015
rect 3358 -6083 3478 -6049
rect 3358 -6117 3401 -6083
rect 3435 -6117 3478 -6083
rect 3358 -6151 3478 -6117
rect 3358 -6185 3401 -6151
rect 3435 -6185 3478 -6151
rect 3358 -6219 3478 -6185
rect 3358 -6253 3401 -6219
rect 3435 -6253 3478 -6219
rect 3358 -6287 3478 -6253
rect 3358 -6321 3401 -6287
rect 3435 -6321 3478 -6287
rect 3358 -6355 3478 -6321
rect 3358 -6389 3401 -6355
rect 3435 -6389 3478 -6355
rect 3358 -6423 3478 -6389
rect 3578 -5607 3698 -5583
rect 3578 -5641 3621 -5607
rect 3655 -5641 3698 -5607
rect 3578 -5675 3698 -5641
rect 3578 -5709 3621 -5675
rect 3655 -5709 3698 -5675
rect 3578 -5743 3698 -5709
rect 3578 -5777 3621 -5743
rect 3655 -5777 3698 -5743
rect 3578 -5811 3698 -5777
rect 3578 -5845 3621 -5811
rect 3655 -5845 3698 -5811
rect 3578 -5879 3698 -5845
rect 3578 -5913 3621 -5879
rect 3655 -5913 3698 -5879
rect 3578 -5947 3698 -5913
rect 3578 -5981 3621 -5947
rect 3655 -5981 3698 -5947
rect 3578 -6015 3698 -5981
rect 3578 -6049 3621 -6015
rect 3655 -6049 3698 -6015
rect 3578 -6083 3698 -6049
rect 3578 -6117 3621 -6083
rect 3655 -6117 3698 -6083
rect 3578 -6151 3698 -6117
rect 3578 -6185 3621 -6151
rect 3655 -6185 3698 -6151
rect 3578 -6219 3698 -6185
rect 3578 -6253 3621 -6219
rect 3655 -6253 3698 -6219
rect 3578 -6287 3698 -6253
rect 3578 -6321 3621 -6287
rect 3655 -6321 3698 -6287
rect 3578 -6355 3698 -6321
rect 3578 -6389 3621 -6355
rect 3655 -6389 3698 -6355
rect 3578 -6423 3698 -6389
rect 3798 -5607 3918 -5583
rect 3798 -5641 3841 -5607
rect 3875 -5641 3918 -5607
rect 3798 -5675 3918 -5641
rect 3798 -5709 3841 -5675
rect 3875 -5709 3918 -5675
rect 3798 -5743 3918 -5709
rect 3798 -5777 3841 -5743
rect 3875 -5777 3918 -5743
rect 3798 -5811 3918 -5777
rect 3798 -5845 3841 -5811
rect 3875 -5845 3918 -5811
rect 3798 -5879 3918 -5845
rect 3798 -5913 3841 -5879
rect 3875 -5913 3918 -5879
rect 3798 -5947 3918 -5913
rect 3798 -5981 3841 -5947
rect 3875 -5981 3918 -5947
rect 3798 -6015 3918 -5981
rect 3798 -6049 3841 -6015
rect 3875 -6049 3918 -6015
rect 3798 -6083 3918 -6049
rect 3798 -6117 3841 -6083
rect 3875 -6117 3918 -6083
rect 3798 -6151 3918 -6117
rect 3798 -6185 3841 -6151
rect 3875 -6185 3918 -6151
rect 3798 -6219 3918 -6185
rect 3798 -6253 3841 -6219
rect 3875 -6253 3918 -6219
rect 3798 -6287 3918 -6253
rect 3798 -6321 3841 -6287
rect 3875 -6321 3918 -6287
rect 3798 -6355 3918 -6321
rect 3798 -6389 3841 -6355
rect 3875 -6389 3918 -6355
rect 3798 -6423 3918 -6389
rect 4492 -5589 4535 -5555
rect 4569 -5589 4612 -5555
rect 4492 -5623 4612 -5589
rect 4492 -5657 4535 -5623
rect 4569 -5657 4612 -5623
rect 4492 -5691 4612 -5657
rect 4492 -5725 4535 -5691
rect 4569 -5725 4612 -5691
rect 4492 -5759 4612 -5725
rect 4492 -5793 4535 -5759
rect 4569 -5793 4612 -5759
rect 4492 -5827 4612 -5793
rect 4492 -5861 4535 -5827
rect 4569 -5861 4612 -5827
rect 4492 -5895 4612 -5861
rect 4492 -5929 4535 -5895
rect 4569 -5929 4612 -5895
rect 4492 -5963 4612 -5929
rect 4492 -5997 4535 -5963
rect 4569 -5997 4612 -5963
rect 4492 -6031 4612 -5997
rect 4492 -6065 4535 -6031
rect 4569 -6065 4612 -6031
rect 4492 -6099 4612 -6065
rect 4492 -6133 4535 -6099
rect 4569 -6133 4612 -6099
rect 4492 -6167 4612 -6133
rect 4492 -6201 4535 -6167
rect 4569 -6201 4612 -6167
rect 4492 -6235 4612 -6201
rect 4492 -6269 4535 -6235
rect 4569 -6269 4612 -6235
rect 4492 -6303 4612 -6269
rect 4492 -6337 4535 -6303
rect 4569 -6337 4612 -6303
rect 4492 -6371 4612 -6337
rect 4492 -6405 4535 -6371
rect 4569 -6405 4612 -6371
rect 4492 -6455 4612 -6405
rect 4712 -5555 4832 -5505
rect 4712 -5589 4755 -5555
rect 4789 -5589 4832 -5555
rect 4712 -5623 4832 -5589
rect 4712 -5657 4755 -5623
rect 4789 -5657 4832 -5623
rect 4712 -5691 4832 -5657
rect 4712 -5725 4755 -5691
rect 4789 -5725 4832 -5691
rect 4712 -5759 4832 -5725
rect 4712 -5793 4755 -5759
rect 4789 -5793 4832 -5759
rect 4712 -5827 4832 -5793
rect 4712 -5861 4755 -5827
rect 4789 -5861 4832 -5827
rect 4712 -5895 4832 -5861
rect 4712 -5929 4755 -5895
rect 4789 -5929 4832 -5895
rect 4712 -5963 4832 -5929
rect 4712 -5997 4755 -5963
rect 4789 -5997 4832 -5963
rect 4712 -6031 4832 -5997
rect 4712 -6065 4755 -6031
rect 4789 -6065 4832 -6031
rect 4712 -6099 4832 -6065
rect 4712 -6133 4755 -6099
rect 4789 -6133 4832 -6099
rect 4712 -6167 4832 -6133
rect 4712 -6201 4755 -6167
rect 4789 -6201 4832 -6167
rect 4712 -6235 4832 -6201
rect 4712 -6269 4755 -6235
rect 4789 -6269 4832 -6235
rect 4712 -6303 4832 -6269
rect 4712 -6337 4755 -6303
rect 4789 -6337 4832 -6303
rect 4712 -6371 4832 -6337
rect 4712 -6405 4755 -6371
rect 4789 -6405 4832 -6371
rect 4712 -6455 4832 -6405
rect 4932 -5555 5052 -5505
rect 4932 -5589 4975 -5555
rect 5009 -5589 5052 -5555
rect 4932 -5623 5052 -5589
rect 4932 -5657 4975 -5623
rect 5009 -5657 5052 -5623
rect 4932 -5691 5052 -5657
rect 4932 -5725 4975 -5691
rect 5009 -5725 5052 -5691
rect 4932 -5759 5052 -5725
rect 4932 -5793 4975 -5759
rect 5009 -5793 5052 -5759
rect 4932 -5827 5052 -5793
rect 4932 -5861 4975 -5827
rect 5009 -5861 5052 -5827
rect 4932 -5895 5052 -5861
rect 4932 -5929 4975 -5895
rect 5009 -5929 5052 -5895
rect 4932 -5963 5052 -5929
rect 4932 -5997 4975 -5963
rect 5009 -5997 5052 -5963
rect 4932 -6031 5052 -5997
rect 4932 -6065 4975 -6031
rect 5009 -6065 5052 -6031
rect 4932 -6099 5052 -6065
rect 4932 -6133 4975 -6099
rect 5009 -6133 5052 -6099
rect 4932 -6167 5052 -6133
rect 4932 -6201 4975 -6167
rect 5009 -6201 5052 -6167
rect 4932 -6235 5052 -6201
rect 4932 -6269 4975 -6235
rect 5009 -6269 5052 -6235
rect 4932 -6303 5052 -6269
rect 4932 -6337 4975 -6303
rect 5009 -6337 5052 -6303
rect 4932 -6371 5052 -6337
rect 4932 -6405 4975 -6371
rect 5009 -6405 5052 -6371
rect 4932 -6455 5052 -6405
rect 5152 -5555 5272 -5505
rect 5152 -5589 5195 -5555
rect 5229 -5589 5272 -5555
rect 5152 -5623 5272 -5589
rect 5152 -5657 5195 -5623
rect 5229 -5657 5272 -5623
rect 5152 -5691 5272 -5657
rect 5152 -5725 5195 -5691
rect 5229 -5725 5272 -5691
rect 5152 -5759 5272 -5725
rect 5152 -5793 5195 -5759
rect 5229 -5793 5272 -5759
rect 5152 -5827 5272 -5793
rect 5152 -5861 5195 -5827
rect 5229 -5861 5272 -5827
rect 5152 -5895 5272 -5861
rect 5152 -5929 5195 -5895
rect 5229 -5929 5272 -5895
rect 5152 -5963 5272 -5929
rect 5152 -5997 5195 -5963
rect 5229 -5997 5272 -5963
rect 5152 -6031 5272 -5997
rect 5152 -6065 5195 -6031
rect 5229 -6065 5272 -6031
rect 5152 -6099 5272 -6065
rect 5152 -6133 5195 -6099
rect 5229 -6133 5272 -6099
rect 5152 -6167 5272 -6133
rect 5152 -6201 5195 -6167
rect 5229 -6201 5272 -6167
rect 5152 -6235 5272 -6201
rect 5152 -6269 5195 -6235
rect 5229 -6269 5272 -6235
rect 5152 -6303 5272 -6269
rect 5152 -6337 5195 -6303
rect 5229 -6337 5272 -6303
rect 5152 -6371 5272 -6337
rect 5152 -6405 5195 -6371
rect 5229 -6405 5272 -6371
rect 5152 -6455 5272 -6405
rect 5372 -5555 5492 -5505
rect 5372 -5589 5415 -5555
rect 5449 -5589 5492 -5555
rect 5372 -5623 5492 -5589
rect 5372 -5657 5415 -5623
rect 5449 -5657 5492 -5623
rect 5372 -5691 5492 -5657
rect 5372 -5725 5415 -5691
rect 5449 -5725 5492 -5691
rect 5372 -5759 5492 -5725
rect 5372 -5793 5415 -5759
rect 5449 -5793 5492 -5759
rect 5372 -5827 5492 -5793
rect 5372 -5861 5415 -5827
rect 5449 -5861 5492 -5827
rect 5372 -5895 5492 -5861
rect 5372 -5929 5415 -5895
rect 5449 -5929 5492 -5895
rect 5372 -5963 5492 -5929
rect 5372 -5997 5415 -5963
rect 5449 -5997 5492 -5963
rect 5372 -6031 5492 -5997
rect 5372 -6065 5415 -6031
rect 5449 -6065 5492 -6031
rect 5372 -6099 5492 -6065
rect 5372 -6133 5415 -6099
rect 5449 -6133 5492 -6099
rect 5372 -6167 5492 -6133
rect 5372 -6201 5415 -6167
rect 5449 -6201 5492 -6167
rect 5372 -6235 5492 -6201
rect 5372 -6269 5415 -6235
rect 5449 -6269 5492 -6235
rect 5372 -6303 5492 -6269
rect 5372 -6337 5415 -6303
rect 5449 -6337 5492 -6303
rect 5372 -6371 5492 -6337
rect 5372 -6405 5415 -6371
rect 5449 -6405 5492 -6371
rect 5372 -6455 5492 -6405
rect 5592 -5555 5712 -5505
rect 5592 -5589 5635 -5555
rect 5669 -5589 5712 -5555
rect 5592 -5623 5712 -5589
rect 5592 -5657 5635 -5623
rect 5669 -5657 5712 -5623
rect 5592 -5691 5712 -5657
rect 5592 -5725 5635 -5691
rect 5669 -5725 5712 -5691
rect 5592 -5759 5712 -5725
rect 5592 -5793 5635 -5759
rect 5669 -5793 5712 -5759
rect 5592 -5827 5712 -5793
rect 5592 -5861 5635 -5827
rect 5669 -5861 5712 -5827
rect 5592 -5895 5712 -5861
rect 5592 -5929 5635 -5895
rect 5669 -5929 5712 -5895
rect 5592 -5963 5712 -5929
rect 5592 -5997 5635 -5963
rect 5669 -5997 5712 -5963
rect 5592 -6031 5712 -5997
rect 5592 -6065 5635 -6031
rect 5669 -6065 5712 -6031
rect 5592 -6099 5712 -6065
rect 5592 -6133 5635 -6099
rect 5669 -6133 5712 -6099
rect 5592 -6167 5712 -6133
rect 5592 -6201 5635 -6167
rect 5669 -6201 5712 -6167
rect 5592 -6235 5712 -6201
rect 5592 -6269 5635 -6235
rect 5669 -6269 5712 -6235
rect 5592 -6303 5712 -6269
rect 5592 -6337 5635 -6303
rect 5669 -6337 5712 -6303
rect 5592 -6371 5712 -6337
rect 5592 -6405 5635 -6371
rect 5669 -6405 5712 -6371
rect 5592 -6455 5712 -6405
rect 5812 -5555 5932 -5505
rect 5812 -5589 5855 -5555
rect 5889 -5589 5932 -5555
rect 5812 -5623 5932 -5589
rect 5812 -5657 5855 -5623
rect 5889 -5657 5932 -5623
rect 5812 -5691 5932 -5657
rect 5812 -5725 5855 -5691
rect 5889 -5725 5932 -5691
rect 5812 -5759 5932 -5725
rect 5812 -5793 5855 -5759
rect 5889 -5793 5932 -5759
rect 5812 -5827 5932 -5793
rect 5812 -5861 5855 -5827
rect 5889 -5861 5932 -5827
rect 5812 -5895 5932 -5861
rect 5812 -5929 5855 -5895
rect 5889 -5929 5932 -5895
rect 5812 -5963 5932 -5929
rect 5812 -5997 5855 -5963
rect 5889 -5997 5932 -5963
rect 5812 -6031 5932 -5997
rect 5812 -6065 5855 -6031
rect 5889 -6065 5932 -6031
rect 5812 -6099 5932 -6065
rect 5812 -6133 5855 -6099
rect 5889 -6133 5932 -6099
rect 5812 -6167 5932 -6133
rect 5812 -6201 5855 -6167
rect 5889 -6201 5932 -6167
rect 5812 -6235 5932 -6201
rect 5812 -6269 5855 -6235
rect 5889 -6269 5932 -6235
rect 5812 -6303 5932 -6269
rect 5812 -6337 5855 -6303
rect 5889 -6337 5932 -6303
rect 5812 -6371 5932 -6337
rect 5812 -6405 5855 -6371
rect 5889 -6405 5932 -6371
rect 5812 -6455 5932 -6405
rect 6032 -5555 6152 -5505
rect 6032 -5589 6075 -5555
rect 6109 -5589 6152 -5555
rect 6032 -5623 6152 -5589
rect 6032 -5657 6075 -5623
rect 6109 -5657 6152 -5623
rect 6032 -5691 6152 -5657
rect 6032 -5725 6075 -5691
rect 6109 -5725 6152 -5691
rect 6032 -5759 6152 -5725
rect 6032 -5793 6075 -5759
rect 6109 -5793 6152 -5759
rect 6032 -5827 6152 -5793
rect 6032 -5861 6075 -5827
rect 6109 -5861 6152 -5827
rect 6032 -5895 6152 -5861
rect 6032 -5929 6075 -5895
rect 6109 -5929 6152 -5895
rect 6032 -5963 6152 -5929
rect 6032 -5997 6075 -5963
rect 6109 -5997 6152 -5963
rect 6032 -6031 6152 -5997
rect 6032 -6065 6075 -6031
rect 6109 -6065 6152 -6031
rect 6032 -6099 6152 -6065
rect 6032 -6133 6075 -6099
rect 6109 -6133 6152 -6099
rect 6032 -6167 6152 -6133
rect 6032 -6201 6075 -6167
rect 6109 -6201 6152 -6167
rect 6032 -6235 6152 -6201
rect 6032 -6269 6075 -6235
rect 6109 -6269 6152 -6235
rect 6032 -6303 6152 -6269
rect 6032 -6337 6075 -6303
rect 6109 -6337 6152 -6303
rect 6032 -6371 6152 -6337
rect 6032 -6405 6075 -6371
rect 6109 -6405 6152 -6371
rect 6032 -6455 6152 -6405
rect 6252 -5555 6372 -5505
rect 6252 -5589 6295 -5555
rect 6329 -5589 6372 -5555
rect 6252 -5623 6372 -5589
rect 6252 -5657 6295 -5623
rect 6329 -5657 6372 -5623
rect 6252 -5691 6372 -5657
rect 6252 -5725 6295 -5691
rect 6329 -5725 6372 -5691
rect 6252 -5759 6372 -5725
rect 6252 -5793 6295 -5759
rect 6329 -5793 6372 -5759
rect 6252 -5827 6372 -5793
rect 6252 -5861 6295 -5827
rect 6329 -5861 6372 -5827
rect 6252 -5895 6372 -5861
rect 6252 -5929 6295 -5895
rect 6329 -5929 6372 -5895
rect 6252 -5963 6372 -5929
rect 6252 -5997 6295 -5963
rect 6329 -5997 6372 -5963
rect 6252 -6031 6372 -5997
rect 6252 -6065 6295 -6031
rect 6329 -6065 6372 -6031
rect 6252 -6099 6372 -6065
rect 6252 -6133 6295 -6099
rect 6329 -6133 6372 -6099
rect 6252 -6167 6372 -6133
rect 6252 -6201 6295 -6167
rect 6329 -6201 6372 -6167
rect 6252 -6235 6372 -6201
rect 6252 -6269 6295 -6235
rect 6329 -6269 6372 -6235
rect 6252 -6303 6372 -6269
rect 6252 -6337 6295 -6303
rect 6329 -6337 6372 -6303
rect 6252 -6371 6372 -6337
rect 6252 -6405 6295 -6371
rect 6329 -6405 6372 -6371
rect 6252 -6455 6372 -6405
rect 6946 -5607 7066 -5583
rect 6946 -5641 6989 -5607
rect 7023 -5641 7066 -5607
rect 6946 -5675 7066 -5641
rect 6946 -5709 6989 -5675
rect 7023 -5709 7066 -5675
rect 6946 -5743 7066 -5709
rect 6946 -5777 6989 -5743
rect 7023 -5777 7066 -5743
rect 6946 -5811 7066 -5777
rect 6946 -5845 6989 -5811
rect 7023 -5845 7066 -5811
rect 6946 -5879 7066 -5845
rect 6946 -5913 6989 -5879
rect 7023 -5913 7066 -5879
rect 6946 -5947 7066 -5913
rect 6946 -5981 6989 -5947
rect 7023 -5981 7066 -5947
rect 6946 -6015 7066 -5981
rect 6946 -6049 6989 -6015
rect 7023 -6049 7066 -6015
rect 6946 -6083 7066 -6049
rect 6946 -6117 6989 -6083
rect 7023 -6117 7066 -6083
rect 6946 -6151 7066 -6117
rect 6946 -6185 6989 -6151
rect 7023 -6185 7066 -6151
rect 6946 -6219 7066 -6185
rect 6946 -6253 6989 -6219
rect 7023 -6253 7066 -6219
rect 6946 -6287 7066 -6253
rect 6946 -6321 6989 -6287
rect 7023 -6321 7066 -6287
rect 6946 -6355 7066 -6321
rect 6946 -6389 6989 -6355
rect 7023 -6389 7066 -6355
rect 6946 -6423 7066 -6389
rect 7166 -5607 7286 -5583
rect 7166 -5641 7209 -5607
rect 7243 -5641 7286 -5607
rect 7166 -5675 7286 -5641
rect 7166 -5709 7209 -5675
rect 7243 -5709 7286 -5675
rect 7166 -5743 7286 -5709
rect 7166 -5777 7209 -5743
rect 7243 -5777 7286 -5743
rect 7166 -5811 7286 -5777
rect 7166 -5845 7209 -5811
rect 7243 -5845 7286 -5811
rect 7166 -5879 7286 -5845
rect 7166 -5913 7209 -5879
rect 7243 -5913 7286 -5879
rect 7166 -5947 7286 -5913
rect 7166 -5981 7209 -5947
rect 7243 -5981 7286 -5947
rect 7166 -6015 7286 -5981
rect 7166 -6049 7209 -6015
rect 7243 -6049 7286 -6015
rect 7166 -6083 7286 -6049
rect 7166 -6117 7209 -6083
rect 7243 -6117 7286 -6083
rect 7166 -6151 7286 -6117
rect 7166 -6185 7209 -6151
rect 7243 -6185 7286 -6151
rect 7166 -6219 7286 -6185
rect 7166 -6253 7209 -6219
rect 7243 -6253 7286 -6219
rect 7166 -6287 7286 -6253
rect 7166 -6321 7209 -6287
rect 7243 -6321 7286 -6287
rect 7166 -6355 7286 -6321
rect 7166 -6389 7209 -6355
rect 7243 -6389 7286 -6355
rect 7166 -6423 7286 -6389
rect 7386 -5607 7506 -5583
rect 7386 -5641 7429 -5607
rect 7463 -5641 7506 -5607
rect 7386 -5675 7506 -5641
rect 7386 -5709 7429 -5675
rect 7463 -5709 7506 -5675
rect 7386 -5743 7506 -5709
rect 7386 -5777 7429 -5743
rect 7463 -5777 7506 -5743
rect 7386 -5811 7506 -5777
rect 7386 -5845 7429 -5811
rect 7463 -5845 7506 -5811
rect 7386 -5879 7506 -5845
rect 7386 -5913 7429 -5879
rect 7463 -5913 7506 -5879
rect 7386 -5947 7506 -5913
rect 7386 -5981 7429 -5947
rect 7463 -5981 7506 -5947
rect 7386 -6015 7506 -5981
rect 7386 -6049 7429 -6015
rect 7463 -6049 7506 -6015
rect 7386 -6083 7506 -6049
rect 7386 -6117 7429 -6083
rect 7463 -6117 7506 -6083
rect 7386 -6151 7506 -6117
rect 7386 -6185 7429 -6151
rect 7463 -6185 7506 -6151
rect 7386 -6219 7506 -6185
rect 7386 -6253 7429 -6219
rect 7463 -6253 7506 -6219
rect 7386 -6287 7506 -6253
rect 7386 -6321 7429 -6287
rect 7463 -6321 7506 -6287
rect 7386 -6355 7506 -6321
rect 7386 -6389 7429 -6355
rect 7463 -6389 7506 -6355
rect 7386 -6423 7506 -6389
rect 7606 -5607 7726 -5583
rect 7606 -5641 7649 -5607
rect 7683 -5641 7726 -5607
rect 7606 -5675 7726 -5641
rect 7606 -5709 7649 -5675
rect 7683 -5709 7726 -5675
rect 7606 -5743 7726 -5709
rect 7606 -5777 7649 -5743
rect 7683 -5777 7726 -5743
rect 7606 -5811 7726 -5777
rect 7606 -5845 7649 -5811
rect 7683 -5845 7726 -5811
rect 7606 -5879 7726 -5845
rect 7606 -5913 7649 -5879
rect 7683 -5913 7726 -5879
rect 7606 -5947 7726 -5913
rect 7606 -5981 7649 -5947
rect 7683 -5981 7726 -5947
rect 7606 -6015 7726 -5981
rect 7606 -6049 7649 -6015
rect 7683 -6049 7726 -6015
rect 7606 -6083 7726 -6049
rect 7606 -6117 7649 -6083
rect 7683 -6117 7726 -6083
rect 7606 -6151 7726 -6117
rect 7606 -6185 7649 -6151
rect 7683 -6185 7726 -6151
rect 7606 -6219 7726 -6185
rect 7606 -6253 7649 -6219
rect 7683 -6253 7726 -6219
rect 7606 -6287 7726 -6253
rect 7606 -6321 7649 -6287
rect 7683 -6321 7726 -6287
rect 7606 -6355 7726 -6321
rect 7606 -6389 7649 -6355
rect 7683 -6389 7726 -6355
rect 7606 -6423 7726 -6389
rect 7826 -5607 7946 -5583
rect 7826 -5641 7869 -5607
rect 7903 -5641 7946 -5607
rect 7826 -5675 7946 -5641
rect 7826 -5709 7869 -5675
rect 7903 -5709 7946 -5675
rect 7826 -5743 7946 -5709
rect 7826 -5777 7869 -5743
rect 7903 -5777 7946 -5743
rect 7826 -5811 7946 -5777
rect 7826 -5845 7869 -5811
rect 7903 -5845 7946 -5811
rect 7826 -5879 7946 -5845
rect 7826 -5913 7869 -5879
rect 7903 -5913 7946 -5879
rect 7826 -5947 7946 -5913
rect 7826 -5981 7869 -5947
rect 7903 -5981 7946 -5947
rect 7826 -6015 7946 -5981
rect 7826 -6049 7869 -6015
rect 7903 -6049 7946 -6015
rect 7826 -6083 7946 -6049
rect 7826 -6117 7869 -6083
rect 7903 -6117 7946 -6083
rect 7826 -6151 7946 -6117
rect 7826 -6185 7869 -6151
rect 7903 -6185 7946 -6151
rect 7826 -6219 7946 -6185
rect 7826 -6253 7869 -6219
rect 7903 -6253 7946 -6219
rect 7826 -6287 7946 -6253
rect 7826 -6321 7869 -6287
rect 7903 -6321 7946 -6287
rect 7826 -6355 7946 -6321
rect 7826 -6389 7869 -6355
rect 7903 -6389 7946 -6355
rect 7826 -6423 7946 -6389
rect 8046 -5607 8166 -5583
rect 8046 -5641 8089 -5607
rect 8123 -5641 8166 -5607
rect 8046 -5675 8166 -5641
rect 8046 -5709 8089 -5675
rect 8123 -5709 8166 -5675
rect 8046 -5743 8166 -5709
rect 8046 -5777 8089 -5743
rect 8123 -5777 8166 -5743
rect 8046 -5811 8166 -5777
rect 8046 -5845 8089 -5811
rect 8123 -5845 8166 -5811
rect 8046 -5879 8166 -5845
rect 8046 -5913 8089 -5879
rect 8123 -5913 8166 -5879
rect 8046 -5947 8166 -5913
rect 8046 -5981 8089 -5947
rect 8123 -5981 8166 -5947
rect 8046 -6015 8166 -5981
rect 8046 -6049 8089 -6015
rect 8123 -6049 8166 -6015
rect 8046 -6083 8166 -6049
rect 8046 -6117 8089 -6083
rect 8123 -6117 8166 -6083
rect 8046 -6151 8166 -6117
rect 8046 -6185 8089 -6151
rect 8123 -6185 8166 -6151
rect 8046 -6219 8166 -6185
rect 8046 -6253 8089 -6219
rect 8123 -6253 8166 -6219
rect 8046 -6287 8166 -6253
rect 8046 -6321 8089 -6287
rect 8123 -6321 8166 -6287
rect 8046 -6355 8166 -6321
rect 8046 -6389 8089 -6355
rect 8123 -6389 8166 -6355
rect 8046 -6423 8166 -6389
rect 8266 -5607 8386 -5583
rect 8266 -5641 8309 -5607
rect 8343 -5641 8386 -5607
rect 8266 -5675 8386 -5641
rect 8266 -5709 8309 -5675
rect 8343 -5709 8386 -5675
rect 8266 -5743 8386 -5709
rect 8266 -5777 8309 -5743
rect 8343 -5777 8386 -5743
rect 8266 -5811 8386 -5777
rect 8266 -5845 8309 -5811
rect 8343 -5845 8386 -5811
rect 8266 -5879 8386 -5845
rect 8266 -5913 8309 -5879
rect 8343 -5913 8386 -5879
rect 8266 -5947 8386 -5913
rect 8266 -5981 8309 -5947
rect 8343 -5981 8386 -5947
rect 8266 -6015 8386 -5981
rect 8266 -6049 8309 -6015
rect 8343 -6049 8386 -6015
rect 8266 -6083 8386 -6049
rect 8266 -6117 8309 -6083
rect 8343 -6117 8386 -6083
rect 8266 -6151 8386 -6117
rect 8266 -6185 8309 -6151
rect 8343 -6185 8386 -6151
rect 8266 -6219 8386 -6185
rect 8266 -6253 8309 -6219
rect 8343 -6253 8386 -6219
rect 8266 -6287 8386 -6253
rect 8266 -6321 8309 -6287
rect 8343 -6321 8386 -6287
rect 8266 -6355 8386 -6321
rect 8266 -6389 8309 -6355
rect 8343 -6389 8386 -6355
rect 8266 -6423 8386 -6389
rect 8486 -5607 8606 -5583
rect 8486 -5641 8529 -5607
rect 8563 -5641 8606 -5607
rect 8486 -5675 8606 -5641
rect 8486 -5709 8529 -5675
rect 8563 -5709 8606 -5675
rect 8486 -5743 8606 -5709
rect 8486 -5777 8529 -5743
rect 8563 -5777 8606 -5743
rect 8486 -5811 8606 -5777
rect 8486 -5845 8529 -5811
rect 8563 -5845 8606 -5811
rect 8486 -5879 8606 -5845
rect 8486 -5913 8529 -5879
rect 8563 -5913 8606 -5879
rect 8486 -5947 8606 -5913
rect 8486 -5981 8529 -5947
rect 8563 -5981 8606 -5947
rect 8486 -6015 8606 -5981
rect 8486 -6049 8529 -6015
rect 8563 -6049 8606 -6015
rect 8486 -6083 8606 -6049
rect 8486 -6117 8529 -6083
rect 8563 -6117 8606 -6083
rect 8486 -6151 8606 -6117
rect 8486 -6185 8529 -6151
rect 8563 -6185 8606 -6151
rect 8486 -6219 8606 -6185
rect 8486 -6253 8529 -6219
rect 8563 -6253 8606 -6219
rect 8486 -6287 8606 -6253
rect 8486 -6321 8529 -6287
rect 8563 -6321 8606 -6287
rect 8486 -6355 8606 -6321
rect 8486 -6389 8529 -6355
rect 8563 -6389 8606 -6355
rect 8486 -6423 8606 -6389
rect 8706 -5607 8826 -5583
rect 8706 -5641 8749 -5607
rect 8783 -5641 8826 -5607
rect 8706 -5675 8826 -5641
rect 8706 -5709 8749 -5675
rect 8783 -5709 8826 -5675
rect 8706 -5743 8826 -5709
rect 8706 -5777 8749 -5743
rect 8783 -5777 8826 -5743
rect 8706 -5811 8826 -5777
rect 8706 -5845 8749 -5811
rect 8783 -5845 8826 -5811
rect 8706 -5879 8826 -5845
rect 8706 -5913 8749 -5879
rect 8783 -5913 8826 -5879
rect 8706 -5947 8826 -5913
rect 8706 -5981 8749 -5947
rect 8783 -5981 8826 -5947
rect 8706 -6015 8826 -5981
rect 8706 -6049 8749 -6015
rect 8783 -6049 8826 -6015
rect 8706 -6083 8826 -6049
rect 8706 -6117 8749 -6083
rect 8783 -6117 8826 -6083
rect 8706 -6151 8826 -6117
rect 8706 -6185 8749 -6151
rect 8783 -6185 8826 -6151
rect 8706 -6219 8826 -6185
rect 8706 -6253 8749 -6219
rect 8783 -6253 8826 -6219
rect 8706 -6287 8826 -6253
rect 8706 -6321 8749 -6287
rect 8783 -6321 8826 -6287
rect 8706 -6355 8826 -6321
rect 8706 -6389 8749 -6355
rect 8783 -6389 8826 -6355
rect 8706 -6423 8826 -6389
<< pdiff >>
rect 4493 -3976 4613 -3900
rect 4493 -4010 4536 -3976
rect 4570 -4010 4613 -3976
rect 4493 -4044 4613 -4010
rect 4493 -4078 4536 -4044
rect 4570 -4078 4613 -4044
rect 4493 -4112 4613 -4078
rect 4493 -4146 4536 -4112
rect 4570 -4146 4613 -4112
rect 4493 -4180 4613 -4146
rect 4493 -4214 4536 -4180
rect 4570 -4214 4613 -4180
rect 4493 -4248 4613 -4214
rect 4493 -4282 4536 -4248
rect 4570 -4282 4613 -4248
rect 4493 -4316 4613 -4282
rect 4493 -4350 4536 -4316
rect 4570 -4350 4613 -4316
rect 4493 -4384 4613 -4350
rect 4493 -4418 4536 -4384
rect 4570 -4418 4613 -4384
rect 4493 -4452 4613 -4418
rect 4493 -4486 4536 -4452
rect 4570 -4486 4613 -4452
rect 4493 -4520 4613 -4486
rect 4493 -4554 4536 -4520
rect 4570 -4554 4613 -4520
rect 4493 -4588 4613 -4554
rect 4493 -4622 4536 -4588
rect 4570 -4622 4613 -4588
rect 4493 -4656 4613 -4622
rect 4493 -4690 4536 -4656
rect 4570 -4690 4613 -4656
rect 4493 -4724 4613 -4690
rect 4493 -4758 4536 -4724
rect 4570 -4758 4613 -4724
rect 4493 -4792 4613 -4758
rect 4493 -4826 4536 -4792
rect 4570 -4826 4613 -4792
rect 4493 -4850 4613 -4826
rect 4713 -3976 4833 -3900
rect 4713 -4010 4756 -3976
rect 4790 -4010 4833 -3976
rect 4713 -4044 4833 -4010
rect 4713 -4078 4756 -4044
rect 4790 -4078 4833 -4044
rect 4713 -4112 4833 -4078
rect 4713 -4146 4756 -4112
rect 4790 -4146 4833 -4112
rect 4713 -4180 4833 -4146
rect 4713 -4214 4756 -4180
rect 4790 -4214 4833 -4180
rect 4713 -4248 4833 -4214
rect 4713 -4282 4756 -4248
rect 4790 -4282 4833 -4248
rect 4713 -4316 4833 -4282
rect 4713 -4350 4756 -4316
rect 4790 -4350 4833 -4316
rect 4713 -4384 4833 -4350
rect 4713 -4418 4756 -4384
rect 4790 -4418 4833 -4384
rect 4713 -4452 4833 -4418
rect 4713 -4486 4756 -4452
rect 4790 -4486 4833 -4452
rect 4713 -4520 4833 -4486
rect 4713 -4554 4756 -4520
rect 4790 -4554 4833 -4520
rect 4713 -4588 4833 -4554
rect 4713 -4622 4756 -4588
rect 4790 -4622 4833 -4588
rect 4713 -4656 4833 -4622
rect 4713 -4690 4756 -4656
rect 4790 -4690 4833 -4656
rect 4713 -4724 4833 -4690
rect 4713 -4758 4756 -4724
rect 4790 -4758 4833 -4724
rect 4713 -4792 4833 -4758
rect 4713 -4826 4756 -4792
rect 4790 -4826 4833 -4792
rect 4713 -4850 4833 -4826
rect 4933 -3976 5053 -3900
rect 4933 -4010 4976 -3976
rect 5010 -4010 5053 -3976
rect 4933 -4044 5053 -4010
rect 4933 -4078 4976 -4044
rect 5010 -4078 5053 -4044
rect 4933 -4112 5053 -4078
rect 4933 -4146 4976 -4112
rect 5010 -4146 5053 -4112
rect 4933 -4180 5053 -4146
rect 4933 -4214 4976 -4180
rect 5010 -4214 5053 -4180
rect 4933 -4248 5053 -4214
rect 4933 -4282 4976 -4248
rect 5010 -4282 5053 -4248
rect 4933 -4316 5053 -4282
rect 4933 -4350 4976 -4316
rect 5010 -4350 5053 -4316
rect 4933 -4384 5053 -4350
rect 4933 -4418 4976 -4384
rect 5010 -4418 5053 -4384
rect 4933 -4452 5053 -4418
rect 4933 -4486 4976 -4452
rect 5010 -4486 5053 -4452
rect 4933 -4520 5053 -4486
rect 4933 -4554 4976 -4520
rect 5010 -4554 5053 -4520
rect 4933 -4588 5053 -4554
rect 4933 -4622 4976 -4588
rect 5010 -4622 5053 -4588
rect 4933 -4656 5053 -4622
rect 4933 -4690 4976 -4656
rect 5010 -4690 5053 -4656
rect 4933 -4724 5053 -4690
rect 4933 -4758 4976 -4724
rect 5010 -4758 5053 -4724
rect 4933 -4792 5053 -4758
rect 4933 -4826 4976 -4792
rect 5010 -4826 5053 -4792
rect 4933 -4850 5053 -4826
rect 5153 -3976 5273 -3900
rect 5153 -4010 5196 -3976
rect 5230 -4010 5273 -3976
rect 5153 -4044 5273 -4010
rect 5153 -4078 5196 -4044
rect 5230 -4078 5273 -4044
rect 5153 -4112 5273 -4078
rect 5153 -4146 5196 -4112
rect 5230 -4146 5273 -4112
rect 5153 -4180 5273 -4146
rect 5153 -4214 5196 -4180
rect 5230 -4214 5273 -4180
rect 5153 -4248 5273 -4214
rect 5153 -4282 5196 -4248
rect 5230 -4282 5273 -4248
rect 5153 -4316 5273 -4282
rect 5153 -4350 5196 -4316
rect 5230 -4350 5273 -4316
rect 5153 -4384 5273 -4350
rect 5153 -4418 5196 -4384
rect 5230 -4418 5273 -4384
rect 5153 -4452 5273 -4418
rect 5153 -4486 5196 -4452
rect 5230 -4486 5273 -4452
rect 5153 -4520 5273 -4486
rect 5153 -4554 5196 -4520
rect 5230 -4554 5273 -4520
rect 5153 -4588 5273 -4554
rect 5153 -4622 5196 -4588
rect 5230 -4622 5273 -4588
rect 5153 -4656 5273 -4622
rect 5153 -4690 5196 -4656
rect 5230 -4690 5273 -4656
rect 5153 -4724 5273 -4690
rect 5153 -4758 5196 -4724
rect 5230 -4758 5273 -4724
rect 5153 -4792 5273 -4758
rect 5153 -4826 5196 -4792
rect 5230 -4826 5273 -4792
rect 5153 -4850 5273 -4826
rect 5373 -3976 5493 -3900
rect 5373 -4010 5416 -3976
rect 5450 -4010 5493 -3976
rect 5373 -4044 5493 -4010
rect 5373 -4078 5416 -4044
rect 5450 -4078 5493 -4044
rect 5373 -4112 5493 -4078
rect 5373 -4146 5416 -4112
rect 5450 -4146 5493 -4112
rect 5373 -4180 5493 -4146
rect 5373 -4214 5416 -4180
rect 5450 -4214 5493 -4180
rect 5373 -4248 5493 -4214
rect 5373 -4282 5416 -4248
rect 5450 -4282 5493 -4248
rect 5373 -4316 5493 -4282
rect 5373 -4350 5416 -4316
rect 5450 -4350 5493 -4316
rect 5373 -4384 5493 -4350
rect 5373 -4418 5416 -4384
rect 5450 -4418 5493 -4384
rect 5373 -4452 5493 -4418
rect 5373 -4486 5416 -4452
rect 5450 -4486 5493 -4452
rect 5373 -4520 5493 -4486
rect 5373 -4554 5416 -4520
rect 5450 -4554 5493 -4520
rect 5373 -4588 5493 -4554
rect 5373 -4622 5416 -4588
rect 5450 -4622 5493 -4588
rect 5373 -4656 5493 -4622
rect 5373 -4690 5416 -4656
rect 5450 -4690 5493 -4656
rect 5373 -4724 5493 -4690
rect 5373 -4758 5416 -4724
rect 5450 -4758 5493 -4724
rect 5373 -4792 5493 -4758
rect 5373 -4826 5416 -4792
rect 5450 -4826 5493 -4792
rect 5373 -4850 5493 -4826
rect 5593 -3976 5713 -3900
rect 5593 -4010 5636 -3976
rect 5670 -4010 5713 -3976
rect 5593 -4044 5713 -4010
rect 5593 -4078 5636 -4044
rect 5670 -4078 5713 -4044
rect 5593 -4112 5713 -4078
rect 5593 -4146 5636 -4112
rect 5670 -4146 5713 -4112
rect 5593 -4180 5713 -4146
rect 5593 -4214 5636 -4180
rect 5670 -4214 5713 -4180
rect 5593 -4248 5713 -4214
rect 5593 -4282 5636 -4248
rect 5670 -4282 5713 -4248
rect 5593 -4316 5713 -4282
rect 5593 -4350 5636 -4316
rect 5670 -4350 5713 -4316
rect 5593 -4384 5713 -4350
rect 5593 -4418 5636 -4384
rect 5670 -4418 5713 -4384
rect 5593 -4452 5713 -4418
rect 5593 -4486 5636 -4452
rect 5670 -4486 5713 -4452
rect 5593 -4520 5713 -4486
rect 5593 -4554 5636 -4520
rect 5670 -4554 5713 -4520
rect 5593 -4588 5713 -4554
rect 5593 -4622 5636 -4588
rect 5670 -4622 5713 -4588
rect 5593 -4656 5713 -4622
rect 5593 -4690 5636 -4656
rect 5670 -4690 5713 -4656
rect 5593 -4724 5713 -4690
rect 5593 -4758 5636 -4724
rect 5670 -4758 5713 -4724
rect 5593 -4792 5713 -4758
rect 5593 -4826 5636 -4792
rect 5670 -4826 5713 -4792
rect 5593 -4850 5713 -4826
rect 5813 -3976 5933 -3900
rect 5813 -4010 5856 -3976
rect 5890 -4010 5933 -3976
rect 5813 -4044 5933 -4010
rect 5813 -4078 5856 -4044
rect 5890 -4078 5933 -4044
rect 5813 -4112 5933 -4078
rect 5813 -4146 5856 -4112
rect 5890 -4146 5933 -4112
rect 5813 -4180 5933 -4146
rect 5813 -4214 5856 -4180
rect 5890 -4214 5933 -4180
rect 5813 -4248 5933 -4214
rect 5813 -4282 5856 -4248
rect 5890 -4282 5933 -4248
rect 5813 -4316 5933 -4282
rect 5813 -4350 5856 -4316
rect 5890 -4350 5933 -4316
rect 5813 -4384 5933 -4350
rect 5813 -4418 5856 -4384
rect 5890 -4418 5933 -4384
rect 5813 -4452 5933 -4418
rect 5813 -4486 5856 -4452
rect 5890 -4486 5933 -4452
rect 5813 -4520 5933 -4486
rect 5813 -4554 5856 -4520
rect 5890 -4554 5933 -4520
rect 5813 -4588 5933 -4554
rect 5813 -4622 5856 -4588
rect 5890 -4622 5933 -4588
rect 5813 -4656 5933 -4622
rect 5813 -4690 5856 -4656
rect 5890 -4690 5933 -4656
rect 5813 -4724 5933 -4690
rect 5813 -4758 5856 -4724
rect 5890 -4758 5933 -4724
rect 5813 -4792 5933 -4758
rect 5813 -4826 5856 -4792
rect 5890 -4826 5933 -4792
rect 5813 -4850 5933 -4826
rect 6033 -3976 6153 -3900
rect 6033 -4010 6076 -3976
rect 6110 -4010 6153 -3976
rect 6033 -4044 6153 -4010
rect 6033 -4078 6076 -4044
rect 6110 -4078 6153 -4044
rect 6033 -4112 6153 -4078
rect 6033 -4146 6076 -4112
rect 6110 -4146 6153 -4112
rect 6033 -4180 6153 -4146
rect 6033 -4214 6076 -4180
rect 6110 -4214 6153 -4180
rect 6033 -4248 6153 -4214
rect 6033 -4282 6076 -4248
rect 6110 -4282 6153 -4248
rect 6033 -4316 6153 -4282
rect 6033 -4350 6076 -4316
rect 6110 -4350 6153 -4316
rect 6033 -4384 6153 -4350
rect 6033 -4418 6076 -4384
rect 6110 -4418 6153 -4384
rect 6033 -4452 6153 -4418
rect 6033 -4486 6076 -4452
rect 6110 -4486 6153 -4452
rect 6033 -4520 6153 -4486
rect 6033 -4554 6076 -4520
rect 6110 -4554 6153 -4520
rect 6033 -4588 6153 -4554
rect 6033 -4622 6076 -4588
rect 6110 -4622 6153 -4588
rect 6033 -4656 6153 -4622
rect 6033 -4690 6076 -4656
rect 6110 -4690 6153 -4656
rect 6033 -4724 6153 -4690
rect 6033 -4758 6076 -4724
rect 6110 -4758 6153 -4724
rect 6033 -4792 6153 -4758
rect 6033 -4826 6076 -4792
rect 6110 -4826 6153 -4792
rect 6033 -4850 6153 -4826
rect 6253 -3976 6373 -3900
rect 6253 -4010 6296 -3976
rect 6330 -4010 6373 -3976
rect 6253 -4044 6373 -4010
rect 6253 -4078 6296 -4044
rect 6330 -4078 6373 -4044
rect 6253 -4112 6373 -4078
rect 6253 -4146 6296 -4112
rect 6330 -4146 6373 -4112
rect 6253 -4180 6373 -4146
rect 6253 -4214 6296 -4180
rect 6330 -4214 6373 -4180
rect 6253 -4248 6373 -4214
rect 6253 -4282 6296 -4248
rect 6330 -4282 6373 -4248
rect 6253 -4316 6373 -4282
rect 6253 -4350 6296 -4316
rect 6330 -4350 6373 -4316
rect 6253 -4384 6373 -4350
rect 6253 -4418 6296 -4384
rect 6330 -4418 6373 -4384
rect 6253 -4452 6373 -4418
rect 6253 -4486 6296 -4452
rect 6330 -4486 6373 -4452
rect 6253 -4520 6373 -4486
rect 6253 -4554 6296 -4520
rect 6330 -4554 6373 -4520
rect 6253 -4588 6373 -4554
rect 6253 -4622 6296 -4588
rect 6330 -4622 6373 -4588
rect 6253 -4656 6373 -4622
rect 6253 -4690 6296 -4656
rect 6330 -4690 6373 -4656
rect 6253 -4724 6373 -4690
rect 6253 -4758 6296 -4724
rect 6330 -4758 6373 -4724
rect 6253 -4792 6373 -4758
rect 6253 -4826 6296 -4792
rect 6330 -4826 6373 -4792
rect 6253 -4850 6373 -4826
<< ndiffc >>
rect 2081 -5641 2115 -5607
rect 2081 -5709 2115 -5675
rect 2081 -5777 2115 -5743
rect 2081 -5845 2115 -5811
rect 2081 -5913 2115 -5879
rect 2081 -5981 2115 -5947
rect 2081 -6049 2115 -6015
rect 2081 -6117 2115 -6083
rect 2081 -6185 2115 -6151
rect 2081 -6253 2115 -6219
rect 2081 -6321 2115 -6287
rect 2081 -6389 2115 -6355
rect 2301 -5641 2335 -5607
rect 2301 -5709 2335 -5675
rect 2301 -5777 2335 -5743
rect 2301 -5845 2335 -5811
rect 2301 -5913 2335 -5879
rect 2301 -5981 2335 -5947
rect 2301 -6049 2335 -6015
rect 2301 -6117 2335 -6083
rect 2301 -6185 2335 -6151
rect 2301 -6253 2335 -6219
rect 2301 -6321 2335 -6287
rect 2301 -6389 2335 -6355
rect 2521 -5641 2555 -5607
rect 2521 -5709 2555 -5675
rect 2521 -5777 2555 -5743
rect 2521 -5845 2555 -5811
rect 2521 -5913 2555 -5879
rect 2521 -5981 2555 -5947
rect 2521 -6049 2555 -6015
rect 2521 -6117 2555 -6083
rect 2521 -6185 2555 -6151
rect 2521 -6253 2555 -6219
rect 2521 -6321 2555 -6287
rect 2521 -6389 2555 -6355
rect 2741 -5641 2775 -5607
rect 2741 -5709 2775 -5675
rect 2741 -5777 2775 -5743
rect 2741 -5845 2775 -5811
rect 2741 -5913 2775 -5879
rect 2741 -5981 2775 -5947
rect 2741 -6049 2775 -6015
rect 2741 -6117 2775 -6083
rect 2741 -6185 2775 -6151
rect 2741 -6253 2775 -6219
rect 2741 -6321 2775 -6287
rect 2741 -6389 2775 -6355
rect 2961 -5641 2995 -5607
rect 2961 -5709 2995 -5675
rect 2961 -5777 2995 -5743
rect 2961 -5845 2995 -5811
rect 2961 -5913 2995 -5879
rect 2961 -5981 2995 -5947
rect 2961 -6049 2995 -6015
rect 2961 -6117 2995 -6083
rect 2961 -6185 2995 -6151
rect 2961 -6253 2995 -6219
rect 2961 -6321 2995 -6287
rect 2961 -6389 2995 -6355
rect 3181 -5641 3215 -5607
rect 3181 -5709 3215 -5675
rect 3181 -5777 3215 -5743
rect 3181 -5845 3215 -5811
rect 3181 -5913 3215 -5879
rect 3181 -5981 3215 -5947
rect 3181 -6049 3215 -6015
rect 3181 -6117 3215 -6083
rect 3181 -6185 3215 -6151
rect 3181 -6253 3215 -6219
rect 3181 -6321 3215 -6287
rect 3181 -6389 3215 -6355
rect 3401 -5641 3435 -5607
rect 3401 -5709 3435 -5675
rect 3401 -5777 3435 -5743
rect 3401 -5845 3435 -5811
rect 3401 -5913 3435 -5879
rect 3401 -5981 3435 -5947
rect 3401 -6049 3435 -6015
rect 3401 -6117 3435 -6083
rect 3401 -6185 3435 -6151
rect 3401 -6253 3435 -6219
rect 3401 -6321 3435 -6287
rect 3401 -6389 3435 -6355
rect 3621 -5641 3655 -5607
rect 3621 -5709 3655 -5675
rect 3621 -5777 3655 -5743
rect 3621 -5845 3655 -5811
rect 3621 -5913 3655 -5879
rect 3621 -5981 3655 -5947
rect 3621 -6049 3655 -6015
rect 3621 -6117 3655 -6083
rect 3621 -6185 3655 -6151
rect 3621 -6253 3655 -6219
rect 3621 -6321 3655 -6287
rect 3621 -6389 3655 -6355
rect 3841 -5641 3875 -5607
rect 3841 -5709 3875 -5675
rect 3841 -5777 3875 -5743
rect 3841 -5845 3875 -5811
rect 3841 -5913 3875 -5879
rect 3841 -5981 3875 -5947
rect 3841 -6049 3875 -6015
rect 3841 -6117 3875 -6083
rect 3841 -6185 3875 -6151
rect 3841 -6253 3875 -6219
rect 3841 -6321 3875 -6287
rect 3841 -6389 3875 -6355
rect 4535 -5589 4569 -5555
rect 4535 -5657 4569 -5623
rect 4535 -5725 4569 -5691
rect 4535 -5793 4569 -5759
rect 4535 -5861 4569 -5827
rect 4535 -5929 4569 -5895
rect 4535 -5997 4569 -5963
rect 4535 -6065 4569 -6031
rect 4535 -6133 4569 -6099
rect 4535 -6201 4569 -6167
rect 4535 -6269 4569 -6235
rect 4535 -6337 4569 -6303
rect 4535 -6405 4569 -6371
rect 4755 -5589 4789 -5555
rect 4755 -5657 4789 -5623
rect 4755 -5725 4789 -5691
rect 4755 -5793 4789 -5759
rect 4755 -5861 4789 -5827
rect 4755 -5929 4789 -5895
rect 4755 -5997 4789 -5963
rect 4755 -6065 4789 -6031
rect 4755 -6133 4789 -6099
rect 4755 -6201 4789 -6167
rect 4755 -6269 4789 -6235
rect 4755 -6337 4789 -6303
rect 4755 -6405 4789 -6371
rect 4975 -5589 5009 -5555
rect 4975 -5657 5009 -5623
rect 4975 -5725 5009 -5691
rect 4975 -5793 5009 -5759
rect 4975 -5861 5009 -5827
rect 4975 -5929 5009 -5895
rect 4975 -5997 5009 -5963
rect 4975 -6065 5009 -6031
rect 4975 -6133 5009 -6099
rect 4975 -6201 5009 -6167
rect 4975 -6269 5009 -6235
rect 4975 -6337 5009 -6303
rect 4975 -6405 5009 -6371
rect 5195 -5589 5229 -5555
rect 5195 -5657 5229 -5623
rect 5195 -5725 5229 -5691
rect 5195 -5793 5229 -5759
rect 5195 -5861 5229 -5827
rect 5195 -5929 5229 -5895
rect 5195 -5997 5229 -5963
rect 5195 -6065 5229 -6031
rect 5195 -6133 5229 -6099
rect 5195 -6201 5229 -6167
rect 5195 -6269 5229 -6235
rect 5195 -6337 5229 -6303
rect 5195 -6405 5229 -6371
rect 5415 -5589 5449 -5555
rect 5415 -5657 5449 -5623
rect 5415 -5725 5449 -5691
rect 5415 -5793 5449 -5759
rect 5415 -5861 5449 -5827
rect 5415 -5929 5449 -5895
rect 5415 -5997 5449 -5963
rect 5415 -6065 5449 -6031
rect 5415 -6133 5449 -6099
rect 5415 -6201 5449 -6167
rect 5415 -6269 5449 -6235
rect 5415 -6337 5449 -6303
rect 5415 -6405 5449 -6371
rect 5635 -5589 5669 -5555
rect 5635 -5657 5669 -5623
rect 5635 -5725 5669 -5691
rect 5635 -5793 5669 -5759
rect 5635 -5861 5669 -5827
rect 5635 -5929 5669 -5895
rect 5635 -5997 5669 -5963
rect 5635 -6065 5669 -6031
rect 5635 -6133 5669 -6099
rect 5635 -6201 5669 -6167
rect 5635 -6269 5669 -6235
rect 5635 -6337 5669 -6303
rect 5635 -6405 5669 -6371
rect 5855 -5589 5889 -5555
rect 5855 -5657 5889 -5623
rect 5855 -5725 5889 -5691
rect 5855 -5793 5889 -5759
rect 5855 -5861 5889 -5827
rect 5855 -5929 5889 -5895
rect 5855 -5997 5889 -5963
rect 5855 -6065 5889 -6031
rect 5855 -6133 5889 -6099
rect 5855 -6201 5889 -6167
rect 5855 -6269 5889 -6235
rect 5855 -6337 5889 -6303
rect 5855 -6405 5889 -6371
rect 6075 -5589 6109 -5555
rect 6075 -5657 6109 -5623
rect 6075 -5725 6109 -5691
rect 6075 -5793 6109 -5759
rect 6075 -5861 6109 -5827
rect 6075 -5929 6109 -5895
rect 6075 -5997 6109 -5963
rect 6075 -6065 6109 -6031
rect 6075 -6133 6109 -6099
rect 6075 -6201 6109 -6167
rect 6075 -6269 6109 -6235
rect 6075 -6337 6109 -6303
rect 6075 -6405 6109 -6371
rect 6295 -5589 6329 -5555
rect 6295 -5657 6329 -5623
rect 6295 -5725 6329 -5691
rect 6295 -5793 6329 -5759
rect 6295 -5861 6329 -5827
rect 6295 -5929 6329 -5895
rect 6295 -5997 6329 -5963
rect 6295 -6065 6329 -6031
rect 6295 -6133 6329 -6099
rect 6295 -6201 6329 -6167
rect 6295 -6269 6329 -6235
rect 6295 -6337 6329 -6303
rect 6295 -6405 6329 -6371
rect 6989 -5641 7023 -5607
rect 6989 -5709 7023 -5675
rect 6989 -5777 7023 -5743
rect 6989 -5845 7023 -5811
rect 6989 -5913 7023 -5879
rect 6989 -5981 7023 -5947
rect 6989 -6049 7023 -6015
rect 6989 -6117 7023 -6083
rect 6989 -6185 7023 -6151
rect 6989 -6253 7023 -6219
rect 6989 -6321 7023 -6287
rect 6989 -6389 7023 -6355
rect 7209 -5641 7243 -5607
rect 7209 -5709 7243 -5675
rect 7209 -5777 7243 -5743
rect 7209 -5845 7243 -5811
rect 7209 -5913 7243 -5879
rect 7209 -5981 7243 -5947
rect 7209 -6049 7243 -6015
rect 7209 -6117 7243 -6083
rect 7209 -6185 7243 -6151
rect 7209 -6253 7243 -6219
rect 7209 -6321 7243 -6287
rect 7209 -6389 7243 -6355
rect 7429 -5641 7463 -5607
rect 7429 -5709 7463 -5675
rect 7429 -5777 7463 -5743
rect 7429 -5845 7463 -5811
rect 7429 -5913 7463 -5879
rect 7429 -5981 7463 -5947
rect 7429 -6049 7463 -6015
rect 7429 -6117 7463 -6083
rect 7429 -6185 7463 -6151
rect 7429 -6253 7463 -6219
rect 7429 -6321 7463 -6287
rect 7429 -6389 7463 -6355
rect 7649 -5641 7683 -5607
rect 7649 -5709 7683 -5675
rect 7649 -5777 7683 -5743
rect 7649 -5845 7683 -5811
rect 7649 -5913 7683 -5879
rect 7649 -5981 7683 -5947
rect 7649 -6049 7683 -6015
rect 7649 -6117 7683 -6083
rect 7649 -6185 7683 -6151
rect 7649 -6253 7683 -6219
rect 7649 -6321 7683 -6287
rect 7649 -6389 7683 -6355
rect 7869 -5641 7903 -5607
rect 7869 -5709 7903 -5675
rect 7869 -5777 7903 -5743
rect 7869 -5845 7903 -5811
rect 7869 -5913 7903 -5879
rect 7869 -5981 7903 -5947
rect 7869 -6049 7903 -6015
rect 7869 -6117 7903 -6083
rect 7869 -6185 7903 -6151
rect 7869 -6253 7903 -6219
rect 7869 -6321 7903 -6287
rect 7869 -6389 7903 -6355
rect 8089 -5641 8123 -5607
rect 8089 -5709 8123 -5675
rect 8089 -5777 8123 -5743
rect 8089 -5845 8123 -5811
rect 8089 -5913 8123 -5879
rect 8089 -5981 8123 -5947
rect 8089 -6049 8123 -6015
rect 8089 -6117 8123 -6083
rect 8089 -6185 8123 -6151
rect 8089 -6253 8123 -6219
rect 8089 -6321 8123 -6287
rect 8089 -6389 8123 -6355
rect 8309 -5641 8343 -5607
rect 8309 -5709 8343 -5675
rect 8309 -5777 8343 -5743
rect 8309 -5845 8343 -5811
rect 8309 -5913 8343 -5879
rect 8309 -5981 8343 -5947
rect 8309 -6049 8343 -6015
rect 8309 -6117 8343 -6083
rect 8309 -6185 8343 -6151
rect 8309 -6253 8343 -6219
rect 8309 -6321 8343 -6287
rect 8309 -6389 8343 -6355
rect 8529 -5641 8563 -5607
rect 8529 -5709 8563 -5675
rect 8529 -5777 8563 -5743
rect 8529 -5845 8563 -5811
rect 8529 -5913 8563 -5879
rect 8529 -5981 8563 -5947
rect 8529 -6049 8563 -6015
rect 8529 -6117 8563 -6083
rect 8529 -6185 8563 -6151
rect 8529 -6253 8563 -6219
rect 8529 -6321 8563 -6287
rect 8529 -6389 8563 -6355
rect 8749 -5641 8783 -5607
rect 8749 -5709 8783 -5675
rect 8749 -5777 8783 -5743
rect 8749 -5845 8783 -5811
rect 8749 -5913 8783 -5879
rect 8749 -5981 8783 -5947
rect 8749 -6049 8783 -6015
rect 8749 -6117 8783 -6083
rect 8749 -6185 8783 -6151
rect 8749 -6253 8783 -6219
rect 8749 -6321 8783 -6287
rect 8749 -6389 8783 -6355
<< pdiffc >>
rect 4536 -4010 4570 -3976
rect 4536 -4078 4570 -4044
rect 4536 -4146 4570 -4112
rect 4536 -4214 4570 -4180
rect 4536 -4282 4570 -4248
rect 4536 -4350 4570 -4316
rect 4536 -4418 4570 -4384
rect 4536 -4486 4570 -4452
rect 4536 -4554 4570 -4520
rect 4536 -4622 4570 -4588
rect 4536 -4690 4570 -4656
rect 4536 -4758 4570 -4724
rect 4536 -4826 4570 -4792
rect 4756 -4010 4790 -3976
rect 4756 -4078 4790 -4044
rect 4756 -4146 4790 -4112
rect 4756 -4214 4790 -4180
rect 4756 -4282 4790 -4248
rect 4756 -4350 4790 -4316
rect 4756 -4418 4790 -4384
rect 4756 -4486 4790 -4452
rect 4756 -4554 4790 -4520
rect 4756 -4622 4790 -4588
rect 4756 -4690 4790 -4656
rect 4756 -4758 4790 -4724
rect 4756 -4826 4790 -4792
rect 4976 -4010 5010 -3976
rect 4976 -4078 5010 -4044
rect 4976 -4146 5010 -4112
rect 4976 -4214 5010 -4180
rect 4976 -4282 5010 -4248
rect 4976 -4350 5010 -4316
rect 4976 -4418 5010 -4384
rect 4976 -4486 5010 -4452
rect 4976 -4554 5010 -4520
rect 4976 -4622 5010 -4588
rect 4976 -4690 5010 -4656
rect 4976 -4758 5010 -4724
rect 4976 -4826 5010 -4792
rect 5196 -4010 5230 -3976
rect 5196 -4078 5230 -4044
rect 5196 -4146 5230 -4112
rect 5196 -4214 5230 -4180
rect 5196 -4282 5230 -4248
rect 5196 -4350 5230 -4316
rect 5196 -4418 5230 -4384
rect 5196 -4486 5230 -4452
rect 5196 -4554 5230 -4520
rect 5196 -4622 5230 -4588
rect 5196 -4690 5230 -4656
rect 5196 -4758 5230 -4724
rect 5196 -4826 5230 -4792
rect 5416 -4010 5450 -3976
rect 5416 -4078 5450 -4044
rect 5416 -4146 5450 -4112
rect 5416 -4214 5450 -4180
rect 5416 -4282 5450 -4248
rect 5416 -4350 5450 -4316
rect 5416 -4418 5450 -4384
rect 5416 -4486 5450 -4452
rect 5416 -4554 5450 -4520
rect 5416 -4622 5450 -4588
rect 5416 -4690 5450 -4656
rect 5416 -4758 5450 -4724
rect 5416 -4826 5450 -4792
rect 5636 -4010 5670 -3976
rect 5636 -4078 5670 -4044
rect 5636 -4146 5670 -4112
rect 5636 -4214 5670 -4180
rect 5636 -4282 5670 -4248
rect 5636 -4350 5670 -4316
rect 5636 -4418 5670 -4384
rect 5636 -4486 5670 -4452
rect 5636 -4554 5670 -4520
rect 5636 -4622 5670 -4588
rect 5636 -4690 5670 -4656
rect 5636 -4758 5670 -4724
rect 5636 -4826 5670 -4792
rect 5856 -4010 5890 -3976
rect 5856 -4078 5890 -4044
rect 5856 -4146 5890 -4112
rect 5856 -4214 5890 -4180
rect 5856 -4282 5890 -4248
rect 5856 -4350 5890 -4316
rect 5856 -4418 5890 -4384
rect 5856 -4486 5890 -4452
rect 5856 -4554 5890 -4520
rect 5856 -4622 5890 -4588
rect 5856 -4690 5890 -4656
rect 5856 -4758 5890 -4724
rect 5856 -4826 5890 -4792
rect 6076 -4010 6110 -3976
rect 6076 -4078 6110 -4044
rect 6076 -4146 6110 -4112
rect 6076 -4214 6110 -4180
rect 6076 -4282 6110 -4248
rect 6076 -4350 6110 -4316
rect 6076 -4418 6110 -4384
rect 6076 -4486 6110 -4452
rect 6076 -4554 6110 -4520
rect 6076 -4622 6110 -4588
rect 6076 -4690 6110 -4656
rect 6076 -4758 6110 -4724
rect 6076 -4826 6110 -4792
rect 6296 -4010 6330 -3976
rect 6296 -4078 6330 -4044
rect 6296 -4146 6330 -4112
rect 6296 -4214 6330 -4180
rect 6296 -4282 6330 -4248
rect 6296 -4350 6330 -4316
rect 6296 -4418 6330 -4384
rect 6296 -4486 6330 -4452
rect 6296 -4554 6330 -4520
rect 6296 -4622 6330 -4588
rect 6296 -4690 6330 -4656
rect 6296 -4758 6330 -4724
rect 6296 -4826 6330 -4792
<< psubdiff >>
rect 4372 -5555 4492 -5505
rect 1918 -5607 2038 -5583
rect 1918 -5641 1961 -5607
rect 1995 -5641 2038 -5607
rect 1918 -5675 2038 -5641
rect 1918 -5709 1961 -5675
rect 1995 -5709 2038 -5675
rect 1918 -5743 2038 -5709
rect 1918 -5777 1961 -5743
rect 1995 -5777 2038 -5743
rect 1918 -5811 2038 -5777
rect 1918 -5845 1961 -5811
rect 1995 -5845 2038 -5811
rect 1918 -5879 2038 -5845
rect 1918 -5913 1961 -5879
rect 1995 -5913 2038 -5879
rect 1918 -5947 2038 -5913
rect 1918 -5981 1961 -5947
rect 1995 -5981 2038 -5947
rect 1918 -6015 2038 -5981
rect 1918 -6049 1961 -6015
rect 1995 -6049 2038 -6015
rect 1918 -6083 2038 -6049
rect 1918 -6117 1961 -6083
rect 1995 -6117 2038 -6083
rect 1918 -6151 2038 -6117
rect 1918 -6185 1961 -6151
rect 1995 -6185 2038 -6151
rect 1918 -6219 2038 -6185
rect 1918 -6253 1961 -6219
rect 1995 -6253 2038 -6219
rect 1918 -6287 2038 -6253
rect 1918 -6321 1961 -6287
rect 1995 -6321 2038 -6287
rect 1918 -6355 2038 -6321
rect 1918 -6389 1961 -6355
rect 1995 -6389 2038 -6355
rect 1918 -6423 2038 -6389
rect 3918 -5607 4038 -5583
rect 3918 -5641 3961 -5607
rect 3995 -5641 4038 -5607
rect 3918 -5675 4038 -5641
rect 3918 -5709 3961 -5675
rect 3995 -5709 4038 -5675
rect 3918 -5743 4038 -5709
rect 3918 -5777 3961 -5743
rect 3995 -5777 4038 -5743
rect 3918 -5811 4038 -5777
rect 3918 -5845 3961 -5811
rect 3995 -5845 4038 -5811
rect 3918 -5879 4038 -5845
rect 3918 -5913 3961 -5879
rect 3995 -5913 4038 -5879
rect 3918 -5947 4038 -5913
rect 3918 -5981 3961 -5947
rect 3995 -5981 4038 -5947
rect 3918 -6015 4038 -5981
rect 3918 -6049 3961 -6015
rect 3995 -6049 4038 -6015
rect 3918 -6083 4038 -6049
rect 3918 -6117 3961 -6083
rect 3995 -6117 4038 -6083
rect 3918 -6151 4038 -6117
rect 3918 -6185 3961 -6151
rect 3995 -6185 4038 -6151
rect 3918 -6219 4038 -6185
rect 3918 -6253 3961 -6219
rect 3995 -6253 4038 -6219
rect 3918 -6287 4038 -6253
rect 3918 -6321 3961 -6287
rect 3995 -6321 4038 -6287
rect 3918 -6355 4038 -6321
rect 3918 -6389 3961 -6355
rect 3995 -6389 4038 -6355
rect 3918 -6423 4038 -6389
rect 4372 -5589 4415 -5555
rect 4449 -5589 4492 -5555
rect 4372 -5623 4492 -5589
rect 4372 -5657 4415 -5623
rect 4449 -5657 4492 -5623
rect 4372 -5691 4492 -5657
rect 4372 -5725 4415 -5691
rect 4449 -5725 4492 -5691
rect 4372 -5759 4492 -5725
rect 4372 -5793 4415 -5759
rect 4449 -5793 4492 -5759
rect 4372 -5827 4492 -5793
rect 4372 -5861 4415 -5827
rect 4449 -5861 4492 -5827
rect 4372 -5895 4492 -5861
rect 4372 -5929 4415 -5895
rect 4449 -5929 4492 -5895
rect 4372 -5963 4492 -5929
rect 4372 -5997 4415 -5963
rect 4449 -5997 4492 -5963
rect 4372 -6031 4492 -5997
rect 4372 -6065 4415 -6031
rect 4449 -6065 4492 -6031
rect 4372 -6099 4492 -6065
rect 4372 -6133 4415 -6099
rect 4449 -6133 4492 -6099
rect 4372 -6167 4492 -6133
rect 4372 -6201 4415 -6167
rect 4449 -6201 4492 -6167
rect 4372 -6235 4492 -6201
rect 4372 -6269 4415 -6235
rect 4449 -6269 4492 -6235
rect 4372 -6303 4492 -6269
rect 4372 -6337 4415 -6303
rect 4449 -6337 4492 -6303
rect 4372 -6371 4492 -6337
rect 4372 -6405 4415 -6371
rect 4449 -6405 4492 -6371
rect 4372 -6455 4492 -6405
rect 6372 -5555 6492 -5505
rect 6372 -5589 6415 -5555
rect 6449 -5589 6492 -5555
rect 6372 -5623 6492 -5589
rect 6372 -5657 6415 -5623
rect 6449 -5657 6492 -5623
rect 6372 -5691 6492 -5657
rect 6372 -5725 6415 -5691
rect 6449 -5725 6492 -5691
rect 6372 -5759 6492 -5725
rect 6372 -5793 6415 -5759
rect 6449 -5793 6492 -5759
rect 6372 -5827 6492 -5793
rect 6372 -5861 6415 -5827
rect 6449 -5861 6492 -5827
rect 6372 -5895 6492 -5861
rect 6372 -5929 6415 -5895
rect 6449 -5929 6492 -5895
rect 6372 -5963 6492 -5929
rect 6372 -5997 6415 -5963
rect 6449 -5997 6492 -5963
rect 6372 -6031 6492 -5997
rect 6372 -6065 6415 -6031
rect 6449 -6065 6492 -6031
rect 6372 -6099 6492 -6065
rect 6372 -6133 6415 -6099
rect 6449 -6133 6492 -6099
rect 6372 -6167 6492 -6133
rect 6372 -6201 6415 -6167
rect 6449 -6201 6492 -6167
rect 6372 -6235 6492 -6201
rect 6372 -6269 6415 -6235
rect 6449 -6269 6492 -6235
rect 6372 -6303 6492 -6269
rect 6372 -6337 6415 -6303
rect 6449 -6337 6492 -6303
rect 6372 -6371 6492 -6337
rect 6372 -6405 6415 -6371
rect 6449 -6405 6492 -6371
rect 6372 -6455 6492 -6405
rect 6826 -5607 6946 -5583
rect 6826 -5641 6869 -5607
rect 6903 -5641 6946 -5607
rect 6826 -5675 6946 -5641
rect 6826 -5709 6869 -5675
rect 6903 -5709 6946 -5675
rect 6826 -5743 6946 -5709
rect 6826 -5777 6869 -5743
rect 6903 -5777 6946 -5743
rect 6826 -5811 6946 -5777
rect 6826 -5845 6869 -5811
rect 6903 -5845 6946 -5811
rect 6826 -5879 6946 -5845
rect 6826 -5913 6869 -5879
rect 6903 -5913 6946 -5879
rect 6826 -5947 6946 -5913
rect 6826 -5981 6869 -5947
rect 6903 -5981 6946 -5947
rect 6826 -6015 6946 -5981
rect 6826 -6049 6869 -6015
rect 6903 -6049 6946 -6015
rect 6826 -6083 6946 -6049
rect 6826 -6117 6869 -6083
rect 6903 -6117 6946 -6083
rect 6826 -6151 6946 -6117
rect 6826 -6185 6869 -6151
rect 6903 -6185 6946 -6151
rect 6826 -6219 6946 -6185
rect 6826 -6253 6869 -6219
rect 6903 -6253 6946 -6219
rect 6826 -6287 6946 -6253
rect 6826 -6321 6869 -6287
rect 6903 -6321 6946 -6287
rect 6826 -6355 6946 -6321
rect 6826 -6389 6869 -6355
rect 6903 -6389 6946 -6355
rect 6826 -6423 6946 -6389
rect 8826 -5607 8946 -5583
rect 8826 -5641 8869 -5607
rect 8903 -5641 8946 -5607
rect 8826 -5675 8946 -5641
rect 8826 -5709 8869 -5675
rect 8903 -5709 8946 -5675
rect 8826 -5743 8946 -5709
rect 8826 -5777 8869 -5743
rect 8903 -5777 8946 -5743
rect 8826 -5811 8946 -5777
rect 8826 -5845 8869 -5811
rect 8903 -5845 8946 -5811
rect 8826 -5879 8946 -5845
rect 8826 -5913 8869 -5879
rect 8903 -5913 8946 -5879
rect 8826 -5947 8946 -5913
rect 8826 -5981 8869 -5947
rect 8903 -5981 8946 -5947
rect 8826 -6015 8946 -5981
rect 8826 -6049 8869 -6015
rect 8903 -6049 8946 -6015
rect 8826 -6083 8946 -6049
rect 8826 -6117 8869 -6083
rect 8903 -6117 8946 -6083
rect 8826 -6151 8946 -6117
rect 8826 -6185 8869 -6151
rect 8903 -6185 8946 -6151
rect 8826 -6219 8946 -6185
rect 8826 -6253 8869 -6219
rect 8903 -6253 8946 -6219
rect 8826 -6287 8946 -6253
rect 8826 -6321 8869 -6287
rect 8903 -6321 8946 -6287
rect 8826 -6355 8946 -6321
rect 8826 -6389 8869 -6355
rect 8903 -6389 8946 -6355
rect 8826 -6423 8946 -6389
<< nsubdiff >>
rect 4373 -3976 4493 -3900
rect 4373 -4010 4416 -3976
rect 4450 -4010 4493 -3976
rect 4373 -4044 4493 -4010
rect 4373 -4078 4416 -4044
rect 4450 -4078 4493 -4044
rect 4373 -4112 4493 -4078
rect 4373 -4146 4416 -4112
rect 4450 -4146 4493 -4112
rect 4373 -4180 4493 -4146
rect 4373 -4214 4416 -4180
rect 4450 -4214 4493 -4180
rect 4373 -4248 4493 -4214
rect 4373 -4282 4416 -4248
rect 4450 -4282 4493 -4248
rect 4373 -4316 4493 -4282
rect 4373 -4350 4416 -4316
rect 4450 -4350 4493 -4316
rect 4373 -4384 4493 -4350
rect 4373 -4418 4416 -4384
rect 4450 -4418 4493 -4384
rect 4373 -4452 4493 -4418
rect 4373 -4486 4416 -4452
rect 4450 -4486 4493 -4452
rect 4373 -4520 4493 -4486
rect 4373 -4554 4416 -4520
rect 4450 -4554 4493 -4520
rect 4373 -4588 4493 -4554
rect 4373 -4622 4416 -4588
rect 4450 -4622 4493 -4588
rect 4373 -4656 4493 -4622
rect 4373 -4690 4416 -4656
rect 4450 -4690 4493 -4656
rect 4373 -4724 4493 -4690
rect 4373 -4758 4416 -4724
rect 4450 -4758 4493 -4724
rect 4373 -4792 4493 -4758
rect 4373 -4826 4416 -4792
rect 4450 -4826 4493 -4792
rect 4373 -4850 4493 -4826
rect 6373 -3976 6493 -3900
rect 6373 -4010 6416 -3976
rect 6450 -4010 6493 -3976
rect 6373 -4044 6493 -4010
rect 6373 -4078 6416 -4044
rect 6450 -4078 6493 -4044
rect 6373 -4112 6493 -4078
rect 6373 -4146 6416 -4112
rect 6450 -4146 6493 -4112
rect 6373 -4180 6493 -4146
rect 6373 -4214 6416 -4180
rect 6450 -4214 6493 -4180
rect 6373 -4248 6493 -4214
rect 6373 -4282 6416 -4248
rect 6450 -4282 6493 -4248
rect 6373 -4316 6493 -4282
rect 6373 -4350 6416 -4316
rect 6450 -4350 6493 -4316
rect 6373 -4384 6493 -4350
rect 6373 -4418 6416 -4384
rect 6450 -4418 6493 -4384
rect 6373 -4452 6493 -4418
rect 6373 -4486 6416 -4452
rect 6450 -4486 6493 -4452
rect 6373 -4520 6493 -4486
rect 6373 -4554 6416 -4520
rect 6450 -4554 6493 -4520
rect 6373 -4588 6493 -4554
rect 6373 -4622 6416 -4588
rect 6450 -4622 6493 -4588
rect 6373 -4656 6493 -4622
rect 6373 -4690 6416 -4656
rect 6450 -4690 6493 -4656
rect 6373 -4724 6493 -4690
rect 6373 -4758 6416 -4724
rect 6450 -4758 6493 -4724
rect 6373 -4792 6493 -4758
rect 6373 -4826 6416 -4792
rect 6450 -4826 6493 -4792
rect 6373 -4850 6493 -4826
<< psubdiffcont >>
rect 1961 -5641 1995 -5607
rect 1961 -5709 1995 -5675
rect 1961 -5777 1995 -5743
rect 1961 -5845 1995 -5811
rect 1961 -5913 1995 -5879
rect 1961 -5981 1995 -5947
rect 1961 -6049 1995 -6015
rect 1961 -6117 1995 -6083
rect 1961 -6185 1995 -6151
rect 1961 -6253 1995 -6219
rect 1961 -6321 1995 -6287
rect 1961 -6389 1995 -6355
rect 3961 -5641 3995 -5607
rect 3961 -5709 3995 -5675
rect 3961 -5777 3995 -5743
rect 3961 -5845 3995 -5811
rect 3961 -5913 3995 -5879
rect 3961 -5981 3995 -5947
rect 3961 -6049 3995 -6015
rect 3961 -6117 3995 -6083
rect 3961 -6185 3995 -6151
rect 3961 -6253 3995 -6219
rect 3961 -6321 3995 -6287
rect 3961 -6389 3995 -6355
rect 4415 -5589 4449 -5555
rect 4415 -5657 4449 -5623
rect 4415 -5725 4449 -5691
rect 4415 -5793 4449 -5759
rect 4415 -5861 4449 -5827
rect 4415 -5929 4449 -5895
rect 4415 -5997 4449 -5963
rect 4415 -6065 4449 -6031
rect 4415 -6133 4449 -6099
rect 4415 -6201 4449 -6167
rect 4415 -6269 4449 -6235
rect 4415 -6337 4449 -6303
rect 4415 -6405 4449 -6371
rect 6415 -5589 6449 -5555
rect 6415 -5657 6449 -5623
rect 6415 -5725 6449 -5691
rect 6415 -5793 6449 -5759
rect 6415 -5861 6449 -5827
rect 6415 -5929 6449 -5895
rect 6415 -5997 6449 -5963
rect 6415 -6065 6449 -6031
rect 6415 -6133 6449 -6099
rect 6415 -6201 6449 -6167
rect 6415 -6269 6449 -6235
rect 6415 -6337 6449 -6303
rect 6415 -6405 6449 -6371
rect 6869 -5641 6903 -5607
rect 6869 -5709 6903 -5675
rect 6869 -5777 6903 -5743
rect 6869 -5845 6903 -5811
rect 6869 -5913 6903 -5879
rect 6869 -5981 6903 -5947
rect 6869 -6049 6903 -6015
rect 6869 -6117 6903 -6083
rect 6869 -6185 6903 -6151
rect 6869 -6253 6903 -6219
rect 6869 -6321 6903 -6287
rect 6869 -6389 6903 -6355
rect 8869 -5641 8903 -5607
rect 8869 -5709 8903 -5675
rect 8869 -5777 8903 -5743
rect 8869 -5845 8903 -5811
rect 8869 -5913 8903 -5879
rect 8869 -5981 8903 -5947
rect 8869 -6049 8903 -6015
rect 8869 -6117 8903 -6083
rect 8869 -6185 8903 -6151
rect 8869 -6253 8903 -6219
rect 8869 -6321 8903 -6287
rect 8869 -6389 8903 -6355
<< nsubdiffcont >>
rect 4416 -4010 4450 -3976
rect 4416 -4078 4450 -4044
rect 4416 -4146 4450 -4112
rect 4416 -4214 4450 -4180
rect 4416 -4282 4450 -4248
rect 4416 -4350 4450 -4316
rect 4416 -4418 4450 -4384
rect 4416 -4486 4450 -4452
rect 4416 -4554 4450 -4520
rect 4416 -4622 4450 -4588
rect 4416 -4690 4450 -4656
rect 4416 -4758 4450 -4724
rect 4416 -4826 4450 -4792
rect 6416 -4010 6450 -3976
rect 6416 -4078 6450 -4044
rect 6416 -4146 6450 -4112
rect 6416 -4214 6450 -4180
rect 6416 -4282 6450 -4248
rect 6416 -4350 6450 -4316
rect 6416 -4418 6450 -4384
rect 6416 -4486 6450 -4452
rect 6416 -4554 6450 -4520
rect 6416 -4622 6450 -4588
rect 6416 -4690 6450 -4656
rect 6416 -4758 6450 -4724
rect 6416 -4826 6450 -4792
<< poly >>
rect 4613 -3743 4761 -3720
rect 4613 -3777 4636 -3743
rect 4670 -3777 4704 -3743
rect 4738 -3777 4761 -3743
rect 4613 -3800 4761 -3777
rect 4613 -3850 6253 -3800
rect 4613 -3900 4713 -3850
rect 4833 -3900 4933 -3850
rect 5053 -3900 5153 -3850
rect 5273 -3900 5373 -3850
rect 5493 -3900 5593 -3850
rect 5713 -3900 5813 -3850
rect 5933 -3900 6033 -3850
rect 6153 -3900 6253 -3850
rect 4613 -4900 4713 -4850
rect 4833 -4900 4933 -4850
rect 5053 -4900 5153 -4850
rect 5273 -4900 5373 -4850
rect 5493 -4900 5593 -4850
rect 5713 -4900 5813 -4850
rect 5933 -4900 6033 -4850
rect 6153 -4900 6253 -4850
rect 2158 -5446 2238 -5423
rect 2158 -5480 2181 -5446
rect 2215 -5480 2238 -5446
rect 2158 -5503 2238 -5480
rect 3038 -5446 3118 -5423
rect 3038 -5480 3061 -5446
rect 3095 -5480 3118 -5446
rect 3038 -5503 3118 -5480
rect 4612 -5455 5372 -5425
rect 2158 -5533 2918 -5503
rect 2158 -5583 2258 -5533
rect 2378 -5583 2478 -5533
rect 2598 -5583 2698 -5533
rect 2818 -5583 2918 -5533
rect 3038 -5533 3798 -5503
rect 4612 -5505 4712 -5455
rect 4832 -5505 4932 -5455
rect 5052 -5505 5152 -5455
rect 5272 -5505 5372 -5455
rect 5492 -5455 6252 -5425
rect 5492 -5505 5592 -5455
rect 5712 -5505 5812 -5455
rect 5932 -5505 6032 -5455
rect 6152 -5505 6252 -5455
rect 3038 -5583 3138 -5533
rect 3258 -5583 3358 -5533
rect 3478 -5583 3578 -5533
rect 3698 -5583 3798 -5533
rect 2158 -6517 2258 -6423
rect 2378 -6453 2478 -6423
rect 2598 -6453 2698 -6423
rect 2818 -6453 2918 -6423
rect 2168 -6540 2248 -6517
rect 2168 -6574 2191 -6540
rect 2225 -6574 2248 -6540
rect 2168 -6597 2248 -6574
rect 3038 -6613 3138 -6423
rect 3258 -6453 3358 -6423
rect 3478 -6453 3578 -6423
rect 3698 -6453 3798 -6423
rect 7066 -5533 7826 -5503
rect 7066 -5583 7166 -5533
rect 7286 -5583 7386 -5533
rect 7506 -5583 7606 -5533
rect 7726 -5583 7826 -5533
rect 7946 -5533 8706 -5503
rect 7946 -5583 8046 -5533
rect 8166 -5583 8266 -5533
rect 8386 -5583 8486 -5533
rect 8606 -5583 8706 -5533
rect 3048 -6622 3128 -6613
rect 3048 -6656 3071 -6622
rect 3105 -6656 3128 -6622
rect 3048 -6679 3128 -6656
rect 4612 -6763 4712 -6455
rect 4832 -6485 4932 -6455
rect 5052 -6485 5152 -6455
rect 5272 -6485 5372 -6455
rect 5492 -6485 5592 -6455
rect 5712 -6485 5812 -6455
rect 5932 -6485 6032 -6455
rect 6152 -6685 6252 -6455
rect 7066 -6599 7166 -6423
rect 7286 -6453 7386 -6423
rect 7506 -6453 7606 -6423
rect 7726 -6453 7826 -6423
rect 7946 -6517 8046 -6423
rect 8166 -6453 8266 -6423
rect 8386 -6453 8486 -6423
rect 8606 -6453 8706 -6423
rect 7953 -6540 8033 -6517
rect 7953 -6574 7976 -6540
rect 8010 -6574 8033 -6540
rect 7953 -6597 8033 -6574
rect 7076 -6622 7156 -6599
rect 7076 -6656 7099 -6622
rect 7133 -6656 7156 -6622
rect 7076 -6679 7156 -6656
rect 6161 -6704 6241 -6685
rect 6161 -6738 6184 -6704
rect 6218 -6738 6241 -6704
rect 6161 -6761 6241 -6738
rect 4622 -6786 4702 -6763
rect 4622 -6820 4645 -6786
rect 4679 -6820 4702 -6786
rect 4622 -6843 4702 -6820
<< polycont >>
rect 4636 -3777 4670 -3743
rect 4704 -3777 4738 -3743
rect 2181 -5480 2215 -5446
rect 3061 -5480 3095 -5446
rect 2191 -6574 2225 -6540
rect 3071 -6656 3105 -6622
rect 7976 -6574 8010 -6540
rect 7099 -6656 7133 -6622
rect 6184 -6738 6218 -6704
rect 4645 -6820 4679 -6786
<< xpolycontact >>
rect 2505 -4455 2575 -4023
rect 2505 -5025 2575 -4593
rect 8291 -4455 8361 -4023
rect 8291 -5025 8361 -4593
<< xpolyres >>
rect 2505 -4593 2575 -4455
rect 8291 -4593 8361 -4455
<< locali >>
rect -101 -3455 10466 -3432
rect -101 -3489 -40 -3455
rect -6 -3489 32 -3455
rect 66 -3489 104 -3455
rect 138 -3489 176 -3455
rect 210 -3489 248 -3455
rect 282 -3489 320 -3455
rect 354 -3489 392 -3455
rect 426 -3489 464 -3455
rect 498 -3489 536 -3455
rect 570 -3489 608 -3455
rect 642 -3489 680 -3455
rect 714 -3489 752 -3455
rect 786 -3489 824 -3455
rect 858 -3489 896 -3455
rect 930 -3489 968 -3455
rect 1002 -3489 1040 -3455
rect 1074 -3489 1112 -3455
rect 1146 -3489 1184 -3455
rect 1218 -3489 1279 -3455
rect 1313 -3489 1351 -3455
rect 1385 -3489 1423 -3455
rect 1457 -3489 1495 -3455
rect 1529 -3489 1567 -3455
rect 1601 -3489 1639 -3455
rect 1673 -3489 1711 -3455
rect 1745 -3489 1783 -3455
rect 1817 -3489 1855 -3455
rect 1889 -3489 1927 -3455
rect 1961 -3489 1999 -3455
rect 2033 -3489 2071 -3455
rect 2105 -3489 2143 -3455
rect 2177 -3489 2215 -3455
rect 2249 -3489 2287 -3455
rect 2321 -3489 2359 -3455
rect 2393 -3489 2431 -3455
rect 2465 -3489 2503 -3455
rect 2537 -3489 2575 -3455
rect 2609 -3489 2647 -3455
rect 2681 -3489 2719 -3455
rect 2753 -3489 2791 -3455
rect 2825 -3489 2863 -3455
rect 2897 -3489 2935 -3455
rect 2969 -3489 3007 -3455
rect 3041 -3489 3079 -3455
rect 3113 -3489 3151 -3455
rect 3185 -3489 3223 -3455
rect 3257 -3489 3295 -3455
rect 3329 -3489 3367 -3455
rect 3401 -3489 3439 -3455
rect 3473 -3489 3511 -3455
rect 3545 -3489 3583 -3455
rect 3617 -3489 3655 -3455
rect 3689 -3489 3727 -3455
rect 3761 -3489 3799 -3455
rect 3833 -3489 3894 -3455
rect 3928 -3489 3966 -3455
rect 4000 -3489 4038 -3455
rect 4072 -3489 4110 -3455
rect 4144 -3489 4182 -3455
rect 4216 -3489 4254 -3455
rect 4288 -3489 4326 -3455
rect 4360 -3489 4398 -3455
rect 4432 -3489 4470 -3455
rect 4504 -3489 4542 -3455
rect 4576 -3489 4614 -3455
rect 4648 -3489 4686 -3455
rect 4720 -3489 4758 -3455
rect 4792 -3489 4830 -3455
rect 4864 -3489 4902 -3455
rect 4936 -3489 4974 -3455
rect 5008 -3489 5046 -3455
rect 5080 -3489 5118 -3455
rect 5152 -3489 5190 -3455
rect 5224 -3489 5262 -3455
rect 5296 -3489 5334 -3455
rect 5368 -3489 5406 -3455
rect 5440 -3489 5478 -3455
rect 5512 -3489 5550 -3455
rect 5584 -3489 5622 -3455
rect 5656 -3489 5694 -3455
rect 5728 -3489 5766 -3455
rect 5800 -3489 5838 -3455
rect 5872 -3489 5910 -3455
rect 5944 -3489 5982 -3455
rect 6016 -3489 6054 -3455
rect 6088 -3489 6126 -3455
rect 6160 -3489 6198 -3455
rect 6232 -3489 6270 -3455
rect 6304 -3489 6342 -3455
rect 6376 -3489 6414 -3455
rect 6448 -3489 6509 -3455
rect 6543 -3489 6581 -3455
rect 6615 -3489 6653 -3455
rect 6687 -3489 6725 -3455
rect 6759 -3489 6797 -3455
rect 6831 -3489 6869 -3455
rect 6903 -3489 6941 -3455
rect 6975 -3489 7013 -3455
rect 7047 -3489 7085 -3455
rect 7119 -3489 7157 -3455
rect 7191 -3489 7229 -3455
rect 7263 -3489 7301 -3455
rect 7335 -3489 7373 -3455
rect 7407 -3489 7445 -3455
rect 7479 -3489 7517 -3455
rect 7551 -3489 7589 -3455
rect 7623 -3489 7661 -3455
rect 7695 -3489 7733 -3455
rect 7767 -3489 7805 -3455
rect 7839 -3489 7877 -3455
rect 7911 -3489 7949 -3455
rect 7983 -3489 8021 -3455
rect 8055 -3489 8093 -3455
rect 8127 -3489 8165 -3455
rect 8199 -3489 8237 -3455
rect 8271 -3489 8309 -3455
rect 8343 -3489 8381 -3455
rect 8415 -3489 8453 -3455
rect 8487 -3489 8525 -3455
rect 8559 -3489 8597 -3455
rect 8631 -3489 8669 -3455
rect 8703 -3489 8741 -3455
rect 8775 -3489 8813 -3455
rect 8847 -3489 8885 -3455
rect 8919 -3489 8957 -3455
rect 8991 -3489 9029 -3455
rect 9063 -3489 9124 -3455
rect 9158 -3489 9196 -3455
rect 9230 -3489 9268 -3455
rect 9302 -3489 9340 -3455
rect 9374 -3489 9412 -3455
rect 9446 -3489 9484 -3455
rect 9518 -3489 9556 -3455
rect 9590 -3489 9628 -3455
rect 9662 -3489 9700 -3455
rect 9734 -3489 9772 -3455
rect 9806 -3489 9844 -3455
rect 9878 -3489 9916 -3455
rect 9950 -3489 9988 -3455
rect 10022 -3489 10060 -3455
rect 10094 -3489 10132 -3455
rect 10166 -3489 10204 -3455
rect 10238 -3489 10276 -3455
rect 10310 -3489 10348 -3455
rect 10382 -3489 10466 -3455
rect -101 -3512 10466 -3489
rect 2184 -3743 4761 -3720
rect 2184 -3777 2207 -3743
rect 2241 -3777 4636 -3743
rect 4670 -3777 4704 -3743
rect 4738 -3777 4761 -3743
rect 2184 -3800 4761 -3777
rect 5360 -3840 5508 -3512
rect 4534 -3880 6333 -3840
rect 4534 -3920 4574 -3880
rect 4973 -3920 5013 -3880
rect 4393 -3976 4593 -3920
rect 4393 -4010 4416 -3976
rect 4450 -4010 4536 -3976
rect 4570 -4010 4593 -3976
rect 4393 -4044 4593 -4010
rect 4393 -4078 4416 -4044
rect 4450 -4078 4536 -4044
rect 4570 -4078 4593 -4044
rect 4393 -4112 4593 -4078
rect 4393 -4146 4416 -4112
rect 4450 -4146 4536 -4112
rect 4570 -4146 4593 -4112
rect 4393 -4180 4593 -4146
rect 4393 -4214 4416 -4180
rect 4450 -4214 4536 -4180
rect 4570 -4214 4593 -4180
rect 4393 -4248 4593 -4214
rect 4393 -4282 4416 -4248
rect 4450 -4282 4536 -4248
rect 4570 -4282 4593 -4248
rect 4393 -4316 4593 -4282
rect 4393 -4350 4416 -4316
rect 4450 -4350 4536 -4316
rect 4570 -4350 4593 -4316
rect 4393 -4384 4593 -4350
rect 4393 -4418 4416 -4384
rect 4450 -4418 4536 -4384
rect 4570 -4418 4593 -4384
rect 4393 -4452 4593 -4418
rect 4393 -4486 4416 -4452
rect 4450 -4486 4536 -4452
rect 4570 -4486 4593 -4452
rect 4393 -4520 4593 -4486
rect 4393 -4554 4416 -4520
rect 4450 -4554 4536 -4520
rect 4570 -4554 4593 -4520
rect 4393 -4588 4593 -4554
rect 4393 -4622 4416 -4588
rect 4450 -4622 4536 -4588
rect 4570 -4622 4593 -4588
rect 4393 -4656 4593 -4622
rect 4393 -4690 4416 -4656
rect 4450 -4690 4536 -4656
rect 4570 -4690 4593 -4656
rect 4393 -4724 4593 -4690
rect 4393 -4758 4416 -4724
rect 4450 -4758 4536 -4724
rect 4570 -4758 4593 -4724
rect 4393 -4792 4593 -4758
rect 4393 -4826 4416 -4792
rect 4450 -4826 4536 -4792
rect 4570 -4826 4593 -4792
rect 4393 -4830 4593 -4826
rect 4733 -3976 4813 -3920
rect 4733 -4010 4756 -3976
rect 4790 -4010 4813 -3976
rect 4733 -4044 4813 -4010
rect 4733 -4078 4756 -4044
rect 4790 -4078 4813 -4044
rect 4733 -4112 4813 -4078
rect 4733 -4146 4756 -4112
rect 4790 -4146 4813 -4112
rect 4733 -4180 4813 -4146
rect 4733 -4214 4756 -4180
rect 4790 -4214 4813 -4180
rect 4733 -4248 4813 -4214
rect 4733 -4282 4756 -4248
rect 4790 -4282 4813 -4248
rect 4733 -4316 4813 -4282
rect 4733 -4350 4756 -4316
rect 4790 -4350 4813 -4316
rect 4733 -4384 4813 -4350
rect 4733 -4418 4756 -4384
rect 4790 -4418 4813 -4384
rect 4733 -4452 4813 -4418
rect 4733 -4486 4756 -4452
rect 4790 -4486 4813 -4452
rect 4733 -4520 4813 -4486
rect 4733 -4554 4756 -4520
rect 4790 -4554 4813 -4520
rect 4733 -4588 4813 -4554
rect 4733 -4622 4756 -4588
rect 4790 -4622 4813 -4588
rect 4733 -4656 4813 -4622
rect 4733 -4690 4756 -4656
rect 4790 -4690 4813 -4656
rect 4733 -4724 4813 -4690
rect 4733 -4758 4756 -4724
rect 4790 -4758 4813 -4724
rect 4733 -4792 4813 -4758
rect 4733 -4826 4756 -4792
rect 4790 -4826 4813 -4792
rect 4733 -4830 4813 -4826
rect 4953 -3976 5033 -3920
rect 4953 -4010 4976 -3976
rect 5010 -4010 5033 -3976
rect 4953 -4044 5033 -4010
rect 4953 -4078 4976 -4044
rect 5010 -4078 5033 -4044
rect 4953 -4112 5033 -4078
rect 4953 -4146 4976 -4112
rect 5010 -4146 5033 -4112
rect 4953 -4180 5033 -4146
rect 4953 -4214 4976 -4180
rect 5010 -4214 5033 -4180
rect 4953 -4248 5033 -4214
rect 4953 -4282 4976 -4248
rect 5010 -4282 5033 -4248
rect 4953 -4316 5033 -4282
rect 4953 -4350 4976 -4316
rect 5010 -4350 5033 -4316
rect 4953 -4384 5033 -4350
rect 4953 -4418 4976 -4384
rect 5010 -4418 5033 -4384
rect 4953 -4452 5033 -4418
rect 4953 -4486 4976 -4452
rect 5010 -4486 5033 -4452
rect 4953 -4520 5033 -4486
rect 4953 -4554 4976 -4520
rect 5010 -4554 5033 -4520
rect 4953 -4588 5033 -4554
rect 4953 -4622 4976 -4588
rect 5010 -4622 5033 -4588
rect 4953 -4656 5033 -4622
rect 4953 -4690 4976 -4656
rect 5010 -4690 5033 -4656
rect 4953 -4724 5033 -4690
rect 4953 -4758 4976 -4724
rect 5010 -4758 5033 -4724
rect 4953 -4792 5033 -4758
rect 4953 -4826 4976 -4792
rect 5010 -4826 5033 -4792
rect 4953 -4830 5033 -4826
rect 5173 -3976 5253 -3920
rect 5360 -3950 5508 -3880
rect 5853 -3920 5893 -3880
rect 6293 -3920 6333 -3880
rect 5173 -4010 5196 -3976
rect 5230 -4010 5253 -3976
rect 5173 -4044 5253 -4010
rect 5173 -4078 5196 -4044
rect 5230 -4078 5253 -4044
rect 5173 -4112 5253 -4078
rect 5173 -4146 5196 -4112
rect 5230 -4146 5253 -4112
rect 5173 -4180 5253 -4146
rect 5173 -4214 5196 -4180
rect 5230 -4214 5253 -4180
rect 5173 -4248 5253 -4214
rect 5173 -4282 5196 -4248
rect 5230 -4282 5253 -4248
rect 5173 -4316 5253 -4282
rect 5173 -4350 5196 -4316
rect 5230 -4350 5253 -4316
rect 5173 -4384 5253 -4350
rect 5173 -4418 5196 -4384
rect 5230 -4418 5253 -4384
rect 5173 -4452 5253 -4418
rect 5173 -4486 5196 -4452
rect 5230 -4486 5253 -4452
rect 5173 -4520 5253 -4486
rect 5173 -4554 5196 -4520
rect 5230 -4554 5253 -4520
rect 5173 -4588 5253 -4554
rect 5173 -4622 5196 -4588
rect 5230 -4622 5253 -4588
rect 5173 -4656 5253 -4622
rect 5173 -4690 5196 -4656
rect 5230 -4690 5253 -4656
rect 5173 -4724 5253 -4690
rect 5173 -4758 5196 -4724
rect 5230 -4758 5253 -4724
rect 5173 -4792 5253 -4758
rect 5173 -4826 5196 -4792
rect 5230 -4826 5253 -4792
rect 5173 -4830 5253 -4826
rect 5393 -3976 5473 -3950
rect 5393 -4010 5416 -3976
rect 5450 -4010 5473 -3976
rect 5393 -4044 5473 -4010
rect 5393 -4078 5416 -4044
rect 5450 -4078 5473 -4044
rect 5393 -4112 5473 -4078
rect 5393 -4146 5416 -4112
rect 5450 -4146 5473 -4112
rect 5393 -4180 5473 -4146
rect 5393 -4214 5416 -4180
rect 5450 -4214 5473 -4180
rect 5393 -4248 5473 -4214
rect 5393 -4282 5416 -4248
rect 5450 -4282 5473 -4248
rect 5393 -4316 5473 -4282
rect 5393 -4350 5416 -4316
rect 5450 -4350 5473 -4316
rect 5393 -4384 5473 -4350
rect 5393 -4418 5416 -4384
rect 5450 -4418 5473 -4384
rect 5393 -4452 5473 -4418
rect 5393 -4486 5416 -4452
rect 5450 -4486 5473 -4452
rect 5393 -4520 5473 -4486
rect 5393 -4554 5416 -4520
rect 5450 -4554 5473 -4520
rect 5393 -4588 5473 -4554
rect 5393 -4622 5416 -4588
rect 5450 -4622 5473 -4588
rect 5393 -4656 5473 -4622
rect 5393 -4690 5416 -4656
rect 5450 -4690 5473 -4656
rect 5393 -4724 5473 -4690
rect 5393 -4758 5416 -4724
rect 5450 -4758 5473 -4724
rect 5393 -4792 5473 -4758
rect 5393 -4826 5416 -4792
rect 5450 -4826 5473 -4792
rect 5393 -4830 5473 -4826
rect 5613 -3976 5693 -3920
rect 5613 -4010 5636 -3976
rect 5670 -4010 5693 -3976
rect 5613 -4044 5693 -4010
rect 5613 -4078 5636 -4044
rect 5670 -4078 5693 -4044
rect 5613 -4112 5693 -4078
rect 5613 -4146 5636 -4112
rect 5670 -4146 5693 -4112
rect 5613 -4180 5693 -4146
rect 5613 -4214 5636 -4180
rect 5670 -4214 5693 -4180
rect 5613 -4248 5693 -4214
rect 5613 -4282 5636 -4248
rect 5670 -4282 5693 -4248
rect 5613 -4316 5693 -4282
rect 5613 -4350 5636 -4316
rect 5670 -4350 5693 -4316
rect 5613 -4384 5693 -4350
rect 5613 -4418 5636 -4384
rect 5670 -4418 5693 -4384
rect 5613 -4452 5693 -4418
rect 5613 -4486 5636 -4452
rect 5670 -4486 5693 -4452
rect 5613 -4520 5693 -4486
rect 5613 -4554 5636 -4520
rect 5670 -4554 5693 -4520
rect 5613 -4588 5693 -4554
rect 5613 -4622 5636 -4588
rect 5670 -4622 5693 -4588
rect 5613 -4656 5693 -4622
rect 5613 -4690 5636 -4656
rect 5670 -4690 5693 -4656
rect 5613 -4724 5693 -4690
rect 5613 -4758 5636 -4724
rect 5670 -4758 5693 -4724
rect 5613 -4792 5693 -4758
rect 5613 -4826 5636 -4792
rect 5670 -4826 5693 -4792
rect 5613 -4830 5693 -4826
rect 5833 -3976 5913 -3920
rect 5833 -4010 5856 -3976
rect 5890 -4010 5913 -3976
rect 5833 -4044 5913 -4010
rect 5833 -4078 5856 -4044
rect 5890 -4078 5913 -4044
rect 5833 -4112 5913 -4078
rect 5833 -4146 5856 -4112
rect 5890 -4146 5913 -4112
rect 5833 -4180 5913 -4146
rect 5833 -4214 5856 -4180
rect 5890 -4214 5913 -4180
rect 5833 -4248 5913 -4214
rect 5833 -4282 5856 -4248
rect 5890 -4282 5913 -4248
rect 5833 -4316 5913 -4282
rect 5833 -4350 5856 -4316
rect 5890 -4350 5913 -4316
rect 5833 -4384 5913 -4350
rect 5833 -4418 5856 -4384
rect 5890 -4418 5913 -4384
rect 5833 -4452 5913 -4418
rect 5833 -4486 5856 -4452
rect 5890 -4486 5913 -4452
rect 5833 -4520 5913 -4486
rect 5833 -4554 5856 -4520
rect 5890 -4554 5913 -4520
rect 5833 -4588 5913 -4554
rect 5833 -4622 5856 -4588
rect 5890 -4622 5913 -4588
rect 5833 -4656 5913 -4622
rect 5833 -4690 5856 -4656
rect 5890 -4690 5913 -4656
rect 5833 -4724 5913 -4690
rect 5833 -4758 5856 -4724
rect 5890 -4758 5913 -4724
rect 5833 -4792 5913 -4758
rect 5833 -4826 5856 -4792
rect 5890 -4826 5913 -4792
rect 5833 -4830 5913 -4826
rect 6053 -3976 6133 -3920
rect 6053 -4010 6076 -3976
rect 6110 -4010 6133 -3976
rect 6053 -4044 6133 -4010
rect 6053 -4078 6076 -4044
rect 6110 -4078 6133 -4044
rect 6053 -4112 6133 -4078
rect 6053 -4146 6076 -4112
rect 6110 -4146 6133 -4112
rect 6053 -4180 6133 -4146
rect 6053 -4214 6076 -4180
rect 6110 -4214 6133 -4180
rect 6053 -4248 6133 -4214
rect 6053 -4282 6076 -4248
rect 6110 -4282 6133 -4248
rect 6053 -4316 6133 -4282
rect 6053 -4350 6076 -4316
rect 6110 -4350 6133 -4316
rect 6053 -4384 6133 -4350
rect 6053 -4418 6076 -4384
rect 6110 -4418 6133 -4384
rect 6053 -4452 6133 -4418
rect 6053 -4486 6076 -4452
rect 6110 -4486 6133 -4452
rect 6053 -4520 6133 -4486
rect 6053 -4554 6076 -4520
rect 6110 -4554 6133 -4520
rect 6053 -4588 6133 -4554
rect 6053 -4622 6076 -4588
rect 6110 -4622 6133 -4588
rect 6053 -4656 6133 -4622
rect 6053 -4690 6076 -4656
rect 6110 -4690 6133 -4656
rect 6053 -4724 6133 -4690
rect 6053 -4758 6076 -4724
rect 6110 -4758 6133 -4724
rect 6053 -4792 6133 -4758
rect 6053 -4826 6076 -4792
rect 6110 -4826 6133 -4792
rect 6053 -4830 6133 -4826
rect 6273 -3976 6473 -3920
rect 6273 -4010 6296 -3976
rect 6330 -4010 6416 -3976
rect 6450 -4010 6473 -3976
rect 6273 -4044 6473 -4010
rect 6273 -4078 6296 -4044
rect 6330 -4078 6416 -4044
rect 6450 -4078 6473 -4044
rect 6273 -4112 6473 -4078
rect 6273 -4146 6296 -4112
rect 6330 -4146 6416 -4112
rect 6450 -4146 6473 -4112
rect 6273 -4180 6473 -4146
rect 6273 -4214 6296 -4180
rect 6330 -4214 6416 -4180
rect 6450 -4214 6473 -4180
rect 6273 -4248 6473 -4214
rect 6273 -4282 6296 -4248
rect 6330 -4282 6416 -4248
rect 6450 -4282 6473 -4248
rect 6273 -4316 6473 -4282
rect 6273 -4350 6296 -4316
rect 6330 -4350 6416 -4316
rect 6450 -4350 6473 -4316
rect 6273 -4384 6473 -4350
rect 6273 -4418 6296 -4384
rect 6330 -4418 6416 -4384
rect 6450 -4418 6473 -4384
rect 6273 -4452 6473 -4418
rect 6273 -4486 6296 -4452
rect 6330 -4486 6416 -4452
rect 6450 -4486 6473 -4452
rect 6273 -4520 6473 -4486
rect 6273 -4554 6296 -4520
rect 6330 -4554 6416 -4520
rect 6450 -4554 6473 -4520
rect 6273 -4588 6473 -4554
rect 6273 -4622 6296 -4588
rect 6330 -4622 6416 -4588
rect 6450 -4622 6473 -4588
rect 6273 -4656 6473 -4622
rect 6273 -4690 6296 -4656
rect 6330 -4690 6416 -4656
rect 6450 -4690 6473 -4656
rect 6273 -4724 6473 -4690
rect 6273 -4758 6296 -4724
rect 6330 -4758 6416 -4724
rect 6450 -4758 6473 -4724
rect 6273 -4792 6473 -4758
rect 6273 -4826 6296 -4792
rect 6330 -4826 6416 -4792
rect 6450 -4826 6473 -4792
rect 6273 -4830 6473 -4826
rect 4753 -4870 4793 -4830
rect 5193 -4870 5233 -4830
rect 4753 -4910 5233 -4870
rect 5633 -4870 5673 -4830
rect 6073 -4870 6113 -4830
rect 5633 -4910 6113 -4870
rect 2505 -5123 2575 -5025
rect 2500 -5146 2580 -5123
rect 2500 -5180 2523 -5146
rect 2557 -5180 2580 -5146
rect 2500 -5203 2580 -5180
rect 2505 -5341 2575 -5203
rect 3578 -5256 3658 -5233
rect 3578 -5290 3601 -5256
rect 3635 -5290 3658 -5256
rect 2500 -5364 2580 -5341
rect 2500 -5398 2523 -5364
rect 2557 -5398 2580 -5364
rect 2500 -5421 2580 -5398
rect 2158 -5446 2238 -5423
rect 2158 -5480 2181 -5446
rect 2215 -5480 2238 -5446
rect 2158 -5503 2238 -5480
rect 2505 -5523 2575 -5421
rect 3038 -5446 3118 -5423
rect 3038 -5480 3061 -5446
rect 3095 -5480 3118 -5446
rect 3038 -5503 3118 -5480
rect 3578 -5523 3658 -5290
rect 4960 -5445 5028 -4910
rect 5839 -5445 5907 -4910
rect 8291 -5233 8361 -5025
rect 8286 -5256 8366 -5233
rect 8286 -5290 8309 -5256
rect 8343 -5290 8366 -5256
rect 8286 -5313 8366 -5290
rect 7206 -5364 7286 -5341
rect 7206 -5398 7229 -5364
rect 7263 -5398 7286 -5364
rect 2298 -5563 2778 -5523
rect 2298 -5603 2338 -5563
rect 2738 -5603 2778 -5563
rect 3178 -5563 3658 -5523
rect 3178 -5603 3218 -5563
rect 3618 -5603 3658 -5563
rect 3841 -5479 5232 -5445
rect 3841 -5603 3875 -5479
rect 4752 -5485 5232 -5479
rect 4752 -5525 4792 -5485
rect 5192 -5525 5232 -5485
rect 5632 -5479 7023 -5445
rect 5632 -5485 6112 -5479
rect 5632 -5525 5672 -5485
rect 6072 -5525 6112 -5485
rect 4392 -5555 4592 -5525
rect 4392 -5589 4415 -5555
rect 4449 -5589 4535 -5555
rect 4569 -5589 4592 -5555
rect 1938 -5607 2018 -5603
rect 1938 -5641 1961 -5607
rect 1995 -5641 2018 -5607
rect 1938 -5675 2018 -5641
rect 1938 -5709 1961 -5675
rect 1995 -5709 2018 -5675
rect 1938 -5743 2018 -5709
rect 1938 -5777 1961 -5743
rect 1995 -5777 2018 -5743
rect 1938 -5811 2018 -5777
rect 1938 -5845 1961 -5811
rect 1995 -5845 2018 -5811
rect 1938 -5879 2018 -5845
rect 1938 -5913 1961 -5879
rect 1995 -5913 2018 -5879
rect 1938 -5947 2018 -5913
rect 1938 -5981 1961 -5947
rect 1995 -5981 2018 -5947
rect 1938 -6015 2018 -5981
rect 1938 -6049 1961 -6015
rect 1995 -6049 2018 -6015
rect 1938 -6083 2018 -6049
rect 1938 -6117 1961 -6083
rect 1995 -6117 2018 -6083
rect 1938 -6151 2018 -6117
rect 1938 -6185 1961 -6151
rect 1995 -6185 2018 -6151
rect 1938 -6219 2018 -6185
rect 1938 -6253 1961 -6219
rect 1995 -6253 2018 -6219
rect 1938 -6287 2018 -6253
rect 1938 -6321 1961 -6287
rect 1995 -6321 2018 -6287
rect 1938 -6355 2018 -6321
rect 1938 -6389 1961 -6355
rect 1995 -6389 2018 -6355
rect 1938 -6968 2018 -6389
rect 2058 -5607 2138 -5603
rect 2058 -5641 2081 -5607
rect 2115 -5641 2138 -5607
rect 2058 -5675 2138 -5641
rect 2058 -5709 2081 -5675
rect 2115 -5709 2138 -5675
rect 2058 -5743 2138 -5709
rect 2058 -5777 2081 -5743
rect 2115 -5777 2138 -5743
rect 2058 -5811 2138 -5777
rect 2058 -5845 2081 -5811
rect 2115 -5845 2138 -5811
rect 2058 -5879 2138 -5845
rect 2058 -5913 2081 -5879
rect 2115 -5913 2138 -5879
rect 2058 -5947 2138 -5913
rect 2058 -5981 2081 -5947
rect 2115 -5981 2138 -5947
rect 2058 -6015 2138 -5981
rect 2058 -6049 2081 -6015
rect 2115 -6049 2138 -6015
rect 2058 -6083 2138 -6049
rect 2058 -6117 2081 -6083
rect 2115 -6117 2138 -6083
rect 2058 -6151 2138 -6117
rect 2058 -6185 2081 -6151
rect 2115 -6185 2138 -6151
rect 2058 -6219 2138 -6185
rect 2058 -6253 2081 -6219
rect 2115 -6253 2138 -6219
rect 2058 -6287 2138 -6253
rect 2058 -6321 2081 -6287
rect 2115 -6321 2138 -6287
rect 2058 -6355 2138 -6321
rect 2058 -6389 2081 -6355
rect 2115 -6389 2138 -6355
rect 2058 -6403 2138 -6389
rect 2278 -5607 2358 -5603
rect 2278 -5641 2301 -5607
rect 2335 -5641 2358 -5607
rect 2278 -5675 2358 -5641
rect 2278 -5709 2301 -5675
rect 2335 -5709 2358 -5675
rect 2278 -5743 2358 -5709
rect 2278 -5777 2301 -5743
rect 2335 -5777 2358 -5743
rect 2278 -5811 2358 -5777
rect 2278 -5845 2301 -5811
rect 2335 -5845 2358 -5811
rect 2278 -5879 2358 -5845
rect 2278 -5913 2301 -5879
rect 2335 -5913 2358 -5879
rect 2278 -5947 2358 -5913
rect 2278 -5981 2301 -5947
rect 2335 -5981 2358 -5947
rect 2278 -6015 2358 -5981
rect 2278 -6049 2301 -6015
rect 2335 -6049 2358 -6015
rect 2278 -6083 2358 -6049
rect 2278 -6117 2301 -6083
rect 2335 -6117 2358 -6083
rect 2278 -6151 2358 -6117
rect 2278 -6185 2301 -6151
rect 2335 -6185 2358 -6151
rect 2278 -6219 2358 -6185
rect 2278 -6253 2301 -6219
rect 2335 -6253 2358 -6219
rect 2278 -6287 2358 -6253
rect 2278 -6321 2301 -6287
rect 2335 -6321 2358 -6287
rect 2278 -6355 2358 -6321
rect 2278 -6389 2301 -6355
rect 2335 -6389 2358 -6355
rect 2278 -6403 2358 -6389
rect 2498 -5607 2578 -5603
rect 2498 -5641 2521 -5607
rect 2555 -5641 2578 -5607
rect 2498 -5675 2578 -5641
rect 2498 -5709 2521 -5675
rect 2555 -5709 2578 -5675
rect 2498 -5743 2578 -5709
rect 2498 -5777 2521 -5743
rect 2555 -5777 2578 -5743
rect 2498 -5811 2578 -5777
rect 2498 -5845 2521 -5811
rect 2555 -5845 2578 -5811
rect 2498 -5879 2578 -5845
rect 2498 -5913 2521 -5879
rect 2555 -5913 2578 -5879
rect 2498 -5947 2578 -5913
rect 2498 -5981 2521 -5947
rect 2555 -5981 2578 -5947
rect 2498 -6015 2578 -5981
rect 2498 -6049 2521 -6015
rect 2555 -6049 2578 -6015
rect 2498 -6083 2578 -6049
rect 2498 -6117 2521 -6083
rect 2555 -6117 2578 -6083
rect 2498 -6151 2578 -6117
rect 2498 -6185 2521 -6151
rect 2555 -6185 2578 -6151
rect 2498 -6219 2578 -6185
rect 2498 -6253 2521 -6219
rect 2555 -6253 2578 -6219
rect 2498 -6287 2578 -6253
rect 2498 -6321 2521 -6287
rect 2555 -6321 2578 -6287
rect 2498 -6355 2578 -6321
rect 2498 -6389 2521 -6355
rect 2555 -6389 2578 -6355
rect 2498 -6403 2578 -6389
rect 2718 -5607 2798 -5603
rect 2718 -5641 2741 -5607
rect 2775 -5641 2798 -5607
rect 2718 -5675 2798 -5641
rect 2718 -5709 2741 -5675
rect 2775 -5709 2798 -5675
rect 2718 -5743 2798 -5709
rect 2718 -5777 2741 -5743
rect 2775 -5777 2798 -5743
rect 2718 -5811 2798 -5777
rect 2718 -5845 2741 -5811
rect 2775 -5845 2798 -5811
rect 2718 -5879 2798 -5845
rect 2718 -5913 2741 -5879
rect 2775 -5913 2798 -5879
rect 2718 -5947 2798 -5913
rect 2718 -5981 2741 -5947
rect 2775 -5981 2798 -5947
rect 2718 -6015 2798 -5981
rect 2718 -6049 2741 -6015
rect 2775 -6049 2798 -6015
rect 2718 -6083 2798 -6049
rect 2718 -6117 2741 -6083
rect 2775 -6117 2798 -6083
rect 2718 -6151 2798 -6117
rect 2718 -6185 2741 -6151
rect 2775 -6185 2798 -6151
rect 2718 -6219 2798 -6185
rect 2718 -6253 2741 -6219
rect 2775 -6253 2798 -6219
rect 2718 -6287 2798 -6253
rect 2718 -6321 2741 -6287
rect 2775 -6321 2798 -6287
rect 2718 -6355 2798 -6321
rect 2718 -6389 2741 -6355
rect 2775 -6389 2798 -6355
rect 2718 -6403 2798 -6389
rect 2938 -5607 3018 -5603
rect 2938 -5641 2961 -5607
rect 2995 -5641 3018 -5607
rect 2938 -5675 3018 -5641
rect 2938 -5709 2961 -5675
rect 2995 -5709 3018 -5675
rect 2938 -5743 3018 -5709
rect 2938 -5777 2961 -5743
rect 2995 -5777 3018 -5743
rect 2938 -5811 3018 -5777
rect 2938 -5845 2961 -5811
rect 2995 -5845 3018 -5811
rect 2938 -5879 3018 -5845
rect 2938 -5913 2961 -5879
rect 2995 -5913 3018 -5879
rect 2938 -5947 3018 -5913
rect 2938 -5981 2961 -5947
rect 2995 -5981 3018 -5947
rect 2938 -6015 3018 -5981
rect 2938 -6049 2961 -6015
rect 2995 -6049 3018 -6015
rect 2938 -6083 3018 -6049
rect 2938 -6117 2961 -6083
rect 2995 -6117 3018 -6083
rect 2938 -6151 3018 -6117
rect 2938 -6185 2961 -6151
rect 2995 -6185 3018 -6151
rect 2938 -6219 3018 -6185
rect 2938 -6253 2961 -6219
rect 2995 -6253 3018 -6219
rect 2938 -6287 3018 -6253
rect 2938 -6321 2961 -6287
rect 2995 -6321 3018 -6287
rect 2938 -6355 3018 -6321
rect 2938 -6389 2961 -6355
rect 2995 -6389 3018 -6355
rect 2938 -6403 3018 -6389
rect 3158 -5607 3238 -5603
rect 3158 -5641 3181 -5607
rect 3215 -5641 3238 -5607
rect 3158 -5675 3238 -5641
rect 3158 -5709 3181 -5675
rect 3215 -5709 3238 -5675
rect 3158 -5743 3238 -5709
rect 3158 -5777 3181 -5743
rect 3215 -5777 3238 -5743
rect 3158 -5811 3238 -5777
rect 3158 -5845 3181 -5811
rect 3215 -5845 3238 -5811
rect 3158 -5879 3238 -5845
rect 3158 -5913 3181 -5879
rect 3215 -5913 3238 -5879
rect 3158 -5947 3238 -5913
rect 3158 -5981 3181 -5947
rect 3215 -5981 3238 -5947
rect 3158 -6015 3238 -5981
rect 3158 -6049 3181 -6015
rect 3215 -6049 3238 -6015
rect 3158 -6083 3238 -6049
rect 3158 -6117 3181 -6083
rect 3215 -6117 3238 -6083
rect 3158 -6151 3238 -6117
rect 3158 -6185 3181 -6151
rect 3215 -6185 3238 -6151
rect 3158 -6219 3238 -6185
rect 3158 -6253 3181 -6219
rect 3215 -6253 3238 -6219
rect 3158 -6287 3238 -6253
rect 3158 -6321 3181 -6287
rect 3215 -6321 3238 -6287
rect 3158 -6355 3238 -6321
rect 3158 -6389 3181 -6355
rect 3215 -6389 3238 -6355
rect 3158 -6403 3238 -6389
rect 3378 -5607 3458 -5603
rect 3378 -5641 3401 -5607
rect 3435 -5641 3458 -5607
rect 3378 -5675 3458 -5641
rect 3378 -5709 3401 -5675
rect 3435 -5709 3458 -5675
rect 3378 -5743 3458 -5709
rect 3378 -5777 3401 -5743
rect 3435 -5777 3458 -5743
rect 3378 -5811 3458 -5777
rect 3378 -5845 3401 -5811
rect 3435 -5845 3458 -5811
rect 3378 -5879 3458 -5845
rect 3378 -5913 3401 -5879
rect 3435 -5913 3458 -5879
rect 3378 -5947 3458 -5913
rect 3378 -5981 3401 -5947
rect 3435 -5981 3458 -5947
rect 3378 -6015 3458 -5981
rect 3378 -6049 3401 -6015
rect 3435 -6049 3458 -6015
rect 3378 -6083 3458 -6049
rect 3378 -6117 3401 -6083
rect 3435 -6117 3458 -6083
rect 3378 -6151 3458 -6117
rect 3378 -6185 3401 -6151
rect 3435 -6185 3458 -6151
rect 3378 -6219 3458 -6185
rect 3378 -6253 3401 -6219
rect 3435 -6253 3458 -6219
rect 3378 -6287 3458 -6253
rect 3378 -6321 3401 -6287
rect 3435 -6321 3458 -6287
rect 3378 -6355 3458 -6321
rect 3378 -6389 3401 -6355
rect 3435 -6389 3458 -6355
rect 3378 -6403 3458 -6389
rect 3598 -5607 3678 -5603
rect 3598 -5641 3621 -5607
rect 3655 -5641 3678 -5607
rect 3598 -5675 3678 -5641
rect 3598 -5709 3621 -5675
rect 3655 -5709 3678 -5675
rect 3598 -5743 3678 -5709
rect 3598 -5777 3621 -5743
rect 3655 -5777 3678 -5743
rect 3598 -5811 3678 -5777
rect 3598 -5845 3621 -5811
rect 3655 -5845 3678 -5811
rect 3598 -5879 3678 -5845
rect 3598 -5913 3621 -5879
rect 3655 -5913 3678 -5879
rect 3598 -5947 3678 -5913
rect 3598 -5981 3621 -5947
rect 3655 -5981 3678 -5947
rect 3598 -6015 3678 -5981
rect 3598 -6049 3621 -6015
rect 3655 -6049 3678 -6015
rect 3598 -6083 3678 -6049
rect 3598 -6117 3621 -6083
rect 3655 -6117 3678 -6083
rect 3598 -6151 3678 -6117
rect 3598 -6185 3621 -6151
rect 3655 -6185 3678 -6151
rect 3598 -6219 3678 -6185
rect 3598 -6253 3621 -6219
rect 3655 -6253 3678 -6219
rect 3598 -6287 3678 -6253
rect 3598 -6321 3621 -6287
rect 3655 -6321 3678 -6287
rect 3598 -6355 3678 -6321
rect 3598 -6389 3621 -6355
rect 3655 -6389 3678 -6355
rect 3598 -6403 3678 -6389
rect 3818 -5607 3898 -5603
rect 3818 -5641 3841 -5607
rect 3875 -5641 3898 -5607
rect 3818 -5675 3898 -5641
rect 3818 -5709 3841 -5675
rect 3875 -5709 3898 -5675
rect 3818 -5743 3898 -5709
rect 3818 -5777 3841 -5743
rect 3875 -5777 3898 -5743
rect 3818 -5811 3898 -5777
rect 3818 -5845 3841 -5811
rect 3875 -5845 3898 -5811
rect 3818 -5879 3898 -5845
rect 3818 -5913 3841 -5879
rect 3875 -5913 3898 -5879
rect 3818 -5947 3898 -5913
rect 3818 -5981 3841 -5947
rect 3875 -5981 3898 -5947
rect 3818 -6015 3898 -5981
rect 3818 -6049 3841 -6015
rect 3875 -6049 3898 -6015
rect 3818 -6083 3898 -6049
rect 3818 -6117 3841 -6083
rect 3875 -6117 3898 -6083
rect 3818 -6151 3898 -6117
rect 3818 -6185 3841 -6151
rect 3875 -6185 3898 -6151
rect 3818 -6219 3898 -6185
rect 3818 -6253 3841 -6219
rect 3875 -6253 3898 -6219
rect 3818 -6287 3898 -6253
rect 3818 -6321 3841 -6287
rect 3875 -6321 3898 -6287
rect 3818 -6355 3898 -6321
rect 3818 -6389 3841 -6355
rect 3875 -6389 3898 -6355
rect 3818 -6403 3898 -6389
rect 3938 -5607 4018 -5603
rect 3938 -5641 3961 -5607
rect 3995 -5641 4018 -5607
rect 3938 -5675 4018 -5641
rect 3938 -5709 3961 -5675
rect 3995 -5709 4018 -5675
rect 3938 -5743 4018 -5709
rect 3938 -5777 3961 -5743
rect 3995 -5777 4018 -5743
rect 3938 -5811 4018 -5777
rect 3938 -5845 3961 -5811
rect 3995 -5845 4018 -5811
rect 3938 -5879 4018 -5845
rect 3938 -5913 3961 -5879
rect 3995 -5913 4018 -5879
rect 3938 -5947 4018 -5913
rect 3938 -5981 3961 -5947
rect 3995 -5981 4018 -5947
rect 3938 -6015 4018 -5981
rect 3938 -6049 3961 -6015
rect 3995 -6049 4018 -6015
rect 3938 -6083 4018 -6049
rect 3938 -6117 3961 -6083
rect 3995 -6117 4018 -6083
rect 3938 -6151 4018 -6117
rect 3938 -6185 3961 -6151
rect 3995 -6185 4018 -6151
rect 3938 -6219 4018 -6185
rect 3938 -6253 3961 -6219
rect 3995 -6253 4018 -6219
rect 3938 -6287 4018 -6253
rect 3938 -6321 3961 -6287
rect 3995 -6321 4018 -6287
rect 3938 -6355 4018 -6321
rect 3938 -6389 3961 -6355
rect 3995 -6389 4018 -6355
rect 2078 -6443 2118 -6403
rect 2518 -6443 2558 -6403
rect 2958 -6443 2998 -6403
rect 3398 -6443 3438 -6403
rect 3838 -6443 3878 -6403
rect 2078 -6483 3878 -6443
rect 2168 -6540 2248 -6517
rect 2168 -6574 2191 -6540
rect 2225 -6574 2248 -6540
rect 2168 -6597 2248 -6574
rect 3048 -6622 3128 -6599
rect 3048 -6656 3071 -6622
rect 3105 -6656 3128 -6622
rect 3048 -6679 3128 -6656
rect 3938 -6968 4018 -6389
rect 4392 -5623 4592 -5589
rect 4392 -5657 4415 -5623
rect 4449 -5657 4535 -5623
rect 4569 -5657 4592 -5623
rect 4392 -5691 4592 -5657
rect 4392 -5725 4415 -5691
rect 4449 -5725 4535 -5691
rect 4569 -5725 4592 -5691
rect 4392 -5759 4592 -5725
rect 4392 -5793 4415 -5759
rect 4449 -5793 4535 -5759
rect 4569 -5793 4592 -5759
rect 4392 -5827 4592 -5793
rect 4392 -5861 4415 -5827
rect 4449 -5861 4535 -5827
rect 4569 -5861 4592 -5827
rect 4392 -5895 4592 -5861
rect 4392 -5929 4415 -5895
rect 4449 -5929 4535 -5895
rect 4569 -5929 4592 -5895
rect 4392 -5963 4592 -5929
rect 4392 -5997 4415 -5963
rect 4449 -5997 4535 -5963
rect 4569 -5997 4592 -5963
rect 4392 -6031 4592 -5997
rect 4392 -6065 4415 -6031
rect 4449 -6065 4535 -6031
rect 4569 -6065 4592 -6031
rect 4392 -6099 4592 -6065
rect 4392 -6133 4415 -6099
rect 4449 -6133 4535 -6099
rect 4569 -6133 4592 -6099
rect 4392 -6167 4592 -6133
rect 4392 -6201 4415 -6167
rect 4449 -6201 4535 -6167
rect 4569 -6201 4592 -6167
rect 4392 -6235 4592 -6201
rect 4392 -6269 4415 -6235
rect 4449 -6269 4535 -6235
rect 4569 -6269 4592 -6235
rect 4392 -6303 4592 -6269
rect 4392 -6337 4415 -6303
rect 4449 -6337 4535 -6303
rect 4569 -6337 4592 -6303
rect 4392 -6371 4592 -6337
rect 4392 -6405 4415 -6371
rect 4449 -6405 4535 -6371
rect 4569 -6405 4592 -6371
rect 4392 -6435 4592 -6405
rect 4732 -5555 4812 -5525
rect 4732 -5589 4755 -5555
rect 4789 -5589 4812 -5555
rect 4732 -5623 4812 -5589
rect 4732 -5657 4755 -5623
rect 4789 -5657 4812 -5623
rect 4732 -5691 4812 -5657
rect 4732 -5725 4755 -5691
rect 4789 -5725 4812 -5691
rect 4732 -5759 4812 -5725
rect 4732 -5793 4755 -5759
rect 4789 -5793 4812 -5759
rect 4732 -5827 4812 -5793
rect 4732 -5861 4755 -5827
rect 4789 -5861 4812 -5827
rect 4732 -5895 4812 -5861
rect 4732 -5929 4755 -5895
rect 4789 -5929 4812 -5895
rect 4732 -5963 4812 -5929
rect 4732 -5997 4755 -5963
rect 4789 -5997 4812 -5963
rect 4732 -6031 4812 -5997
rect 4732 -6065 4755 -6031
rect 4789 -6065 4812 -6031
rect 4732 -6099 4812 -6065
rect 4732 -6133 4755 -6099
rect 4789 -6133 4812 -6099
rect 4732 -6167 4812 -6133
rect 4732 -6201 4755 -6167
rect 4789 -6201 4812 -6167
rect 4732 -6235 4812 -6201
rect 4732 -6269 4755 -6235
rect 4789 -6269 4812 -6235
rect 4732 -6303 4812 -6269
rect 4732 -6337 4755 -6303
rect 4789 -6337 4812 -6303
rect 4732 -6371 4812 -6337
rect 4732 -6405 4755 -6371
rect 4789 -6405 4812 -6371
rect 4732 -6435 4812 -6405
rect 4952 -5555 5032 -5525
rect 4952 -5589 4975 -5555
rect 5009 -5589 5032 -5555
rect 4952 -5623 5032 -5589
rect 4952 -5657 4975 -5623
rect 5009 -5657 5032 -5623
rect 4952 -5691 5032 -5657
rect 4952 -5725 4975 -5691
rect 5009 -5725 5032 -5691
rect 4952 -5759 5032 -5725
rect 4952 -5793 4975 -5759
rect 5009 -5793 5032 -5759
rect 4952 -5827 5032 -5793
rect 4952 -5861 4975 -5827
rect 5009 -5861 5032 -5827
rect 4952 -5895 5032 -5861
rect 4952 -5929 4975 -5895
rect 5009 -5929 5032 -5895
rect 4952 -5963 5032 -5929
rect 4952 -5997 4975 -5963
rect 5009 -5997 5032 -5963
rect 4952 -6031 5032 -5997
rect 4952 -6065 4975 -6031
rect 5009 -6065 5032 -6031
rect 4952 -6099 5032 -6065
rect 4952 -6133 4975 -6099
rect 5009 -6133 5032 -6099
rect 4952 -6167 5032 -6133
rect 4952 -6201 4975 -6167
rect 5009 -6201 5032 -6167
rect 4952 -6235 5032 -6201
rect 4952 -6269 4975 -6235
rect 5009 -6269 5032 -6235
rect 4952 -6303 5032 -6269
rect 4952 -6337 4975 -6303
rect 5009 -6337 5032 -6303
rect 4952 -6371 5032 -6337
rect 4952 -6405 4975 -6371
rect 5009 -6405 5032 -6371
rect 4952 -6435 5032 -6405
rect 5172 -5555 5252 -5525
rect 5172 -5589 5195 -5555
rect 5229 -5589 5252 -5555
rect 5172 -5623 5252 -5589
rect 5172 -5657 5195 -5623
rect 5229 -5657 5252 -5623
rect 5172 -5691 5252 -5657
rect 5172 -5725 5195 -5691
rect 5229 -5725 5252 -5691
rect 5172 -5759 5252 -5725
rect 5172 -5793 5195 -5759
rect 5229 -5793 5252 -5759
rect 5172 -5827 5252 -5793
rect 5172 -5861 5195 -5827
rect 5229 -5861 5252 -5827
rect 5172 -5895 5252 -5861
rect 5172 -5929 5195 -5895
rect 5229 -5929 5252 -5895
rect 5172 -5963 5252 -5929
rect 5172 -5997 5195 -5963
rect 5229 -5997 5252 -5963
rect 5172 -6031 5252 -5997
rect 5172 -6065 5195 -6031
rect 5229 -6065 5252 -6031
rect 5172 -6099 5252 -6065
rect 5172 -6133 5195 -6099
rect 5229 -6133 5252 -6099
rect 5172 -6167 5252 -6133
rect 5172 -6201 5195 -6167
rect 5229 -6201 5252 -6167
rect 5172 -6235 5252 -6201
rect 5172 -6269 5195 -6235
rect 5229 -6269 5252 -6235
rect 5172 -6303 5252 -6269
rect 5172 -6337 5195 -6303
rect 5229 -6337 5252 -6303
rect 5172 -6371 5252 -6337
rect 5172 -6405 5195 -6371
rect 5229 -6405 5252 -6371
rect 5172 -6435 5252 -6405
rect 5392 -5555 5472 -5525
rect 5392 -5589 5415 -5555
rect 5449 -5589 5472 -5555
rect 5392 -5623 5472 -5589
rect 5392 -5657 5415 -5623
rect 5449 -5657 5472 -5623
rect 5392 -5691 5472 -5657
rect 5392 -5725 5415 -5691
rect 5449 -5725 5472 -5691
rect 5392 -5759 5472 -5725
rect 5392 -5793 5415 -5759
rect 5449 -5793 5472 -5759
rect 5392 -5827 5472 -5793
rect 5392 -5861 5415 -5827
rect 5449 -5861 5472 -5827
rect 5392 -5895 5472 -5861
rect 5392 -5929 5415 -5895
rect 5449 -5929 5472 -5895
rect 5392 -5963 5472 -5929
rect 5392 -5997 5415 -5963
rect 5449 -5997 5472 -5963
rect 5392 -6031 5472 -5997
rect 5392 -6065 5415 -6031
rect 5449 -6065 5472 -6031
rect 5392 -6099 5472 -6065
rect 5392 -6133 5415 -6099
rect 5449 -6133 5472 -6099
rect 5392 -6167 5472 -6133
rect 5392 -6201 5415 -6167
rect 5449 -6201 5472 -6167
rect 5392 -6235 5472 -6201
rect 5392 -6269 5415 -6235
rect 5449 -6269 5472 -6235
rect 5392 -6303 5472 -6269
rect 5392 -6337 5415 -6303
rect 5449 -6337 5472 -6303
rect 5392 -6371 5472 -6337
rect 5392 -6405 5415 -6371
rect 5449 -6405 5472 -6371
rect 5392 -6435 5472 -6405
rect 5612 -5555 5692 -5525
rect 5612 -5589 5635 -5555
rect 5669 -5589 5692 -5555
rect 5612 -5623 5692 -5589
rect 5612 -5657 5635 -5623
rect 5669 -5657 5692 -5623
rect 5612 -5691 5692 -5657
rect 5612 -5725 5635 -5691
rect 5669 -5725 5692 -5691
rect 5612 -5759 5692 -5725
rect 5612 -5793 5635 -5759
rect 5669 -5793 5692 -5759
rect 5612 -5827 5692 -5793
rect 5612 -5861 5635 -5827
rect 5669 -5861 5692 -5827
rect 5612 -5895 5692 -5861
rect 5612 -5929 5635 -5895
rect 5669 -5929 5692 -5895
rect 5612 -5963 5692 -5929
rect 5612 -5997 5635 -5963
rect 5669 -5997 5692 -5963
rect 5612 -6031 5692 -5997
rect 5612 -6065 5635 -6031
rect 5669 -6065 5692 -6031
rect 5612 -6099 5692 -6065
rect 5612 -6133 5635 -6099
rect 5669 -6133 5692 -6099
rect 5612 -6167 5692 -6133
rect 5612 -6201 5635 -6167
rect 5669 -6201 5692 -6167
rect 5612 -6235 5692 -6201
rect 5612 -6269 5635 -6235
rect 5669 -6269 5692 -6235
rect 5612 -6303 5692 -6269
rect 5612 -6337 5635 -6303
rect 5669 -6337 5692 -6303
rect 5612 -6371 5692 -6337
rect 5612 -6405 5635 -6371
rect 5669 -6405 5692 -6371
rect 5612 -6435 5692 -6405
rect 5832 -5555 5912 -5525
rect 5832 -5589 5855 -5555
rect 5889 -5589 5912 -5555
rect 5832 -5623 5912 -5589
rect 5832 -5657 5855 -5623
rect 5889 -5657 5912 -5623
rect 5832 -5691 5912 -5657
rect 5832 -5725 5855 -5691
rect 5889 -5725 5912 -5691
rect 5832 -5759 5912 -5725
rect 5832 -5793 5855 -5759
rect 5889 -5793 5912 -5759
rect 5832 -5827 5912 -5793
rect 5832 -5861 5855 -5827
rect 5889 -5861 5912 -5827
rect 5832 -5895 5912 -5861
rect 5832 -5929 5855 -5895
rect 5889 -5929 5912 -5895
rect 5832 -5963 5912 -5929
rect 5832 -5997 5855 -5963
rect 5889 -5997 5912 -5963
rect 5832 -6031 5912 -5997
rect 5832 -6065 5855 -6031
rect 5889 -6065 5912 -6031
rect 5832 -6099 5912 -6065
rect 5832 -6133 5855 -6099
rect 5889 -6133 5912 -6099
rect 5832 -6167 5912 -6133
rect 5832 -6201 5855 -6167
rect 5889 -6201 5912 -6167
rect 5832 -6235 5912 -6201
rect 5832 -6269 5855 -6235
rect 5889 -6269 5912 -6235
rect 5832 -6303 5912 -6269
rect 5832 -6337 5855 -6303
rect 5889 -6337 5912 -6303
rect 5832 -6371 5912 -6337
rect 5832 -6405 5855 -6371
rect 5889 -6405 5912 -6371
rect 5832 -6435 5912 -6405
rect 6052 -5555 6132 -5525
rect 6052 -5589 6075 -5555
rect 6109 -5589 6132 -5555
rect 6052 -5623 6132 -5589
rect 6052 -5657 6075 -5623
rect 6109 -5657 6132 -5623
rect 6052 -5691 6132 -5657
rect 6052 -5725 6075 -5691
rect 6109 -5725 6132 -5691
rect 6052 -5759 6132 -5725
rect 6052 -5793 6075 -5759
rect 6109 -5793 6132 -5759
rect 6052 -5827 6132 -5793
rect 6052 -5861 6075 -5827
rect 6109 -5861 6132 -5827
rect 6052 -5895 6132 -5861
rect 6052 -5929 6075 -5895
rect 6109 -5929 6132 -5895
rect 6052 -5963 6132 -5929
rect 6052 -5997 6075 -5963
rect 6109 -5997 6132 -5963
rect 6052 -6031 6132 -5997
rect 6052 -6065 6075 -6031
rect 6109 -6065 6132 -6031
rect 6052 -6099 6132 -6065
rect 6052 -6133 6075 -6099
rect 6109 -6133 6132 -6099
rect 6052 -6167 6132 -6133
rect 6052 -6201 6075 -6167
rect 6109 -6201 6132 -6167
rect 6052 -6235 6132 -6201
rect 6052 -6269 6075 -6235
rect 6109 -6269 6132 -6235
rect 6052 -6303 6132 -6269
rect 6052 -6337 6075 -6303
rect 6109 -6337 6132 -6303
rect 6052 -6371 6132 -6337
rect 6052 -6405 6075 -6371
rect 6109 -6405 6132 -6371
rect 6052 -6435 6132 -6405
rect 6272 -5555 6472 -5525
rect 6272 -5589 6295 -5555
rect 6329 -5589 6415 -5555
rect 6449 -5589 6472 -5555
rect 6272 -5623 6472 -5589
rect 6989 -5603 7023 -5479
rect 7206 -5523 7286 -5398
rect 8291 -5523 8361 -5313
rect 7206 -5563 7686 -5523
rect 7206 -5603 7246 -5563
rect 7646 -5603 7686 -5563
rect 8086 -5563 8566 -5523
rect 8086 -5603 8126 -5563
rect 8526 -5603 8566 -5563
rect 6272 -5657 6295 -5623
rect 6329 -5657 6415 -5623
rect 6449 -5657 6472 -5623
rect 6272 -5691 6472 -5657
rect 6272 -5725 6295 -5691
rect 6329 -5725 6415 -5691
rect 6449 -5725 6472 -5691
rect 6272 -5759 6472 -5725
rect 6272 -5793 6295 -5759
rect 6329 -5793 6415 -5759
rect 6449 -5793 6472 -5759
rect 6272 -5827 6472 -5793
rect 6272 -5861 6295 -5827
rect 6329 -5861 6415 -5827
rect 6449 -5861 6472 -5827
rect 6272 -5895 6472 -5861
rect 6272 -5929 6295 -5895
rect 6329 -5929 6415 -5895
rect 6449 -5929 6472 -5895
rect 6272 -5963 6472 -5929
rect 6272 -5997 6295 -5963
rect 6329 -5997 6415 -5963
rect 6449 -5997 6472 -5963
rect 6272 -6031 6472 -5997
rect 6272 -6065 6295 -6031
rect 6329 -6065 6415 -6031
rect 6449 -6065 6472 -6031
rect 6272 -6099 6472 -6065
rect 6272 -6133 6295 -6099
rect 6329 -6133 6415 -6099
rect 6449 -6133 6472 -6099
rect 6272 -6167 6472 -6133
rect 6272 -6201 6295 -6167
rect 6329 -6201 6415 -6167
rect 6449 -6201 6472 -6167
rect 6272 -6235 6472 -6201
rect 6272 -6269 6295 -6235
rect 6329 -6269 6415 -6235
rect 6449 -6269 6472 -6235
rect 6272 -6303 6472 -6269
rect 6272 -6337 6295 -6303
rect 6329 -6337 6415 -6303
rect 6449 -6337 6472 -6303
rect 6272 -6371 6472 -6337
rect 6272 -6405 6295 -6371
rect 6329 -6405 6415 -6371
rect 6449 -6405 6472 -6371
rect 6272 -6435 6472 -6405
rect 6846 -5607 6926 -5603
rect 6846 -5641 6869 -5607
rect 6903 -5641 6926 -5607
rect 6846 -5675 6926 -5641
rect 6846 -5709 6869 -5675
rect 6903 -5709 6926 -5675
rect 6846 -5743 6926 -5709
rect 6846 -5777 6869 -5743
rect 6903 -5777 6926 -5743
rect 6846 -5811 6926 -5777
rect 6846 -5845 6869 -5811
rect 6903 -5845 6926 -5811
rect 6846 -5879 6926 -5845
rect 6846 -5913 6869 -5879
rect 6903 -5913 6926 -5879
rect 6846 -5947 6926 -5913
rect 6846 -5981 6869 -5947
rect 6903 -5981 6926 -5947
rect 6846 -6015 6926 -5981
rect 6846 -6049 6869 -6015
rect 6903 -6049 6926 -6015
rect 6846 -6083 6926 -6049
rect 6846 -6117 6869 -6083
rect 6903 -6117 6926 -6083
rect 6846 -6151 6926 -6117
rect 6846 -6185 6869 -6151
rect 6903 -6185 6926 -6151
rect 6846 -6219 6926 -6185
rect 6846 -6253 6869 -6219
rect 6903 -6253 6926 -6219
rect 6846 -6287 6926 -6253
rect 6846 -6321 6869 -6287
rect 6903 -6321 6926 -6287
rect 6846 -6355 6926 -6321
rect 6846 -6389 6869 -6355
rect 6903 -6389 6926 -6355
rect 4532 -6475 4572 -6435
rect 4972 -6475 5012 -6435
rect 5412 -6475 5452 -6435
rect 5852 -6475 5892 -6435
rect 6292 -6475 6332 -6435
rect 4532 -6515 6332 -6475
rect 4622 -6786 4702 -6763
rect 4622 -6820 4645 -6786
rect 4679 -6820 4702 -6786
rect 4622 -6843 4702 -6820
rect 5034 -6968 5834 -6515
rect 6161 -6704 6241 -6681
rect 6161 -6738 6184 -6704
rect 6218 -6738 6241 -6704
rect 6161 -6761 6241 -6738
rect 6846 -6968 6926 -6389
rect 6966 -5607 7046 -5603
rect 6966 -5641 6989 -5607
rect 7023 -5641 7046 -5607
rect 6966 -5675 7046 -5641
rect 6966 -5709 6989 -5675
rect 7023 -5709 7046 -5675
rect 6966 -5743 7046 -5709
rect 6966 -5777 6989 -5743
rect 7023 -5777 7046 -5743
rect 6966 -5811 7046 -5777
rect 6966 -5845 6989 -5811
rect 7023 -5845 7046 -5811
rect 6966 -5879 7046 -5845
rect 6966 -5913 6989 -5879
rect 7023 -5913 7046 -5879
rect 6966 -5947 7046 -5913
rect 6966 -5981 6989 -5947
rect 7023 -5981 7046 -5947
rect 6966 -6015 7046 -5981
rect 6966 -6049 6989 -6015
rect 7023 -6049 7046 -6015
rect 6966 -6083 7046 -6049
rect 6966 -6117 6989 -6083
rect 7023 -6117 7046 -6083
rect 6966 -6151 7046 -6117
rect 6966 -6185 6989 -6151
rect 7023 -6185 7046 -6151
rect 6966 -6219 7046 -6185
rect 6966 -6253 6989 -6219
rect 7023 -6253 7046 -6219
rect 6966 -6287 7046 -6253
rect 6966 -6321 6989 -6287
rect 7023 -6321 7046 -6287
rect 6966 -6355 7046 -6321
rect 6966 -6389 6989 -6355
rect 7023 -6389 7046 -6355
rect 6966 -6403 7046 -6389
rect 7186 -5607 7266 -5603
rect 7186 -5641 7209 -5607
rect 7243 -5641 7266 -5607
rect 7186 -5675 7266 -5641
rect 7186 -5709 7209 -5675
rect 7243 -5709 7266 -5675
rect 7186 -5743 7266 -5709
rect 7186 -5777 7209 -5743
rect 7243 -5777 7266 -5743
rect 7186 -5811 7266 -5777
rect 7186 -5845 7209 -5811
rect 7243 -5845 7266 -5811
rect 7186 -5879 7266 -5845
rect 7186 -5913 7209 -5879
rect 7243 -5913 7266 -5879
rect 7186 -5947 7266 -5913
rect 7186 -5981 7209 -5947
rect 7243 -5981 7266 -5947
rect 7186 -6015 7266 -5981
rect 7186 -6049 7209 -6015
rect 7243 -6049 7266 -6015
rect 7186 -6083 7266 -6049
rect 7186 -6117 7209 -6083
rect 7243 -6117 7266 -6083
rect 7186 -6151 7266 -6117
rect 7186 -6185 7209 -6151
rect 7243 -6185 7266 -6151
rect 7186 -6219 7266 -6185
rect 7186 -6253 7209 -6219
rect 7243 -6253 7266 -6219
rect 7186 -6287 7266 -6253
rect 7186 -6321 7209 -6287
rect 7243 -6321 7266 -6287
rect 7186 -6355 7266 -6321
rect 7186 -6389 7209 -6355
rect 7243 -6389 7266 -6355
rect 7186 -6403 7266 -6389
rect 7406 -5607 7486 -5603
rect 7406 -5641 7429 -5607
rect 7463 -5641 7486 -5607
rect 7406 -5675 7486 -5641
rect 7406 -5709 7429 -5675
rect 7463 -5709 7486 -5675
rect 7406 -5743 7486 -5709
rect 7406 -5777 7429 -5743
rect 7463 -5777 7486 -5743
rect 7406 -5811 7486 -5777
rect 7406 -5845 7429 -5811
rect 7463 -5845 7486 -5811
rect 7406 -5879 7486 -5845
rect 7406 -5913 7429 -5879
rect 7463 -5913 7486 -5879
rect 7406 -5947 7486 -5913
rect 7406 -5981 7429 -5947
rect 7463 -5981 7486 -5947
rect 7406 -6015 7486 -5981
rect 7406 -6049 7429 -6015
rect 7463 -6049 7486 -6015
rect 7406 -6083 7486 -6049
rect 7406 -6117 7429 -6083
rect 7463 -6117 7486 -6083
rect 7406 -6151 7486 -6117
rect 7406 -6185 7429 -6151
rect 7463 -6185 7486 -6151
rect 7406 -6219 7486 -6185
rect 7406 -6253 7429 -6219
rect 7463 -6253 7486 -6219
rect 7406 -6287 7486 -6253
rect 7406 -6321 7429 -6287
rect 7463 -6321 7486 -6287
rect 7406 -6355 7486 -6321
rect 7406 -6389 7429 -6355
rect 7463 -6389 7486 -6355
rect 7406 -6403 7486 -6389
rect 7626 -5607 7706 -5603
rect 7626 -5641 7649 -5607
rect 7683 -5641 7706 -5607
rect 7626 -5675 7706 -5641
rect 7626 -5709 7649 -5675
rect 7683 -5709 7706 -5675
rect 7626 -5743 7706 -5709
rect 7626 -5777 7649 -5743
rect 7683 -5777 7706 -5743
rect 7626 -5811 7706 -5777
rect 7626 -5845 7649 -5811
rect 7683 -5845 7706 -5811
rect 7626 -5879 7706 -5845
rect 7626 -5913 7649 -5879
rect 7683 -5913 7706 -5879
rect 7626 -5947 7706 -5913
rect 7626 -5981 7649 -5947
rect 7683 -5981 7706 -5947
rect 7626 -6015 7706 -5981
rect 7626 -6049 7649 -6015
rect 7683 -6049 7706 -6015
rect 7626 -6083 7706 -6049
rect 7626 -6117 7649 -6083
rect 7683 -6117 7706 -6083
rect 7626 -6151 7706 -6117
rect 7626 -6185 7649 -6151
rect 7683 -6185 7706 -6151
rect 7626 -6219 7706 -6185
rect 7626 -6253 7649 -6219
rect 7683 -6253 7706 -6219
rect 7626 -6287 7706 -6253
rect 7626 -6321 7649 -6287
rect 7683 -6321 7706 -6287
rect 7626 -6355 7706 -6321
rect 7626 -6389 7649 -6355
rect 7683 -6389 7706 -6355
rect 7626 -6403 7706 -6389
rect 7846 -5607 7926 -5603
rect 7846 -5641 7869 -5607
rect 7903 -5641 7926 -5607
rect 7846 -5675 7926 -5641
rect 7846 -5709 7869 -5675
rect 7903 -5709 7926 -5675
rect 7846 -5743 7926 -5709
rect 7846 -5777 7869 -5743
rect 7903 -5777 7926 -5743
rect 7846 -5811 7926 -5777
rect 7846 -5845 7869 -5811
rect 7903 -5845 7926 -5811
rect 7846 -5879 7926 -5845
rect 7846 -5913 7869 -5879
rect 7903 -5913 7926 -5879
rect 7846 -5947 7926 -5913
rect 7846 -5981 7869 -5947
rect 7903 -5981 7926 -5947
rect 7846 -6015 7926 -5981
rect 7846 -6049 7869 -6015
rect 7903 -6049 7926 -6015
rect 7846 -6083 7926 -6049
rect 7846 -6117 7869 -6083
rect 7903 -6117 7926 -6083
rect 7846 -6151 7926 -6117
rect 7846 -6185 7869 -6151
rect 7903 -6185 7926 -6151
rect 7846 -6219 7926 -6185
rect 7846 -6253 7869 -6219
rect 7903 -6253 7926 -6219
rect 7846 -6287 7926 -6253
rect 7846 -6321 7869 -6287
rect 7903 -6321 7926 -6287
rect 7846 -6355 7926 -6321
rect 7846 -6389 7869 -6355
rect 7903 -6389 7926 -6355
rect 7846 -6403 7926 -6389
rect 8066 -5607 8146 -5603
rect 8066 -5641 8089 -5607
rect 8123 -5641 8146 -5607
rect 8066 -5675 8146 -5641
rect 8066 -5709 8089 -5675
rect 8123 -5709 8146 -5675
rect 8066 -5743 8146 -5709
rect 8066 -5777 8089 -5743
rect 8123 -5777 8146 -5743
rect 8066 -5811 8146 -5777
rect 8066 -5845 8089 -5811
rect 8123 -5845 8146 -5811
rect 8066 -5879 8146 -5845
rect 8066 -5913 8089 -5879
rect 8123 -5913 8146 -5879
rect 8066 -5947 8146 -5913
rect 8066 -5981 8089 -5947
rect 8123 -5981 8146 -5947
rect 8066 -6015 8146 -5981
rect 8066 -6049 8089 -6015
rect 8123 -6049 8146 -6015
rect 8066 -6083 8146 -6049
rect 8066 -6117 8089 -6083
rect 8123 -6117 8146 -6083
rect 8066 -6151 8146 -6117
rect 8066 -6185 8089 -6151
rect 8123 -6185 8146 -6151
rect 8066 -6219 8146 -6185
rect 8066 -6253 8089 -6219
rect 8123 -6253 8146 -6219
rect 8066 -6287 8146 -6253
rect 8066 -6321 8089 -6287
rect 8123 -6321 8146 -6287
rect 8066 -6355 8146 -6321
rect 8066 -6389 8089 -6355
rect 8123 -6389 8146 -6355
rect 8066 -6403 8146 -6389
rect 8286 -5607 8366 -5603
rect 8286 -5641 8309 -5607
rect 8343 -5641 8366 -5607
rect 8286 -5675 8366 -5641
rect 8286 -5709 8309 -5675
rect 8343 -5709 8366 -5675
rect 8286 -5743 8366 -5709
rect 8286 -5777 8309 -5743
rect 8343 -5777 8366 -5743
rect 8286 -5811 8366 -5777
rect 8286 -5845 8309 -5811
rect 8343 -5845 8366 -5811
rect 8286 -5879 8366 -5845
rect 8286 -5913 8309 -5879
rect 8343 -5913 8366 -5879
rect 8286 -5947 8366 -5913
rect 8286 -5981 8309 -5947
rect 8343 -5981 8366 -5947
rect 8286 -6015 8366 -5981
rect 8286 -6049 8309 -6015
rect 8343 -6049 8366 -6015
rect 8286 -6083 8366 -6049
rect 8286 -6117 8309 -6083
rect 8343 -6117 8366 -6083
rect 8286 -6151 8366 -6117
rect 8286 -6185 8309 -6151
rect 8343 -6185 8366 -6151
rect 8286 -6219 8366 -6185
rect 8286 -6253 8309 -6219
rect 8343 -6253 8366 -6219
rect 8286 -6287 8366 -6253
rect 8286 -6321 8309 -6287
rect 8343 -6321 8366 -6287
rect 8286 -6355 8366 -6321
rect 8286 -6389 8309 -6355
rect 8343 -6389 8366 -6355
rect 8286 -6403 8366 -6389
rect 8506 -5607 8586 -5603
rect 8506 -5641 8529 -5607
rect 8563 -5641 8586 -5607
rect 8506 -5675 8586 -5641
rect 8506 -5709 8529 -5675
rect 8563 -5709 8586 -5675
rect 8506 -5743 8586 -5709
rect 8506 -5777 8529 -5743
rect 8563 -5777 8586 -5743
rect 8506 -5811 8586 -5777
rect 8506 -5845 8529 -5811
rect 8563 -5845 8586 -5811
rect 8506 -5879 8586 -5845
rect 8506 -5913 8529 -5879
rect 8563 -5913 8586 -5879
rect 8506 -5947 8586 -5913
rect 8506 -5981 8529 -5947
rect 8563 -5981 8586 -5947
rect 8506 -6015 8586 -5981
rect 8506 -6049 8529 -6015
rect 8563 -6049 8586 -6015
rect 8506 -6083 8586 -6049
rect 8506 -6117 8529 -6083
rect 8563 -6117 8586 -6083
rect 8506 -6151 8586 -6117
rect 8506 -6185 8529 -6151
rect 8563 -6185 8586 -6151
rect 8506 -6219 8586 -6185
rect 8506 -6253 8529 -6219
rect 8563 -6253 8586 -6219
rect 8506 -6287 8586 -6253
rect 8506 -6321 8529 -6287
rect 8563 -6321 8586 -6287
rect 8506 -6355 8586 -6321
rect 8506 -6389 8529 -6355
rect 8563 -6389 8586 -6355
rect 8506 -6403 8586 -6389
rect 8726 -5607 8806 -5603
rect 8726 -5641 8749 -5607
rect 8783 -5641 8806 -5607
rect 8726 -5675 8806 -5641
rect 8726 -5709 8749 -5675
rect 8783 -5709 8806 -5675
rect 8726 -5743 8806 -5709
rect 8726 -5777 8749 -5743
rect 8783 -5777 8806 -5743
rect 8726 -5811 8806 -5777
rect 8726 -5845 8749 -5811
rect 8783 -5845 8806 -5811
rect 8726 -5879 8806 -5845
rect 8726 -5913 8749 -5879
rect 8783 -5913 8806 -5879
rect 8726 -5947 8806 -5913
rect 8726 -5981 8749 -5947
rect 8783 -5981 8806 -5947
rect 8726 -6015 8806 -5981
rect 8726 -6049 8749 -6015
rect 8783 -6049 8806 -6015
rect 8726 -6083 8806 -6049
rect 8726 -6117 8749 -6083
rect 8783 -6117 8806 -6083
rect 8726 -6151 8806 -6117
rect 8726 -6185 8749 -6151
rect 8783 -6185 8806 -6151
rect 8726 -6219 8806 -6185
rect 8726 -6253 8749 -6219
rect 8783 -6253 8806 -6219
rect 8726 -6287 8806 -6253
rect 8726 -6321 8749 -6287
rect 8783 -6321 8806 -6287
rect 8726 -6355 8806 -6321
rect 8726 -6389 8749 -6355
rect 8783 -6389 8806 -6355
rect 8726 -6403 8806 -6389
rect 8846 -5607 8926 -5603
rect 8846 -5641 8869 -5607
rect 8903 -5641 8926 -5607
rect 8846 -5675 8926 -5641
rect 8846 -5709 8869 -5675
rect 8903 -5709 8926 -5675
rect 8846 -5743 8926 -5709
rect 8846 -5777 8869 -5743
rect 8903 -5777 8926 -5743
rect 8846 -5811 8926 -5777
rect 8846 -5845 8869 -5811
rect 8903 -5845 8926 -5811
rect 8846 -5879 8926 -5845
rect 8846 -5913 8869 -5879
rect 8903 -5913 8926 -5879
rect 8846 -5947 8926 -5913
rect 8846 -5981 8869 -5947
rect 8903 -5981 8926 -5947
rect 8846 -6015 8926 -5981
rect 8846 -6049 8869 -6015
rect 8903 -6049 8926 -6015
rect 8846 -6083 8926 -6049
rect 8846 -6117 8869 -6083
rect 8903 -6117 8926 -6083
rect 8846 -6151 8926 -6117
rect 8846 -6185 8869 -6151
rect 8903 -6185 8926 -6151
rect 8846 -6219 8926 -6185
rect 8846 -6253 8869 -6219
rect 8903 -6253 8926 -6219
rect 8846 -6287 8926 -6253
rect 8846 -6321 8869 -6287
rect 8903 -6321 8926 -6287
rect 8846 -6355 8926 -6321
rect 8846 -6389 8869 -6355
rect 8903 -6389 8926 -6355
rect 6986 -6443 7026 -6403
rect 7426 -6443 7466 -6403
rect 7866 -6443 7906 -6403
rect 8306 -6443 8346 -6403
rect 8746 -6443 8786 -6403
rect 6986 -6483 8786 -6443
rect 7953 -6540 8033 -6517
rect 7953 -6574 7976 -6540
rect 8010 -6574 8033 -6540
rect 7953 -6597 8033 -6574
rect 7076 -6622 7156 -6599
rect 7076 -6656 7099 -6622
rect 7133 -6656 7156 -6622
rect 7076 -6679 7156 -6656
rect 8846 -6968 8926 -6389
rect -102 -6991 10465 -6968
rect -102 -7025 -41 -6991
rect -7 -7025 31 -6991
rect 65 -7025 103 -6991
rect 137 -7025 175 -6991
rect 209 -7025 247 -6991
rect 281 -7025 319 -6991
rect 353 -7025 391 -6991
rect 425 -7025 463 -6991
rect 497 -7025 535 -6991
rect 569 -7025 607 -6991
rect 641 -7025 679 -6991
rect 713 -7025 751 -6991
rect 785 -7025 823 -6991
rect 857 -7025 895 -6991
rect 929 -7025 967 -6991
rect 1001 -7025 1039 -6991
rect 1073 -7025 1111 -6991
rect 1145 -7025 1183 -6991
rect 1217 -7025 1278 -6991
rect 1312 -7025 1350 -6991
rect 1384 -7025 1422 -6991
rect 1456 -7025 1494 -6991
rect 1528 -7025 1566 -6991
rect 1600 -7025 1638 -6991
rect 1672 -7025 1710 -6991
rect 1744 -7025 1782 -6991
rect 1816 -7025 1854 -6991
rect 1888 -7025 1926 -6991
rect 1960 -7025 1998 -6991
rect 2032 -7025 2070 -6991
rect 2104 -7025 2142 -6991
rect 2176 -7025 2214 -6991
rect 2248 -7025 2286 -6991
rect 2320 -7025 2358 -6991
rect 2392 -7025 2430 -6991
rect 2464 -7025 2502 -6991
rect 2536 -7025 2574 -6991
rect 2608 -7025 2646 -6991
rect 2680 -7025 2718 -6991
rect 2752 -7025 2790 -6991
rect 2824 -7025 2862 -6991
rect 2896 -7025 2934 -6991
rect 2968 -7025 3006 -6991
rect 3040 -7025 3078 -6991
rect 3112 -7025 3150 -6991
rect 3184 -7025 3222 -6991
rect 3256 -7025 3294 -6991
rect 3328 -7025 3366 -6991
rect 3400 -7025 3438 -6991
rect 3472 -7025 3510 -6991
rect 3544 -7025 3582 -6991
rect 3616 -7025 3654 -6991
rect 3688 -7025 3726 -6991
rect 3760 -7025 3798 -6991
rect 3832 -7025 3893 -6991
rect 3927 -7025 3965 -6991
rect 3999 -7025 4037 -6991
rect 4071 -7025 4109 -6991
rect 4143 -7025 4181 -6991
rect 4215 -7025 4253 -6991
rect 4287 -7025 4325 -6991
rect 4359 -7025 4397 -6991
rect 4431 -7025 4469 -6991
rect 4503 -7025 4541 -6991
rect 4575 -7025 4613 -6991
rect 4647 -7025 4685 -6991
rect 4719 -7025 4757 -6991
rect 4791 -7025 4829 -6991
rect 4863 -7025 4901 -6991
rect 4935 -7025 4973 -6991
rect 5007 -7025 5045 -6991
rect 5079 -7025 5117 -6991
rect 5151 -7025 5189 -6991
rect 5223 -7025 5261 -6991
rect 5295 -7025 5333 -6991
rect 5367 -7025 5405 -6991
rect 5439 -7025 5477 -6991
rect 5511 -7025 5549 -6991
rect 5583 -7025 5621 -6991
rect 5655 -7025 5693 -6991
rect 5727 -7025 5765 -6991
rect 5799 -7025 5837 -6991
rect 5871 -7025 5909 -6991
rect 5943 -7025 5981 -6991
rect 6015 -7025 6053 -6991
rect 6087 -7025 6125 -6991
rect 6159 -7025 6197 -6991
rect 6231 -7025 6269 -6991
rect 6303 -7025 6341 -6991
rect 6375 -7025 6413 -6991
rect 6447 -7025 6508 -6991
rect 6542 -7025 6580 -6991
rect 6614 -7025 6652 -6991
rect 6686 -7025 6724 -6991
rect 6758 -7025 6796 -6991
rect 6830 -7025 6868 -6991
rect 6902 -7025 6940 -6991
rect 6974 -7025 7012 -6991
rect 7046 -7025 7084 -6991
rect 7118 -7025 7156 -6991
rect 7190 -7025 7228 -6991
rect 7262 -7025 7300 -6991
rect 7334 -7025 7372 -6991
rect 7406 -7025 7444 -6991
rect 7478 -7025 7516 -6991
rect 7550 -7025 7588 -6991
rect 7622 -7025 7660 -6991
rect 7694 -7025 7732 -6991
rect 7766 -7025 7804 -6991
rect 7838 -7025 7876 -6991
rect 7910 -7025 7948 -6991
rect 7982 -7025 8020 -6991
rect 8054 -7025 8092 -6991
rect 8126 -7025 8164 -6991
rect 8198 -7025 8236 -6991
rect 8270 -7025 8308 -6991
rect 8342 -7025 8380 -6991
rect 8414 -7025 8452 -6991
rect 8486 -7025 8524 -6991
rect 8558 -7025 8596 -6991
rect 8630 -7025 8668 -6991
rect 8702 -7025 8740 -6991
rect 8774 -7025 8812 -6991
rect 8846 -7025 8884 -6991
rect 8918 -7025 8956 -6991
rect 8990 -7025 9028 -6991
rect 9062 -7025 9123 -6991
rect 9157 -7025 9195 -6991
rect 9229 -7025 9267 -6991
rect 9301 -7025 9339 -6991
rect 9373 -7025 9411 -6991
rect 9445 -7025 9483 -6991
rect 9517 -7025 9555 -6991
rect 9589 -7025 9627 -6991
rect 9661 -7025 9699 -6991
rect 9733 -7025 9771 -6991
rect 9805 -7025 9843 -6991
rect 9877 -7025 9915 -6991
rect 9949 -7025 9987 -6991
rect 10021 -7025 10059 -6991
rect 10093 -7025 10131 -6991
rect 10165 -7025 10203 -6991
rect 10237 -7025 10275 -6991
rect 10309 -7025 10347 -6991
rect 10381 -7025 10465 -6991
rect -102 -7048 10465 -7025
<< viali >>
rect -40 -3489 -6 -3455
rect 32 -3489 66 -3455
rect 104 -3489 138 -3455
rect 176 -3489 210 -3455
rect 248 -3489 282 -3455
rect 320 -3489 354 -3455
rect 392 -3489 426 -3455
rect 464 -3489 498 -3455
rect 536 -3489 570 -3455
rect 608 -3489 642 -3455
rect 680 -3489 714 -3455
rect 752 -3489 786 -3455
rect 824 -3489 858 -3455
rect 896 -3489 930 -3455
rect 968 -3489 1002 -3455
rect 1040 -3489 1074 -3455
rect 1112 -3489 1146 -3455
rect 1184 -3489 1218 -3455
rect 1279 -3489 1313 -3455
rect 1351 -3489 1385 -3455
rect 1423 -3489 1457 -3455
rect 1495 -3489 1529 -3455
rect 1567 -3489 1601 -3455
rect 1639 -3489 1673 -3455
rect 1711 -3489 1745 -3455
rect 1783 -3489 1817 -3455
rect 1855 -3489 1889 -3455
rect 1927 -3489 1961 -3455
rect 1999 -3489 2033 -3455
rect 2071 -3489 2105 -3455
rect 2143 -3489 2177 -3455
rect 2215 -3489 2249 -3455
rect 2287 -3489 2321 -3455
rect 2359 -3489 2393 -3455
rect 2431 -3489 2465 -3455
rect 2503 -3489 2537 -3455
rect 2575 -3489 2609 -3455
rect 2647 -3489 2681 -3455
rect 2719 -3489 2753 -3455
rect 2791 -3489 2825 -3455
rect 2863 -3489 2897 -3455
rect 2935 -3489 2969 -3455
rect 3007 -3489 3041 -3455
rect 3079 -3489 3113 -3455
rect 3151 -3489 3185 -3455
rect 3223 -3489 3257 -3455
rect 3295 -3489 3329 -3455
rect 3367 -3489 3401 -3455
rect 3439 -3489 3473 -3455
rect 3511 -3489 3545 -3455
rect 3583 -3489 3617 -3455
rect 3655 -3489 3689 -3455
rect 3727 -3489 3761 -3455
rect 3799 -3489 3833 -3455
rect 3894 -3489 3928 -3455
rect 3966 -3489 4000 -3455
rect 4038 -3489 4072 -3455
rect 4110 -3489 4144 -3455
rect 4182 -3489 4216 -3455
rect 4254 -3489 4288 -3455
rect 4326 -3489 4360 -3455
rect 4398 -3489 4432 -3455
rect 4470 -3489 4504 -3455
rect 4542 -3489 4576 -3455
rect 4614 -3489 4648 -3455
rect 4686 -3489 4720 -3455
rect 4758 -3489 4792 -3455
rect 4830 -3489 4864 -3455
rect 4902 -3489 4936 -3455
rect 4974 -3489 5008 -3455
rect 5046 -3489 5080 -3455
rect 5118 -3489 5152 -3455
rect 5190 -3489 5224 -3455
rect 5262 -3489 5296 -3455
rect 5334 -3489 5368 -3455
rect 5406 -3489 5440 -3455
rect 5478 -3489 5512 -3455
rect 5550 -3489 5584 -3455
rect 5622 -3489 5656 -3455
rect 5694 -3489 5728 -3455
rect 5766 -3489 5800 -3455
rect 5838 -3489 5872 -3455
rect 5910 -3489 5944 -3455
rect 5982 -3489 6016 -3455
rect 6054 -3489 6088 -3455
rect 6126 -3489 6160 -3455
rect 6198 -3489 6232 -3455
rect 6270 -3489 6304 -3455
rect 6342 -3489 6376 -3455
rect 6414 -3489 6448 -3455
rect 6509 -3489 6543 -3455
rect 6581 -3489 6615 -3455
rect 6653 -3489 6687 -3455
rect 6725 -3489 6759 -3455
rect 6797 -3489 6831 -3455
rect 6869 -3489 6903 -3455
rect 6941 -3489 6975 -3455
rect 7013 -3489 7047 -3455
rect 7085 -3489 7119 -3455
rect 7157 -3489 7191 -3455
rect 7229 -3489 7263 -3455
rect 7301 -3489 7335 -3455
rect 7373 -3489 7407 -3455
rect 7445 -3489 7479 -3455
rect 7517 -3489 7551 -3455
rect 7589 -3489 7623 -3455
rect 7661 -3489 7695 -3455
rect 7733 -3489 7767 -3455
rect 7805 -3489 7839 -3455
rect 7877 -3489 7911 -3455
rect 7949 -3489 7983 -3455
rect 8021 -3489 8055 -3455
rect 8093 -3489 8127 -3455
rect 8165 -3489 8199 -3455
rect 8237 -3489 8271 -3455
rect 8309 -3489 8343 -3455
rect 8381 -3489 8415 -3455
rect 8453 -3489 8487 -3455
rect 8525 -3489 8559 -3455
rect 8597 -3489 8631 -3455
rect 8669 -3489 8703 -3455
rect 8741 -3489 8775 -3455
rect 8813 -3489 8847 -3455
rect 8885 -3489 8919 -3455
rect 8957 -3489 8991 -3455
rect 9029 -3489 9063 -3455
rect 9124 -3489 9158 -3455
rect 9196 -3489 9230 -3455
rect 9268 -3489 9302 -3455
rect 9340 -3489 9374 -3455
rect 9412 -3489 9446 -3455
rect 9484 -3489 9518 -3455
rect 9556 -3489 9590 -3455
rect 9628 -3489 9662 -3455
rect 9700 -3489 9734 -3455
rect 9772 -3489 9806 -3455
rect 9844 -3489 9878 -3455
rect 9916 -3489 9950 -3455
rect 9988 -3489 10022 -3455
rect 10060 -3489 10094 -3455
rect 10132 -3489 10166 -3455
rect 10204 -3489 10238 -3455
rect 10276 -3489 10310 -3455
rect 10348 -3489 10382 -3455
rect 2207 -3777 2241 -3743
rect 2523 -4077 2557 -4043
rect 2523 -4149 2557 -4115
rect 2523 -4221 2557 -4187
rect 2523 -4293 2557 -4259
rect 2523 -4365 2557 -4331
rect 2523 -4437 2557 -4403
rect 2523 -4646 2557 -4612
rect 2523 -4718 2557 -4684
rect 2523 -4790 2557 -4756
rect 2523 -4862 2557 -4828
rect 8309 -4077 8343 -4043
rect 8309 -4149 8343 -4115
rect 8309 -4221 8343 -4187
rect 8309 -4293 8343 -4259
rect 8309 -4365 8343 -4331
rect 8309 -4437 8343 -4403
rect 8309 -4646 8343 -4612
rect 8309 -4718 8343 -4684
rect 8309 -4790 8343 -4756
rect 2523 -4934 2557 -4900
rect 8309 -4862 8343 -4828
rect 2523 -5006 2557 -4972
rect 2523 -5180 2557 -5146
rect 3601 -5290 3635 -5256
rect 2523 -5398 2557 -5364
rect 2181 -5480 2215 -5446
rect 3061 -5480 3095 -5446
rect 8309 -4934 8343 -4900
rect 8309 -5006 8343 -4972
rect 8309 -5290 8343 -5256
rect 7229 -5398 7263 -5364
rect 2191 -6574 2225 -6540
rect 3071 -6656 3105 -6622
rect 4645 -6820 4679 -6786
rect 6184 -6738 6218 -6704
rect 7976 -6574 8010 -6540
rect 7099 -6656 7133 -6622
rect -41 -7025 -7 -6991
rect 31 -7025 65 -6991
rect 103 -7025 137 -6991
rect 175 -7025 209 -6991
rect 247 -7025 281 -6991
rect 319 -7025 353 -6991
rect 391 -7025 425 -6991
rect 463 -7025 497 -6991
rect 535 -7025 569 -6991
rect 607 -7025 641 -6991
rect 679 -7025 713 -6991
rect 751 -7025 785 -6991
rect 823 -7025 857 -6991
rect 895 -7025 929 -6991
rect 967 -7025 1001 -6991
rect 1039 -7025 1073 -6991
rect 1111 -7025 1145 -6991
rect 1183 -7025 1217 -6991
rect 1278 -7025 1312 -6991
rect 1350 -7025 1384 -6991
rect 1422 -7025 1456 -6991
rect 1494 -7025 1528 -6991
rect 1566 -7025 1600 -6991
rect 1638 -7025 1672 -6991
rect 1710 -7025 1744 -6991
rect 1782 -7025 1816 -6991
rect 1854 -7025 1888 -6991
rect 1926 -7025 1960 -6991
rect 1998 -7025 2032 -6991
rect 2070 -7025 2104 -6991
rect 2142 -7025 2176 -6991
rect 2214 -7025 2248 -6991
rect 2286 -7025 2320 -6991
rect 2358 -7025 2392 -6991
rect 2430 -7025 2464 -6991
rect 2502 -7025 2536 -6991
rect 2574 -7025 2608 -6991
rect 2646 -7025 2680 -6991
rect 2718 -7025 2752 -6991
rect 2790 -7025 2824 -6991
rect 2862 -7025 2896 -6991
rect 2934 -7025 2968 -6991
rect 3006 -7025 3040 -6991
rect 3078 -7025 3112 -6991
rect 3150 -7025 3184 -6991
rect 3222 -7025 3256 -6991
rect 3294 -7025 3328 -6991
rect 3366 -7025 3400 -6991
rect 3438 -7025 3472 -6991
rect 3510 -7025 3544 -6991
rect 3582 -7025 3616 -6991
rect 3654 -7025 3688 -6991
rect 3726 -7025 3760 -6991
rect 3798 -7025 3832 -6991
rect 3893 -7025 3927 -6991
rect 3965 -7025 3999 -6991
rect 4037 -7025 4071 -6991
rect 4109 -7025 4143 -6991
rect 4181 -7025 4215 -6991
rect 4253 -7025 4287 -6991
rect 4325 -7025 4359 -6991
rect 4397 -7025 4431 -6991
rect 4469 -7025 4503 -6991
rect 4541 -7025 4575 -6991
rect 4613 -7025 4647 -6991
rect 4685 -7025 4719 -6991
rect 4757 -7025 4791 -6991
rect 4829 -7025 4863 -6991
rect 4901 -7025 4935 -6991
rect 4973 -7025 5007 -6991
rect 5045 -7025 5079 -6991
rect 5117 -7025 5151 -6991
rect 5189 -7025 5223 -6991
rect 5261 -7025 5295 -6991
rect 5333 -7025 5367 -6991
rect 5405 -7025 5439 -6991
rect 5477 -7025 5511 -6991
rect 5549 -7025 5583 -6991
rect 5621 -7025 5655 -6991
rect 5693 -7025 5727 -6991
rect 5765 -7025 5799 -6991
rect 5837 -7025 5871 -6991
rect 5909 -7025 5943 -6991
rect 5981 -7025 6015 -6991
rect 6053 -7025 6087 -6991
rect 6125 -7025 6159 -6991
rect 6197 -7025 6231 -6991
rect 6269 -7025 6303 -6991
rect 6341 -7025 6375 -6991
rect 6413 -7025 6447 -6991
rect 6508 -7025 6542 -6991
rect 6580 -7025 6614 -6991
rect 6652 -7025 6686 -6991
rect 6724 -7025 6758 -6991
rect 6796 -7025 6830 -6991
rect 6868 -7025 6902 -6991
rect 6940 -7025 6974 -6991
rect 7012 -7025 7046 -6991
rect 7084 -7025 7118 -6991
rect 7156 -7025 7190 -6991
rect 7228 -7025 7262 -6991
rect 7300 -7025 7334 -6991
rect 7372 -7025 7406 -6991
rect 7444 -7025 7478 -6991
rect 7516 -7025 7550 -6991
rect 7588 -7025 7622 -6991
rect 7660 -7025 7694 -6991
rect 7732 -7025 7766 -6991
rect 7804 -7025 7838 -6991
rect 7876 -7025 7910 -6991
rect 7948 -7025 7982 -6991
rect 8020 -7025 8054 -6991
rect 8092 -7025 8126 -6991
rect 8164 -7025 8198 -6991
rect 8236 -7025 8270 -6991
rect 8308 -7025 8342 -6991
rect 8380 -7025 8414 -6991
rect 8452 -7025 8486 -6991
rect 8524 -7025 8558 -6991
rect 8596 -7025 8630 -6991
rect 8668 -7025 8702 -6991
rect 8740 -7025 8774 -6991
rect 8812 -7025 8846 -6991
rect 8884 -7025 8918 -6991
rect 8956 -7025 8990 -6991
rect 9028 -7025 9062 -6991
rect 9123 -7025 9157 -6991
rect 9195 -7025 9229 -6991
rect 9267 -7025 9301 -6991
rect 9339 -7025 9373 -6991
rect 9411 -7025 9445 -6991
rect 9483 -7025 9517 -6991
rect 9555 -7025 9589 -6991
rect 9627 -7025 9661 -6991
rect 9699 -7025 9733 -6991
rect 9771 -7025 9805 -6991
rect 9843 -7025 9877 -6991
rect 9915 -7025 9949 -6991
rect 9987 -7025 10021 -6991
rect 10059 -7025 10093 -6991
rect 10131 -7025 10165 -6991
rect 10203 -7025 10237 -6991
rect 10275 -7025 10309 -6991
rect 10347 -7025 10381 -6991
<< metal1 >>
rect -101 -3455 10466 -3422
rect -101 -3489 -40 -3455
rect -6 -3489 32 -3455
rect 66 -3489 104 -3455
rect 138 -3489 176 -3455
rect 210 -3489 248 -3455
rect 282 -3489 320 -3455
rect 354 -3489 392 -3455
rect 426 -3489 464 -3455
rect 498 -3489 536 -3455
rect 570 -3489 608 -3455
rect 642 -3489 680 -3455
rect 714 -3489 752 -3455
rect 786 -3489 824 -3455
rect 858 -3489 896 -3455
rect 930 -3489 968 -3455
rect 1002 -3489 1040 -3455
rect 1074 -3489 1112 -3455
rect 1146 -3489 1184 -3455
rect 1218 -3489 1279 -3455
rect 1313 -3489 1351 -3455
rect 1385 -3489 1423 -3455
rect 1457 -3489 1495 -3455
rect 1529 -3489 1567 -3455
rect 1601 -3489 1639 -3455
rect 1673 -3489 1711 -3455
rect 1745 -3489 1783 -3455
rect 1817 -3489 1855 -3455
rect 1889 -3489 1927 -3455
rect 1961 -3489 1999 -3455
rect 2033 -3489 2071 -3455
rect 2105 -3489 2143 -3455
rect 2177 -3489 2215 -3455
rect 2249 -3489 2287 -3455
rect 2321 -3489 2359 -3455
rect 2393 -3489 2431 -3455
rect 2465 -3489 2503 -3455
rect 2537 -3489 2575 -3455
rect 2609 -3489 2647 -3455
rect 2681 -3489 2719 -3455
rect 2753 -3489 2791 -3455
rect 2825 -3489 2863 -3455
rect 2897 -3489 2935 -3455
rect 2969 -3489 3007 -3455
rect 3041 -3489 3079 -3455
rect 3113 -3489 3151 -3455
rect 3185 -3489 3223 -3455
rect 3257 -3489 3295 -3455
rect 3329 -3489 3367 -3455
rect 3401 -3489 3439 -3455
rect 3473 -3489 3511 -3455
rect 3545 -3489 3583 -3455
rect 3617 -3489 3655 -3455
rect 3689 -3489 3727 -3455
rect 3761 -3489 3799 -3455
rect 3833 -3489 3894 -3455
rect 3928 -3489 3966 -3455
rect 4000 -3489 4038 -3455
rect 4072 -3489 4110 -3455
rect 4144 -3489 4182 -3455
rect 4216 -3489 4254 -3455
rect 4288 -3489 4326 -3455
rect 4360 -3489 4398 -3455
rect 4432 -3489 4470 -3455
rect 4504 -3489 4542 -3455
rect 4576 -3489 4614 -3455
rect 4648 -3489 4686 -3455
rect 4720 -3489 4758 -3455
rect 4792 -3489 4830 -3455
rect 4864 -3489 4902 -3455
rect 4936 -3489 4974 -3455
rect 5008 -3489 5046 -3455
rect 5080 -3489 5118 -3455
rect 5152 -3489 5190 -3455
rect 5224 -3489 5262 -3455
rect 5296 -3489 5334 -3455
rect 5368 -3489 5406 -3455
rect 5440 -3489 5478 -3455
rect 5512 -3489 5550 -3455
rect 5584 -3489 5622 -3455
rect 5656 -3489 5694 -3455
rect 5728 -3489 5766 -3455
rect 5800 -3489 5838 -3455
rect 5872 -3489 5910 -3455
rect 5944 -3489 5982 -3455
rect 6016 -3489 6054 -3455
rect 6088 -3489 6126 -3455
rect 6160 -3489 6198 -3455
rect 6232 -3489 6270 -3455
rect 6304 -3489 6342 -3455
rect 6376 -3489 6414 -3455
rect 6448 -3489 6509 -3455
rect 6543 -3489 6581 -3455
rect 6615 -3489 6653 -3455
rect 6687 -3489 6725 -3455
rect 6759 -3489 6797 -3455
rect 6831 -3489 6869 -3455
rect 6903 -3489 6941 -3455
rect 6975 -3489 7013 -3455
rect 7047 -3489 7085 -3455
rect 7119 -3489 7157 -3455
rect 7191 -3489 7229 -3455
rect 7263 -3489 7301 -3455
rect 7335 -3489 7373 -3455
rect 7407 -3489 7445 -3455
rect 7479 -3489 7517 -3455
rect 7551 -3489 7589 -3455
rect 7623 -3489 7661 -3455
rect 7695 -3489 7733 -3455
rect 7767 -3489 7805 -3455
rect 7839 -3489 7877 -3455
rect 7911 -3489 7949 -3455
rect 7983 -3489 8021 -3455
rect 8055 -3489 8093 -3455
rect 8127 -3489 8165 -3455
rect 8199 -3489 8237 -3455
rect 8271 -3489 8309 -3455
rect 8343 -3489 8381 -3455
rect 8415 -3489 8453 -3455
rect 8487 -3489 8525 -3455
rect 8559 -3489 8597 -3455
rect 8631 -3489 8669 -3455
rect 8703 -3489 8741 -3455
rect 8775 -3489 8813 -3455
rect 8847 -3489 8885 -3455
rect 8919 -3489 8957 -3455
rect 8991 -3489 9029 -3455
rect 9063 -3489 9124 -3455
rect 9158 -3489 9196 -3455
rect 9230 -3489 9268 -3455
rect 9302 -3489 9340 -3455
rect 9374 -3489 9412 -3455
rect 9446 -3489 9484 -3455
rect 9518 -3489 9556 -3455
rect 9590 -3489 9628 -3455
rect 9662 -3489 9700 -3455
rect 9734 -3489 9772 -3455
rect 9806 -3489 9844 -3455
rect 9878 -3489 9916 -3455
rect 9950 -3489 9988 -3455
rect 10022 -3489 10060 -3455
rect 10094 -3489 10132 -3455
rect 10166 -3489 10204 -3455
rect 10238 -3489 10276 -3455
rect 10310 -3489 10348 -3455
rect 10382 -3489 10466 -3455
rect -101 -3522 10466 -3489
rect 2184 -3743 2264 -3720
rect 2184 -3746 2207 -3743
rect 1802 -3774 2207 -3746
rect 2184 -3777 2207 -3774
rect 2241 -3777 2264 -3743
rect 2184 -3800 2264 -3777
rect 2515 -4043 2565 -3522
rect 2515 -4077 2523 -4043
rect 2557 -4077 2565 -4043
rect 2515 -4115 2565 -4077
rect 2515 -4149 2523 -4115
rect 2557 -4149 2565 -4115
rect 2515 -4187 2565 -4149
rect 2515 -4221 2523 -4187
rect 2557 -4221 2565 -4187
rect 2515 -4259 2565 -4221
rect 2515 -4293 2523 -4259
rect 2557 -4293 2565 -4259
rect 2515 -4331 2565 -4293
rect 2515 -4365 2523 -4331
rect 2557 -4365 2565 -4331
rect 2515 -4403 2565 -4365
rect 2515 -4437 2523 -4403
rect 2557 -4437 2565 -4403
rect 2515 -4450 2565 -4437
rect 8301 -4043 8351 -3522
rect 8301 -4077 8309 -4043
rect 8343 -4077 8351 -4043
rect 8301 -4115 8351 -4077
rect 8301 -4149 8309 -4115
rect 8343 -4149 8351 -4115
rect 8301 -4187 8351 -4149
rect 8301 -4221 8309 -4187
rect 8343 -4221 8351 -4187
rect 8301 -4259 8351 -4221
rect 8301 -4293 8309 -4259
rect 8343 -4293 8351 -4259
rect 8301 -4331 8351 -4293
rect 8301 -4365 8309 -4331
rect 8343 -4365 8351 -4331
rect 8301 -4403 8351 -4365
rect 8301 -4437 8309 -4403
rect 8343 -4437 8351 -4403
rect 8301 -4450 8351 -4437
rect 2515 -4612 2565 -4598
rect 2515 -4646 2523 -4612
rect 2557 -4646 2565 -4612
rect 2515 -4684 2565 -4646
rect 2515 -4718 2523 -4684
rect 2557 -4718 2565 -4684
rect 2515 -4756 2565 -4718
rect 2515 -4790 2523 -4756
rect 2557 -4790 2565 -4756
rect 2515 -4828 2565 -4790
rect 2515 -4862 2523 -4828
rect 2557 -4862 2565 -4828
rect 2515 -4900 2565 -4862
rect 2515 -4934 2523 -4900
rect 2557 -4934 2565 -4900
rect 2515 -4972 2565 -4934
rect 2515 -5006 2523 -4972
rect 2557 -5006 2565 -4972
rect 2515 -5019 2565 -5006
rect 8301 -4612 8351 -4598
rect 8301 -4646 8309 -4612
rect 8343 -4646 8351 -4612
rect 8301 -4684 8351 -4646
rect 8301 -4718 8309 -4684
rect 8343 -4718 8351 -4684
rect 8301 -4756 8351 -4718
rect 8301 -4790 8309 -4756
rect 8343 -4790 8351 -4756
rect 8301 -4828 8351 -4790
rect 8301 -4862 8309 -4828
rect 8343 -4862 8351 -4828
rect 8301 -4900 8351 -4862
rect 8301 -4934 8309 -4900
rect 8343 -4934 8351 -4900
rect 8301 -4972 8351 -4934
rect 8301 -5006 8309 -4972
rect 8343 -5006 8351 -4972
rect 8301 -5019 8351 -5006
rect 2500 -5137 2580 -5123
rect 2500 -5189 2514 -5137
rect 2566 -5189 2580 -5137
rect 2500 -5203 2580 -5189
rect 3578 -5256 3658 -5233
rect 3578 -5290 3601 -5256
rect 3635 -5260 3658 -5256
rect 8286 -5247 8366 -5233
rect 8286 -5260 8300 -5247
rect 3635 -5288 8300 -5260
rect 3635 -5290 3658 -5288
rect 3578 -5313 3658 -5290
rect 8286 -5299 8300 -5288
rect 8352 -5299 8366 -5247
rect 8286 -5313 8366 -5299
rect 2500 -5364 2580 -5341
rect 1802 -5395 2294 -5367
rect 2158 -5446 2238 -5423
rect 2158 -5450 2181 -5446
rect 1802 -5478 2181 -5450
rect 2158 -5480 2181 -5478
rect 2215 -5480 2238 -5446
rect 2266 -5451 2294 -5395
rect 2500 -5398 2523 -5364
rect 2557 -5367 2580 -5364
rect 7206 -5364 7286 -5341
rect 7206 -5367 7229 -5364
rect 2557 -5395 7229 -5367
rect 2557 -5398 2580 -5395
rect 2500 -5421 2580 -5398
rect 7206 -5398 7229 -5395
rect 7263 -5398 7286 -5364
rect 7206 -5421 7286 -5398
rect 3038 -5446 3118 -5423
rect 3038 -5451 3061 -5446
rect 2266 -5479 3061 -5451
rect 2158 -5503 2238 -5480
rect 3038 -5480 3061 -5479
rect 3095 -5480 3118 -5446
rect 3038 -5503 3118 -5480
rect 2168 -6540 2248 -6517
rect 2168 -6574 2191 -6540
rect 2225 -6543 2248 -6540
rect 7953 -6540 8033 -6517
rect 7953 -6543 7976 -6540
rect 2225 -6571 7976 -6543
rect 2225 -6574 2248 -6571
rect 2168 -6597 2248 -6574
rect 7953 -6574 7976 -6571
rect 8010 -6574 8033 -6540
rect 7953 -6597 8033 -6574
rect 3048 -6622 3128 -6599
rect 3048 -6656 3071 -6622
rect 3105 -6625 3128 -6622
rect 7076 -6622 7156 -6599
rect 7076 -6625 7099 -6622
rect 3105 -6653 7099 -6625
rect 3105 -6656 3128 -6653
rect 3048 -6679 3128 -6656
rect 7076 -6656 7099 -6653
rect 7133 -6656 7156 -6622
rect 7076 -6679 7156 -6656
rect 6161 -6704 6241 -6681
rect 6161 -6707 6184 -6704
rect 1802 -6735 6184 -6707
rect 6161 -6738 6184 -6735
rect 6218 -6738 6241 -6704
rect 6161 -6761 6241 -6738
rect 4622 -6786 4702 -6763
rect 4622 -6790 4645 -6786
rect 1802 -6818 4645 -6790
rect 4622 -6820 4645 -6818
rect 4679 -6820 4702 -6786
rect 4622 -6843 4702 -6820
rect -102 -6991 10465 -6958
rect -102 -7025 -41 -6991
rect -7 -7025 31 -6991
rect 65 -7025 103 -6991
rect 137 -7025 175 -6991
rect 209 -7025 247 -6991
rect 281 -7025 319 -6991
rect 353 -7025 391 -6991
rect 425 -7025 463 -6991
rect 497 -7025 535 -6991
rect 569 -7025 607 -6991
rect 641 -7025 679 -6991
rect 713 -7025 751 -6991
rect 785 -7025 823 -6991
rect 857 -7025 895 -6991
rect 929 -7025 967 -6991
rect 1001 -7025 1039 -6991
rect 1073 -7025 1111 -6991
rect 1145 -7025 1183 -6991
rect 1217 -7025 1278 -6991
rect 1312 -7025 1350 -6991
rect 1384 -7025 1422 -6991
rect 1456 -7025 1494 -6991
rect 1528 -7025 1566 -6991
rect 1600 -7025 1638 -6991
rect 1672 -7025 1710 -6991
rect 1744 -7025 1782 -6991
rect 1816 -7025 1854 -6991
rect 1888 -7025 1926 -6991
rect 1960 -7025 1998 -6991
rect 2032 -7025 2070 -6991
rect 2104 -7025 2142 -6991
rect 2176 -7025 2214 -6991
rect 2248 -7025 2286 -6991
rect 2320 -7025 2358 -6991
rect 2392 -7025 2430 -6991
rect 2464 -7025 2502 -6991
rect 2536 -7025 2574 -6991
rect 2608 -7025 2646 -6991
rect 2680 -7025 2718 -6991
rect 2752 -7025 2790 -6991
rect 2824 -7025 2862 -6991
rect 2896 -7025 2934 -6991
rect 2968 -7025 3006 -6991
rect 3040 -7025 3078 -6991
rect 3112 -7025 3150 -6991
rect 3184 -7025 3222 -6991
rect 3256 -7025 3294 -6991
rect 3328 -7025 3366 -6991
rect 3400 -7025 3438 -6991
rect 3472 -7025 3510 -6991
rect 3544 -7025 3582 -6991
rect 3616 -7025 3654 -6991
rect 3688 -7025 3726 -6991
rect 3760 -7025 3798 -6991
rect 3832 -7025 3893 -6991
rect 3927 -7025 3965 -6991
rect 3999 -7025 4037 -6991
rect 4071 -7025 4109 -6991
rect 4143 -7025 4181 -6991
rect 4215 -7025 4253 -6991
rect 4287 -7025 4325 -6991
rect 4359 -7025 4397 -6991
rect 4431 -7025 4469 -6991
rect 4503 -7025 4541 -6991
rect 4575 -7025 4613 -6991
rect 4647 -7025 4685 -6991
rect 4719 -7025 4757 -6991
rect 4791 -7025 4829 -6991
rect 4863 -7025 4901 -6991
rect 4935 -7025 4973 -6991
rect 5007 -7025 5045 -6991
rect 5079 -7025 5117 -6991
rect 5151 -7025 5189 -6991
rect 5223 -7025 5261 -6991
rect 5295 -7025 5333 -6991
rect 5367 -7025 5405 -6991
rect 5439 -7025 5477 -6991
rect 5511 -7025 5549 -6991
rect 5583 -7025 5621 -6991
rect 5655 -7025 5693 -6991
rect 5727 -7025 5765 -6991
rect 5799 -7025 5837 -6991
rect 5871 -7025 5909 -6991
rect 5943 -7025 5981 -6991
rect 6015 -7025 6053 -6991
rect 6087 -7025 6125 -6991
rect 6159 -7025 6197 -6991
rect 6231 -7025 6269 -6991
rect 6303 -7025 6341 -6991
rect 6375 -7025 6413 -6991
rect 6447 -7025 6508 -6991
rect 6542 -7025 6580 -6991
rect 6614 -7025 6652 -6991
rect 6686 -7025 6724 -6991
rect 6758 -7025 6796 -6991
rect 6830 -7025 6868 -6991
rect 6902 -7025 6940 -6991
rect 6974 -7025 7012 -6991
rect 7046 -7025 7084 -6991
rect 7118 -7025 7156 -6991
rect 7190 -7025 7228 -6991
rect 7262 -7025 7300 -6991
rect 7334 -7025 7372 -6991
rect 7406 -7025 7444 -6991
rect 7478 -7025 7516 -6991
rect 7550 -7025 7588 -6991
rect 7622 -7025 7660 -6991
rect 7694 -7025 7732 -6991
rect 7766 -7025 7804 -6991
rect 7838 -7025 7876 -6991
rect 7910 -7025 7948 -6991
rect 7982 -7025 8020 -6991
rect 8054 -7025 8092 -6991
rect 8126 -7025 8164 -6991
rect 8198 -7025 8236 -6991
rect 8270 -7025 8308 -6991
rect 8342 -7025 8380 -6991
rect 8414 -7025 8452 -6991
rect 8486 -7025 8524 -6991
rect 8558 -7025 8596 -6991
rect 8630 -7025 8668 -6991
rect 8702 -7025 8740 -6991
rect 8774 -7025 8812 -6991
rect 8846 -7025 8884 -6991
rect 8918 -7025 8956 -6991
rect 8990 -7025 9028 -6991
rect 9062 -7025 9123 -6991
rect 9157 -7025 9195 -6991
rect 9229 -7025 9267 -6991
rect 9301 -7025 9339 -6991
rect 9373 -7025 9411 -6991
rect 9445 -7025 9483 -6991
rect 9517 -7025 9555 -6991
rect 9589 -7025 9627 -6991
rect 9661 -7025 9699 -6991
rect 9733 -7025 9771 -6991
rect 9805 -7025 9843 -6991
rect 9877 -7025 9915 -6991
rect 9949 -7025 9987 -6991
rect 10021 -7025 10059 -6991
rect 10093 -7025 10131 -6991
rect 10165 -7025 10203 -6991
rect 10237 -7025 10275 -6991
rect 10309 -7025 10347 -6991
rect 10381 -7025 10465 -6991
rect -102 -7058 10465 -7025
<< via1 >>
rect 2514 -5146 2566 -5137
rect 2514 -5180 2523 -5146
rect 2523 -5180 2557 -5146
rect 2557 -5180 2566 -5146
rect 2514 -5189 2566 -5180
rect 8300 -5256 8352 -5247
rect 8300 -5290 8309 -5256
rect 8309 -5290 8343 -5256
rect 8343 -5290 8352 -5256
rect 8300 -5299 8352 -5290
<< metal2 >>
rect 2332 -5149 2360 -3364
rect 2500 -5137 2580 -5123
rect 2500 -5149 2514 -5137
rect 2332 -5177 2514 -5149
rect 2500 -5189 2514 -5177
rect 2566 -5189 2580 -5137
rect 2500 -5203 2580 -5189
rect 8286 -5247 8366 -5233
rect 8286 -5299 8300 -5247
rect 8352 -5259 8366 -5247
rect 8506 -5259 8534 -3364
rect 8352 -5287 8534 -5259
rect 8352 -5299 8366 -5287
rect 8286 -5313 8366 -5299
<< labels >>
flabel metal1 s 1815 -3768 1830 -3755 2 FreeSans 100000 0 0 0 v_bias_p
port 1 nsew
flabel metal1 s 5333 -7025 5512 -6991 2 FreeSans 100000 0 0 0 Ground
port 2 nsew
flabel metal1 s 5368 -3489 5406 -3455 2 FreeSans 100000 0 0 0 VDD
port 3 nsew
flabel metal1 s 1811 -6812 1826 -6796 2 FreeSans 100000 0 0 0 RFP
port 4 nsew
flabel metal1 s 1811 -6729 1826 -6713 2 FreeSans 100000 0 0 0 RFN
port 5 nsew
flabel metal1 s 1815 -5473 1833 -5456 2 FreeSans 100000 0 0 0 LOP
port 6 nsew
flabel metal1 s 1816 -5390 1834 -5373 2 FreeSans 100000 0 0 0 LON
port 7 nsew
flabel metal2 s 2381 -5169 2397 -5156 2 FreeSans 100000 0 0 0 VoutP
port 8 nsew
flabel metal2 s 8448 -5281 8467 -5264 2 FreeSans 100000 0 0 0 VoutN
port 9 nsew
<< properties >>
string path 18.780 -3.635 18.780 5.750 
<< end >>
