magic
tech sky130A
timestamp 1662343253
<< nwell >>
rect -1260 650 -1025 1000
<< nmos >>
rect -1120 465 -1105 615
<< pmos >>
rect -1120 675 -1105 975
<< ndiff >>
rect -1180 600 -1120 615
rect -1180 480 -1165 600
rect -1135 480 -1120 600
rect -1180 465 -1120 480
rect -1105 600 -1045 615
rect -1105 480 -1090 600
rect -1060 480 -1045 600
rect -1105 465 -1045 480
<< pdiff >>
rect -1180 960 -1120 975
rect -1180 690 -1165 960
rect -1135 690 -1120 960
rect -1180 675 -1120 690
rect -1105 960 -1045 975
rect -1105 690 -1090 960
rect -1060 690 -1045 960
rect -1105 675 -1045 690
<< ndiffc >>
rect -1165 480 -1135 600
rect -1090 480 -1060 600
<< pdiffc >>
rect -1165 690 -1135 960
rect -1090 690 -1060 960
<< psubdiff >>
rect -1240 600 -1180 615
rect -1240 480 -1225 600
rect -1195 480 -1180 600
rect -1240 465 -1180 480
<< nsubdiff >>
rect -1240 960 -1180 975
rect -1240 690 -1225 960
rect -1195 690 -1180 960
rect -1240 675 -1180 690
<< psubdiffcont >>
rect -1225 480 -1195 600
<< nsubdiffcont >>
rect -1225 690 -1195 960
<< poly >>
rect -1120 975 -1105 990
rect -1120 615 -1105 675
rect -1120 450 -1105 465
rect -1145 440 -1105 450
rect -1145 420 -1135 440
rect -1115 420 -1105 440
rect -1145 410 -1105 420
<< polycont >>
rect -1135 420 -1115 440
<< locali >>
rect -1235 960 -1125 970
rect -1235 690 -1225 960
rect -1195 690 -1165 960
rect -1135 690 -1125 960
rect -1235 680 -1125 690
rect -1100 960 -1050 965
rect -1100 690 -1090 960
rect -1060 690 -1050 960
rect -1100 680 -1050 690
rect -1075 610 -1050 680
rect -1235 600 -1125 610
rect -1235 480 -1225 600
rect -1195 480 -1165 600
rect -1135 480 -1125 600
rect -1235 470 -1125 480
rect -1100 600 -1050 610
rect -1100 480 -1090 600
rect -1060 480 -1050 600
rect -1100 470 -1050 480
rect -1075 450 -1050 470
rect -1260 440 -1105 450
rect -1260 430 -1135 440
rect -1145 420 -1135 430
rect -1115 420 -1105 440
rect -1075 430 -1025 450
rect -1145 410 -1105 420
<< viali >>
rect -1225 690 -1195 960
rect -1165 690 -1135 960
rect -1225 480 -1195 600
rect -1165 480 -1135 600
<< metal1 >>
rect -1260 960 -1125 970
rect -1260 690 -1225 960
rect -1195 690 -1165 960
rect -1135 690 -1125 960
rect -1260 680 -1125 690
rect -1260 600 -1125 610
rect -1260 480 -1225 600
rect -1195 480 -1165 600
rect -1135 480 -1125 600
rect -1260 470 -1125 480
<< labels >>
rlabel locali -1025 440 -1025 440 3 OUT
port 3 e
rlabel metal1 -1260 810 -1260 810 7 VP
port 1 w
rlabel metal1 -1260 535 -1260 535 7 VN
port 4 w
rlabel locali -1260 440 -1260 440 7 A
port 2 w
<< end >>
