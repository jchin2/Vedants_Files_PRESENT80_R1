magic
tech sky130A
magscale 1 2
timestamp 1671058898
<< poly >>
rect -44 226 44 242
rect -44 192 -17 226
rect 17 192 44 226
rect -44 169 44 192
rect -44 -192 44 -169
rect -44 -226 -17 -192
rect 17 -226 44 -192
rect -44 -242 44 -226
<< polycont >>
rect -17 192 17 226
rect -17 -226 17 -192
<< npolyres >>
rect -44 -169 44 169
<< locali >>
rect -44 192 -17 226
rect 17 192 44 226
rect -28 189 -17 192
rect 17 189 28 192
rect -28 186 28 189
rect -28 -189 28 -186
rect -28 -192 -17 -189
rect 17 -192 28 -189
rect -44 -226 -17 -192
rect 17 -226 44 -192
<< viali >>
rect -17 192 17 223
rect -17 189 17 192
rect -17 -192 17 -189
rect -17 -223 17 -192
<< metal1 >>
rect -40 223 40 232
rect -40 189 -17 223
rect 17 189 40 223
rect -40 180 40 189
rect -40 -189 40 -180
rect -40 -223 -17 -189
rect 17 -223 40 -189
rect -40 -232 40 -223
<< end >>
