* NGSPICE file created from EESPFAL_Sbox_flat.ext - technology: sky130A

.subckt EESPFAL_Sbox_flat GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar Dis1 Dis2 Dis3
+ s0 s0_bar s1_bar s1 s2 s2_bar s3_bar s3 CLK1 CLK2 CLK3
X0 CLK2.t52 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t5 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 CLK2.t51 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B Dis1.t0 GND.t229 GND.t204 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X2 CLK2.t21 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar GND.t97 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X3 GND.t309 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t3 GND.t85 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 CLK1.t56 x1.t0 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B GND.t163 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X5 CLK1.t151 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t5 CLK1.t150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_1170_n10570# x3_bar.t0 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t0 GND.t162 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t4 Dis1.t1 GND.t228 GND.t187 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t3 Dis2.t0 GND.t149 GND.t148 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 CLK2.t30 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_6859_n7070# GND.t121 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X10 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A x0.t0 a_3070_n7070# GND.t59 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X11 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t6 CLK1.t42 CLK1.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 GND.t86 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar GND.t85 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_1510_n7070# x1.t1 CLK1.t55 GND.t161 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X14 CLK3.t27 s0.t6 s0_bar.t3 CLK3.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 CLK2.t91 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t6 a_6800_n10570# GND.t140 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X16 CLK1.t101 x1_bar.t0 a_1170_n2029# GND.t91 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X17 CLK3.t17 s2_bar.t5 s2.t3 CLK3.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 CLK3.t42 s1.t7 s1_bar.t3 CLK3.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar x1.t2 CLK1.t58 GND.t39 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X20 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t0 x3.t0 a_3030_n2029# GND.t164 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X21 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar GND.t254 GND.t132 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X22 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar Dis2.t1 GND.t151 GND.t150 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X23 s0.t0 Dis3.t0 GND.t31 GND.t30 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X24 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar CLK1.t79 CLK1.t78 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X25 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar Dis1.t2 GND.t226 GND.t200 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X26 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar x0.t1 a_1510_n7070# GND.t63 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X27 a_1470_n2029# x1.t3 CLK1.t62 GND.t165 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X28 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t5 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t6 CLK1.t185 CLK1.t184 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X29 a_2730_791# x1_bar.t1 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B GND.t110 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X30 s2_bar.t4 s2.t7 CLK3.t37 CLK3.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X31 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t6 CLK2.t50 CLK2.t49 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X32 CLK2.t62 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t3 CLK2.t61 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X33 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t0 Dis2.t2 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X34 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t2 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t7 CLK2.t90 GND.t50 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X35 CLK2.t48 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t5 GND.t154 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X36 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t5 Dis1.t3 GND.t227 GND.t198 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X37 CLK1.t131 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t6 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t4 CLK1.t130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X38 CLK2.t22 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t4 GND.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X39 CLK1.t15 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B CLK1.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X40 a_1170_n9890# x0_bar.t0 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t0 GND.t162 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X41 CLK2.t38 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B CLK2.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X42 CLK1.t99 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar CLK1.t98 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X43 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/B CLK1.t46 CLK1.t45 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X44 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar x0.t2 CLK1.t24 GND.t46 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X45 CLK1.t93 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t6 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t4 CLK1.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X46 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t4 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t6 CLK2.t12 GND.t79 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X47 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t6 GND.t89 GND.t88 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X48 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t6 CLK1.t30 CLK1.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X49 a_3030_n9890# x1_bar.t2 CLK1.t186 GND.t106 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X50 CLK1.t33 x2_bar.t0 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X51 CLK2.t68 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t5 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 CLK2.t67 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X52 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar Dis1.t4 GND.t225 GND.t150 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X53 CLK1.t26 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t6 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t5 CLK1.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X54 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B CLK1.t176 CLK1.t175 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X55 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar GND.t172 GND.t171 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X56 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t3 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t6 CLK1.t89 CLK1.t88 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X57 s0_bar.t1 s0.t7 GND.t65 GND.t64 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X58 a_2770_n7750# x2_bar.t1 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t1 GND.t62 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X59 CLK1.t187 x1_bar.t3 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar GND.t288 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X60 GND.t224 Dis1.t5 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t4 GND.t192 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X61 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B CLK1.t11 CLK1.t10 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X62 GND.t105 s1_bar.t5 s1.t1 GND.t104 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X63 GND.t109 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t7 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t3 GND.t108 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X64 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t0 x3.t1 a_3030_1471# GND.t170 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X65 CLK1.t60 x1.t4 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar GND.t55 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X66 GND.t223 Dis1.t6 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t5 GND.t206 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X67 GND.t222 Dis1.t7 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t4 GND.t183 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X68 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar Dis2.t3 GND.t18 GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X69 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar Dis1.t8 GND.t221 GND.t220 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X70 GND.t5 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar GND.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X71 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t0 x3.t2 a_1470_1471# GND.t80 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X72 CLK2.t87 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT CLK2.t86 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X73 CLK1.t180 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t7 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t5 CLK1.t179 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X74 CLK1.t9 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar CLK1.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X75 CLK2.t110 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t5 CLK2.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X76 GND.t136 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_INV4_2/A_bar GND.t135 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.6e+12p ps=1.68e+07u w=1.5e+06u l=150000u
X77 CLK1.t134 x3_bar.t1 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B GND.t163 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X78 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A CLK1.t97 CLK1.t96 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X79 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar Dis1.t9 GND.t219 GND.t213 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X80 GND.t218 Dis1.t10 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B GND.t211 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X81 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar GND.t235 GND.t152 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X82 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t5 CLK2.t114 CLK2.t113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X83 s1_bar.t1 s1.t8 GND.t314 GND.t313 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X84 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t7 GND.t74 GND.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X85 a_7190_n4930# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar a_7040_n4930# GND.t130 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X86 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar CLK2.t79 GND.t252 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X87 CLK1.t61 x1.t5 a_2730_n9890# GND.t56 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X88 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar GND.t102 GND.t101 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X89 GND.t124 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar GND.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X90 CLK1.t170 x3_bar.t2 a_3070_n4929# GND.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X91 s3_bar.t3 s3.t7 CLK3.t46 CLK3.t45 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X92 CLK1.t161 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar EESPFAL_s3_0/EESPFAL_INV4_0/A CLK1.t160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X93 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t1 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 GND.t299 GND.t298 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X94 CLK1.t27 x2_bar.t2 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B GND.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X95 GND.t217 Dis1.t11 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B GND.t194 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X96 CLK2.t25 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t6 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 CLK2.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X97 a_2730_n1349# x0_bar.t1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t3 GND.t113 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X98 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar CLK1.t167 CLK1.t166 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X99 CLK3.t38 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t6 a_7190_n4930# GND.t40 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X100 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NOR_v3_0/B CLK2.t100 CLK2.t99 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X101 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t8 CLK1.t140 CLK1.t139 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X102 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT CLK2.t3 CLK2.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X103 CLK1.t6 x1_bar.t4 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar GND.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X104 s0.t1 s0_bar.t5 CLK3.t21 CLK3.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X105 GND.t283 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X106 s1.t3 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t7 CLK3.t15 GND.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X107 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t0 x0.t3 a_1470_n1349# GND.t47 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X108 CLK2.t18 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar CLK2.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X109 s2.t0 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT CLK3.t0 GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X110 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar x3_bar.t3 CLK1.t171 GND.t142 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X111 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar Dis1.t12 GND.t216 GND.t215 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X112 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT CLK2.t108 CLK2.t107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X113 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar x3.t3 CLK1.t183 GND.t284 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X114 CLK1.t178 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t8 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t5 CLK1.t177 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X115 EESPFAL_s3_0/EESPFAL_INV4_0/A EESPFAL_s3_0/EESPFAL_INV4_0/A_bar GND.t251 GND.t250 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X116 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar GND.t129 GND.t128 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X117 CLK2.t80 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar GND.t147 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X118 CLK3.t10 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT s0.t4 GND.t115 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X119 GND.t33 Dis3.t1 s2_bar.t0 GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X120 s3.t1 s3_bar.t5 CLK3.t8 CLK3.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X121 CLK2.t7 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t2 CLK2.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X122 a_1210_n7070# x0_bar.t2 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar GND.t72 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X123 CLK1.t157 EESPFAL_s3_0/EESPFAL_INV4_0/A EESPFAL_s3_0/EESPFAL_INV4_0/A_bar CLK1.t156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X124 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t6 CLK2.t14 CLK2.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X125 CLK2.t78 EESPFAL_s3_0/EESPFAL_INV4_0/A EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t4 GND.t249 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X126 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar Dis2.t4 GND.t270 GND.t269 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X127 a_2730_1471# x3_bar.t4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t2 GND.t110 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X128 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t7 CLK2.t115 GND.t144 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X129 CLK3.t33 s1_bar.t6 s1.t5 CLK3.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X130 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t2 Dis1.t13 GND.t214 GND.t213 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X131 a_6859_n7070# EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B GND.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X132 a_3070_n7070# x1_bar.t5 CLK1.t7 GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X133 GND.t232 Dis3.t2 s3_bar.t0 GND.t231 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X134 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t0 x3.t4 a_3030_n10570# GND.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X135 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar EESPFAL_s1_0/EESPFAL_INV4_0/A CLK1.t138 CLK1.t137 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X136 CLK1.t31 x1_bar.t6 a_1210_n7070# GND.t60 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X137 a_1170_n2029# x3_bar.t5 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t1 GND.t111 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X138 s2.t2 s2_bar.t6 CLK3.t3 CLK3.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X139 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar CLK2.t95 CLK2.t94 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X140 CLK2.t53 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t7 a_5050_791# GND.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X141 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar CLK1.t146 CLK1.t145 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X142 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar CLK2.t66 CLK2.t65 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X143 CLK3.t23 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar a_7070_791# GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X144 CLK3.t14 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t6 a_6971_n12711# GND.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X145 s1_bar.t2 s1.t9 CLK3.t44 CLK3.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X146 GND.t212 Dis1.t14 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B GND.t211 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X147 s0_bar.t2 s0.t8 CLK3.t25 CLK3.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X148 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar EESPFAL_s3_0/EESPFAL_INV4_0/A CLK1.t155 CLK1.t154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X149 a_2731_n12710# x3.t5 EESPFAL_s3_0/EESPFAL_INV4_0/A GND.t70 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X150 a_3030_n2029# x1_bar.t7 CLK1.t32 GND.t61 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X151 a_7070_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT GND.t139 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X152 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t3 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t7 CLK1.t124 CLK1.t123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X153 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar Dis2.t5 GND.t271 GND.t30 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X154 GND.t28 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar GND.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X155 CLK3.t9 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT s3.t2 GND.t84 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X156 GND.t114 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar GND.t82 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X157 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t7 GND.t107 GND.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X158 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar x2.t0 CLK1.t66 GND.t90 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X159 CLK1.t21 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t6 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t0 CLK1.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X160 CLK2.t93 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT CLK2.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X161 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/B CLK1.t111 CLK1.t110 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X162 CLK1.t144 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B CLK1.t143 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X163 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/B CLK1.t3 CLK1.t2 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X164 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_1/B CLK1.t19 CLK1.t18 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X165 GND.t49 s3_bar.t6 s3.t0 GND.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X166 CLK1.t75 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/B CLK1.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X167 CLK1.t194 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t8 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t5 CLK1.t193 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X168 CLK2.t104 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar CLK2.t103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X169 CLK2.t20 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t1 GND.t97 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X170 a_6971_n12711# EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar a_6821_n12711# GND.t262 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X171 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B x1.t6 CLK1.t57 GND.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X172 CLK1.t59 x1.t7 a_2770_n7070# GND.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X173 GND.t208 Dis1.t15 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t5 GND.t181 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X174 GND.t138 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar GND.t137 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X175 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t8 CLK1.t52 CLK1.t51 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X176 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar GND.t297 GND.t171 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X177 GND.t78 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar GND.t77 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X178 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t6 GND.t287 GND.t273 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X179 CLK1.t64 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t8 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t1 CLK1.t63 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X180 CLK1.t147 x2.t1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar GND.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X181 a_3790_1471# x1_bar.t8 CLK1.t117 GND.t147 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X182 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT CLK2.t16 CLK2.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X183 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar CLK1.t13 CLK1.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X184 GND.t210 Dis1.t16 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar GND.t179 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X185 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar CLK2.t36 CLK2.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X186 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar x2.t2 a_3790_1471# GND.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X187 GND.t117 Dis2.t6 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT GND.t116 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X188 GND.t58 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t7 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t1 GND.t57 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X189 CLK1.t53 x1.t8 a_2730_n2029# GND.t41 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X190 a_2730_n10570# x3_bar.t6 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t1 GND.t73 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X191 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar x3_bar.t7 CLK1.t116 GND.t143 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X192 a_6800_n1349# EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT GND.t3 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X193 CLK1.t172 x3_bar.t8 a_2881_n4169# GND.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X194 GND.t119 Dis2.t7 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT GND.t118 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X195 GND.t36 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t8 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t3 GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X196 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t1 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 GND.t100 GND.t99 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X197 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t1 x3.t6 a_1470_n10570# GND.t160 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X198 CLK2.t106 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t9 a_6859_n7750# GND.t121 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X199 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t0 x2.t3 a_3070_n7750# GND.t59 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X200 GND.t207 Dis1.t17 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B GND.t206 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X201 GND.t159 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar GND.t77 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X202 GND.t281 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar GND.t137 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X203 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar Dis1.t18 GND.t209 GND.t173 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X204 s1.t4 Dis3.t3 GND.t234 GND.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X205 a_1510_n7750# x3.t7 CLK1.t129 GND.t161 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X206 CLK2.t89 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t9 a_6800_n1349# GND.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X207 CLK1.t95 x2.t4 a_2730_791# GND.t93 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X208 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t1 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t7 GND.t38 GND.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X209 CLK2.t43 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t3 GND.t134 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X210 GND.t276 Dis2.t8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t0 GND.t275 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X211 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar Dis1.t19 GND.t205 GND.t204 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X212 GND.t203 Dis1.t20 EESPFAL_s1_0/EESPFAL_INV4_0/A GND.t202 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X213 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar GND.t96 GND.t95 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X214 GND.t125 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar GND.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X215 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t5 Dis1.t21 GND.t201 GND.t200 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X216 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t0 x2.t5 a_1510_n7750# GND.t63 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X217 CLK3.t4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t7 a_6971_n4170# GND.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X218 a_7040_n4930# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 s2_bar.t1 GND.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X219 CLK1.t28 x2_bar.t3 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar GND.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X220 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t7 CLK1.t133 CLK1.t132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X221 a_2730_n9890# x0_bar.t3 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t2 GND.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X222 s1.t0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT CLK3.t1 GND.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X223 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t8 CLK2.t10 GND.t50 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X224 a_2881_n4169# x1.t9 a_2731_n4169# GND.t145 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X225 CLK1.t67 x2_bar.t4 a_1170_n1349# GND.t91 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X226 CLK1.t68 x2_bar.t5 a_1170_n10570# GND.t92 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X227 a_3070_n4929# x1.t10 a_2920_n4929# GND.t146 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X228 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t2 x0.t4 a_1470_n9890# GND.t160 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X229 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t3 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 GND.t243 GND.t242 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X230 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t7 CLK1.t5 CLK1.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X231 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t2 x0.t5 a_3030_n1349# GND.t164 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X232 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar GND.t261 GND.t260 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X233 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar x0_bar.t4 CLK1.t114 GND.t141 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X234 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar x3.t8 CLK1.t198 GND.t239 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X235 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar Dis2.t9 GND.t277 GND.t148 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X236 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t8 CLK2.t112 CLK2.t111 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X237 CLK1.t17 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar CLK1.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X238 CLK3.t11 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT s1.t2 GND.t123 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X239 a_1470_n1349# x2.t6 CLK1.t168 GND.t165 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X240 GND.t20 s2_bar.t7 s2.t1 GND.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X241 CLK1.t71 x0.t6 a_2730_1471# GND.t93 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X242 CLK2.t42 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t9 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT CLK2.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X243 CLK2.t58 EESPFAL_s1_0/EESPFAL_INV4_0/A EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t2 GND.t168 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X244 GND.t305 Dis2.t10 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B GND.t196 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X245 GND.t307 Dis2.t11 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t4 GND.t306 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X246 CLK1.t77 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/B CLK1.t76 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X247 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_INV4_2/A_bar CLK1.t182 CLK1.t86 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X248 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar x2.t7 CLK1.t22 GND.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X249 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t1 Dis1.t22 GND.t199 GND.t198 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X250 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT CLK2.t29 CLK2.t28 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X251 s2_bar.t2 s2.t8 GND.t127 GND.t126 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X252 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t9 CLK1.t153 CLK1.t152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X253 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar x2_bar.t6 CLK1.t49 GND.t80 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X254 CLK2.t27 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar CLK2.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X255 CLK2.t8 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar GND.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X256 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B CLK1.t105 CLK1.t104 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X257 CLK1.t181 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar EESPFAL_s2_0/EESPFAL_INV4_2/A CLK1.t84 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X258 a_2920_n4929# x0.t7 a_2770_n4929# GND.t94 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X259 a_6800_n10570# EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT GND.t76 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X260 s1.t6 s1_bar.t7 CLK3.t35 CLK3.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X261 CLK2.t9 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t8 a_7070_1471# GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X262 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar GND.t240 GND.t64 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X263 CLK1.t109 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar CLK1.t108 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X264 CLK1.t37 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar EESPFAL_s1_0/EESPFAL_INV4_0/A CLK1.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X265 CLK1.t1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar CLK1.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X266 CLK2.t105 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar GND.t115 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X267 CLK2.t69 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar GND.t154 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X268 GND.t294 Dis2.t12 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t0 GND.t293 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X269 GND.t296 Dis2.t13 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT GND.t295 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X270 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar CLK1.t191 CLK1.t190 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X271 CLK1.t44 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar CLK1.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X272 CLK1.t39 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t9 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t4 CLK1.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X273 CLK1.t103 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar CLK1.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X274 CLK2.t34 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar CLK2.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X275 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar CLK1.t83 CLK1.t82 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X276 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t9 CLK2.t88 GND.t265 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X277 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar GND.t153 GND.t152 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X278 a_1170_1471# x3_bar.t9 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t1 GND.t259 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X279 CLK1.t165 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_1/B CLK1.t164 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X280 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t2 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 CLK2.t117 CLK2.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X281 CLK1.t128 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar CLK1.t127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X282 CLK1.t142 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t8 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t3 CLK1.t141 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X283 CLK2.t98 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar CLK2.t97 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X284 CLK2.t83 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t7 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT CLK2.t82 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X285 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar CLK2.t23 GND.t79 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X286 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar GND.t103 GND.t88 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X287 GND.t197 Dis1.t23 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B GND.t196 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X288 GND.t255 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t8 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t2 GND.t108 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X289 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t3 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t8 CLK1.t113 CLK1.t112 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X290 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t0 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 CLK2.t77 CLK2.t76 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X291 CLK1.t118 x1_bar.t9 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B GND.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X292 GND.t195 Dis1.t24 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B GND.t194 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X293 GND.t24 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B GND.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X294 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar CLK1.t73 CLK1.t72 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X295 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B CLK2.t102 CLK2.t101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X296 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t7 GND.t289 GND.t260 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X297 a_2770_n7070# x0_bar.t5 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A GND.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X298 GND.t193 Dis1.t25 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A GND.t192 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X299 GND.t1 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t0 GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X300 EESPFAL_s3_0/EESPFAL_INV4_0/A EESPFAL_s3_0/EESPFAL_INV4_0/A_bar CLK1.t159 CLK1.t158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X301 GND.t7 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t7 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X302 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t8 GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X303 CLK1.t50 x2_bar.t7 a_2881_n12710# GND.t81 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X304 CLK2.t75 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t1 CLK2.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X305 GND.t14 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t0 GND.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X306 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B GND.t263 GND.t101 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X307 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT CLK2.t32 CLK2.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X308 a_6800_n9890# EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT GND.t76 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X309 GND.t290 Dis2.t14 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT GND.t266 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X310 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 Dis2.t15 GND.t292 GND.t291 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X311 GND.t83 s0_bar.t6 s0.t2 GND.t82 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X312 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t8 GND.t301 GND.t128 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X313 a_2730_n2029# x3_bar.t10 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t4 GND.t113 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X314 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t9 CLK1.t48 CLK1.t47 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X315 CLK3.t6 s3.t8 s3_bar.t2 CLK3.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X316 a_1210_n7750# x2_bar.t8 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t4 GND.t72 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X317 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t0 x3.t9 a_1470_n2029# GND.t47 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X318 CLK3.t13 s2.t9 s2_bar.t3 CLK3.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X319 CLK2.t44 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t9 a_6800_n9890# GND.t140 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X320 CLK2.t64 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NOR_v3_0/B CLK2.t63 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X321 GND.t237 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t7 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 GND.t236 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X322 a_6859_n7750# EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT GND.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X323 a_3070_n7750# x3_bar.t11 CLK1.t94 GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X324 GND.t167 EESPFAL_s1_0/EESPFAL_INV4_0/A EESPFAL_s1_0/EESPFAL_INV4_0/A_bar GND.t166 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X325 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B x2_bar.t9 CLK1.t115 GND.t142 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X326 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar Dis1.t26 GND.t191 GND.t185 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X327 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar CLK2.t85 CLK2.t84 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X328 CLK1.t169 x3_bar.t12 a_1210_n7750# GND.t60 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X329 s3_bar.t1 s3.t9 GND.t286 GND.t285 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X330 a_3030_n10570# x2_bar.t10 CLK1.t90 GND.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X331 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t3 Dis2.t16 GND.t302 GND.t269 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X332 GND.t190 Dis1.t27 EESPFAL_s3_0/EESPFAL_INV4_0/A GND.t189 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X333 EESPFAL_s1_0/EESPFAL_INV4_0/A EESPFAL_s1_0/EESPFAL_INV4_0/A_bar GND.t68 GND.t67 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X334 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t5 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t9 CLK2.t45 GND.t144 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X335 CLK1.t148 x1_bar.t10 a_1170_n9890# GND.t92 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X336 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar CLK1.t87 CLK1.t86 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X337 CLK3.t31 s3_bar.t7 s3.t5 CLK3.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X338 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar GND.t98 GND.t95 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X339 CLK1.t70 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t9 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t3 CLK1.t69 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X340 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t5 x0.t8 a_3030_n9890# GND.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X341 a_1170_n1349# x0_bar.t6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t2 GND.t111 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X342 a_2731_n4169# x0_bar.t7 EESPFAL_s1_0/EESPFAL_INV4_0/A GND.t300 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X343 GND.t315 Dis3.t4 s0_bar.t4 GND.t295 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X344 CLK1.t174 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar CLK1.t173 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X345 a_1470_n9890# x1.t11 CLK1.t54 GND.t87 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X346 CLK1.t85 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A CLK1.t84 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X347 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar CLK2.t96 GND.t280 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X348 GND.t156 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t8 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 GND.t155 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X349 CLK1.t196 x0_bar.t8 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar GND.t310 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X350 CLK1.t162 x3.t10 a_2770_n7750# GND.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X351 a_3030_n1349# x2_bar.t11 CLK1.t91 GND.t61 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X352 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar x3.t11 CLK1.t163 GND.t253 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X353 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar CLK2.t73 CLK2.t72 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X354 s3.t3 Dis3.t5 GND.t317 GND.t316 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X355 s2.t4 Dis3.t6 GND.t43 GND.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X356 GND.t248 EESPFAL_s3_0/EESPFAL_INV4_0/A EESPFAL_s3_0/EESPFAL_INV4_0/A_bar GND.t247 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X357 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 Dis2.t17 GND.t304 GND.t303 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X358 a_2881_n12710# x0.t9 a_2731_n12710# GND.t112 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X359 CLK2.t71 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT CLK2.t70 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X360 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t1 Dis1.t28 GND.t188 GND.t187 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X361 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar CLK1.t122 CLK1.t121 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X362 CLK1.t107 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_INV4_2/A_bar CLK1.t98 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X363 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t8 CLK2.t47 CLK2.t46 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X364 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_INV4_2/A_bar GND.t279 GND.t278 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X365 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar Dis1.t29 GND.t186 GND.t185 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X366 GND.t184 Dis1.t30 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t5 GND.t183 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X367 s3.t4 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t8 CLK3.t40 GND.t312 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X368 a_6821_n4170# EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 s1_bar.t4 GND.t241 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X369 GND.t45 Dis3.t7 s1_bar.t0 GND.t44 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X370 GND.t182 Dis1.t31 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t4 GND.t181 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X371 CLK1.t189 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/B CLK1.t188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X372 CLK1.t81 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/B CLK1.t80 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X373 CLK1.t136 EESPFAL_s1_0/EESPFAL_INV4_0/A EESPFAL_s1_0/EESPFAL_INV4_0/A_bar CLK1.t135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X374 GND.t264 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t9 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t3 GND.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X375 CLK1.t192 x3.t12 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B GND.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X376 a_3030_1471# x0_bar.t9 CLK1.t197 GND.t311 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X377 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar x1_bar.t11 CLK1.t149 GND.t239 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X378 GND.t180 Dis1.t32 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B GND.t179 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X379 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar GND.t274 GND.t273 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X380 a_5050_791# EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s0_0/EESPFAL_NOR_v3_0/B GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X381 CLK1.t100 x0_bar.t10 a_1170_1471# GND.t122 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X382 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar Dis1.t33 GND.t178 GND.t177 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X383 CLK1.t120 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B CLK1.t119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X384 a_2770_n4929# x2.t8 EESPFAL_s2_0/EESPFAL_INV4_2/A GND.t131 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X385 a_7070_791# EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar s0_bar.t0 GND.t139 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X386 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t10 GND.t133 GND.t132 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X387 CLK2.t55 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t9 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT CLK2.t54 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X388 GND.t176 Dis1.t34 EESPFAL_s2_0/EESPFAL_INV4_2/A GND.t175 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X389 CLK3.t19 s0_bar.t7 s0.t3 CLK3.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X390 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar Dis1.t35 GND.t174 GND.t173 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X391 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 Dis2.t18 GND.t245 GND.t244 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X392 a_1470_1471# x0.t10 CLK1.t40 GND.t55 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X393 a_6971_n4170# EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar a_6821_n4170# GND.t272 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X394 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar CLK2.t11 GND.t66 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X395 CLK1.t23 x2.t9 a_2730_n1349# GND.t41 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X396 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t2 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 CLK2.t40 CLK2.t39 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X397 CLK2.t1 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t1 CLK2.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X398 a_1470_n10570# x2.t10 CLK1.t65 GND.t87 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X399 EESPFAL_s1_0/EESPFAL_INV4_0/A EESPFAL_s1_0/EESPFAL_INV4_0/A_bar CLK1.t35 CLK1.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X400 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT CLK2.t5 CLK2.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X401 CLK3.t29 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B s2.t6 GND.t282 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X402 a_6800_n2029# EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT GND.t3 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X403 GND.t246 Dis2.t19 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT GND.t118 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X404 GND.t267 Dis2.t20 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT GND.t266 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X405 s3.t6 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT CLK3.t39 GND.t308 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X406 GND.t169 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t9 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t3 GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X407 GND.t22 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar GND.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X408 CLK1.t195 x2.t11 a_2730_n10570# GND.t56 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X409 CLK2.t60 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t4 CLK2.t59 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X410 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar EESPFAL_s2_0/EESPFAL_INV4_2/A CLK1.t106 CLK1.t96 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X411 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t10 CLK2.t19 GND.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X412 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/B CLK1.t126 CLK1.t125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X413 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t9 CLK2.t57 CLK2.t56 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X414 s0.t5 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B CLK3.t28 GND.t265 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X415 GND.t120 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar GND.t57 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X416 GND.t268 Dis2.t21 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B GND.t116 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X417 a_6821_n12711# EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 s3_bar.t4 GND.t158 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X418 s2.t5 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t8 CLK3.t22 GND.t230 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X419 CLK2.t81 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t9 a_6800_n2029# GND.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
R0 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t5 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t6 819.4
R1 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t7 775.706
R2 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t5 514.133
R3 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t8 305.266
R4 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n1 166.734
R5 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n7 163.511
R6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n5 102.4
R7 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n6 88.255
R8 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t2 81.939
R9 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n2 76
R10 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n3 57.6
R11 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n0 51.537
R12 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t1 39.4
R13 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t0 39.4
R14 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t4 24
R15 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t3 24
R16 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n4 6.4
R17 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_s1_0/EESPFAL_INV4_0/OUT_bar 3.2
R18 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 819.4
R19 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 506.1
R20 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 313.3
R21 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 305.997
R22 EESPFAL_s1_0/EESPFAL_INV4_0/OUT EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 206.179
R23 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 187.539
R24 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 128.334
R25 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 115.2
R26 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 57.937
R27 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 57.6
R28 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 41.6
R29 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 39.4
R30 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 39.4
R31 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 24
R32 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 24
R33 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 8.764
R34 EESPFAL_s1_0/EESPFAL_INV4_0/OUT EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 4.65
R35 CLK2.n311 CLK2.n137 407.048
R36 CLK2.n357 CLK2.n117 407.048
R37 CLK2.n251 CLK2.n250 407.048
R38 CLK2.n292 CLK2.n291 407.048
R39 CLK2.n207 CLK2.n206 407.048
R40 CLK2.n240 CLK2.n239 407.048
R41 CLK2.n319 CLK2.n137 400
R42 CLK2.n320 CLK2.n319 400
R43 CLK2.n356 CLK2.n355 400
R44 CLK2.n357 CLK2.n356 400
R45 CLK2.n252 CLK2.n168 400
R46 CLK2.n252 CLK2.n251 400
R47 CLK2.n291 CLK2.n290 400
R48 CLK2.n290 CLK2.n148 400
R49 CLK2.n321 CLK2.n320 366.379
R50 CLK2.n355 CLK2.n118 366.379
R51 CLK2.n260 CLK2.n168 366.379
R52 CLK2.n282 CLK2.n148 366.379
R53 CLK2.n208 CLK2.n207 366.379
R54 CLK2.n239 CLK2.n238 366.379
R55 CLK2.n321 CLK2.n131 131.034
R56 CLK2.n330 CLK2.n131 131.034
R57 CLK2.n333 CLK2.n331 131.034
R58 CLK2.n342 CLK2.n341 131.034
R59 CLK2.n344 CLK2.n343 131.034
R60 CLK2.n343 CLK2.n118 131.034
R61 CLK2.n282 CLK2.n281 131.034
R62 CLK2.n281 CLK2.n280 131.034
R63 CLK2.n272 CLK2.n161 131.034
R64 CLK2.n270 CLK2.n162 131.034
R65 CLK2.n262 CLK2.n261 131.034
R66 CLK2.n261 CLK2.n260 131.034
R67 CLK2.n238 CLK2.n182 131.034
R68 CLK2.n229 CLK2.n182 131.034
R69 CLK2.n228 CLK2.n227 131.034
R70 CLK2.n219 CLK2.n218 131.034
R71 CLK2.n217 CLK2.n195 131.034
R72 CLK2.n208 CLK2.n195 131.034
R73 CLK2.t46 CLK2.n332 122.844
R74 CLK2.n332 CLK2.t109 122.844
R75 CLK2.t84 CLK2.n271 122.844
R76 CLK2.n271 CLK2.t17 122.844
R77 CLK2.n194 CLK2.t116 122.844
R78 CLK2.t67 CLK2.n194 122.844
R79 CLK2.n331 CLK2.t54 106.465
R80 CLK2.t107 CLK2.n342 106.465
R81 CLK2.n161 CLK2.t86 106.465
R82 CLK2.t15 CLK2.n162 106.465
R83 CLK2.t61 CLK2.n228 106.465
R84 CLK2.n218 CLK2.t13 106.465
R85 CLK2.n858 CLK2.n857 104.32
R86 CLK2.n312 CLK2.n138 96
R87 CLK2.n318 CLK2.n138 96
R88 CLK2.n318 CLK2.n136 96
R89 CLK2.n322 CLK2.n136 96
R90 CLK2.n322 CLK2.n132 96
R91 CLK2.n329 CLK2.n132 96
R92 CLK2.n329 CLK2.n130 96
R93 CLK2.n334 CLK2.n130 96
R94 CLK2.n334 CLK2.n125 96
R95 CLK2.n340 CLK2.n125 96
R96 CLK2.n340 CLK2.n124 96
R97 CLK2.n345 CLK2.n124 96
R98 CLK2.n345 CLK2.n119 96
R99 CLK2.n353 CLK2.n119 96
R100 CLK2.n354 CLK2.n353 96
R101 CLK2.n354 CLK2.n114 96
R102 CLK2.n358 CLK2.n114 96
R103 CLK2.n359 CLK2.n358 96
R104 CLK2.n293 CLK2.n147 96
R105 CLK2.n289 CLK2.n147 96
R106 CLK2.n289 CLK2.n149 96
R107 CLK2.n283 CLK2.n149 96
R108 CLK2.n283 CLK2.n153 96
R109 CLK2.n279 CLK2.n153 96
R110 CLK2.n279 CLK2.n154 96
R111 CLK2.n273 CLK2.n154 96
R112 CLK2.n273 CLK2.n160 96
R113 CLK2.n269 CLK2.n160 96
R114 CLK2.n269 CLK2.n163 96
R115 CLK2.n263 CLK2.n163 96
R116 CLK2.n263 CLK2.n167 96
R117 CLK2.n259 CLK2.n167 96
R118 CLK2.n259 CLK2.n169 96
R119 CLK2.n253 CLK2.n169 96
R120 CLK2.n253 CLK2.n175 96
R121 CLK2.n249 CLK2.n175 96
R122 CLK2.n241 CLK2.n181 96
R123 CLK2.n237 CLK2.n181 96
R124 CLK2.n237 CLK2.n183 96
R125 CLK2.n230 CLK2.n183 96
R126 CLK2.n230 CLK2.n187 96
R127 CLK2.n226 CLK2.n187 96
R128 CLK2.n226 CLK2.n188 96
R129 CLK2.n220 CLK2.n188 96
R130 CLK2.n220 CLK2.n193 96
R131 CLK2.n216 CLK2.n193 96
R132 CLK2.n216 CLK2.n196 96
R133 CLK2.n209 CLK2.n196 96
R134 CLK2.n209 CLK2.n200 96
R135 CLK2.n205 CLK2.n200 96
R136 CLK2.n361 CLK2.n117 88
R137 CLK2.n292 CLK2.n144 85.261
R138 CLK2.n250 CLK2.n176 85.261
R139 CLK2.n240 CLK2.n178 85.261
R140 CLK2.n206 CLK2.n201 85.261
R141 CLK2.n311 CLK2.n310 85.261
R142 CLK2.n745 CLK2.t93 44.338
R143 CLK2.n716 CLK2.t32 44.338
R144 CLK2.n596 CLK2.t60 44.338
R145 CLK2.n567 CLK2.t114 44.338
R146 CLK2.n156 CLK2.t87 44.338
R147 CLK2.n165 CLK2.t16 44.338
R148 CLK2.n427 CLK2.t83 44.338
R149 CLK2.n398 CLK2.t3 44.338
R150 CLK2.n915 CLK2.t64 44.338
R151 CLK2.n886 CLK2.t100 44.338
R152 CLK2.n836 CLK2.t5 44.337
R153 CLK2.n809 CLK2.t42 44.337
R154 CLK2.n642 CLK2.t50 44.337
R155 CLK2.n671 CLK2.t75 44.337
R156 CLK2.n520 CLK2.t102 44.337
R157 CLK2.n491 CLK2.t38 44.337
R158 CLK2.n348 CLK2.t108 44.337
R159 CLK2.n326 CLK2.t55 44.337
R160 CLK2.n213 CLK2.t14 44.337
R161 CLK2.n233 CLK2.t62 44.337
R162 CLK2.n56 CLK2.t29 44.337
R163 CLK2.n27 CLK2.t71 44.337
R164 CLK2.n859 CLK2.t66 39.4
R165 CLK2.n859 CLK2.t98 39.4
R166 CLK2.n83 CLK2.t112 39.4
R167 CLK2.n83 CLK2.t7 39.4
R168 CLK2.n89 CLK2.t95 39.4
R169 CLK2.n89 CLK2.t34 39.4
R170 CLK2.n623 CLK2.t77 39.4
R171 CLK2.n623 CLK2.t52 39.4
R172 CLK2.n548 CLK2.t40 39.4
R173 CLK2.n548 CLK2.t25 39.4
R174 CLK2.n101 CLK2.t36 39.4
R175 CLK2.n101 CLK2.t104 39.4
R176 CLK2.n105 CLK2.t57 39.4
R177 CLK2.n105 CLK2.t1 39.4
R178 CLK2.n127 CLK2.t47 39.4
R179 CLK2.n127 CLK2.t110 39.4
R180 CLK2.n157 CLK2.t85 39.4
R181 CLK2.n157 CLK2.t18 39.4
R182 CLK2.n190 CLK2.t117 39.4
R183 CLK2.n190 CLK2.t68 39.4
R184 CLK2.n0 CLK2.t73 39.4
R185 CLK2.n0 CLK2.t27 39.4
R186 CLK2.n2 CLK2.t9 30.775
R187 CLK2.n550 CLK2.t96 29.713
R188 CLK2.n625 CLK2.t11 29.712
R189 CLK2.n202 CLK2.t79 29.712
R190 CLK2.n244 CLK2.t78 29.712
R191 CLK2.n911 CLK2.t63 24.568
R192 CLK2.n887 CLK2.t99 24.568
R193 CLK2.n810 CLK2.t41 24.568
R194 CLK2.n832 CLK2.t4 24.568
R195 CLK2.n741 CLK2.t92 24.568
R196 CLK2.n717 CLK2.t31 24.568
R197 CLK2.n667 CLK2.t74 24.568
R198 CLK2.n643 CLK2.t49 24.568
R199 CLK2.n592 CLK2.t59 24.568
R200 CLK2.n568 CLK2.t113 24.568
R201 CLK2.n492 CLK2.t37 24.568
R202 CLK2.n516 CLK2.t101 24.568
R203 CLK2.n423 CLK2.t82 24.568
R204 CLK2.n399 CLK2.t2 24.568
R205 CLK2.t54 CLK2.n330 24.568
R206 CLK2.n344 CLK2.t107 24.568
R207 CLK2.n280 CLK2.t86 24.568
R208 CLK2.n262 CLK2.t15 24.568
R209 CLK2.n229 CLK2.t61 24.568
R210 CLK2.t13 CLK2.n217 24.568
R211 CLK2.n28 CLK2.t70 24.568
R212 CLK2.n52 CLK2.t28 24.568
R213 CLK2.n945 CLK2.t53 24
R214 CLK2.n80 CLK2.t45 24
R215 CLK2.n80 CLK2.t22 24
R216 CLK2.n774 CLK2.t81 24
R217 CLK2.n90 CLK2.t115 24
R218 CLK2.n90 CLK2.t8 24
R219 CLK2.n96 CLK2.t43 24
R220 CLK2.n100 CLK2.t23 24
R221 CLK2.n100 CLK2.t69 24
R222 CLK2.n462 CLK2.t30 24
R223 CLK2.n456 CLK2.t106 24
R224 CLK2.n116 CLK2.t90 24
R225 CLK2.n116 CLK2.t20 24
R226 CLK2.n299 CLK2.t91 24
R227 CLK2.n172 CLK2.t10 24
R228 CLK2.n172 CLK2.t21 24
R229 CLK2.n303 CLK2.t44 24
R230 CLK2.n372 CLK2.t12 24
R231 CLK2.n372 CLK2.t48 24
R232 CLK2.n93 CLK2.t58 24
R233 CLK2.n84 CLK2.t89 24
R234 CLK2.n860 CLK2.t19 24
R235 CLK2.n860 CLK2.t80 24
R236 CLK2.n949 CLK2.t88 24
R237 CLK2.n949 CLK2.t105 24
R238 CLK2.n731 CLK2.n728 12.8
R239 CLK2.n657 CLK2.n654 12.8
R240 CLK2.n582 CLK2.n579 12.8
R241 CLK2.n510 CLK2.n507 12.8
R242 CLK2.n413 CLK2.n410 12.8
R243 CLK2.n313 CLK2.n310 12.8
R244 CLK2.n313 CLK2.n139 12.8
R245 CLK2.n317 CLK2.n139 12.8
R246 CLK2.n317 CLK2.n135 12.8
R247 CLK2.n323 CLK2.n135 12.8
R248 CLK2.n323 CLK2.n133 12.8
R249 CLK2.n328 CLK2.n133 12.8
R250 CLK2.n328 CLK2.n129 12.8
R251 CLK2.n335 CLK2.n129 12.8
R252 CLK2.n335 CLK2.n126 12.8
R253 CLK2.n339 CLK2.n126 12.8
R254 CLK2.n339 CLK2.n123 12.8
R255 CLK2.n346 CLK2.n123 12.8
R256 CLK2.n346 CLK2.n120 12.8
R257 CLK2.n352 CLK2.n120 12.8
R258 CLK2.n365 CLK2.n115 12.8
R259 CLK2.n360 CLK2.n115 12.8
R260 CLK2.n298 CLK2.n143 12.8
R261 CLK2.n294 CLK2.n144 12.8
R262 CLK2.n294 CLK2.n146 12.8
R263 CLK2.n288 CLK2.n146 12.8
R264 CLK2.n288 CLK2.n150 12.8
R265 CLK2.n284 CLK2.n150 12.8
R266 CLK2.n284 CLK2.n152 12.8
R267 CLK2.n278 CLK2.n152 12.8
R268 CLK2.n278 CLK2.n155 12.8
R269 CLK2.n274 CLK2.n155 12.8
R270 CLK2.n274 CLK2.n159 12.8
R271 CLK2.n268 CLK2.n159 12.8
R272 CLK2.n268 CLK2.n164 12.8
R273 CLK2.n264 CLK2.n164 12.8
R274 CLK2.n264 CLK2.n166 12.8
R275 CLK2.n258 CLK2.n166 12.8
R276 CLK2.n258 CLK2.n170 12.8
R277 CLK2.n254 CLK2.n170 12.8
R278 CLK2.n254 CLK2.n174 12.8
R279 CLK2.n248 CLK2.n174 12.8
R280 CLK2.n248 CLK2.n176 12.8
R281 CLK2.n242 CLK2.n178 12.8
R282 CLK2.n242 CLK2.n180 12.8
R283 CLK2.n236 CLK2.n180 12.8
R284 CLK2.n236 CLK2.n184 12.8
R285 CLK2.n231 CLK2.n184 12.8
R286 CLK2.n231 CLK2.n186 12.8
R287 CLK2.n225 CLK2.n186 12.8
R288 CLK2.n225 CLK2.n189 12.8
R289 CLK2.n221 CLK2.n189 12.8
R290 CLK2.n221 CLK2.n192 12.8
R291 CLK2.n215 CLK2.n192 12.8
R292 CLK2.n215 CLK2.n197 12.8
R293 CLK2.n210 CLK2.n197 12.8
R294 CLK2.n210 CLK2.n199 12.8
R295 CLK2.n204 CLK2.n199 12.8
R296 CLK2.n204 CLK2.n201 12.8
R297 CLK2.n305 CLK2.n304 12.8
R298 CLK2.n826 CLK2.n823 12.8
R299 CLK2.n901 CLK2.n898 12.8
R300 CLK2.n46 CLK2.n43 12.8
R301 CLK2.n366 CLK2.n365 11.84
R302 CLK2.n352 CLK2.n121 11.04
R303 CLK2.n350 CLK2.n121 9.3
R304 CLK2.n113 CLK2.n112 9.3
R305 CLK2.n768 CLK2.n767 8.855
R306 CLK2.n686 CLK2.n685 8.855
R307 CLK2.n612 CLK2.n611 8.855
R308 CLK2.n469 CLK2.n468 8.855
R309 CLK2.n108 CLK2.n107 8.855
R310 CLK2.n358 CLK2.n115 8.855
R311 CLK2.n358 CLK2.n357 8.855
R312 CLK2.n313 CLK2.n312 8.855
R313 CLK2.n299 CLK2.n298 8.855
R314 CLK2.n294 CLK2.n293 8.855
R315 CLK2.n242 CLK2.n241 8.855
R316 CLK2.n181 CLK2.n180 8.855
R317 CLK2.n239 CLK2.n181 8.855
R318 CLK2.n237 CLK2.n236 8.855
R319 CLK2.n238 CLK2.n237 8.855
R320 CLK2.n184 CLK2.n183 8.855
R321 CLK2.n183 CLK2.n182 8.855
R322 CLK2.n231 CLK2.n230 8.855
R323 CLK2.n230 CLK2.n229 8.855
R324 CLK2.n187 CLK2.n186 8.855
R325 CLK2.n228 CLK2.n187 8.855
R326 CLK2.n226 CLK2.n225 8.855
R327 CLK2.n227 CLK2.n226 8.855
R328 CLK2.n189 CLK2.n188 8.855
R329 CLK2.n194 CLK2.n188 8.855
R330 CLK2.n221 CLK2.n220 8.855
R331 CLK2.n220 CLK2.n219 8.855
R332 CLK2.n193 CLK2.n192 8.855
R333 CLK2.n218 CLK2.n193 8.855
R334 CLK2.n216 CLK2.n215 8.855
R335 CLK2.n217 CLK2.n216 8.855
R336 CLK2.n197 CLK2.n196 8.855
R337 CLK2.n196 CLK2.n195 8.855
R338 CLK2.n210 CLK2.n209 8.855
R339 CLK2.n209 CLK2.n208 8.855
R340 CLK2.n200 CLK2.n199 8.855
R341 CLK2.n207 CLK2.n200 8.855
R342 CLK2.n205 CLK2.n204 8.855
R343 CLK2.n147 CLK2.n146 8.855
R344 CLK2.n291 CLK2.n147 8.855
R345 CLK2.n289 CLK2.n288 8.855
R346 CLK2.n290 CLK2.n289 8.855
R347 CLK2.n150 CLK2.n149 8.855
R348 CLK2.n149 CLK2.n148 8.855
R349 CLK2.n284 CLK2.n283 8.855
R350 CLK2.n283 CLK2.n282 8.855
R351 CLK2.n153 CLK2.n152 8.855
R352 CLK2.n281 CLK2.n153 8.855
R353 CLK2.n279 CLK2.n278 8.855
R354 CLK2.n280 CLK2.n279 8.855
R355 CLK2.n155 CLK2.n154 8.855
R356 CLK2.n161 CLK2.n154 8.855
R357 CLK2.n274 CLK2.n273 8.855
R358 CLK2.n273 CLK2.n272 8.855
R359 CLK2.n160 CLK2.n159 8.855
R360 CLK2.n271 CLK2.n160 8.855
R361 CLK2.n269 CLK2.n268 8.855
R362 CLK2.n270 CLK2.n269 8.855
R363 CLK2.n164 CLK2.n163 8.855
R364 CLK2.n163 CLK2.n162 8.855
R365 CLK2.n264 CLK2.n263 8.855
R366 CLK2.n263 CLK2.n262 8.855
R367 CLK2.n167 CLK2.n166 8.855
R368 CLK2.n261 CLK2.n167 8.855
R369 CLK2.n259 CLK2.n258 8.855
R370 CLK2.n260 CLK2.n259 8.855
R371 CLK2.n170 CLK2.n169 8.855
R372 CLK2.n169 CLK2.n168 8.855
R373 CLK2.n254 CLK2.n253 8.855
R374 CLK2.n253 CLK2.n252 8.855
R375 CLK2.n175 CLK2.n174 8.855
R376 CLK2.n251 CLK2.n175 8.855
R377 CLK2.n249 CLK2.n248 8.855
R378 CLK2.n304 CLK2.n303 8.855
R379 CLK2.n360 CLK2.n359 8.855
R380 CLK2.n139 CLK2.n138 8.855
R381 CLK2.n138 CLK2.n137 8.855
R382 CLK2.n318 CLK2.n317 8.855
R383 CLK2.n319 CLK2.n318 8.855
R384 CLK2.n136 CLK2.n135 8.855
R385 CLK2.n320 CLK2.n136 8.855
R386 CLK2.n323 CLK2.n322 8.855
R387 CLK2.n322 CLK2.n321 8.855
R388 CLK2.n133 CLK2.n132 8.855
R389 CLK2.n132 CLK2.n131 8.855
R390 CLK2.n329 CLK2.n328 8.855
R391 CLK2.n330 CLK2.n329 8.855
R392 CLK2.n130 CLK2.n129 8.855
R393 CLK2.n331 CLK2.n130 8.855
R394 CLK2.n335 CLK2.n334 8.855
R395 CLK2.n334 CLK2.n333 8.855
R396 CLK2.n126 CLK2.n125 8.855
R397 CLK2.n332 CLK2.n125 8.855
R398 CLK2.n340 CLK2.n339 8.855
R399 CLK2.n341 CLK2.n340 8.855
R400 CLK2.n124 CLK2.n123 8.855
R401 CLK2.n342 CLK2.n124 8.855
R402 CLK2.n346 CLK2.n345 8.855
R403 CLK2.n345 CLK2.n344 8.855
R404 CLK2.n120 CLK2.n119 8.855
R405 CLK2.n343 CLK2.n119 8.855
R406 CLK2.n353 CLK2.n352 8.855
R407 CLK2.n353 CLK2.n118 8.855
R408 CLK2.n354 CLK2.n113 8.855
R409 CLK2.n355 CLK2.n354 8.855
R410 CLK2.n365 CLK2.n114 8.855
R411 CLK2.n356 CLK2.n114 8.855
R412 CLK2.n450 CLK2.n449 8.855
R413 CLK2.n446 CLK2.n445 8.855
R414 CLK2.n445 CLK2.n444 8.855
R415 CLK2.n442 CLK2.n441 8.855
R416 CLK2.n441 CLK2.n440 8.855
R417 CLK2.n438 CLK2.n437 8.855
R418 CLK2.n437 CLK2.n436 8.855
R419 CLK2.n434 CLK2.n433 8.855
R420 CLK2.n433 CLK2.n432 8.855
R421 CLK2.n430 CLK2.n429 8.855
R422 CLK2.n429 CLK2.n428 8.855
R423 CLK2.n425 CLK2.n424 8.855
R424 CLK2.n424 CLK2.n423 8.855
R425 CLK2.n421 CLK2.n420 8.855
R426 CLK2.n420 CLK2.n419 8.855
R427 CLK2.n417 CLK2.n416 8.855
R428 CLK2.n416 CLK2.n415 8.855
R429 CLK2.n413 CLK2.n412 8.855
R430 CLK2.n412 CLK2.n411 8.855
R431 CLK2.n410 CLK2.n409 8.855
R432 CLK2.n409 CLK2.n408 8.855
R433 CLK2.n405 CLK2.n404 8.855
R434 CLK2.n404 CLK2.n403 8.855
R435 CLK2.n401 CLK2.n400 8.855
R436 CLK2.n400 CLK2.n399 8.855
R437 CLK2.n396 CLK2.n395 8.855
R438 CLK2.n395 CLK2.n394 8.855
R439 CLK2.n392 CLK2.n391 8.855
R440 CLK2.n391 CLK2.n390 8.855
R441 CLK2.n107 CLK2.n106 8.855
R442 CLK2.n385 CLK2.n384 8.855
R443 CLK2.n384 CLK2.n383 8.855
R444 CLK2.n379 CLK2.n378 8.855
R445 CLK2.n378 CLK2.n377 8.855
R446 CLK2.n375 CLK2.n374 8.855
R447 CLK2.n473 CLK2.n472 8.855
R448 CLK2.n472 CLK2.n471 8.855
R449 CLK2.n477 CLK2.n476 8.855
R450 CLK2.n476 CLK2.n475 8.855
R451 CLK2.n481 CLK2.n480 8.855
R452 CLK2.n480 CLK2.n479 8.855
R453 CLK2.n485 CLK2.n484 8.855
R454 CLK2.n484 CLK2.n483 8.855
R455 CLK2.n489 CLK2.n488 8.855
R456 CLK2.n488 CLK2.n487 8.855
R457 CLK2.n494 CLK2.n493 8.855
R458 CLK2.n493 CLK2.n492 8.855
R459 CLK2.n498 CLK2.n497 8.855
R460 CLK2.n497 CLK2.n496 8.855
R461 CLK2.n502 CLK2.n501 8.855
R462 CLK2.n501 CLK2.n500 8.855
R463 CLK2.n507 CLK2.n506 8.855
R464 CLK2.n506 CLK2.n505 8.855
R465 CLK2.n510 CLK2.n509 8.855
R466 CLK2.n509 CLK2.n508 8.855
R467 CLK2.n514 CLK2.n513 8.855
R468 CLK2.n513 CLK2.n512 8.855
R469 CLK2.n518 CLK2.n517 8.855
R470 CLK2.n517 CLK2.n516 8.855
R471 CLK2.n523 CLK2.n522 8.855
R472 CLK2.n522 CLK2.n521 8.855
R473 CLK2.n527 CLK2.n526 8.855
R474 CLK2.n526 CLK2.n525 8.855
R475 CLK2.n531 CLK2.n530 8.855
R476 CLK2.n530 CLK2.n529 8.855
R477 CLK2.n535 CLK2.n534 8.855
R478 CLK2.n534 CLK2.n533 8.855
R479 CLK2.n540 CLK2.n539 8.855
R480 CLK2.n539 CLK2.n538 8.855
R481 CLK2.n544 CLK2.n543 8.855
R482 CLK2.n607 CLK2.n606 8.855
R483 CLK2.n606 CLK2.n605 8.855
R484 CLK2.n603 CLK2.n602 8.855
R485 CLK2.n602 CLK2.n601 8.855
R486 CLK2.n599 CLK2.n598 8.855
R487 CLK2.n598 CLK2.n597 8.855
R488 CLK2.n594 CLK2.n593 8.855
R489 CLK2.n593 CLK2.n592 8.855
R490 CLK2.n590 CLK2.n589 8.855
R491 CLK2.n589 CLK2.n588 8.855
R492 CLK2.n586 CLK2.n585 8.855
R493 CLK2.n585 CLK2.n584 8.855
R494 CLK2.n582 CLK2.n581 8.855
R495 CLK2.n581 CLK2.n580 8.855
R496 CLK2.n579 CLK2.n578 8.855
R497 CLK2.n578 CLK2.n577 8.855
R498 CLK2.n574 CLK2.n573 8.855
R499 CLK2.n573 CLK2.n572 8.855
R500 CLK2.n570 CLK2.n569 8.855
R501 CLK2.n569 CLK2.n568 8.855
R502 CLK2.n565 CLK2.n564 8.855
R503 CLK2.n564 CLK2.n563 8.855
R504 CLK2.n561 CLK2.n560 8.855
R505 CLK2.n560 CLK2.n559 8.855
R506 CLK2.n557 CLK2.n556 8.855
R507 CLK2.n556 CLK2.n555 8.855
R508 CLK2.n553 CLK2.n552 8.855
R509 CLK2.n682 CLK2.n681 8.855
R510 CLK2.n681 CLK2.n680 8.855
R511 CLK2.n678 CLK2.n677 8.855
R512 CLK2.n677 CLK2.n676 8.855
R513 CLK2.n674 CLK2.n673 8.855
R514 CLK2.n673 CLK2.n672 8.855
R515 CLK2.n669 CLK2.n668 8.855
R516 CLK2.n668 CLK2.n667 8.855
R517 CLK2.n665 CLK2.n664 8.855
R518 CLK2.n664 CLK2.n663 8.855
R519 CLK2.n661 CLK2.n660 8.855
R520 CLK2.n660 CLK2.n659 8.855
R521 CLK2.n657 CLK2.n656 8.855
R522 CLK2.n656 CLK2.n655 8.855
R523 CLK2.n654 CLK2.n653 8.855
R524 CLK2.n653 CLK2.n652 8.855
R525 CLK2.n649 CLK2.n648 8.855
R526 CLK2.n648 CLK2.n647 8.855
R527 CLK2.n645 CLK2.n644 8.855
R528 CLK2.n644 CLK2.n643 8.855
R529 CLK2.n640 CLK2.n639 8.855
R530 CLK2.n639 CLK2.n638 8.855
R531 CLK2.n636 CLK2.n635 8.855
R532 CLK2.n635 CLK2.n634 8.855
R533 CLK2.n632 CLK2.n631 8.855
R534 CLK2.n631 CLK2.n630 8.855
R535 CLK2.n628 CLK2.n627 8.855
R536 CLK2.n764 CLK2.n763 8.855
R537 CLK2.n763 CLK2.n762 8.855
R538 CLK2.n760 CLK2.n759 8.855
R539 CLK2.n759 CLK2.n758 8.855
R540 CLK2.n756 CLK2.n755 8.855
R541 CLK2.n755 CLK2.n754 8.855
R542 CLK2.n752 CLK2.n751 8.855
R543 CLK2.n751 CLK2.n750 8.855
R544 CLK2.n748 CLK2.n747 8.855
R545 CLK2.n747 CLK2.n746 8.855
R546 CLK2.n743 CLK2.n742 8.855
R547 CLK2.n742 CLK2.n741 8.855
R548 CLK2.n739 CLK2.n738 8.855
R549 CLK2.n738 CLK2.n737 8.855
R550 CLK2.n735 CLK2.n734 8.855
R551 CLK2.n734 CLK2.n733 8.855
R552 CLK2.n731 CLK2.n730 8.855
R553 CLK2.n730 CLK2.n729 8.855
R554 CLK2.n728 CLK2.n727 8.855
R555 CLK2.n727 CLK2.n726 8.855
R556 CLK2.n723 CLK2.n722 8.855
R557 CLK2.n722 CLK2.n721 8.855
R558 CLK2.n719 CLK2.n718 8.855
R559 CLK2.n718 CLK2.n717 8.855
R560 CLK2.n714 CLK2.n713 8.855
R561 CLK2.n713 CLK2.n712 8.855
R562 CLK2.n710 CLK2.n709 8.855
R563 CLK2.n709 CLK2.n708 8.855
R564 CLK2.n706 CLK2.n705 8.855
R565 CLK2.n705 CLK2.n704 8.855
R566 CLK2.n702 CLK2.n701 8.855
R567 CLK2.n701 CLK2.n700 8.855
R568 CLK2.n697 CLK2.n696 8.855
R569 CLK2.n696 CLK2.n695 8.855
R570 CLK2.n693 CLK2.n692 8.855
R571 CLK2.n787 CLK2.n786 8.855
R572 CLK2.n791 CLK2.n790 8.855
R573 CLK2.n790 CLK2.n789 8.855
R574 CLK2.n795 CLK2.n794 8.855
R575 CLK2.n794 CLK2.n793 8.855
R576 CLK2.n799 CLK2.n798 8.855
R577 CLK2.n798 CLK2.n797 8.855
R578 CLK2.n803 CLK2.n802 8.855
R579 CLK2.n802 CLK2.n801 8.855
R580 CLK2.n807 CLK2.n806 8.855
R581 CLK2.n806 CLK2.n805 8.855
R582 CLK2.n812 CLK2.n811 8.855
R583 CLK2.n811 CLK2.n810 8.855
R584 CLK2.n816 CLK2.n815 8.855
R585 CLK2.n815 CLK2.n814 8.855
R586 CLK2.n820 CLK2.n819 8.855
R587 CLK2.n819 CLK2.n818 8.855
R588 CLK2.n823 CLK2.n82 8.855
R589 CLK2.n82 CLK2.n81 8.855
R590 CLK2.n826 CLK2.n825 8.855
R591 CLK2.n825 CLK2.n824 8.855
R592 CLK2.n830 CLK2.n829 8.855
R593 CLK2.n829 CLK2.n828 8.855
R594 CLK2.n834 CLK2.n833 8.855
R595 CLK2.n833 CLK2.n832 8.855
R596 CLK2.n839 CLK2.n838 8.855
R597 CLK2.n838 CLK2.n837 8.855
R598 CLK2.n843 CLK2.n842 8.855
R599 CLK2.n842 CLK2.n841 8.855
R600 CLK2.n847 CLK2.n846 8.855
R601 CLK2.n846 CLK2.n845 8.855
R602 CLK2.n851 CLK2.n850 8.855
R603 CLK2.n850 CLK2.n849 8.855
R604 CLK2.n77 CLK2.n76 8.855
R605 CLK2.n76 CLK2.n75 8.855
R606 CLK2.n856 CLK2.n79 8.855
R607 CLK2.n938 CLK2.n937 8.855
R608 CLK2.n934 CLK2.n933 8.855
R609 CLK2.n933 CLK2.n932 8.855
R610 CLK2.n930 CLK2.n929 8.855
R611 CLK2.n929 CLK2.n928 8.855
R612 CLK2.n926 CLK2.n925 8.855
R613 CLK2.n925 CLK2.n924 8.855
R614 CLK2.n922 CLK2.n921 8.855
R615 CLK2.n921 CLK2.n920 8.855
R616 CLK2.n918 CLK2.n917 8.855
R617 CLK2.n917 CLK2.n916 8.855
R618 CLK2.n913 CLK2.n912 8.855
R619 CLK2.n912 CLK2.n911 8.855
R620 CLK2.n909 CLK2.n908 8.855
R621 CLK2.n908 CLK2.n907 8.855
R622 CLK2.n905 CLK2.n904 8.855
R623 CLK2.n904 CLK2.n903 8.855
R624 CLK2.n901 CLK2.n900 8.855
R625 CLK2.n900 CLK2.n899 8.855
R626 CLK2.n898 CLK2.n897 8.855
R627 CLK2.n897 CLK2.n896 8.855
R628 CLK2.n893 CLK2.n892 8.855
R629 CLK2.n892 CLK2.n891 8.855
R630 CLK2.n889 CLK2.n888 8.855
R631 CLK2.n888 CLK2.n887 8.855
R632 CLK2.n884 CLK2.n883 8.855
R633 CLK2.n883 CLK2.n882 8.855
R634 CLK2.n880 CLK2.n879 8.855
R635 CLK2.n879 CLK2.n878 8.855
R636 CLK2.n876 CLK2.n875 8.855
R637 CLK2.n875 CLK2.n874 8.855
R638 CLK2.n872 CLK2.n871 8.855
R639 CLK2.n871 CLK2.n870 8.855
R640 CLK2.n867 CLK2.n866 8.855
R641 CLK2.n866 CLK2.n865 8.855
R642 CLK2.n863 CLK2.n862 8.855
R643 CLK2.n5 CLK2.n4 8.855
R644 CLK2.n9 CLK2.n8 8.855
R645 CLK2.n8 CLK2.n7 8.855
R646 CLK2.n13 CLK2.n12 8.855
R647 CLK2.n12 CLK2.n11 8.855
R648 CLK2.n17 CLK2.n16 8.855
R649 CLK2.n16 CLK2.n15 8.855
R650 CLK2.n21 CLK2.n20 8.855
R651 CLK2.n20 CLK2.n19 8.855
R652 CLK2.n25 CLK2.n24 8.855
R653 CLK2.n24 CLK2.n23 8.855
R654 CLK2.n30 CLK2.n29 8.855
R655 CLK2.n29 CLK2.n28 8.855
R656 CLK2.n34 CLK2.n33 8.855
R657 CLK2.n33 CLK2.n32 8.855
R658 CLK2.n38 CLK2.n37 8.855
R659 CLK2.n37 CLK2.n36 8.855
R660 CLK2.n43 CLK2.n42 8.855
R661 CLK2.n42 CLK2.n41 8.855
R662 CLK2.n46 CLK2.n45 8.855
R663 CLK2.n45 CLK2.n44 8.855
R664 CLK2.n50 CLK2.n49 8.855
R665 CLK2.n49 CLK2.n48 8.855
R666 CLK2.n54 CLK2.n53 8.855
R667 CLK2.n53 CLK2.n52 8.855
R668 CLK2.n59 CLK2.n58 8.855
R669 CLK2.n58 CLK2.n57 8.855
R670 CLK2.n63 CLK2.n62 8.855
R671 CLK2.n62 CLK2.n61 8.855
R672 CLK2.n67 CLK2.n66 8.855
R673 CLK2.n66 CLK2.n65 8.855
R674 CLK2.n71 CLK2.n70 8.855
R675 CLK2.n70 CLK2.n69 8.855
R676 CLK2.n962 CLK2.n960 8.855
R677 CLK2.n960 CLK2.n959 8.855
R678 CLK2.n956 CLK2.n955 8.855
R679 CLK2.n464 CLK2.n463 8.365
R680 CLK2.n307 CLK2.n141 8.365
R681 CLK2.n622 CLK2.n94 8.365
R682 CLK2.n780 CLK2.n85 8.365
R683 CLK2.n947 CLK2.n946 8.365
R684 CLK2.n903 CLK2.t65 8.189
R685 CLK2.n896 CLK2.t97 8.189
R686 CLK2.n818 CLK2.t111 8.189
R687 CLK2.n824 CLK2.t6 8.189
R688 CLK2.n733 CLK2.t94 8.189
R689 CLK2.n726 CLK2.t33 8.189
R690 CLK2.n659 CLK2.t76 8.189
R691 CLK2.n652 CLK2.t51 8.189
R692 CLK2.n584 CLK2.t39 8.189
R693 CLK2.n577 CLK2.t24 8.189
R694 CLK2.n500 CLK2.t35 8.189
R695 CLK2.n508 CLK2.t103 8.189
R696 CLK2.n415 CLK2.t56 8.189
R697 CLK2.n408 CLK2.t0 8.189
R698 CLK2.n333 CLK2.t46 8.189
R699 CLK2.n341 CLK2.t109 8.189
R700 CLK2.n272 CLK2.t84 8.189
R701 CLK2.t17 CLK2.n270 8.189
R702 CLK2.n227 CLK2.t116 8.189
R703 CLK2.n219 CLK2.t67 8.189
R704 CLK2.n36 CLK2.t72 8.189
R705 CLK2.n44 CLK2.t26 8.189
R706 CLK2.n948 CLK2.n947 7.422
R707 CLK2.n853 CLK2.n80 6.776
R708 CLK2.n699 CLK2.n90 6.776
R709 CLK2.n537 CLK2.n100 6.776
R710 CLK2.n363 CLK2.n116 6.776
R711 CLK2.n173 CLK2.n172 6.776
R712 CLK2.n381 CLK2.n372 6.776
R713 CLK2.n869 CLK2.n860 6.776
R714 CLK2.n618 CLK2.n97 6.755
R715 CLK2.n301 CLK2.n300 6.754
R716 CLK2.n776 CLK2.n775 6.754
R717 CLK2.n458 CLK2.n457 6.754
R718 CLK2.n857 CLK2.n856 6.72
R719 CLK2.n857 CLK2.n77 6.08
R720 CLK2.n902 CLK2.n859 4.938
R721 CLK2.n822 CLK2.n83 4.938
R722 CLK2.n732 CLK2.n89 4.938
R723 CLK2.n658 CLK2.n623 4.938
R724 CLK2.n583 CLK2.n548 4.938
R725 CLK2.n504 CLK2.n101 4.938
R726 CLK2.n414 CLK2.n105 4.938
R727 CLK2.n337 CLK2.n127 4.938
R728 CLK2.n158 CLK2.n157 4.938
R729 CLK2.n223 CLK2.n190 4.938
R730 CLK2.n40 CLK2.n0 4.938
R731 CLK2.n296 CLK2.n144 4.675
R732 CLK2.n452 CLK2.n104 4.675
R733 CLK2.n466 CLK2.n465 4.675
R734 CLK2.n770 CLK2.n88 4.675
R735 CLK2.n940 CLK2.n858 4.675
R736 CLK2.n2 CLK2.n1 4.675
R737 CLK2.n202 CLK2.n201 4.662
R738 CLK2.n614 CLK2.n99 4.662
R739 CLK2.n550 CLK2.n549 4.662
R740 CLK2.n625 CLK2.n624 4.662
R741 CLK2.n243 CLK2.n242 4.65
R742 CLK2.n180 CLK2.n179 4.65
R743 CLK2.n236 CLK2.n235 4.65
R744 CLK2.n234 CLK2.n184 4.65
R745 CLK2.n232 CLK2.n231 4.65
R746 CLK2.n186 CLK2.n185 4.65
R747 CLK2.n225 CLK2.n224 4.65
R748 CLK2.n223 CLK2.n189 4.65
R749 CLK2.n222 CLK2.n221 4.65
R750 CLK2.n192 CLK2.n191 4.65
R751 CLK2.n215 CLK2.n214 4.65
R752 CLK2.n212 CLK2.n197 4.65
R753 CLK2.n211 CLK2.n210 4.65
R754 CLK2.n199 CLK2.n198 4.65
R755 CLK2.n204 CLK2.n203 4.65
R756 CLK2.n245 CLK2.n178 4.65
R757 CLK2.n246 CLK2.n176 4.65
R758 CLK2.n295 CLK2.n294 4.65
R759 CLK2.n146 CLK2.n145 4.65
R760 CLK2.n288 CLK2.n287 4.65
R761 CLK2.n286 CLK2.n150 4.65
R762 CLK2.n285 CLK2.n284 4.65
R763 CLK2.n152 CLK2.n151 4.65
R764 CLK2.n278 CLK2.n277 4.65
R765 CLK2.n276 CLK2.n155 4.65
R766 CLK2.n275 CLK2.n274 4.65
R767 CLK2.n159 CLK2.n158 4.65
R768 CLK2.n268 CLK2.n267 4.65
R769 CLK2.n266 CLK2.n164 4.65
R770 CLK2.n265 CLK2.n264 4.65
R771 CLK2.n171 CLK2.n166 4.65
R772 CLK2.n258 CLK2.n257 4.65
R773 CLK2.n256 CLK2.n170 4.65
R774 CLK2.n255 CLK2.n254 4.65
R775 CLK2.n177 CLK2.n174 4.65
R776 CLK2.n248 CLK2.n247 4.65
R777 CLK2.n143 CLK2.n142 4.65
R778 CLK2.n298 CLK2.n297 4.65
R779 CLK2.n306 CLK2.n305 4.65
R780 CLK2.n314 CLK2.n313 4.65
R781 CLK2.n362 CLK2.n115 4.65
R782 CLK2.n315 CLK2.n139 4.65
R783 CLK2.n317 CLK2.n316 4.65
R784 CLK2.n135 CLK2.n134 4.65
R785 CLK2.n324 CLK2.n323 4.65
R786 CLK2.n325 CLK2.n133 4.65
R787 CLK2.n328 CLK2.n327 4.65
R788 CLK2.n129 CLK2.n128 4.65
R789 CLK2.n336 CLK2.n335 4.65
R790 CLK2.n337 CLK2.n126 4.65
R791 CLK2.n339 CLK2.n338 4.65
R792 CLK2.n123 CLK2.n122 4.65
R793 CLK2.n347 CLK2.n346 4.65
R794 CLK2.n349 CLK2.n120 4.65
R795 CLK2.n352 CLK2.n351 4.65
R796 CLK2.n365 CLK2.n364 4.65
R797 CLK2.n389 CLK2.n108 4.65
R798 CLK2.n451 CLK2.n450 4.65
R799 CLK2.n447 CLK2.n446 4.65
R800 CLK2.n443 CLK2.n442 4.65
R801 CLK2.n439 CLK2.n438 4.65
R802 CLK2.n435 CLK2.n434 4.65
R803 CLK2.n431 CLK2.n430 4.65
R804 CLK2.n426 CLK2.n425 4.65
R805 CLK2.n422 CLK2.n421 4.65
R806 CLK2.n418 CLK2.n417 4.65
R807 CLK2.n414 CLK2.n413 4.65
R808 CLK2.n410 CLK2.n407 4.65
R809 CLK2.n406 CLK2.n405 4.65
R810 CLK2.n402 CLK2.n401 4.65
R811 CLK2.n397 CLK2.n396 4.65
R812 CLK2.n393 CLK2.n392 4.65
R813 CLK2.n380 CLK2.n379 4.65
R814 CLK2.n455 CLK2.n103 4.65
R815 CLK2.n454 CLK2.n453 4.65
R816 CLK2.n461 CLK2.n460 4.65
R817 CLK2.n547 CLK2.n546 4.65
R818 CLK2.n470 CLK2.n469 4.65
R819 CLK2.n474 CLK2.n473 4.65
R820 CLK2.n478 CLK2.n477 4.65
R821 CLK2.n482 CLK2.n481 4.65
R822 CLK2.n486 CLK2.n485 4.65
R823 CLK2.n490 CLK2.n489 4.65
R824 CLK2.n495 CLK2.n494 4.65
R825 CLK2.n499 CLK2.n498 4.65
R826 CLK2.n503 CLK2.n502 4.65
R827 CLK2.n507 CLK2.n504 4.65
R828 CLK2.n511 CLK2.n510 4.65
R829 CLK2.n515 CLK2.n514 4.65
R830 CLK2.n519 CLK2.n518 4.65
R831 CLK2.n524 CLK2.n523 4.65
R832 CLK2.n528 CLK2.n527 4.65
R833 CLK2.n532 CLK2.n531 4.65
R834 CLK2.n536 CLK2.n535 4.65
R835 CLK2.n541 CLK2.n540 4.65
R836 CLK2.n545 CLK2.n544 4.65
R837 CLK2.n613 CLK2.n612 4.65
R838 CLK2.n608 CLK2.n607 4.65
R839 CLK2.n604 CLK2.n603 4.65
R840 CLK2.n600 CLK2.n599 4.65
R841 CLK2.n595 CLK2.n594 4.65
R842 CLK2.n591 CLK2.n590 4.65
R843 CLK2.n587 CLK2.n586 4.65
R844 CLK2.n583 CLK2.n582 4.65
R845 CLK2.n579 CLK2.n576 4.65
R846 CLK2.n575 CLK2.n574 4.65
R847 CLK2.n571 CLK2.n570 4.65
R848 CLK2.n566 CLK2.n565 4.65
R849 CLK2.n562 CLK2.n561 4.65
R850 CLK2.n558 CLK2.n557 4.65
R851 CLK2.n554 CLK2.n553 4.65
R852 CLK2.n617 CLK2.n98 4.65
R853 CLK2.n616 CLK2.n615 4.65
R854 CLK2.n621 CLK2.n620 4.65
R855 CLK2.n687 CLK2.n686 4.65
R856 CLK2.n683 CLK2.n682 4.65
R857 CLK2.n679 CLK2.n678 4.65
R858 CLK2.n675 CLK2.n674 4.65
R859 CLK2.n670 CLK2.n669 4.65
R860 CLK2.n666 CLK2.n665 4.65
R861 CLK2.n662 CLK2.n661 4.65
R862 CLK2.n658 CLK2.n657 4.65
R863 CLK2.n654 CLK2.n651 4.65
R864 CLK2.n650 CLK2.n649 4.65
R865 CLK2.n646 CLK2.n645 4.65
R866 CLK2.n641 CLK2.n640 4.65
R867 CLK2.n637 CLK2.n636 4.65
R868 CLK2.n633 CLK2.n632 4.65
R869 CLK2.n629 CLK2.n628 4.65
R870 CLK2.n689 CLK2.n92 4.65
R871 CLK2.n690 CLK2.n91 4.65
R872 CLK2.n769 CLK2.n768 4.65
R873 CLK2.n765 CLK2.n764 4.65
R874 CLK2.n761 CLK2.n760 4.65
R875 CLK2.n757 CLK2.n756 4.65
R876 CLK2.n753 CLK2.n752 4.65
R877 CLK2.n749 CLK2.n748 4.65
R878 CLK2.n744 CLK2.n743 4.65
R879 CLK2.n740 CLK2.n739 4.65
R880 CLK2.n736 CLK2.n735 4.65
R881 CLK2.n732 CLK2.n731 4.65
R882 CLK2.n728 CLK2.n725 4.65
R883 CLK2.n724 CLK2.n723 4.65
R884 CLK2.n720 CLK2.n719 4.65
R885 CLK2.n715 CLK2.n714 4.65
R886 CLK2.n711 CLK2.n710 4.65
R887 CLK2.n707 CLK2.n706 4.65
R888 CLK2.n703 CLK2.n702 4.65
R889 CLK2.n698 CLK2.n697 4.65
R890 CLK2.n694 CLK2.n693 4.65
R891 CLK2.n773 CLK2.n87 4.65
R892 CLK2.n772 CLK2.n771 4.65
R893 CLK2.n779 CLK2.n778 4.65
R894 CLK2.n788 CLK2.n787 4.65
R895 CLK2.n792 CLK2.n791 4.65
R896 CLK2.n796 CLK2.n795 4.65
R897 CLK2.n800 CLK2.n799 4.65
R898 CLK2.n804 CLK2.n803 4.65
R899 CLK2.n808 CLK2.n807 4.65
R900 CLK2.n813 CLK2.n812 4.65
R901 CLK2.n817 CLK2.n816 4.65
R902 CLK2.n821 CLK2.n820 4.65
R903 CLK2.n823 CLK2.n822 4.65
R904 CLK2.n827 CLK2.n826 4.65
R905 CLK2.n831 CLK2.n830 4.65
R906 CLK2.n835 CLK2.n834 4.65
R907 CLK2.n840 CLK2.n839 4.65
R908 CLK2.n844 CLK2.n843 4.65
R909 CLK2.n848 CLK2.n847 4.65
R910 CLK2.n852 CLK2.n851 4.65
R911 CLK2.n939 CLK2.n938 4.65
R912 CLK2.n935 CLK2.n934 4.65
R913 CLK2.n931 CLK2.n930 4.65
R914 CLK2.n927 CLK2.n926 4.65
R915 CLK2.n923 CLK2.n922 4.65
R916 CLK2.n919 CLK2.n918 4.65
R917 CLK2.n914 CLK2.n913 4.65
R918 CLK2.n910 CLK2.n909 4.65
R919 CLK2.n906 CLK2.n905 4.65
R920 CLK2.n902 CLK2.n901 4.65
R921 CLK2.n898 CLK2.n895 4.65
R922 CLK2.n894 CLK2.n893 4.65
R923 CLK2.n890 CLK2.n889 4.65
R924 CLK2.n885 CLK2.n884 4.65
R925 CLK2.n881 CLK2.n880 4.65
R926 CLK2.n877 CLK2.n876 4.65
R927 CLK2.n873 CLK2.n872 4.65
R928 CLK2.n868 CLK2.n867 4.65
R929 CLK2.n944 CLK2.n943 4.65
R930 CLK2.n942 CLK2.n941 4.65
R931 CLK2.n953 CLK2.n74 4.65
R932 CLK2.n952 CLK2.n951 4.65
R933 CLK2.n6 CLK2.n5 4.65
R934 CLK2.n10 CLK2.n9 4.65
R935 CLK2.n14 CLK2.n13 4.65
R936 CLK2.n18 CLK2.n17 4.65
R937 CLK2.n22 CLK2.n21 4.65
R938 CLK2.n26 CLK2.n25 4.65
R939 CLK2.n31 CLK2.n30 4.65
R940 CLK2.n35 CLK2.n34 4.65
R941 CLK2.n39 CLK2.n38 4.65
R942 CLK2.n43 CLK2.n40 4.65
R943 CLK2.n47 CLK2.n46 4.65
R944 CLK2.n51 CLK2.n50 4.65
R945 CLK2.n55 CLK2.n54 4.65
R946 CLK2.n60 CLK2.n59 4.65
R947 CLK2.n64 CLK2.n63 4.65
R948 CLK2.n68 CLK2.n67 4.65
R949 CLK2.n72 CLK2.n71 4.65
R950 CLK2 CLK2.n964 4.52
R951 CLK2.n784 EESPFAL_s1_0/CLK2 4.509
R952 EESPFAL_s3_0/CLK2 CLK2.n140 4.509
R953 CLK2.n367 CLK2.n366 4.5
R954 CLK2.n369 CLK2.n111 4.5
R955 CLK2.n300 CLK2.n143 3.715
R956 CLK2.n305 CLK2.n141 3.715
R957 CLK2.n951 CLK2.n950 3.715
R958 CLK2.n304 CLK2.n302 3.039
R959 CLK2.n619 CLK2.n95 3.039
R960 CLK2.n777 CLK2.n86 3.039
R961 CLK2.n459 CLK2.n102 3.039
R962 CLK2.n310 CLK2.n309 3.033
R963 CLK2.n386 CLK2.n385 3.033
R964 CLK2.n783 CLK2.n782 3.033
R965 CLK2.n963 CLK2.n962 3.033
R966 CLK2.n962 CLK2.n961 2.72
R967 CLK2.n361 CLK2.n360 2.682
R968 CLK2.n376 CLK2.n375 2.682
R969 CLK2.n856 CLK2.n855 2.682
R970 CLK2.n864 CLK2.n863 2.682
R971 CLK2.n957 CLK2.n956 2.682
R972 CLK2.n619 CLK2.n618 2.6
R973 CLK2.n775 CLK2.n774 2.57
R974 CLK2.n97 CLK2.n96 2.57
R975 CLK2.n463 CLK2.n462 2.57
R976 CLK2.n457 CLK2.n456 2.57
R977 CLK2.n300 CLK2.n299 2.57
R978 CLK2.n303 CLK2.n141 2.57
R979 CLK2.n94 CLK2.n93 2.57
R980 CLK2.n85 CLK2.n84 2.57
R981 CLK2.n946 CLK2.n945 2.57
R982 CLK2.n950 CLK2.n949 2.57
R983 CLK2.n370 CLK2.n110 2.251
R984 CLK2.n369 CLK2.n368 2.246
R985 CLK2.n965 CLK2.n73 2.246
R986 CLK2.n459 CLK2.n458 2.224
R987 CLK2.n302 CLK2.n301 2.224
R988 CLK2.n777 CLK2.n776 2.224
R989 CLK2.n297 CLK2.n296 2.203
R990 CLK2.n308 CLK2.n307 2.203
R991 CLK2.n454 CLK2.n452 2.203
R992 CLK2.n466 CLK2.n464 2.203
R993 CLK2.n772 CLK2.n770 2.203
R994 CLK2.n781 CLK2.n780 2.203
R995 CLK2.n942 CLK2.n940 2.203
R996 CLK2.n964 CLK2.n953 2.203
R997 CLK2.n121 CLK2.n113 1.76
R998 CLK2.n79 CLK2.n78 1.656
R999 CLK2.n449 CLK2.n448 1.655
R1000 CLK2.n4 CLK2.n3 1.655
R1001 CLK2.n767 CLK2.n766 1.655
R1002 CLK2.n685 CLK2.n684 1.655
R1003 CLK2.n611 CLK2.n610 1.655
R1004 CLK2.n468 CLK2.n467 1.655
R1005 CLK2.n312 CLK2.n311 1.655
R1006 CLK2.n293 CLK2.n292 1.655
R1007 CLK2.n241 CLK2.n240 1.655
R1008 CLK2.n206 CLK2.n205 1.655
R1009 CLK2.n250 CLK2.n249 1.655
R1010 CLK2.n359 CLK2.n117 1.655
R1011 CLK2.n374 CLK2.n373 1.655
R1012 CLK2.n543 CLK2.n542 1.655
R1013 CLK2.n552 CLK2.n551 1.655
R1014 CLK2.n627 CLK2.n626 1.655
R1015 CLK2.n692 CLK2.n691 1.655
R1016 CLK2.n786 CLK2.n785 1.655
R1017 CLK2.n937 CLK2.n936 1.655
R1018 CLK2.n862 CLK2.n861 1.655
R1019 CLK2.n955 CLK2.n954 1.655
R1020 CLK2.n387 CLK2.n371 1.497
R1021 CLK2.n616 CLK2.n614 1.14
R1022 CLK2.n688 CLK2.n622 1.14
R1023 CLK2.n362 CLK2.n361 1.095
R1024 CLK2.n380 CLK2.n376 1.095
R1025 CLK2.n855 CLK2.n854 1.095
R1026 CLK2.n868 CLK2.n864 1.095
R1027 CLK2.n958 CLK2.n957 1.073
R1028 CLK2.n246 CLK2.n245 1.047
R1029 CLK2.n690 CLK2.n689 1.047
R1030 CLK2.n609 CLK2.n547 1.046
R1031 CLK2.n366 CLK2.n113 0.96
R1032 EESPFAL_s1_0/CLK2 CLK2.n783 0.928
R1033 CLK2.n309 EESPFAL_s3_0/CLK2 0.927
R1034 EESPFAL_s2_0/CLK2 CLK2.n370 0.648
R1035 CLK2.n297 CLK2.n142 0.125
R1036 CLK2.n307 CLK2.n306 0.125
R1037 CLK2.n455 CLK2.n454 0.125
R1038 CLK2.n464 CLK2.n461 0.125
R1039 CLK2.n617 CLK2.n616 0.125
R1040 CLK2.n622 CLK2.n621 0.125
R1041 CLK2.n773 CLK2.n772 0.125
R1042 CLK2.n780 CLK2.n779 0.125
R1043 CLK2.n944 CLK2.n942 0.125
R1044 CLK2.n953 CLK2.n952 0.125
R1045 CLK2.n952 CLK2.n948 0.125
R1046 CLK2.n306 CLK2.n302 0.12
R1047 CLK2.n621 CLK2.n619 0.12
R1048 CLK2.n779 CLK2.n777 0.12
R1049 CLK2.n461 CLK2.n459 0.119
R1050 CLK2.n618 CLK2.n617 0.119
R1051 CLK2.n301 CLK2.n142 0.119
R1052 CLK2.n776 CLK2.n773 0.119
R1053 CLK2.n458 CLK2.n455 0.117
R1054 CLK2.n243 CLK2.n179 0.1
R1055 CLK2.n235 CLK2.n179 0.1
R1056 CLK2.n235 CLK2.n234 0.1
R1057 CLK2.n232 CLK2.n185 0.1
R1058 CLK2.n224 CLK2.n185 0.1
R1059 CLK2.n224 CLK2.n223 0.1
R1060 CLK2.n222 CLK2.n191 0.1
R1061 CLK2.n214 CLK2.n191 0.1
R1062 CLK2.n212 CLK2.n211 0.1
R1063 CLK2.n211 CLK2.n198 0.1
R1064 CLK2.n203 CLK2.n198 0.1
R1065 CLK2.n295 CLK2.n145 0.1
R1066 CLK2.n287 CLK2.n145 0.1
R1067 CLK2.n287 CLK2.n286 0.1
R1068 CLK2.n286 CLK2.n285 0.1
R1069 CLK2.n285 CLK2.n151 0.1
R1070 CLK2.n277 CLK2.n276 0.1
R1071 CLK2.n276 CLK2.n275 0.1
R1072 CLK2.n275 CLK2.n158 0.1
R1073 CLK2.n267 CLK2.n266 0.1
R1074 CLK2.n266 CLK2.n265 0.1
R1075 CLK2.n257 CLK2.n171 0.1
R1076 CLK2.n257 CLK2.n256 0.1
R1077 CLK2.n256 CLK2.n255 0.1
R1078 CLK2.n247 CLK2.n177 0.1
R1079 CLK2.n247 CLK2.n246 0.1
R1080 CLK2.n315 CLK2.n314 0.1
R1081 CLK2.n316 CLK2.n315 0.1
R1082 CLK2.n316 CLK2.n134 0.1
R1083 CLK2.n324 CLK2.n134 0.1
R1084 CLK2.n325 CLK2.n324 0.1
R1085 CLK2.n327 CLK2.n128 0.1
R1086 CLK2.n336 CLK2.n128 0.1
R1087 CLK2.n337 CLK2.n336 0.1
R1088 CLK2.n338 CLK2.n122 0.1
R1089 CLK2.n347 CLK2.n122 0.1
R1090 CLK2.n351 CLK2.n349 0.1
R1091 CLK2.n451 CLK2.n447 0.1
R1092 CLK2.n447 CLK2.n443 0.1
R1093 CLK2.n443 CLK2.n439 0.1
R1094 CLK2.n439 CLK2.n435 0.1
R1095 CLK2.n435 CLK2.n431 0.1
R1096 CLK2.n426 CLK2.n422 0.1
R1097 CLK2.n422 CLK2.n418 0.1
R1098 CLK2.n418 CLK2.n414 0.1
R1099 CLK2.n407 CLK2.n406 0.1
R1100 CLK2.n406 CLK2.n402 0.1
R1101 CLK2.n397 CLK2.n393 0.1
R1102 CLK2.n393 CLK2.n389 0.1
R1103 CLK2.n474 CLK2.n470 0.1
R1104 CLK2.n478 CLK2.n474 0.1
R1105 CLK2.n482 CLK2.n478 0.1
R1106 CLK2.n486 CLK2.n482 0.1
R1107 CLK2.n490 CLK2.n486 0.1
R1108 CLK2.n499 CLK2.n495 0.1
R1109 CLK2.n503 CLK2.n499 0.1
R1110 CLK2.n504 CLK2.n503 0.1
R1111 CLK2.n515 CLK2.n511 0.1
R1112 CLK2.n519 CLK2.n515 0.1
R1113 CLK2.n528 CLK2.n524 0.1
R1114 CLK2.n532 CLK2.n528 0.1
R1115 CLK2.n536 CLK2.n532 0.1
R1116 CLK2.n545 CLK2.n541 0.1
R1117 CLK2.n547 CLK2.n545 0.1
R1118 CLK2.n608 CLK2.n604 0.1
R1119 CLK2.n604 CLK2.n600 0.1
R1120 CLK2.n595 CLK2.n591 0.1
R1121 CLK2.n591 CLK2.n587 0.1
R1122 CLK2.n587 CLK2.n583 0.1
R1123 CLK2.n576 CLK2.n575 0.1
R1124 CLK2.n575 CLK2.n571 0.1
R1125 CLK2.n566 CLK2.n562 0.1
R1126 CLK2.n562 CLK2.n558 0.1
R1127 CLK2.n558 CLK2.n554 0.1
R1128 CLK2.n687 CLK2.n683 0.1
R1129 CLK2.n683 CLK2.n679 0.1
R1130 CLK2.n679 CLK2.n675 0.1
R1131 CLK2.n670 CLK2.n666 0.1
R1132 CLK2.n666 CLK2.n662 0.1
R1133 CLK2.n662 CLK2.n658 0.1
R1134 CLK2.n651 CLK2.n650 0.1
R1135 CLK2.n650 CLK2.n646 0.1
R1136 CLK2.n641 CLK2.n637 0.1
R1137 CLK2.n637 CLK2.n633 0.1
R1138 CLK2.n633 CLK2.n629 0.1
R1139 CLK2.n769 CLK2.n765 0.1
R1140 CLK2.n765 CLK2.n761 0.1
R1141 CLK2.n761 CLK2.n757 0.1
R1142 CLK2.n757 CLK2.n753 0.1
R1143 CLK2.n753 CLK2.n749 0.1
R1144 CLK2.n744 CLK2.n740 0.1
R1145 CLK2.n740 CLK2.n736 0.1
R1146 CLK2.n736 CLK2.n732 0.1
R1147 CLK2.n725 CLK2.n724 0.1
R1148 CLK2.n724 CLK2.n720 0.1
R1149 CLK2.n715 CLK2.n711 0.1
R1150 CLK2.n711 CLK2.n707 0.1
R1151 CLK2.n707 CLK2.n703 0.1
R1152 CLK2.n698 CLK2.n694 0.1
R1153 CLK2.n694 CLK2.n690 0.1
R1154 CLK2.n792 CLK2.n788 0.1
R1155 CLK2.n796 CLK2.n792 0.1
R1156 CLK2.n800 CLK2.n796 0.1
R1157 CLK2.n804 CLK2.n800 0.1
R1158 CLK2.n808 CLK2.n804 0.1
R1159 CLK2.n817 CLK2.n813 0.1
R1160 CLK2.n821 CLK2.n817 0.1
R1161 CLK2.n822 CLK2.n821 0.1
R1162 CLK2.n831 CLK2.n827 0.1
R1163 CLK2.n835 CLK2.n831 0.1
R1164 CLK2.n844 CLK2.n840 0.1
R1165 CLK2.n848 CLK2.n844 0.1
R1166 CLK2.n852 CLK2.n848 0.1
R1167 CLK2.n939 CLK2.n935 0.1
R1168 CLK2.n935 CLK2.n931 0.1
R1169 CLK2.n931 CLK2.n927 0.1
R1170 CLK2.n927 CLK2.n923 0.1
R1171 CLK2.n923 CLK2.n919 0.1
R1172 CLK2.n914 CLK2.n910 0.1
R1173 CLK2.n910 CLK2.n906 0.1
R1174 CLK2.n906 CLK2.n902 0.1
R1175 CLK2.n895 CLK2.n894 0.1
R1176 CLK2.n894 CLK2.n890 0.1
R1177 CLK2.n885 CLK2.n881 0.1
R1178 CLK2.n881 CLK2.n877 0.1
R1179 CLK2.n877 CLK2.n873 0.1
R1180 CLK2.n10 CLK2.n6 0.1
R1181 CLK2.n14 CLK2.n10 0.1
R1182 CLK2.n18 CLK2.n14 0.1
R1183 CLK2.n22 CLK2.n18 0.1
R1184 CLK2.n26 CLK2.n22 0.1
R1185 CLK2.n35 CLK2.n31 0.1
R1186 CLK2.n39 CLK2.n35 0.1
R1187 CLK2.n40 CLK2.n39 0.1
R1188 CLK2.n51 CLK2.n47 0.1
R1189 CLK2.n55 CLK2.n51 0.1
R1190 CLK2.n64 CLK2.n60 0.1
R1191 CLK2.n68 CLK2.n64 0.1
R1192 CLK2.n72 CLK2.n68 0.1
R1193 CLK2.n244 CLK2.n243 0.087
R1194 CLK2.n203 CLK2.n202 0.087
R1195 CLK2.n255 CLK2.n173 0.087
R1196 CLK2.n364 CLK2.n363 0.087
R1197 CLK2.n537 CLK2.n536 0.087
R1198 CLK2.n614 CLK2.n613 0.087
R1199 CLK2.n554 CLK2.n550 0.087
R1200 CLK2.n688 CLK2.n687 0.087
R1201 CLK2.n629 CLK2.n625 0.087
R1202 CLK2.n703 CLK2.n699 0.087
R1203 CLK2.n853 CLK2.n852 0.087
R1204 CLK2.n873 CLK2.n869 0.087
R1205 CLK2.n351 CLK2.n350 0.086
R1206 CLK2.n73 CLK2.n72 0.077
R1207 CLK2.n233 CLK2.n232 0.075
R1208 EESPFAL_s3_0/EESPFAL_INV4_0/CLK CLK2.n222 0.075
R1209 CLK2.n214 CLK2.n213 0.075
R1210 CLK2.n296 CLK2.n295 0.075
R1211 CLK2.n277 CLK2.n156 0.075
R1212 CLK2.n267 EESPFAL_s3_0/EESPFAL_NAND_v3_1/CLK 0.075
R1213 CLK2.n265 CLK2.n165 0.075
R1214 CLK2.n327 CLK2.n326 0.075
R1215 CLK2.n338 EESPFAL_s3_0/EESPFAL_NAND_v3_0/CLK 0.075
R1216 CLK2.n348 CLK2.n347 0.075
R1217 CLK2.n452 CLK2.n451 0.075
R1218 CLK2.n427 CLK2.n426 0.075
R1219 CLK2.n407 EESPFAL_s2_0/EESPFAL_NAND_v3_1/CLK 0.075
R1220 CLK2.n402 CLK2.n398 0.075
R1221 CLK2.n470 CLK2.n466 0.075
R1222 CLK2.n495 CLK2.n491 0.075
R1223 CLK2.n511 EESPFAL_s2_0/EESPFAL_NAND_v3_0/CLK 0.075
R1224 CLK2.n520 CLK2.n519 0.075
R1225 CLK2.n613 CLK2.n609 0.075
R1226 CLK2.n596 CLK2.n595 0.075
R1227 CLK2.n576 EESPFAL_s2_0/EESPFAL_INV4_2/CLK 0.075
R1228 CLK2.n571 CLK2.n567 0.075
R1229 CLK2.n671 CLK2.n670 0.075
R1230 CLK2.n651 EESPFAL_s1_0/EESPFAL_INV4_0/CLK 0.075
R1231 CLK2.n646 CLK2.n642 0.075
R1232 CLK2.n770 CLK2.n769 0.075
R1233 CLK2.n745 CLK2.n744 0.075
R1234 CLK2.n725 EESPFAL_s1_0/EESPFAL_NAND_v3_1/CLK 0.075
R1235 CLK2.n720 CLK2.n716 0.075
R1236 CLK2.n813 CLK2.n809 0.075
R1237 CLK2.n827 EESPFAL_s1_0/EESPFAL_NAND_v3_0/CLK 0.075
R1238 CLK2.n836 CLK2.n835 0.075
R1239 CLK2.n940 CLK2.n939 0.075
R1240 CLK2.n915 CLK2.n914 0.075
R1241 CLK2.n895 EESPFAL_s0_0/EESPFAL_NAND_v3_1/CLK 0.075
R1242 CLK2.n890 CLK2.n886 0.075
R1243 CLK2.n6 CLK2.n2 0.075
R1244 CLK2.n31 CLK2.n27 0.075
R1245 CLK2.n47 CLK2 0.075
R1246 CLK2.n56 CLK2.n55 0.075
R1247 CLK2.n382 CLK2.n381 0.074
R1248 CLK2.n314 CLK2.n140 0.072
R1249 CLK2.n389 CLK2.n388 0.072
R1250 CLK2.n788 CLK2.n784 0.072
R1251 CLK2.n947 CLK2.n944 0.062
R1252 CLK2.n364 CLK2.n111 0.06
R1253 CLK2.n371 EESPFAL_s2_0/CLK2 0.042
R1254 CLK2.n388 CLK2.n387 0.026
R1255 CLK2.n234 CLK2.n233 0.025
R1256 CLK2.n223 EESPFAL_s3_0/EESPFAL_INV4_0/CLK 0.025
R1257 CLK2.n213 CLK2.n212 0.025
R1258 CLK2.n156 CLK2.n151 0.025
R1259 EESPFAL_s3_0/EESPFAL_NAND_v3_1/CLK CLK2.n158 0.025
R1260 CLK2.n171 CLK2.n165 0.025
R1261 CLK2.n309 CLK2.n308 0.025
R1262 CLK2.n326 CLK2.n325 0.025
R1263 EESPFAL_s3_0/EESPFAL_NAND_v3_0/CLK CLK2.n337 0.025
R1264 CLK2.n349 CLK2.n348 0.025
R1265 CLK2.n431 CLK2.n427 0.025
R1266 CLK2.n414 EESPFAL_s2_0/EESPFAL_NAND_v3_1/CLK 0.025
R1267 CLK2.n398 CLK2.n397 0.025
R1268 CLK2.n491 CLK2.n490 0.025
R1269 CLK2.n504 EESPFAL_s2_0/EESPFAL_NAND_v3_0/CLK 0.025
R1270 CLK2.n524 CLK2.n520 0.025
R1271 CLK2.n609 CLK2.n608 0.025
R1272 CLK2.n600 CLK2.n596 0.025
R1273 CLK2.n583 EESPFAL_s2_0/EESPFAL_INV4_2/CLK 0.025
R1274 CLK2.n567 CLK2.n566 0.025
R1275 CLK2.n675 CLK2.n671 0.025
R1276 CLK2.n658 EESPFAL_s1_0/EESPFAL_INV4_0/CLK 0.025
R1277 CLK2.n642 CLK2.n641 0.025
R1278 CLK2.n749 CLK2.n745 0.025
R1279 CLK2.n732 EESPFAL_s1_0/EESPFAL_NAND_v3_1/CLK 0.025
R1280 CLK2.n716 CLK2.n715 0.025
R1281 CLK2.n783 CLK2.n781 0.025
R1282 CLK2.n809 CLK2.n808 0.025
R1283 CLK2.n822 EESPFAL_s1_0/EESPFAL_NAND_v3_0/CLK 0.025
R1284 CLK2.n840 CLK2.n836 0.025
R1285 CLK2.n919 CLK2.n915 0.025
R1286 CLK2.n902 EESPFAL_s0_0/EESPFAL_NAND_v3_1/CLK 0.025
R1287 CLK2.n886 CLK2.n885 0.025
R1288 CLK2.n27 CLK2.n26 0.025
R1289 CLK2.n40 CLK2 0.025
R1290 CLK2.n60 CLK2.n56 0.025
R1291 EESPFAL_s0_0/CLK2 CLK2.n965 0.023
R1292 CLK2.n963 CLK2.n958 0.021
R1293 CLK2.n370 CLK2.n369 0.017
R1294 CLK2.n111 CLK2.n110 0.015
R1295 CLK2.n965 CLK2 0.014
R1296 CLK2.n386 CLK2.n382 0.013
R1297 CLK2.n350 CLK2.n112 0.013
R1298 CLK2.n371 CLK2.n109 0.012
R1299 CLK2.n245 CLK2.n244 0.012
R1300 CLK2.n177 CLK2.n173 0.012
R1301 CLK2.n363 CLK2.n362 0.012
R1302 CLK2.n381 CLK2.n380 0.012
R1303 CLK2.n541 CLK2.n537 0.012
R1304 CLK2.n689 CLK2.n688 0.012
R1305 CLK2.n699 CLK2.n698 0.012
R1306 CLK2.n854 CLK2.n853 0.012
R1307 CLK2.n869 CLK2.n868 0.012
R1308 CLK2.n964 CLK2.n963 0.012
R1309 CLK2.n964 CLK2.n73 0.01
R1310 CLK2.n368 CLK2.n367 0.009
R1311 CLK2.n368 CLK2.n110 0.009
R1312 CLK2.n367 CLK2.n112 0.007
R1313 CLK2.n308 CLK2.n140 0.002
R1314 CLK2.n784 CLK2.n781 0.002
R1315 CLK2.n387 CLK2.n386 0.001
R1316 Dis1.n1 Dis1 598.4
R1317 Dis1.n18 EESPFAL_s2_0/EESPFAL_INV4_0/Dis 563.2
R1318 Dis1.n14 EESPFAL_s2_0/EESPFAL_INV4_1/Dis 563.2
R1319 Dis1.n29 EESPFAL_s1_0/EESPFAL_INV4_2/Dis 556.8
R1320 Dis1.n25 EESPFAL_s1_0/EESPFAL_INV4_1/Dis 556.8
R1321 Dis1.n10 EESPFAL_s3_0/EESPFAL_INV4_2/Dis 556.8
R1322 Dis1.n6 EESPFAL_s3_0/EESPFAL_INV4_1/Dis 556.8
R1323 Dis1.n0 Dis1.t23 504.5
R1324 Dis1.n32 Dis1.t17 504.5
R1325 Dis1.n28 Dis1.t32 504.5
R1326 Dis1.n24 Dis1.t16 504.5
R1327 Dis1.n21 Dis1.t34 504.5
R1328 Dis1.n17 Dis1.t11 504.5
R1329 Dis1.n13 Dis1.t24 504.5
R1330 Dis1.n9 Dis1.t10 504.5
R1331 Dis1.n5 Dis1.t14 504.5
R1332 Dis1.n4 Dis1.t27 504.5
R1333 Dis1.n3 Dis1.t20 504.5
R1334 Dis1.n2 Dis1.t13 389.3
R1335 Dis1.n1 Dis1.t6 389.3
R1336 Dis1.n0 Dis1.t4 389.3
R1337 Dis1.n32 Dis1.t9 389.3
R1338 Dis1.n30 Dis1.t22 389.3
R1339 Dis1.n29 Dis1.t31 389.3
R1340 Dis1.n28 Dis1.t19 389.3
R1341 Dis1.n26 Dis1.t3 389.3
R1342 Dis1.n25 Dis1.t15 389.3
R1343 Dis1.n24 Dis1.t0 389.3
R1344 Dis1.n21 Dis1.t12 389.3
R1345 Dis1.n19 Dis1.t2 389.3
R1346 Dis1.n18 Dis1.t25 389.3
R1347 Dis1.n17 Dis1.t18 389.3
R1348 Dis1.n15 Dis1.t21 389.3
R1349 Dis1.n14 Dis1.t5 389.3
R1350 Dis1.n13 Dis1.t35 389.3
R1351 Dis1.n11 Dis1.t28 389.3
R1352 Dis1.n10 Dis1.t7 389.3
R1353 Dis1.n9 Dis1.t26 389.3
R1354 Dis1.n7 Dis1.t1 389.3
R1355 Dis1.n6 Dis1.t30 389.3
R1356 Dis1.n5 Dis1.t29 389.3
R1357 Dis1.n4 Dis1.t33 389.3
R1358 Dis1.n3 Dis1.t8 389.3
R1359 Dis1.n22 EESPFAL_s2_0/EESPFAL_4in_NAND_0/Dis 281.856
R1360 Dis1.n33 EESPFAL_s0_0/EESPFAL_NAND_v3_2/Dis 241.216
R1361 Dis1.n34 EESPFAL_s0_0/EESPFAL_XOR_v3_0/Dis 240.897
R1362 Dis1.n8 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/Dis 235.714
R1363 Dis1.n23 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/Dis 227.781
R1364 Dis1.n31 EESPFAL_s1_0/EESPFAL_XOR_v3_0/Dis 227.456
R1365 Dis1.n27 EESPFAL_s1_0/EESPFAL_XOR_v3_1/Dis 227.456
R1366 Dis1.n12 EESPFAL_s3_0/EESPFAL_XOR_v3_0/Dis 227.456
R1367 Dis1.n8 EESPFAL_s3_0/EESPFAL_XOR_v3_1/Dis 227.456
R1368 Dis1.n20 EESPFAL_s2_0/EESPFAL_XOR_v3_1/Dis 137.536
R1369 Dis1.n16 EESPFAL_s2_0/EESPFAL_XOR_v3_0/Dis 137.536
R1370 Dis1.n2 Dis1.n1 115.2
R1371 Dis1.n30 Dis1.n29 115.2
R1372 Dis1.n26 Dis1.n25 115.2
R1373 Dis1.n19 Dis1.n18 115.2
R1374 Dis1.n15 Dis1.n14 115.2
R1375 Dis1.n11 Dis1.n10 115.2
R1376 Dis1.n7 Dis1.n6 115.2
R1377 Dis1.n22 Dis1.n20 9.213
R1378 Dis1.n27 Dis1.n23 7.933
R1379 Dis1.n33 EESPFAL_s1_0/Dis1 4.681
R1380 Dis1.n16 EESPFAL_s2_0/Dis1 3.351
R1381 EESPFAL_s1_0/Dis1 Dis1.n31 3.266
R1382 EESPFAL_s3_0/Dis1 Dis1.n12 3.266
R1383 Dis1 Dis1.n0 3.2
R1384 EESPFAL_s0_0/EESPFAL_XOR_v3_0/Dis Dis1.n2 3.2
R1385 EESPFAL_s0_0/EESPFAL_NAND_v3_2/Dis Dis1.n32 3.2
R1386 EESPFAL_s1_0/EESPFAL_INV4_2/Dis Dis1.n28 3.2
R1387 EESPFAL_s1_0/EESPFAL_XOR_v3_0/Dis Dis1.n30 3.2
R1388 EESPFAL_s1_0/EESPFAL_INV4_1/Dis Dis1.n24 3.2
R1389 EESPFAL_s1_0/EESPFAL_XOR_v3_1/Dis Dis1.n26 3.2
R1390 EESPFAL_s2_0/EESPFAL_4in_NAND_0/Dis Dis1.n21 3.2
R1391 EESPFAL_s2_0/EESPFAL_INV4_0/Dis Dis1.n17 3.2
R1392 EESPFAL_s2_0/EESPFAL_XOR_v3_1/Dis Dis1.n19 3.2
R1393 EESPFAL_s2_0/EESPFAL_INV4_1/Dis Dis1.n13 3.2
R1394 EESPFAL_s2_0/EESPFAL_XOR_v3_0/Dis Dis1.n15 3.2
R1395 EESPFAL_s3_0/EESPFAL_INV4_2/Dis Dis1.n9 3.2
R1396 EESPFAL_s3_0/EESPFAL_XOR_v3_0/Dis Dis1.n11 3.2
R1397 EESPFAL_s3_0/EESPFAL_INV4_1/Dis Dis1.n5 3.2
R1398 EESPFAL_s3_0/EESPFAL_XOR_v3_1/Dis Dis1.n7 3.2
R1399 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/Dis Dis1.n4 3.2
R1400 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/Dis Dis1.n3 3.2
R1401 Dis1 Dis1.n34 3.049
R1402 EESPFAL_s2_0/Dis1 EESPFAL_s3_0/Dis1 2.199
R1403 Dis1.n23 Dis1.n22 1.174
R1404 Dis1.n12 Dis1.n8 0.627
R1405 Dis1.n20 Dis1.n16 0.627
R1406 Dis1.n31 Dis1.n27 0.627
R1407 Dis1.n34 Dis1.n33 0.625
R1408 EESPFAL_s0_0/Dis1 Dis1 0.2
R1409 GND.n1755 GND.n1400 16794.9
R1410 GND.n1659 GND.n1460 14060
R1411 GND.n1455 GND.n1454 6512
R1412 GND.n1400 GND.n1399 4190.48
R1413 GND.n1399 GND.t257 3724.87
R1414 GND.n1530 GND.n1526 3616.44
R1415 GND.n1659 GND.n1459 3616.44
R1416 GND.t291 GND.t280 3300
R1417 GND.n1526 GND.t40 3214.61
R1418 GND.n1459 GND.t15 3214.61
R1419 GND.n1454 GND.t275 2910
R1420 GND.t275 GND.t99 1500
R1421 GND.t99 GND.t236 1500
R1422 GND.n1709 GND.t291 1250
R1423 GND.n1454 GND.t134 968
R1424 GND.n1460 GND.n1455 880
R1425 GND.n1214 GND.n1213 594.594
R1426 GND.n1216 GND.n1214 594.594
R1427 GND.n1216 GND.n1215 594.594
R1428 GND.n1226 GND.n1225 594.594
R1429 GND.n1236 GND.n1095 594.594
R1430 GND.n1238 GND.n1237 594.594
R1431 GND.n1238 GND.n1089 594.594
R1432 GND.n1246 GND.n1089 594.594
R1433 GND.n1149 GND.n1148 594.594
R1434 GND.n1151 GND.n1150 594.594
R1435 GND.n1160 GND.n1159 594.594
R1436 GND.n1162 GND.n1160 594.594
R1437 GND.n1162 GND.n1161 594.594
R1438 GND.n1172 GND.n1171 594.594
R1439 GND.n1182 GND.n1124 594.594
R1440 GND.n1184 GND.n1183 594.594
R1441 GND.n1184 GND.n1118 594.594
R1442 GND.n1192 GND.n1118 594.594
R1443 GND.n1194 GND.n1193 594.594
R1444 GND.n1202 GND.n1112 594.594
R1445 GND.n1258 GND.n1257 594.594
R1446 GND.n1260 GND.n1259 594.594
R1447 GND.n1269 GND.n1268 594.594
R1448 GND.n1271 GND.n1269 594.594
R1449 GND.n1271 GND.n1270 594.594
R1450 GND.n1281 GND.n1280 594.594
R1451 GND.n1291 GND.n1067 594.594
R1452 GND.n1293 GND.n1292 594.594
R1453 GND.n1293 GND.n1061 594.594
R1454 GND.n1301 GND.n1061 594.594
R1455 GND.n1303 GND.n1302 594.594
R1456 GND.n1312 GND.n1055 594.594
R1457 GND.n1213 GND.t249 557.432
R1458 GND.n1227 GND.t298 557.432
R1459 GND.n1227 GND.t6 557.432
R1460 GND.t252 GND.n1246 557.432
R1461 GND.n1159 GND.t158 557.432
R1462 GND.n1173 GND.t285 557.432
R1463 GND.n1173 GND.t48 557.432
R1464 GND.t312 GND.n1192 557.432
R1465 GND.n1268 GND.t70 557.432
R1466 GND.n1282 GND.t250 557.432
R1467 GND.n1282 GND.t247 557.432
R1468 GND.t90 GND.n1301 557.432
R1469 GND.n1755 GND.n1754 523.031
R1470 GND.t66 GND.n1753 490.341
R1471 GND.n1225 GND.t293 483.108
R1472 GND.t303 GND.n1236 483.108
R1473 GND.n1151 GND.t262 483.108
R1474 GND.n1171 GND.t231 483.108
R1475 GND.t316 GND.n1182 483.108
R1476 GND.n1194 GND.t84 483.108
R1477 GND.n1260 GND.t112 483.108
R1478 GND.n1280 GND.t189 483.108
R1479 GND.t177 GND.n1291 483.108
R1480 GND.n1303 GND.t310 483.108
R1481 GND.n1148 GND.t71 408.783
R1482 GND.t308 GND.n1202 408.783
R1483 GND.n1257 GND.t81 408.783
R1484 GND.t143 GND.n1312 408.783
R1485 GND.n942 GND.n941 341.085
R1486 GND.n944 GND.n942 341.085
R1487 GND.n944 GND.n943 341.085
R1488 GND.n954 GND.n953 341.085
R1489 GND.n964 GND.n837 341.085
R1490 GND.n966 GND.n965 341.085
R1491 GND.n966 GND.n831 341.085
R1492 GND.n974 GND.n831 341.085
R1493 GND.n888 GND.n887 341.085
R1494 GND.n889 GND.n874 341.085
R1495 GND.n898 GND.n874 341.085
R1496 GND.n899 GND.n898 341.085
R1497 GND.n901 GND.n900 341.085
R1498 GND.n911 GND.n910 341.085
R1499 GND.n920 GND.n861 341.085
R1500 GND.n921 GND.n920 341.085
R1501 GND.n922 GND.n921 341.085
R1502 GND.n930 GND.n855 341.085
R1503 GND.n982 GND.n981 341.085
R1504 GND.n990 GND.n822 341.085
R1505 GND.n992 GND.n991 341.085
R1506 GND.n1001 GND.n816 341.085
R1507 GND.n1002 GND.n1001 341.085
R1508 GND.n1003 GND.n1002 341.085
R1509 GND.n1014 GND.n810 341.085
R1510 GND.n1017 GND.n1016 341.085
R1511 GND.n1027 GND.n1026 341.085
R1512 GND.n1029 GND.n1027 341.085
R1513 GND.n1029 GND.n1028 341.085
R1514 GND.n1038 GND.n1037 341.085
R1515 GND.n1040 GND.n1039 341.085
R1516 GND.n1050 GND.n1049 341.085
R1517 GND.n683 GND.n682 341.085
R1518 GND.n685 GND.n683 341.085
R1519 GND.n685 GND.n684 341.085
R1520 GND.n695 GND.n694 341.085
R1521 GND.n705 GND.n578 341.085
R1522 GND.n707 GND.n706 341.085
R1523 GND.n707 GND.n572 341.085
R1524 GND.n715 GND.n572 341.085
R1525 GND.n629 GND.n628 341.085
R1526 GND.n630 GND.n615 341.085
R1527 GND.n639 GND.n615 341.085
R1528 GND.n640 GND.n639 341.085
R1529 GND.n642 GND.n641 341.085
R1530 GND.n652 GND.n651 341.085
R1531 GND.n661 GND.n602 341.085
R1532 GND.n662 GND.n661 341.085
R1533 GND.n663 GND.n662 341.085
R1534 GND.n671 GND.n596 341.085
R1535 GND.n723 GND.n722 341.085
R1536 GND.n731 GND.n563 341.085
R1537 GND.n733 GND.n732 341.085
R1538 GND.n742 GND.n557 341.085
R1539 GND.n743 GND.n742 341.085
R1540 GND.n744 GND.n743 341.085
R1541 GND.n755 GND.n551 341.085
R1542 GND.n758 GND.n757 341.085
R1543 GND.n768 GND.n767 341.085
R1544 GND.n770 GND.n768 341.085
R1545 GND.n770 GND.n769 341.085
R1546 GND.n779 GND.n778 341.085
R1547 GND.n781 GND.n780 341.085
R1548 GND.n791 GND.n790 341.085
R1549 GND.n941 GND.t163 319.767
R1550 GND.n955 GND.t95 319.767
R1551 GND.n955 GND.t77 319.767
R1552 GND.t239 GND.n974 319.767
R1553 GND.n889 GND.t76 319.767
R1554 GND.n909 GND.t260 319.767
R1555 GND.t85 GND.n909 319.767
R1556 GND.n922 GND.t50 319.767
R1557 GND.t73 GND.n816 319.767
R1558 GND.n1015 GND.t37 319.767
R1559 GND.t35 GND.n1015 319.767
R1560 GND.n1028 GND.t160 319.767
R1561 GND.n682 GND.t53 319.767
R1562 GND.n696 GND.t152 319.767
R1563 GND.n696 GND.t21 319.767
R1564 GND.t39 GND.n715 319.767
R1565 GND.n630 GND.t23 319.767
R1566 GND.n650 GND.t128 319.767
R1567 GND.t0 GND.n650 319.767
R1568 GND.n663 GND.t79 319.767
R1569 GND.t62 GND.n557 319.767
R1570 GND.n756 GND.t88 319.767
R1571 GND.t57 GND.n756 319.767
R1572 GND.n769 GND.t63 319.767
R1573 GND.n953 GND.t211 277.131
R1574 GND.t185 GND.n964 277.131
R1575 GND.n887 GND.t140 277.131
R1576 GND.n901 GND.t266 277.131
R1577 GND.n911 GND.t16 277.131
R1578 GND.t97 GND.n930 277.131
R1579 GND.n991 GND.t56 277.131
R1580 GND.t183 GND.n810 277.131
R1581 GND.n1016 GND.t187 277.131
R1582 GND.t87 GND.n1038 277.131
R1583 GND.n694 GND.t194 277.131
R1584 GND.t173 GND.n705 277.131
R1585 GND.n628 GND.t121 277.131
R1586 GND.n642 GND.t116 277.131
R1587 GND.n652 GND.t148 277.131
R1588 GND.t154 GND.n671 277.131
R1589 GND.n732 GND.t52 277.131
R1590 GND.t192 GND.n551 277.131
R1591 GND.n757 GND.t200 277.131
R1592 GND.t161 GND.n779 277.131
R1593 GND.n273 GND.t259 269.289
R1594 GND.n171 GND.t170 269.289
R1595 GND.n1675 GND.n1449 261.515
R1596 GND.n1676 GND.n1675 261.515
R1597 GND.n1677 GND.n1676 261.515
R1598 GND.n1686 GND.n1443 261.515
R1599 GND.n1687 GND.n1686 261.515
R1600 GND.n1688 GND.n1687 261.515
R1601 GND.n1688 GND.n1437 261.515
R1602 GND.n1697 GND.n1437 261.515
R1603 GND.n1698 GND.n1697 261.515
R1604 GND.n1699 GND.n1698 261.515
R1605 GND.n1707 GND.n1430 261.515
R1606 GND.n1708 GND.n1707 261.515
R1607 GND.n1718 GND.n1423 261.515
R1608 GND.n1719 GND.n1718 261.515
R1609 GND.n1720 GND.n1417 261.515
R1610 GND.n1729 GND.n1417 261.515
R1611 GND.n1730 GND.n1729 261.515
R1612 GND.n1731 GND.n1411 261.515
R1613 GND.n1740 GND.n1411 261.515
R1614 GND.n1741 GND.n1740 261.515
R1615 GND.n1742 GND.n1741 261.515
R1616 GND.n1742 GND.n1404 261.515
R1617 GND.n1753 GND.n1404 261.515
R1618 GND.n1709 GND.t236 250
R1619 GND.n1460 GND.n1449 235.364
R1620 GND.t106 GND.n822 234.496
R1621 GND.n1039 GND.t92 234.496
R1622 GND.t12 GND.n563 234.496
R1623 GND.n780 GND.t60 234.496
R1624 GND.n1561 GND.n1515 233.453
R1625 GND.n1563 GND.n1562 233.453
R1626 GND.n1572 GND.n1509 233.453
R1627 GND.n1582 GND.n1503 233.453
R1628 GND.n1592 GND.n1496 233.453
R1629 GND.n1594 GND.n1593 233.453
R1630 GND.n1602 GND.n1489 233.453
R1631 GND.n1612 GND.n1484 233.453
R1632 GND.n1623 GND.n1478 233.453
R1633 GND.n1625 GND.n1624 233.453
R1634 GND.n1633 GND.n1472 233.453
R1635 GND.t168 GND.n1443 228.826
R1636 GND.t242 GND.n1423 228.826
R1637 GND.t155 GND.n1719 228.826
R1638 GND.n1540 GND.n1526 221.582
R1639 GND.n1646 GND.n1459 221.582
R1640 GND.n1551 GND.t34 217.625
R1641 GND.n1635 GND.t2 217.625
R1642 GND.n1553 GND.t75 213.669
R1643 GND.n1584 GND.t126 213.669
R1644 GND.t104 GND.n1603 213.669
R1645 GND.t157 GND.n1634 213.669
R1646 GND.n1203 GND.t308 192.984
R1647 GND.n1250 GND.t81 192.984
R1648 GND.n1143 GND.t71 192.984
R1649 GND.n1313 GND.t143 192.984
R1650 GND.n981 GND.t69 191.86
R1651 GND.t162 GND.n1050 191.86
R1652 GND.n722 GND.t59 191.86
R1653 GND.t72 GND.n791 191.86
R1654 GND.n1543 GND.t130 174.1
R1655 GND.n1574 GND.t32 174.1
R1656 GND.t233 GND.n1613 174.1
R1657 GND.t123 GND.n1645 174.1
R1658 GND.t306 GND.n1430 163.447
R1659 GND.t244 GND.n1730 163.447
R1660 GND.n1897 GND.n1896 163.19
R1661 GND.n1772 GND.n1771 162.23
R1662 GND.n1782 GND.n1781 162.23
R1663 GND.n1792 GND.n1791 162.23
R1664 GND.n1802 GND.n1801 162.23
R1665 GND.n1803 GND.n1370 162.23
R1666 GND.n1814 GND.n1813 162.23
R1667 GND.n1824 GND.n1823 162.23
R1668 GND.n1835 GND.n1350 162.23
R1669 GND.n1845 GND.n1344 162.23
R1670 GND.n1856 GND.n1855 162.23
R1671 GND.n1857 GND.n1338 162.23
R1672 GND.n1867 GND.n1332 162.23
R1673 GND.n1877 GND.n1326 162.23
R1674 GND.n1887 GND.n1319 162.23
R1675 GND.n433 GND.t164 158.378
R1676 GND.n533 GND.t111 158.378
R1677 GND.t69 GND.n980 158.378
R1678 GND.n1051 GND.t162 158.378
R1679 GND.t59 GND.n721 158.378
R1680 GND.n792 GND.t72 158.378
R1681 GND.n1756 GND.n1403 157.6
R1682 GND.n1532 GND.n1527 157.6
R1683 GND.n1212 GND.n1107 157.6
R1684 GND.n1212 GND.n1106 157.6
R1685 GND.n1217 GND.n1106 157.6
R1686 GND.n1217 GND.n1102 157.6
R1687 GND.n1224 GND.n1102 157.6
R1688 GND.n1224 GND.n1101 157.6
R1689 GND.n1228 GND.n1101 157.6
R1690 GND.n1228 GND.n1096 157.6
R1691 GND.n1235 GND.n1096 157.6
R1692 GND.n1235 GND.n1094 157.6
R1693 GND.n1239 GND.n1094 157.6
R1694 GND.n1239 GND.n1090 157.6
R1695 GND.n1245 GND.n1090 157.6
R1696 GND.n1245 GND.n1088 157.6
R1697 GND.n1147 GND.n1141 157.6
R1698 GND.n1147 GND.n1140 157.6
R1699 GND.n1152 GND.n1140 157.6
R1700 GND.n1152 GND.n1136 157.6
R1701 GND.n1158 GND.n1136 157.6
R1702 GND.n1158 GND.n1135 157.6
R1703 GND.n1163 GND.n1135 157.6
R1704 GND.n1163 GND.n1131 157.6
R1705 GND.n1170 GND.n1131 157.6
R1706 GND.n1170 GND.n1130 157.6
R1707 GND.n1174 GND.n1130 157.6
R1708 GND.n1174 GND.n1125 157.6
R1709 GND.n1181 GND.n1125 157.6
R1710 GND.n1181 GND.n1123 157.6
R1711 GND.n1185 GND.n1123 157.6
R1712 GND.n1185 GND.n1119 157.6
R1713 GND.n1191 GND.n1119 157.6
R1714 GND.n1191 GND.n1117 157.6
R1715 GND.n1195 GND.n1117 157.6
R1716 GND.n1195 GND.n1113 157.6
R1717 GND.n1201 GND.n1113 157.6
R1718 GND.n1201 GND.n1111 157.6
R1719 GND.n1256 GND.n1084 157.6
R1720 GND.n1256 GND.n1083 157.6
R1721 GND.n1261 GND.n1083 157.6
R1722 GND.n1261 GND.n1079 157.6
R1723 GND.n1267 GND.n1079 157.6
R1724 GND.n1267 GND.n1078 157.6
R1725 GND.n1272 GND.n1078 157.6
R1726 GND.n1272 GND.n1074 157.6
R1727 GND.n1279 GND.n1074 157.6
R1728 GND.n1279 GND.n1073 157.6
R1729 GND.n1283 GND.n1073 157.6
R1730 GND.n1283 GND.n1068 157.6
R1731 GND.n1290 GND.n1068 157.6
R1732 GND.n1290 GND.n1066 157.6
R1733 GND.n1294 GND.n1066 157.6
R1734 GND.n1294 GND.n1062 157.6
R1735 GND.n1300 GND.n1062 157.6
R1736 GND.n1300 GND.n1060 157.6
R1737 GND.n1304 GND.n1060 157.6
R1738 GND.n1304 GND.n1056 157.6
R1739 GND.n1311 GND.n1056 157.6
R1740 GND.n1311 GND.n1054 157.6
R1741 GND.n940 GND.n850 157.6
R1742 GND.n940 GND.n849 157.6
R1743 GND.n945 GND.n849 157.6
R1744 GND.n945 GND.n845 157.6
R1745 GND.n952 GND.n845 157.6
R1746 GND.n952 GND.n844 157.6
R1747 GND.n956 GND.n844 157.6
R1748 GND.n956 GND.n838 157.6
R1749 GND.n963 GND.n838 157.6
R1750 GND.n963 GND.n836 157.6
R1751 GND.n967 GND.n836 157.6
R1752 GND.n967 GND.n832 157.6
R1753 GND.n973 GND.n832 157.6
R1754 GND.n973 GND.n830 157.6
R1755 GND.n886 GND.n880 157.6
R1756 GND.n886 GND.n879 157.6
R1757 GND.n890 GND.n879 157.6
R1758 GND.n890 GND.n875 157.6
R1759 GND.n897 GND.n875 157.6
R1760 GND.n897 GND.n873 157.6
R1761 GND.n902 GND.n873 157.6
R1762 GND.n902 GND.n867 157.6
R1763 GND.n908 GND.n867 157.6
R1764 GND.n908 GND.n866 157.6
R1765 GND.n912 GND.n866 157.6
R1766 GND.n912 GND.n862 157.6
R1767 GND.n919 GND.n862 157.6
R1768 GND.n919 GND.n860 157.6
R1769 GND.n923 GND.n860 157.6
R1770 GND.n923 GND.n856 157.6
R1771 GND.n929 GND.n856 157.6
R1772 GND.n929 GND.n854 157.6
R1773 GND.n980 GND.n827 157.6
R1774 GND.n983 GND.n827 157.6
R1775 GND.n983 GND.n823 157.6
R1776 GND.n989 GND.n823 157.6
R1777 GND.n989 GND.n821 157.6
R1778 GND.n993 GND.n821 157.6
R1779 GND.n993 GND.n817 157.6
R1780 GND.n1000 GND.n817 157.6
R1781 GND.n1000 GND.n815 157.6
R1782 GND.n1004 GND.n815 157.6
R1783 GND.n1004 GND.n811 157.6
R1784 GND.n1013 GND.n811 157.6
R1785 GND.n1013 GND.n809 157.6
R1786 GND.n1018 GND.n809 157.6
R1787 GND.n1018 GND.n806 157.6
R1788 GND.n1025 GND.n806 157.6
R1789 GND.n1025 GND.n805 157.6
R1790 GND.n1030 GND.n805 157.6
R1791 GND.n1030 GND.n801 157.6
R1792 GND.n1036 GND.n801 157.6
R1793 GND.n1036 GND.n800 157.6
R1794 GND.n1041 GND.n800 157.6
R1795 GND.n1041 GND.n796 157.6
R1796 GND.n1048 GND.n796 157.6
R1797 GND.n1048 GND.n795 157.6
R1798 GND.n1051 GND.n795 157.6
R1799 GND.n681 GND.n591 157.6
R1800 GND.n681 GND.n590 157.6
R1801 GND.n686 GND.n590 157.6
R1802 GND.n686 GND.n586 157.6
R1803 GND.n693 GND.n586 157.6
R1804 GND.n693 GND.n585 157.6
R1805 GND.n697 GND.n585 157.6
R1806 GND.n697 GND.n579 157.6
R1807 GND.n704 GND.n579 157.6
R1808 GND.n704 GND.n577 157.6
R1809 GND.n708 GND.n577 157.6
R1810 GND.n708 GND.n573 157.6
R1811 GND.n714 GND.n573 157.6
R1812 GND.n714 GND.n571 157.6
R1813 GND.n627 GND.n621 157.6
R1814 GND.n627 GND.n620 157.6
R1815 GND.n631 GND.n620 157.6
R1816 GND.n631 GND.n616 157.6
R1817 GND.n638 GND.n616 157.6
R1818 GND.n638 GND.n614 157.6
R1819 GND.n643 GND.n614 157.6
R1820 GND.n643 GND.n608 157.6
R1821 GND.n649 GND.n608 157.6
R1822 GND.n649 GND.n607 157.6
R1823 GND.n653 GND.n607 157.6
R1824 GND.n653 GND.n603 157.6
R1825 GND.n660 GND.n603 157.6
R1826 GND.n660 GND.n601 157.6
R1827 GND.n664 GND.n601 157.6
R1828 GND.n664 GND.n597 157.6
R1829 GND.n670 GND.n597 157.6
R1830 GND.n670 GND.n595 157.6
R1831 GND.n721 GND.n568 157.6
R1832 GND.n724 GND.n568 157.6
R1833 GND.n724 GND.n564 157.6
R1834 GND.n730 GND.n564 157.6
R1835 GND.n730 GND.n562 157.6
R1836 GND.n734 GND.n562 157.6
R1837 GND.n734 GND.n558 157.6
R1838 GND.n741 GND.n558 157.6
R1839 GND.n741 GND.n556 157.6
R1840 GND.n745 GND.n556 157.6
R1841 GND.n745 GND.n552 157.6
R1842 GND.n754 GND.n552 157.6
R1843 GND.n754 GND.n550 157.6
R1844 GND.n759 GND.n550 157.6
R1845 GND.n759 GND.n547 157.6
R1846 GND.n766 GND.n547 157.6
R1847 GND.n766 GND.n546 157.6
R1848 GND.n771 GND.n546 157.6
R1849 GND.n771 GND.n542 157.6
R1850 GND.n777 GND.n542 157.6
R1851 GND.n777 GND.n541 157.6
R1852 GND.n782 GND.n541 157.6
R1853 GND.n782 GND.n537 157.6
R1854 GND.n789 GND.n537 157.6
R1855 GND.n789 GND.n536 157.6
R1856 GND.n792 GND.n536 157.6
R1857 GND.n1763 GND.n1395 156.724
R1858 GND.n1771 GND.n1394 154.316
R1859 GND.n1781 GND.n1388 154.316
R1860 GND.n1791 GND.n1382 154.316
R1861 GND.n1801 GND.n1376 154.316
R1862 GND.n1803 GND.n1802 154.316
R1863 GND.n1813 GND.n1370 154.316
R1864 GND.n1823 GND.n1364 154.316
R1865 GND.n1833 GND.n1356 154.316
R1866 GND.n1843 GND.n1350 154.316
R1867 GND.n1855 GND.n1344 154.316
R1868 GND.n1857 GND.n1856 154.316
R1869 GND.n1865 GND.n1338 154.316
R1870 GND.n1875 GND.n1332 154.316
R1871 GND.n1885 GND.n1326 154.316
R1872 GND.n1895 GND.n1319 154.316
R1873 GND.n1752 GND.n1403 148.783
R1874 GND.n1667 GND.n1450 148.783
R1875 GND.n1896 GND.t54 147.437
R1876 GND.t300 GND.n1376 142.446
R1877 GND.t67 GND.n1356 142.446
R1878 GND.t135 GND.n1833 142.446
R1879 GND.t284 GND.n1865 142.446
R1880 GND.n1144 GND.n1143 135.387
R1881 GND.n1793 GND.t131 134.532
R1882 GND.n1825 GND.t278 134.532
R1883 GND.t166 GND.n1834 134.532
R1884 GND.t253 GND.n1866 134.532
R1885 GND.n268 GND.t122 133.857
R1886 GND.n178 GND.t311 133.857
R1887 GND.n1207 GND.n1206 132.648
R1888 GND.n1314 GND.n1313 132.648
R1889 GND.n1248 GND.n1247 132.647
R1890 GND.n1204 GND.n1203 132.647
R1891 GND.n1251 GND.n1250 132.647
R1892 GND.n1709 GND.n1708 130.757
R1893 GND.n1710 GND.n1709 130.757
R1894 GND.n1658 GND.n1458 122.642
R1895 GND.n883 GND.n882 118.662
R1896 GND.n624 GND.n623 118.662
R1897 GND.n935 GND.n934 115.922
R1898 GND.n676 GND.n675 115.922
R1899 GND.n976 GND.n975 115.922
R1900 GND.n932 GND.n931 115.922
R1901 GND.n717 GND.n716 115.922
R1902 GND.n673 GND.n672 115.922
R1903 GND.n1215 GND.t293 111.486
R1904 GND.n1237 GND.t303 111.486
R1905 GND.t262 GND.n1149 111.486
R1906 GND.n1161 GND.t231 111.486
R1907 GND.n1183 GND.t316 111.486
R1908 GND.t84 GND.n1112 111.486
R1909 GND.t112 GND.n1258 111.486
R1910 GND.n1270 GND.t189 111.486
R1911 GND.n1292 GND.t177 111.486
R1912 GND.t310 GND.n1055 111.486
R1913 GND.n440 GND.t61 106.589
R1914 GND.n528 GND.t91 106.589
R1915 GND.n982 GND.t106 106.589
R1916 GND.n1049 GND.t92 106.589
R1917 GND.n723 GND.t12 106.589
R1918 GND.n790 GND.t60 106.589
R1919 GND.t145 GND.n1382 102.877
R1920 GND.t202 GND.n1364 102.877
R1921 GND.t215 GND.n1843 102.877
R1922 GND.t11 GND.n1875 102.877
R1923 GND.t146 GND.n1772 98.92
R1924 GND.n1773 GND.t258 98.92
R1925 GND.n1886 GND.t141 98.92
R1926 GND.n1887 GND.t46 98.92
R1927 GND.n1699 GND.t306 98.068
R1928 GND.n1731 GND.t244 98.068
R1929 GND.n1783 GND.t94 94.964
R1930 GND.n1815 GND.t175 94.964
R1931 GND.t220 GND.n1844 94.964
R1932 GND.t288 GND.n1876 94.964
R1933 GND.n1541 GND.n1540 83.093
R1934 GND.n1543 GND.n1542 83.093
R1935 GND.n1552 GND.n1551 83.093
R1936 GND.n1562 GND.n1561 83.093
R1937 GND.n1573 GND.n1572 83.093
R1938 GND.n1574 GND.n1503 83.093
R1939 GND.n1583 GND.n1582 83.093
R1940 GND.n1604 GND.n1484 83.093
R1941 GND.n1613 GND.n1612 83.093
R1942 GND.n1614 GND.n1478 83.093
R1943 GND.n1625 GND.n1472 83.093
R1944 GND.n1636 GND.n1635 83.093
R1945 GND.n1645 GND.n1644 83.093
R1946 GND.n1647 GND.n1646 83.093
R1947 GND.n1657 GND.n1461 81.207
R1948 GND.n1539 GND.n1527 81.207
R1949 GND.n9 GND.t29 70.155
R1950 GND.n83 GND.t115 70.155
R1951 GND.n91 GND.t51 70.155
R1952 GND.n165 GND.t147 70.155
R1953 GND.n363 GND.t25 70.155
R1954 GND.n931 GND.t97 70.155
R1955 GND.n672 GND.t154 70.155
R1956 GND.n291 GND.t256 70.155
R1957 GND.n882 GND.t140 70.155
R1958 GND.n623 GND.t121 70.155
R1959 GND.n1399 GND.n1394 67.266
R1960 GND.n1544 GND.n1525 64.572
R1961 GND.n1550 GND.n1521 64.572
R1962 GND.n1554 GND.n1520 64.572
R1963 GND.n1560 GND.n1516 64.572
R1964 GND.n1564 GND.n1514 64.572
R1965 GND.n1571 GND.n1510 64.572
R1966 GND.n1575 GND.n1508 64.572
R1967 GND.n1581 GND.n1504 64.572
R1968 GND.n1585 GND.n1502 64.572
R1969 GND.n1591 GND.n1497 64.572
R1970 GND.n1595 GND.n1495 64.572
R1971 GND.n1601 GND.n1490 64.572
R1972 GND.n1605 GND.n1488 64.572
R1973 GND.n1611 GND.n1485 64.572
R1974 GND.n1615 GND.n1483 64.572
R1975 GND.n1622 GND.n1479 64.572
R1976 GND.n1626 GND.n1477 64.572
R1977 GND.n1632 GND.n1473 64.572
R1978 GND.n1637 GND.n1471 64.572
R1979 GND.n1643 GND.n1467 64.572
R1980 GND.n1648 GND.n1466 64.572
R1981 GND.n186 GND.t93 63.953
R1982 GND.n211 GND.t206 63.953
R1983 GND.n235 GND.t213 63.953
R1984 GND.n260 GND.t55 63.953
R1985 GND.n34 GND.t295 63.953
R1986 GND.n58 GND.t30 63.953
R1987 GND.n116 GND.t196 63.953
R1988 GND.n140 GND.t150 63.953
R1989 GND.n388 GND.t179 63.953
R1990 GND.n410 GND.t204 63.953
R1991 GND.n316 GND.t118 63.953
R1992 GND.n338 GND.t269 63.953
R1993 GND.n448 GND.t41 63.953
R1994 GND.n473 GND.t181 63.953
R1995 GND.n495 GND.t198 63.953
R1996 GND.n520 GND.t165 63.953
R1997 GND.n943 GND.t211 63.953
R1998 GND.n965 GND.t185 63.953
R1999 GND.t266 GND.n899 63.953
R2000 GND.t16 GND.n861 63.953
R2001 GND.t56 GND.n990 63.953
R2002 GND.n1003 GND.t183 63.953
R2003 GND.n1026 GND.t187 63.953
R2004 GND.n1040 GND.t87 63.953
R2005 GND.n684 GND.t194 63.953
R2006 GND.n706 GND.t173 63.953
R2007 GND.t116 GND.n640 63.953
R2008 GND.t148 GND.n602 63.953
R2009 GND.t52 GND.n731 63.953
R2010 GND.n744 GND.t192 63.953
R2011 GND.n767 GND.t200 63.953
R2012 GND.n781 GND.t161 63.953
R2013 GND.t241 GND.n1509 63.309
R2014 GND.t19 GND.n1592 63.309
R2015 GND.t313 GND.n1489 63.309
R2016 GND.t230 GND.n1623 63.309
R2017 GND.t258 GND.n1388 63.309
R2018 GND.t141 GND.n1885 63.309
R2019 GND.t130 GND.n1541 59.352
R2020 GND.n1553 GND.t272 59.352
R2021 GND.t32 GND.n1573 59.352
R2022 GND.n1584 GND.t44 59.352
R2023 GND.n1603 GND.t42 59.352
R2024 GND.n1614 GND.t233 59.352
R2025 GND.n1634 GND.t282 59.352
R2026 GND.n1647 GND.t123 59.352
R2027 GND.t94 GND.n1782 59.352
R2028 GND.n1783 GND.t145 59.352
R2029 GND.t175 GND.n1814 59.352
R2030 GND.n1815 GND.t202 59.352
R2031 GND.n1844 GND.t215 59.352
R2032 GND.n1845 GND.t220 59.352
R2033 GND.n1876 GND.t11 59.352
R2034 GND.n1877 GND.t288 59.352
R2035 GND.n1773 GND.t146 55.395
R2036 GND.t46 GND.n1886 55.395
R2037 EESPFAL_s3_0/GND GND.n1314 48.86
R2038 GND.n1894 GND.n1318 45.747
R2039 GND.n1770 GND.n1393 44.872
R2040 GND.n1774 GND.n1389 44.872
R2041 GND.n1780 GND.n1387 44.872
R2042 GND.n1784 GND.n1383 44.872
R2043 GND.n1790 GND.n1381 44.872
R2044 GND.n1794 GND.n1377 44.872
R2045 GND.n1800 GND.n1375 44.872
R2046 GND.n1804 GND.n1371 44.872
R2047 GND.n1812 GND.n1369 44.872
R2048 GND.n1816 GND.n1365 44.872
R2049 GND.n1822 GND.n1363 44.872
R2050 GND.n1826 GND.n1357 44.872
R2051 GND.n1832 GND.n1355 44.872
R2052 GND.n1836 GND.n1351 44.872
R2053 GND.n1842 GND.n1349 44.872
R2054 GND.n1846 GND.n1345 44.872
R2055 GND.n1854 GND.n1343 44.872
R2056 GND.n1858 GND.n1339 44.872
R2057 GND.n1864 GND.n1337 44.872
R2058 GND.n1868 GND.n1333 44.872
R2059 GND.n1874 GND.n1331 44.872
R2060 GND.n1878 GND.n1327 44.872
R2061 GND.n1884 GND.n1325 44.872
R2062 GND.n1888 GND.n1320 44.872
R2063 GND.n1247 GND.t252 44.336
R2064 GND.n1206 GND.t249 44.336
R2065 GND.n1674 GND.n1450 43.535
R2066 GND.n1674 GND.n1448 43.535
R2067 GND.n1678 GND.n1448 43.535
R2068 GND.n1678 GND.n1444 43.535
R2069 GND.n1685 GND.n1444 43.535
R2070 GND.n1685 GND.n1442 43.535
R2071 GND.n1689 GND.n1442 43.535
R2072 GND.n1689 GND.n1438 43.535
R2073 GND.n1696 GND.n1438 43.535
R2074 GND.n1696 GND.n1436 43.535
R2075 GND.n1700 GND.n1436 43.535
R2076 GND.n1700 GND.n1431 43.535
R2077 GND.n1706 GND.n1431 43.535
R2078 GND.n1706 GND.n1429 43.535
R2079 GND.n1711 GND.n1429 43.535
R2080 GND.n1711 GND.n1424 43.535
R2081 GND.n1717 GND.n1424 43.535
R2082 GND.n1717 GND.n1422 43.535
R2083 GND.n1721 GND.n1422 43.535
R2084 GND.n1721 GND.n1418 43.535
R2085 GND.n1728 GND.n1418 43.535
R2086 GND.n1728 GND.n1416 43.535
R2087 GND.n1732 GND.n1416 43.535
R2088 GND.n1732 GND.n1412 43.535
R2089 GND.n1739 GND.n1412 43.535
R2090 GND.n1739 GND.n1410 43.535
R2091 GND.n1743 GND.n1410 43.535
R2092 GND.n1743 GND.n1405 43.535
R2093 GND.n1752 GND.n1405 43.535
R2094 GND.n1770 GND.n1395 42.683
R2095 GND.n1774 GND.n1393 42.683
R2096 GND.n1780 GND.n1389 42.683
R2097 GND.n1784 GND.n1387 42.683
R2098 GND.n1790 GND.n1383 42.683
R2099 GND.n1794 GND.n1381 42.683
R2100 GND.n1800 GND.n1377 42.683
R2101 GND.n1804 GND.n1375 42.683
R2102 GND.n1812 GND.n1371 42.683
R2103 GND.n1816 GND.n1369 42.683
R2104 GND.n1822 GND.n1365 42.683
R2105 GND.n1826 GND.n1363 42.683
R2106 GND.n1832 GND.n1357 42.683
R2107 GND.n1836 GND.n1355 42.683
R2108 GND.n1842 GND.n1351 42.683
R2109 GND.n1846 GND.n1349 42.683
R2110 GND.n1854 GND.n1345 42.683
R2111 GND.n1858 GND.n1343 42.683
R2112 GND.n1864 GND.n1339 42.683
R2113 GND.n1868 GND.n1337 42.683
R2114 GND.n1874 GND.n1333 42.683
R2115 GND.n1878 GND.n1331 42.683
R2116 GND.n1884 GND.n1327 42.683
R2117 GND.n1888 GND.n1325 42.683
R2118 GND.n1894 GND.n1320 42.683
R2119 GND.n1316 GND.n793 37.93
R2120 GND.t298 GND.n1226 37.162
R2121 GND.t6 GND.n1095 37.162
R2122 GND.n1150 GND.t158 37.162
R2123 GND.t285 GND.n1172 37.162
R2124 GND.t48 GND.n1124 37.162
R2125 GND.n1193 GND.t312 37.162
R2126 GND.n1259 GND.t70 37.162
R2127 GND.t250 GND.n1281 37.162
R2128 GND.t247 GND.n1067 37.162
R2129 GND.n1302 GND.t90 37.162
R2130 GND.n1677 GND.t168 32.689
R2131 GND.n1710 GND.t242 32.689
R2132 GND.n1720 GND.t155 32.689
R2133 GND.n1754 GND.t66 32.689
R2134 GND.n275 GND.n274 31.53
R2135 GND.n1899 GND.n534 31.53
R2136 GND.n1315 GND.n1052 31.53
R2137 GND.n33 GND.t296 29.103
R2138 GND.n62 GND.t271 29.103
R2139 GND.n115 GND.t197 29.103
R2140 GND.n144 GND.t225 29.103
R2141 GND.n210 GND.t223 29.103
R2142 GND.n239 GND.t214 29.103
R2143 GND.n315 GND.t119 29.103
R2144 GND.n342 GND.t302 29.103
R2145 GND.n387 GND.t180 29.103
R2146 GND.n414 GND.t205 29.103
R2147 GND.n472 GND.t182 29.103
R2148 GND.n499 GND.t199 29.103
R2149 GND.n1809 GND.t203 29.103
R2150 GND.n1851 GND.t221 29.103
R2151 GND.n1693 GND.t307 29.103
R2152 GND.n1736 GND.t245 29.103
R2153 GND.n1500 GND.t45 29.103
R2154 GND.n1619 GND.t234 29.103
R2155 GND.n1166 GND.t232 29.103
R2156 GND.n1121 GND.t317 29.103
R2157 GND.n1220 GND.t294 29.103
R2158 GND.n1092 GND.t304 29.103
R2159 GND.n1275 GND.t190 29.103
R2160 GND.n1064 GND.t178 29.103
R2161 GND.n894 GND.t290 29.103
R2162 GND.n916 GND.t17 29.103
R2163 GND.n948 GND.t218 29.103
R2164 GND.n834 GND.t191 29.103
R2165 GND.n813 GND.t222 29.103
R2166 GND.n1022 GND.t188 29.103
R2167 GND.n635 GND.t268 29.103
R2168 GND.n657 GND.t277 29.103
R2169 GND.n689 GND.t217 29.103
R2170 GND.n575 GND.t209 29.103
R2171 GND.n554 GND.t193 29.103
R2172 GND.n763 GND.t226 29.103
R2173 GND.n33 GND.t315 29.102
R2174 GND.n62 GND.t31 29.102
R2175 GND.n115 GND.t305 29.102
R2176 GND.n144 GND.t151 29.102
R2177 GND.n210 GND.t207 29.102
R2178 GND.n239 GND.t219 29.102
R2179 GND.n315 GND.t246 29.102
R2180 GND.n342 GND.t270 29.102
R2181 GND.n387 GND.t210 29.102
R2182 GND.n414 GND.t229 29.102
R2183 GND.n472 GND.t208 29.102
R2184 GND.n499 GND.t227 29.102
R2185 GND.n1849 GND.t216 29.102
R2186 GND.n1808 GND.t176 29.102
R2187 GND.n1724 GND.t292 29.102
R2188 GND.n1682 GND.t276 29.102
R2189 GND.n1607 GND.t43 29.102
R2190 GND.n1568 GND.t33 29.102
R2191 GND.n894 GND.t267 29.102
R2192 GND.n916 GND.t18 29.102
R2193 GND.n948 GND.t212 29.102
R2194 GND.n834 GND.t186 29.102
R2195 GND.n813 GND.t184 29.102
R2196 GND.n1022 GND.t228 29.102
R2197 GND.n635 GND.t117 29.102
R2198 GND.n657 GND.t149 29.102
R2199 GND.n689 GND.t195 29.102
R2200 GND.n575 GND.t174 29.102
R2201 GND.n554 GND.t224 29.102
R2202 GND.n763 GND.t201 29.102
R2203 GND.n427 GND.t142 27.519
R2204 GND.n975 GND.t239 27.519
R2205 GND.n716 GND.t39 27.519
R2206 GND.n371 GND.t238 27.519
R2207 GND.n934 GND.t163 27.519
R2208 GND.n675 GND.t53 27.519
R2209 GND.n4 GND.t254 24
R2210 GND.n4 GND.t28 24
R2211 GND.n3 GND.t133 24
R2212 GND.n3 GND.t264 24
R2213 GND.n8 GND.t65 24
R2214 GND.n8 GND.t83 24
R2215 GND.n7 GND.t240 24
R2216 GND.n7 GND.t114 24
R2217 GND.n6 GND.t172 24
R2218 GND.n6 GND.t281 24
R2219 GND.n5 GND.t297 24
R2220 GND.n5 GND.t138 24
R2221 GND.n282 GND.t10 24
R2222 GND.n282 GND.t255 24
R2223 GND.n281 GND.t74 24
R2224 GND.n281 GND.t109 24
R2225 GND.n286 GND.t263 24
R2226 GND.n286 GND.t24 24
R2227 GND.n285 GND.t102 24
R2228 GND.n285 GND.t5 24
R2229 GND.n290 GND.t274 24
R2230 GND.n290 GND.t124 24
R2231 GND.n289 GND.t287 24
R2232 GND.n289 GND.t14 24
R2233 GND.n1360 GND.t279 24
R2234 GND.n1360 GND.t136 24
R2235 GND.n1359 GND.t68 24
R2236 GND.n1359 GND.t167 24
R2237 GND.n1433 GND.t100 24
R2238 GND.n1433 GND.t237 24
R2239 GND.n1426 GND.t243 24
R2240 GND.n1426 GND.t156 24
R2241 GND.n1499 GND.t127 24
R2242 GND.n1499 GND.t20 24
R2243 GND.n1492 GND.t314 24
R2244 GND.n1492 GND.t105 24
R2245 GND.n1070 GND.t251 24
R2246 GND.n1070 GND.t248 24
R2247 GND.n1098 GND.t299 24
R2248 GND.n1098 GND.t7 24
R2249 GND.n1127 GND.t286 24
R2250 GND.n1127 GND.t49 24
R2251 GND.n1009 GND.t107 24
R2252 GND.n1009 GND.t169 24
R2253 GND.n1008 GND.t38 24
R2254 GND.n1008 GND.t36 24
R2255 GND.n841 GND.t98 24
R2256 GND.n841 GND.t78 24
R2257 GND.n840 GND.t96 24
R2258 GND.n840 GND.t159 24
R2259 GND.n870 GND.t261 24
R2260 GND.n870 GND.t86 24
R2261 GND.n869 GND.t289 24
R2262 GND.n869 GND.t309 24
R2263 GND.n750 GND.t89 24
R2264 GND.n750 GND.t58 24
R2265 GND.n749 GND.t103 24
R2266 GND.n749 GND.t120 24
R2267 GND.n582 GND.t153 24
R2268 GND.n582 GND.t22 24
R2269 GND.n581 GND.t235 24
R2270 GND.n581 GND.t125 24
R2271 GND.n611 GND.t301 24
R2272 GND.n611 GND.t1 24
R2273 GND.n610 GND.t129 24
R2274 GND.n610 GND.t283 24
R2275 GND.t272 GND.n1515 23.741
R2276 GND.t44 GND.n1496 23.741
R2277 GND.t42 GND.n1602 23.741
R2278 GND.t282 GND.n1633 23.741
R2279 GND.t54 GND.n1895 23.741
R2280 GND.n1539 GND.n1525 22.983
R2281 GND.n1544 GND.n1521 22.983
R2282 GND.n1550 GND.n1520 22.983
R2283 GND.n1554 GND.n1516 22.983
R2284 GND.n1560 GND.n1514 22.983
R2285 GND.n1564 GND.n1510 22.983
R2286 GND.n1571 GND.n1508 22.983
R2287 GND.n1575 GND.n1504 22.983
R2288 GND.n1581 GND.n1502 22.983
R2289 GND.n1585 GND.n1497 22.983
R2290 GND.n1591 GND.n1495 22.983
R2291 GND.n1595 GND.n1490 22.983
R2292 GND.n1601 GND.n1488 22.983
R2293 GND.n1605 GND.n1485 22.983
R2294 GND.n1611 GND.n1483 22.983
R2295 GND.n1615 GND.n1479 22.983
R2296 GND.n1622 GND.n1477 22.983
R2297 GND.n1626 GND.n1473 22.983
R2298 GND.n1632 GND.n1471 22.983
R2299 GND.n1637 GND.n1467 22.983
R2300 GND.n1643 GND.n1466 22.983
R2301 GND.n1648 GND.n1461 22.983
R2302 GND.n194 GND.t110 21.317
R2303 GND.n219 GND.t132 21.317
R2304 GND.n227 GND.t27 21.317
R2305 GND.n252 GND.t80 21.317
R2306 GND.n17 GND.t139 21.317
R2307 GND.n42 GND.t64 21.317
R2308 GND.n50 GND.t82 21.317
R2309 GND.n75 GND.t265 21.317
R2310 GND.n99 GND.t26 21.317
R2311 GND.n124 GND.t171 21.317
R2312 GND.n132 GND.t137 21.317
R2313 GND.n157 GND.t8 21.317
R2314 GND.n396 GND.t101 21.317
R2315 GND.n402 GND.t4 21.317
R2316 GND.n299 GND.t3 21.317
R2317 GND.n324 GND.t273 21.317
R2318 GND.n330 GND.t13 21.317
R2319 GND.n355 GND.t144 21.317
R2320 GND.n456 GND.t113 21.317
R2321 GND.n481 GND.t9 21.317
R2322 GND.n487 GND.t108 21.317
R2323 GND.n512 GND.t47 21.317
R2324 GND.t95 GND.n954 21.317
R2325 GND.t77 GND.n837 21.317
R2326 GND.t76 GND.n888 21.317
R2327 GND.n900 GND.t260 21.317
R2328 GND.n910 GND.t85 21.317
R2329 GND.t50 GND.n855 21.317
R2330 GND.n992 GND.t73 21.317
R2331 GND.t37 GND.n1014 21.317
R2332 GND.n1017 GND.t35 21.317
R2333 GND.n1037 GND.t160 21.317
R2334 GND.t152 GND.n695 21.317
R2335 GND.t21 GND.n578 21.317
R2336 GND.t23 GND.n629 21.317
R2337 GND.n641 GND.t128 21.317
R2338 GND.n651 GND.t0 21.317
R2339 GND.t79 GND.n596 21.317
R2340 GND.n733 GND.t62 21.317
R2341 GND.t88 GND.n755 21.317
R2342 GND.n758 GND.t57 21.317
R2343 GND.n778 GND.t63 21.317
R2344 GND.t75 GND.n1552 19.784
R2345 GND.n1563 GND.t241 19.784
R2346 GND.t126 GND.n1583 19.784
R2347 GND.n1593 GND.t19 19.784
R2348 GND.n1594 GND.t313 19.784
R2349 GND.n1604 GND.t104 19.784
R2350 GND.n1624 GND.t230 19.784
R2351 GND.n1636 GND.t157 19.784
R2352 GND.t131 GND.n1792 19.784
R2353 GND.n1793 GND.t300 19.784
R2354 GND.t278 GND.n1824 19.784
R2355 GND.n1825 GND.t67 19.784
R2356 GND.n1834 GND.t135 19.784
R2357 GND.n1835 GND.t166 19.784
R2358 GND.n1866 GND.t284 19.784
R2359 GND.n1867 GND.t253 19.784
R2360 GND.n1531 GND.n1529 19.462
R2361 GND.n1762 GND.n1761 17.358
R2362 GND.n1666 GND.n1665 17.357
R2363 GND.n1661 GND.n1660 17.35
R2364 GND.n1542 GND.t34 15.827
R2365 GND.n1644 GND.t2 15.827
R2366 GND.n52 GND.n49 12.8
R2367 GND.n134 GND.n131 12.8
R2368 GND.n229 GND.n226 12.8
R2369 GND.n404 GND.n401 12.8
R2370 GND.n332 GND.n329 12.8
R2371 GND.n489 GND.n486 12.8
R2372 GND.n1207 GND.n1108 12.8
R2373 GND.n1211 GND.n1108 12.8
R2374 GND.n1211 GND.n1105 12.8
R2375 GND.n1218 GND.n1105 12.8
R2376 GND.n1218 GND.n1103 12.8
R2377 GND.n1223 GND.n1103 12.8
R2378 GND.n1223 GND.n1100 12.8
R2379 GND.n1229 GND.n1100 12.8
R2380 GND.n1229 GND.n1097 12.8
R2381 GND.n1234 GND.n1097 12.8
R2382 GND.n1234 GND.n1093 12.8
R2383 GND.n1240 GND.n1093 12.8
R2384 GND.n1240 GND.n1091 12.8
R2385 GND.n1244 GND.n1091 12.8
R2386 GND.n1244 GND.n1087 12.8
R2387 GND.n1248 GND.n1087 12.8
R2388 GND.n1146 GND.n1142 12.8
R2389 GND.n1146 GND.n1139 12.8
R2390 GND.n1153 GND.n1139 12.8
R2391 GND.n1153 GND.n1137 12.8
R2392 GND.n1157 GND.n1137 12.8
R2393 GND.n1157 GND.n1134 12.8
R2394 GND.n1164 GND.n1134 12.8
R2395 GND.n1164 GND.n1132 12.8
R2396 GND.n1169 GND.n1132 12.8
R2397 GND.n1169 GND.n1129 12.8
R2398 GND.n1175 GND.n1129 12.8
R2399 GND.n1175 GND.n1126 12.8
R2400 GND.n1180 GND.n1126 12.8
R2401 GND.n1180 GND.n1122 12.8
R2402 GND.n1186 GND.n1122 12.8
R2403 GND.n1186 GND.n1120 12.8
R2404 GND.n1190 GND.n1120 12.8
R2405 GND.n1190 GND.n1116 12.8
R2406 GND.n1196 GND.n1116 12.8
R2407 GND.n1196 GND.n1114 12.8
R2408 GND.n1200 GND.n1114 12.8
R2409 GND.n1200 GND.n1110 12.8
R2410 GND.n1204 GND.n1110 12.8
R2411 GND.n1251 GND.n1085 12.8
R2412 GND.n1255 GND.n1085 12.8
R2413 GND.n1255 GND.n1082 12.8
R2414 GND.n1262 GND.n1082 12.8
R2415 GND.n1262 GND.n1080 12.8
R2416 GND.n1266 GND.n1080 12.8
R2417 GND.n1266 GND.n1077 12.8
R2418 GND.n1273 GND.n1077 12.8
R2419 GND.n1273 GND.n1075 12.8
R2420 GND.n1278 GND.n1075 12.8
R2421 GND.n1278 GND.n1072 12.8
R2422 GND.n1284 GND.n1072 12.8
R2423 GND.n1284 GND.n1069 12.8
R2424 GND.n1289 GND.n1069 12.8
R2425 GND.n1289 GND.n1065 12.8
R2426 GND.n1295 GND.n1065 12.8
R2427 GND.n1295 GND.n1063 12.8
R2428 GND.n1299 GND.n1063 12.8
R2429 GND.n1299 GND.n1059 12.8
R2430 GND.n1305 GND.n1059 12.8
R2431 GND.n1305 GND.n1057 12.8
R2432 GND.n1310 GND.n1057 12.8
R2433 GND.n1310 GND.n1309 12.8
R2434 GND.n935 GND.n851 12.8
R2435 GND.n939 GND.n851 12.8
R2436 GND.n939 GND.n848 12.8
R2437 GND.n946 GND.n848 12.8
R2438 GND.n946 GND.n846 12.8
R2439 GND.n951 GND.n846 12.8
R2440 GND.n951 GND.n843 12.8
R2441 GND.n957 GND.n843 12.8
R2442 GND.n957 GND.n839 12.8
R2443 GND.n962 GND.n839 12.8
R2444 GND.n962 GND.n835 12.8
R2445 GND.n968 GND.n835 12.8
R2446 GND.n968 GND.n833 12.8
R2447 GND.n972 GND.n833 12.8
R2448 GND.n972 GND.n829 12.8
R2449 GND.n976 GND.n829 12.8
R2450 GND.n885 GND.n881 12.8
R2451 GND.n885 GND.n878 12.8
R2452 GND.n891 GND.n878 12.8
R2453 GND.n891 GND.n876 12.8
R2454 GND.n896 GND.n876 12.8
R2455 GND.n896 GND.n872 12.8
R2456 GND.n903 GND.n872 12.8
R2457 GND.n903 GND.n868 12.8
R2458 GND.n907 GND.n868 12.8
R2459 GND.n907 GND.n865 12.8
R2460 GND.n913 GND.n865 12.8
R2461 GND.n913 GND.n863 12.8
R2462 GND.n918 GND.n863 12.8
R2463 GND.n918 GND.n859 12.8
R2464 GND.n924 GND.n859 12.8
R2465 GND.n924 GND.n857 12.8
R2466 GND.n928 GND.n857 12.8
R2467 GND.n928 GND.n853 12.8
R2468 GND.n932 GND.n853 12.8
R2469 GND.n979 GND.n826 12.8
R2470 GND.n984 GND.n826 12.8
R2471 GND.n984 GND.n824 12.8
R2472 GND.n988 GND.n824 12.8
R2473 GND.n988 GND.n820 12.8
R2474 GND.n994 GND.n820 12.8
R2475 GND.n994 GND.n818 12.8
R2476 GND.n999 GND.n818 12.8
R2477 GND.n999 GND.n814 12.8
R2478 GND.n1005 GND.n814 12.8
R2479 GND.n1005 GND.n812 12.8
R2480 GND.n1012 GND.n812 12.8
R2481 GND.n1012 GND.n808 12.8
R2482 GND.n1019 GND.n808 12.8
R2483 GND.n1019 GND.n807 12.8
R2484 GND.n1024 GND.n807 12.8
R2485 GND.n1024 GND.n804 12.8
R2486 GND.n1031 GND.n804 12.8
R2487 GND.n1031 GND.n802 12.8
R2488 GND.n1035 GND.n802 12.8
R2489 GND.n1035 GND.n799 12.8
R2490 GND.n1042 GND.n799 12.8
R2491 GND.n1042 GND.n797 12.8
R2492 GND.n1047 GND.n797 12.8
R2493 GND.n1047 GND.n1046 12.8
R2494 GND.n676 GND.n592 12.8
R2495 GND.n680 GND.n592 12.8
R2496 GND.n680 GND.n589 12.8
R2497 GND.n687 GND.n589 12.8
R2498 GND.n687 GND.n587 12.8
R2499 GND.n692 GND.n587 12.8
R2500 GND.n692 GND.n584 12.8
R2501 GND.n698 GND.n584 12.8
R2502 GND.n698 GND.n580 12.8
R2503 GND.n703 GND.n580 12.8
R2504 GND.n703 GND.n576 12.8
R2505 GND.n709 GND.n576 12.8
R2506 GND.n709 GND.n574 12.8
R2507 GND.n713 GND.n574 12.8
R2508 GND.n713 GND.n570 12.8
R2509 GND.n717 GND.n570 12.8
R2510 GND.n626 GND.n622 12.8
R2511 GND.n626 GND.n619 12.8
R2512 GND.n632 GND.n619 12.8
R2513 GND.n632 GND.n617 12.8
R2514 GND.n637 GND.n617 12.8
R2515 GND.n637 GND.n613 12.8
R2516 GND.n644 GND.n613 12.8
R2517 GND.n644 GND.n609 12.8
R2518 GND.n648 GND.n609 12.8
R2519 GND.n648 GND.n606 12.8
R2520 GND.n654 GND.n606 12.8
R2521 GND.n654 GND.n604 12.8
R2522 GND.n659 GND.n604 12.8
R2523 GND.n659 GND.n600 12.8
R2524 GND.n665 GND.n600 12.8
R2525 GND.n665 GND.n598 12.8
R2526 GND.n669 GND.n598 12.8
R2527 GND.n669 GND.n594 12.8
R2528 GND.n673 GND.n594 12.8
R2529 GND.n720 GND.n567 12.8
R2530 GND.n725 GND.n567 12.8
R2531 GND.n725 GND.n565 12.8
R2532 GND.n729 GND.n565 12.8
R2533 GND.n729 GND.n561 12.8
R2534 GND.n735 GND.n561 12.8
R2535 GND.n735 GND.n559 12.8
R2536 GND.n740 GND.n559 12.8
R2537 GND.n740 GND.n555 12.8
R2538 GND.n746 GND.n555 12.8
R2539 GND.n746 GND.n553 12.8
R2540 GND.n753 GND.n553 12.8
R2541 GND.n753 GND.n549 12.8
R2542 GND.n760 GND.n549 12.8
R2543 GND.n760 GND.n548 12.8
R2544 GND.n765 GND.n548 12.8
R2545 GND.n765 GND.n545 12.8
R2546 GND.n772 GND.n545 12.8
R2547 GND.n772 GND.n543 12.8
R2548 GND.n776 GND.n543 12.8
R2549 GND.n776 GND.n540 12.8
R2550 GND.n783 GND.n540 12.8
R2551 GND.n783 GND.n538 12.8
R2552 GND.n788 GND.n538 12.8
R2553 GND.n788 GND.n787 12.8
R2554 GND.n1898 GND.n1897 12.475
R2555 GND.n11 GND.n10 9.154
R2556 GND.n93 GND.n92 9.154
R2557 GND.n97 GND.n96 9.154
R2558 GND.n96 GND.n95 9.154
R2559 GND.n101 GND.n100 9.154
R2560 GND.n100 GND.n99 9.154
R2561 GND.n105 GND.n104 9.154
R2562 GND.n104 GND.n103 9.154
R2563 GND.n109 GND.n108 9.154
R2564 GND.n108 GND.n107 9.154
R2565 GND.n113 GND.n112 9.154
R2566 GND.n112 GND.n111 9.154
R2567 GND.n118 GND.n117 9.154
R2568 GND.n117 GND.n116 9.154
R2569 GND.n122 GND.n121 9.154
R2570 GND.n121 GND.n120 9.154
R2571 GND.n126 GND.n125 9.154
R2572 GND.n125 GND.n124 9.154
R2573 GND.n131 GND.n130 9.154
R2574 GND.n130 GND.n129 9.154
R2575 GND.n134 GND.n133 9.154
R2576 GND.n133 GND.n132 9.154
R2577 GND.n138 GND.n137 9.154
R2578 GND.n137 GND.n136 9.154
R2579 GND.n142 GND.n141 9.154
R2580 GND.n141 GND.n140 9.154
R2581 GND.n147 GND.n146 9.154
R2582 GND.n146 GND.n145 9.154
R2583 GND.n151 GND.n150 9.154
R2584 GND.n150 GND.n149 9.154
R2585 GND.n155 GND.n154 9.154
R2586 GND.n154 GND.n153 9.154
R2587 GND.n159 GND.n158 9.154
R2588 GND.n158 GND.n157 9.154
R2589 GND.n163 GND.n162 9.154
R2590 GND.n162 GND.n161 9.154
R2591 GND.n167 GND.n166 9.154
R2592 GND.n15 GND.n14 9.154
R2593 GND.n14 GND.n13 9.154
R2594 GND.n19 GND.n18 9.154
R2595 GND.n18 GND.n17 9.154
R2596 GND.n23 GND.n22 9.154
R2597 GND.n22 GND.n21 9.154
R2598 GND.n27 GND.n26 9.154
R2599 GND.n26 GND.n25 9.154
R2600 GND.n31 GND.n30 9.154
R2601 GND.n30 GND.n29 9.154
R2602 GND.n36 GND.n35 9.154
R2603 GND.n35 GND.n34 9.154
R2604 GND.n40 GND.n39 9.154
R2605 GND.n39 GND.n38 9.154
R2606 GND.n44 GND.n43 9.154
R2607 GND.n43 GND.n42 9.154
R2608 GND.n49 GND.n48 9.154
R2609 GND.n48 GND.n47 9.154
R2610 GND.n52 GND.n51 9.154
R2611 GND.n51 GND.n50 9.154
R2612 GND.n56 GND.n55 9.154
R2613 GND.n55 GND.n54 9.154
R2614 GND.n60 GND.n59 9.154
R2615 GND.n59 GND.n58 9.154
R2616 GND.n65 GND.n64 9.154
R2617 GND.n64 GND.n63 9.154
R2618 GND.n69 GND.n68 9.154
R2619 GND.n68 GND.n67 9.154
R2620 GND.n73 GND.n72 9.154
R2621 GND.n72 GND.n71 9.154
R2622 GND.n77 GND.n76 9.154
R2623 GND.n76 GND.n75 9.154
R2624 GND.n81 GND.n80 9.154
R2625 GND.n80 GND.n79 9.154
R2626 GND.n85 GND.n84 9.154
R2627 GND.n176 GND.n175 9.154
R2628 GND.n175 GND.n174 9.154
R2629 GND.n180 GND.n179 9.154
R2630 GND.n179 GND.n178 9.154
R2631 GND.n184 GND.n183 9.154
R2632 GND.n183 GND.n182 9.154
R2633 GND.n188 GND.n187 9.154
R2634 GND.n187 GND.n186 9.154
R2635 GND.n192 GND.n191 9.154
R2636 GND.n191 GND.n190 9.154
R2637 GND.n196 GND.n195 9.154
R2638 GND.n195 GND.n194 9.154
R2639 GND.n200 GND.n199 9.154
R2640 GND.n199 GND.n198 9.154
R2641 GND.n204 GND.n203 9.154
R2642 GND.n203 GND.n202 9.154
R2643 GND.n208 GND.n207 9.154
R2644 GND.n207 GND.n206 9.154
R2645 GND.n213 GND.n212 9.154
R2646 GND.n212 GND.n211 9.154
R2647 GND.n217 GND.n216 9.154
R2648 GND.n216 GND.n215 9.154
R2649 GND.n221 GND.n220 9.154
R2650 GND.n220 GND.n219 9.154
R2651 GND.n226 GND.n225 9.154
R2652 GND.n225 GND.n224 9.154
R2653 GND.n229 GND.n228 9.154
R2654 GND.n228 GND.n227 9.154
R2655 GND.n233 GND.n232 9.154
R2656 GND.n232 GND.n231 9.154
R2657 GND.n237 GND.n236 9.154
R2658 GND.n236 GND.n235 9.154
R2659 GND.n242 GND.n241 9.154
R2660 GND.n241 GND.n240 9.154
R2661 GND.n246 GND.n245 9.154
R2662 GND.n245 GND.n244 9.154
R2663 GND.n250 GND.n249 9.154
R2664 GND.n249 GND.n248 9.154
R2665 GND.n254 GND.n253 9.154
R2666 GND.n253 GND.n252 9.154
R2667 GND.n258 GND.n257 9.154
R2668 GND.n257 GND.n256 9.154
R2669 GND.n262 GND.n261 9.154
R2670 GND.n261 GND.n260 9.154
R2671 GND.n266 GND.n265 9.154
R2672 GND.n265 GND.n264 9.154
R2673 GND.n270 GND.n269 9.154
R2674 GND.n269 GND.n268 9.154
R2675 GND.n2 GND.n1 9.154
R2676 GND.n1 GND.n0 9.154
R2677 GND.n274 GND.n273 9.154
R2678 GND.n172 GND.n171 9.154
R2679 GND.n293 GND.n292 9.154
R2680 GND.n297 GND.n296 9.154
R2681 GND.n296 GND.n295 9.154
R2682 GND.n301 GND.n300 9.154
R2683 GND.n300 GND.n299 9.154
R2684 GND.n305 GND.n304 9.154
R2685 GND.n304 GND.n303 9.154
R2686 GND.n309 GND.n308 9.154
R2687 GND.n308 GND.n307 9.154
R2688 GND.n313 GND.n312 9.154
R2689 GND.n312 GND.n311 9.154
R2690 GND.n318 GND.n317 9.154
R2691 GND.n317 GND.n316 9.154
R2692 GND.n322 GND.n321 9.154
R2693 GND.n321 GND.n320 9.154
R2694 GND.n326 GND.n325 9.154
R2695 GND.n325 GND.n324 9.154
R2696 GND.n329 GND.n288 9.154
R2697 GND.n288 GND.n287 9.154
R2698 GND.n332 GND.n331 9.154
R2699 GND.n331 GND.n330 9.154
R2700 GND.n336 GND.n335 9.154
R2701 GND.n335 GND.n334 9.154
R2702 GND.n340 GND.n339 9.154
R2703 GND.n339 GND.n338 9.154
R2704 GND.n345 GND.n344 9.154
R2705 GND.n344 GND.n343 9.154
R2706 GND.n349 GND.n348 9.154
R2707 GND.n348 GND.n347 9.154
R2708 GND.n353 GND.n352 9.154
R2709 GND.n352 GND.n351 9.154
R2710 GND.n357 GND.n356 9.154
R2711 GND.n356 GND.n355 9.154
R2712 GND.n361 GND.n360 9.154
R2713 GND.n360 GND.n359 9.154
R2714 GND.n365 GND.n364 9.154
R2715 GND.n373 GND.n372 9.154
R2716 GND.n377 GND.n376 9.154
R2717 GND.n376 GND.n375 9.154
R2718 GND.n381 GND.n380 9.154
R2719 GND.n380 GND.n379 9.154
R2720 GND.n385 GND.n384 9.154
R2721 GND.n384 GND.n383 9.154
R2722 GND.n390 GND.n389 9.154
R2723 GND.n389 GND.n388 9.154
R2724 GND.n394 GND.n393 9.154
R2725 GND.n393 GND.n392 9.154
R2726 GND.n398 GND.n397 9.154
R2727 GND.n397 GND.n396 9.154
R2728 GND.n401 GND.n284 9.154
R2729 GND.n284 GND.n283 9.154
R2730 GND.n404 GND.n403 9.154
R2731 GND.n403 GND.n402 9.154
R2732 GND.n408 GND.n407 9.154
R2733 GND.n407 GND.n406 9.154
R2734 GND.n412 GND.n411 9.154
R2735 GND.n411 GND.n410 9.154
R2736 GND.n417 GND.n416 9.154
R2737 GND.n416 GND.n415 9.154
R2738 GND.n421 GND.n420 9.154
R2739 GND.n420 GND.n419 9.154
R2740 GND.n425 GND.n424 9.154
R2741 GND.n424 GND.n423 9.154
R2742 GND.n429 GND.n428 9.154
R2743 GND.n534 GND.n533 9.154
R2744 GND.n434 GND.n433 9.154
R2745 GND.n438 GND.n437 9.154
R2746 GND.n437 GND.n436 9.154
R2747 GND.n442 GND.n441 9.154
R2748 GND.n441 GND.n440 9.154
R2749 GND.n446 GND.n445 9.154
R2750 GND.n445 GND.n444 9.154
R2751 GND.n450 GND.n449 9.154
R2752 GND.n449 GND.n448 9.154
R2753 GND.n454 GND.n453 9.154
R2754 GND.n453 GND.n452 9.154
R2755 GND.n458 GND.n457 9.154
R2756 GND.n457 GND.n456 9.154
R2757 GND.n462 GND.n461 9.154
R2758 GND.n461 GND.n460 9.154
R2759 GND.n466 GND.n465 9.154
R2760 GND.n465 GND.n464 9.154
R2761 GND.n470 GND.n469 9.154
R2762 GND.n469 GND.n468 9.154
R2763 GND.n475 GND.n474 9.154
R2764 GND.n474 GND.n473 9.154
R2765 GND.n479 GND.n478 9.154
R2766 GND.n478 GND.n477 9.154
R2767 GND.n483 GND.n482 9.154
R2768 GND.n482 GND.n481 9.154
R2769 GND.n486 GND.n280 9.154
R2770 GND.n280 GND.n279 9.154
R2771 GND.n489 GND.n488 9.154
R2772 GND.n488 GND.n487 9.154
R2773 GND.n493 GND.n492 9.154
R2774 GND.n492 GND.n491 9.154
R2775 GND.n497 GND.n496 9.154
R2776 GND.n496 GND.n495 9.154
R2777 GND.n502 GND.n501 9.154
R2778 GND.n501 GND.n500 9.154
R2779 GND.n506 GND.n505 9.154
R2780 GND.n505 GND.n504 9.154
R2781 GND.n510 GND.n509 9.154
R2782 GND.n509 GND.n508 9.154
R2783 GND.n514 GND.n513 9.154
R2784 GND.n513 GND.n512 9.154
R2785 GND.n518 GND.n517 9.154
R2786 GND.n517 GND.n516 9.154
R2787 GND.n522 GND.n521 9.154
R2788 GND.n521 GND.n520 9.154
R2789 GND.n526 GND.n525 9.154
R2790 GND.n525 GND.n524 9.154
R2791 GND.n530 GND.n529 9.154
R2792 GND.n529 GND.n528 9.154
R2793 GND.n278 GND.n277 9.154
R2794 GND.n277 GND.n276 9.154
R2795 GND.n1533 GND.n1532 9.154
R2796 GND.n1528 GND.n1527 9.154
R2797 GND.n1530 GND.n1527 9.154
R2798 GND.n1539 GND.n1538 9.154
R2799 GND.n1540 GND.n1539 9.154
R2800 GND.n1545 GND.n1544 9.154
R2801 GND.n1544 GND.n1543 9.154
R2802 GND.n1550 GND.n1549 9.154
R2803 GND.n1551 GND.n1550 9.154
R2804 GND.n1555 GND.n1554 9.154
R2805 GND.n1554 GND.n1553 9.154
R2806 GND.n1560 GND.n1559 9.154
R2807 GND.n1561 GND.n1560 9.154
R2808 GND.n1565 GND.n1564 9.154
R2809 GND.n1564 GND.n1563 9.154
R2810 GND.n1571 GND.n1570 9.154
R2811 GND.n1572 GND.n1571 9.154
R2812 GND.n1576 GND.n1575 9.154
R2813 GND.n1575 GND.n1574 9.154
R2814 GND.n1581 GND.n1580 9.154
R2815 GND.n1582 GND.n1581 9.154
R2816 GND.n1586 GND.n1585 9.154
R2817 GND.n1585 GND.n1584 9.154
R2818 GND.n1591 GND.n1590 9.154
R2819 GND.n1592 GND.n1591 9.154
R2820 GND.n1596 GND.n1595 9.154
R2821 GND.n1595 GND.n1594 9.154
R2822 GND.n1601 GND.n1600 9.154
R2823 GND.n1602 GND.n1601 9.154
R2824 GND.n1606 GND.n1605 9.154
R2825 GND.n1605 GND.n1604 9.154
R2826 GND.n1611 GND.n1610 9.154
R2827 GND.n1612 GND.n1611 9.154
R2828 GND.n1616 GND.n1615 9.154
R2829 GND.n1615 GND.n1614 9.154
R2830 GND.n1622 GND.n1621 9.154
R2831 GND.n1623 GND.n1622 9.154
R2832 GND.n1627 GND.n1626 9.154
R2833 GND.n1626 GND.n1625 9.154
R2834 GND.n1632 GND.n1631 9.154
R2835 GND.n1633 GND.n1632 9.154
R2836 GND.n1638 GND.n1637 9.154
R2837 GND.n1637 GND.n1636 9.154
R2838 GND.n1643 GND.n1642 9.154
R2839 GND.n1644 GND.n1643 9.154
R2840 GND.n1649 GND.n1648 9.154
R2841 GND.n1648 GND.n1647 9.154
R2842 GND.n1525 GND.n1524 9.154
R2843 GND.n1541 GND.n1525 9.154
R2844 GND.n1522 GND.n1521 9.154
R2845 GND.n1542 GND.n1521 9.154
R2846 GND.n1520 GND.n1519 9.154
R2847 GND.n1552 GND.n1520 9.154
R2848 GND.n1517 GND.n1516 9.154
R2849 GND.n1516 GND.n1515 9.154
R2850 GND.n1514 GND.n1513 9.154
R2851 GND.n1562 GND.n1514 9.154
R2852 GND.n1511 GND.n1510 9.154
R2853 GND.n1510 GND.n1509 9.154
R2854 GND.n1508 GND.n1507 9.154
R2855 GND.n1573 GND.n1508 9.154
R2856 GND.n1505 GND.n1504 9.154
R2857 GND.n1504 GND.n1503 9.154
R2858 GND.n1502 GND.n1501 9.154
R2859 GND.n1583 GND.n1502 9.154
R2860 GND.n1498 GND.n1497 9.154
R2861 GND.n1497 GND.n1496 9.154
R2862 GND.n1495 GND.n1494 9.154
R2863 GND.n1593 GND.n1495 9.154
R2864 GND.n1491 GND.n1490 9.154
R2865 GND.n1490 GND.n1489 9.154
R2866 GND.n1488 GND.n1487 9.154
R2867 GND.n1603 GND.n1488 9.154
R2868 GND.n1486 GND.n1485 9.154
R2869 GND.n1485 GND.n1484 9.154
R2870 GND.n1483 GND.n1482 9.154
R2871 GND.n1613 GND.n1483 9.154
R2872 GND.n1480 GND.n1479 9.154
R2873 GND.n1479 GND.n1478 9.154
R2874 GND.n1477 GND.n1476 9.154
R2875 GND.n1624 GND.n1477 9.154
R2876 GND.n1474 GND.n1473 9.154
R2877 GND.n1473 GND.n1472 9.154
R2878 GND.n1471 GND.n1470 9.154
R2879 GND.n1634 GND.n1471 9.154
R2880 GND.n1468 GND.n1467 9.154
R2881 GND.n1635 GND.n1467 9.154
R2882 GND.n1466 GND.n1465 9.154
R2883 GND.n1645 GND.n1466 9.154
R2884 GND.n1462 GND.n1461 9.154
R2885 GND.n1646 GND.n1461 9.154
R2886 GND.n1657 GND.n1656 9.154
R2887 GND.n1652 GND.n1458 9.154
R2888 GND.n1668 GND.n1667 9.154
R2889 GND.n1679 GND.n1678 9.154
R2890 GND.n1678 GND.n1677 9.154
R2891 GND.n1685 GND.n1684 9.154
R2892 GND.n1686 GND.n1685 9.154
R2893 GND.n1690 GND.n1689 9.154
R2894 GND.n1689 GND.n1688 9.154
R2895 GND.n1696 GND.n1695 9.154
R2896 GND.n1697 GND.n1696 9.154
R2897 GND.n1701 GND.n1700 9.154
R2898 GND.n1700 GND.n1699 9.154
R2899 GND.n1706 GND.n1705 9.154
R2900 GND.n1707 GND.n1706 9.154
R2901 GND.n1712 GND.n1711 9.154
R2902 GND.n1711 GND.n1710 9.154
R2903 GND.n1717 GND.n1716 9.154
R2904 GND.n1718 GND.n1717 9.154
R2905 GND.n1722 GND.n1721 9.154
R2906 GND.n1721 GND.n1720 9.154
R2907 GND.n1728 GND.n1727 9.154
R2908 GND.n1729 GND.n1728 9.154
R2909 GND.n1733 GND.n1732 9.154
R2910 GND.n1732 GND.n1731 9.154
R2911 GND.n1739 GND.n1738 9.154
R2912 GND.n1740 GND.n1739 9.154
R2913 GND.n1744 GND.n1743 9.154
R2914 GND.n1743 GND.n1742 9.154
R2915 GND.n1752 GND.n1751 9.154
R2916 GND.n1753 GND.n1752 9.154
R2917 GND.n1747 GND.n1403 9.154
R2918 GND.n1754 GND.n1403 9.154
R2919 GND.n1757 GND.n1756 9.154
R2920 GND.n1756 GND.n1755 9.154
R2921 GND.n1674 GND.n1673 9.154
R2922 GND.n1675 GND.n1674 9.154
R2923 GND.n1451 GND.n1450 9.154
R2924 GND.n1450 GND.n1449 9.154
R2925 GND.n1448 GND.n1447 9.154
R2926 GND.n1676 GND.n1448 9.154
R2927 GND.n1445 GND.n1444 9.154
R2928 GND.n1444 GND.n1443 9.154
R2929 GND.n1442 GND.n1441 9.154
R2930 GND.n1687 GND.n1442 9.154
R2931 GND.n1439 GND.n1438 9.154
R2932 GND.n1438 GND.n1437 9.154
R2933 GND.n1436 GND.n1435 9.154
R2934 GND.n1698 GND.n1436 9.154
R2935 GND.n1432 GND.n1431 9.154
R2936 GND.n1431 GND.n1430 9.154
R2937 GND.n1429 GND.n1428 9.154
R2938 GND.n1708 GND.n1429 9.154
R2939 GND.n1425 GND.n1424 9.154
R2940 GND.n1424 GND.n1423 9.154
R2941 GND.n1422 GND.n1421 9.154
R2942 GND.n1719 GND.n1422 9.154
R2943 GND.n1419 GND.n1418 9.154
R2944 GND.n1418 GND.n1417 9.154
R2945 GND.n1416 GND.n1415 9.154
R2946 GND.n1730 GND.n1416 9.154
R2947 GND.n1413 GND.n1412 9.154
R2948 GND.n1412 GND.n1411 9.154
R2949 GND.n1410 GND.n1409 9.154
R2950 GND.n1741 GND.n1410 9.154
R2951 GND.n1406 GND.n1405 9.154
R2952 GND.n1405 GND.n1404 9.154
R2953 GND.n1770 GND.n1769 9.154
R2954 GND.n1771 GND.n1770 9.154
R2955 GND.n1775 GND.n1774 9.154
R2956 GND.n1774 GND.n1773 9.154
R2957 GND.n1780 GND.n1779 9.154
R2958 GND.n1781 GND.n1780 9.154
R2959 GND.n1785 GND.n1784 9.154
R2960 GND.n1784 GND.n1783 9.154
R2961 GND.n1790 GND.n1789 9.154
R2962 GND.n1791 GND.n1790 9.154
R2963 GND.n1795 GND.n1794 9.154
R2964 GND.n1794 GND.n1793 9.154
R2965 GND.n1800 GND.n1799 9.154
R2966 GND.n1801 GND.n1800 9.154
R2967 GND.n1805 GND.n1804 9.154
R2968 GND.n1804 GND.n1803 9.154
R2969 GND.n1812 GND.n1811 9.154
R2970 GND.n1813 GND.n1812 9.154
R2971 GND.n1817 GND.n1816 9.154
R2972 GND.n1816 GND.n1815 9.154
R2973 GND.n1822 GND.n1821 9.154
R2974 GND.n1823 GND.n1822 9.154
R2975 GND.n1827 GND.n1826 9.154
R2976 GND.n1826 GND.n1825 9.154
R2977 GND.n1832 GND.n1831 9.154
R2978 GND.n1833 GND.n1832 9.154
R2979 GND.n1837 GND.n1836 9.154
R2980 GND.n1836 GND.n1835 9.154
R2981 GND.n1842 GND.n1841 9.154
R2982 GND.n1843 GND.n1842 9.154
R2983 GND.n1847 GND.n1846 9.154
R2984 GND.n1846 GND.n1845 9.154
R2985 GND.n1854 GND.n1853 9.154
R2986 GND.n1855 GND.n1854 9.154
R2987 GND.n1859 GND.n1858 9.154
R2988 GND.n1858 GND.n1857 9.154
R2989 GND.n1864 GND.n1863 9.154
R2990 GND.n1865 GND.n1864 9.154
R2991 GND.n1869 GND.n1868 9.154
R2992 GND.n1868 GND.n1867 9.154
R2993 GND.n1874 GND.n1873 9.154
R2994 GND.n1875 GND.n1874 9.154
R2995 GND.n1879 GND.n1878 9.154
R2996 GND.n1878 GND.n1877 9.154
R2997 GND.n1884 GND.n1883 9.154
R2998 GND.n1885 GND.n1884 9.154
R2999 GND.n1889 GND.n1888 9.154
R3000 GND.n1888 GND.n1887 9.154
R3001 GND.n1894 GND.n1893 9.154
R3002 GND.n1895 GND.n1894 9.154
R3003 GND.n1764 GND.n1763 9.154
R3004 GND.n1396 GND.n1395 9.154
R3005 GND.n1395 GND.n1394 9.154
R3006 GND.n1393 GND.n1392 9.154
R3007 GND.n1772 GND.n1393 9.154
R3008 GND.n1390 GND.n1389 9.154
R3009 GND.n1389 GND.n1388 9.154
R3010 GND.n1387 GND.n1386 9.154
R3011 GND.n1782 GND.n1387 9.154
R3012 GND.n1384 GND.n1383 9.154
R3013 GND.n1383 GND.n1382 9.154
R3014 GND.n1381 GND.n1380 9.154
R3015 GND.n1792 GND.n1381 9.154
R3016 GND.n1378 GND.n1377 9.154
R3017 GND.n1377 GND.n1376 9.154
R3018 GND.n1375 GND.n1374 9.154
R3019 GND.n1802 GND.n1375 9.154
R3020 GND.n1372 GND.n1371 9.154
R3021 GND.n1371 GND.n1370 9.154
R3022 GND.n1369 GND.n1368 9.154
R3023 GND.n1814 GND.n1369 9.154
R3024 GND.n1366 GND.n1365 9.154
R3025 GND.n1365 GND.n1364 9.154
R3026 GND.n1363 GND.n1362 9.154
R3027 GND.n1824 GND.n1363 9.154
R3028 GND.n1358 GND.n1357 9.154
R3029 GND.n1357 GND.n1356 9.154
R3030 GND.n1355 GND.n1354 9.154
R3031 GND.n1834 GND.n1355 9.154
R3032 GND.n1352 GND.n1351 9.154
R3033 GND.n1351 GND.n1350 9.154
R3034 GND.n1349 GND.n1348 9.154
R3035 GND.n1844 GND.n1349 9.154
R3036 GND.n1346 GND.n1345 9.154
R3037 GND.n1345 GND.n1344 9.154
R3038 GND.n1343 GND.n1342 9.154
R3039 GND.n1856 GND.n1343 9.154
R3040 GND.n1340 GND.n1339 9.154
R3041 GND.n1339 GND.n1338 9.154
R3042 GND.n1337 GND.n1336 9.154
R3043 GND.n1866 GND.n1337 9.154
R3044 GND.n1334 GND.n1333 9.154
R3045 GND.n1333 GND.n1332 9.154
R3046 GND.n1331 GND.n1330 9.154
R3047 GND.n1876 GND.n1331 9.154
R3048 GND.n1328 GND.n1327 9.154
R3049 GND.n1327 GND.n1326 9.154
R3050 GND.n1325 GND.n1324 9.154
R3051 GND.n1886 GND.n1325 9.154
R3052 GND.n1321 GND.n1320 9.154
R3053 GND.n1320 GND.n1319 9.154
R3054 GND.n1322 GND.n1318 9.154
R3055 GND.n1142 GND.n1141 9.154
R3056 GND.n1147 GND.n1146 9.154
R3057 GND.n1148 GND.n1147 9.154
R3058 GND.n1140 GND.n1139 9.154
R3059 GND.n1149 GND.n1140 9.154
R3060 GND.n1153 GND.n1152 9.154
R3061 GND.n1152 GND.n1151 9.154
R3062 GND.n1137 GND.n1136 9.154
R3063 GND.n1150 GND.n1136 9.154
R3064 GND.n1158 GND.n1157 9.154
R3065 GND.n1159 GND.n1158 9.154
R3066 GND.n1135 GND.n1134 9.154
R3067 GND.n1160 GND.n1135 9.154
R3068 GND.n1164 GND.n1163 9.154
R3069 GND.n1163 GND.n1162 9.154
R3070 GND.n1132 GND.n1131 9.154
R3071 GND.n1161 GND.n1131 9.154
R3072 GND.n1170 GND.n1169 9.154
R3073 GND.n1171 GND.n1170 9.154
R3074 GND.n1130 GND.n1129 9.154
R3075 GND.n1172 GND.n1130 9.154
R3076 GND.n1175 GND.n1174 9.154
R3077 GND.n1174 GND.n1173 9.154
R3078 GND.n1126 GND.n1125 9.154
R3079 GND.n1125 GND.n1124 9.154
R3080 GND.n1181 GND.n1180 9.154
R3081 GND.n1182 GND.n1181 9.154
R3082 GND.n1123 GND.n1122 9.154
R3083 GND.n1183 GND.n1123 9.154
R3084 GND.n1186 GND.n1185 9.154
R3085 GND.n1185 GND.n1184 9.154
R3086 GND.n1120 GND.n1119 9.154
R3087 GND.n1119 GND.n1118 9.154
R3088 GND.n1191 GND.n1190 9.154
R3089 GND.n1192 GND.n1191 9.154
R3090 GND.n1117 GND.n1116 9.154
R3091 GND.n1193 GND.n1117 9.154
R3092 GND.n1196 GND.n1195 9.154
R3093 GND.n1195 GND.n1194 9.154
R3094 GND.n1114 GND.n1113 9.154
R3095 GND.n1113 GND.n1112 9.154
R3096 GND.n1201 GND.n1200 9.154
R3097 GND.n1202 GND.n1201 9.154
R3098 GND.n1111 GND.n1110 9.154
R3099 GND.n1108 GND.n1107 9.154
R3100 GND.n1212 GND.n1211 9.154
R3101 GND.n1213 GND.n1212 9.154
R3102 GND.n1106 GND.n1105 9.154
R3103 GND.n1214 GND.n1106 9.154
R3104 GND.n1218 GND.n1217 9.154
R3105 GND.n1217 GND.n1216 9.154
R3106 GND.n1103 GND.n1102 9.154
R3107 GND.n1215 GND.n1102 9.154
R3108 GND.n1224 GND.n1223 9.154
R3109 GND.n1225 GND.n1224 9.154
R3110 GND.n1101 GND.n1100 9.154
R3111 GND.n1226 GND.n1101 9.154
R3112 GND.n1229 GND.n1228 9.154
R3113 GND.n1228 GND.n1227 9.154
R3114 GND.n1097 GND.n1096 9.154
R3115 GND.n1096 GND.n1095 9.154
R3116 GND.n1235 GND.n1234 9.154
R3117 GND.n1236 GND.n1235 9.154
R3118 GND.n1094 GND.n1093 9.154
R3119 GND.n1237 GND.n1094 9.154
R3120 GND.n1240 GND.n1239 9.154
R3121 GND.n1239 GND.n1238 9.154
R3122 GND.n1091 GND.n1090 9.154
R3123 GND.n1090 GND.n1089 9.154
R3124 GND.n1245 GND.n1244 9.154
R3125 GND.n1246 GND.n1245 9.154
R3126 GND.n1088 GND.n1087 9.154
R3127 GND.n1085 GND.n1084 9.154
R3128 GND.n1256 GND.n1255 9.154
R3129 GND.n1257 GND.n1256 9.154
R3130 GND.n1083 GND.n1082 9.154
R3131 GND.n1258 GND.n1083 9.154
R3132 GND.n1262 GND.n1261 9.154
R3133 GND.n1261 GND.n1260 9.154
R3134 GND.n1080 GND.n1079 9.154
R3135 GND.n1259 GND.n1079 9.154
R3136 GND.n1267 GND.n1266 9.154
R3137 GND.n1268 GND.n1267 9.154
R3138 GND.n1078 GND.n1077 9.154
R3139 GND.n1269 GND.n1078 9.154
R3140 GND.n1273 GND.n1272 9.154
R3141 GND.n1272 GND.n1271 9.154
R3142 GND.n1075 GND.n1074 9.154
R3143 GND.n1270 GND.n1074 9.154
R3144 GND.n1279 GND.n1278 9.154
R3145 GND.n1280 GND.n1279 9.154
R3146 GND.n1073 GND.n1072 9.154
R3147 GND.n1281 GND.n1073 9.154
R3148 GND.n1284 GND.n1283 9.154
R3149 GND.n1283 GND.n1282 9.154
R3150 GND.n1069 GND.n1068 9.154
R3151 GND.n1068 GND.n1067 9.154
R3152 GND.n1290 GND.n1289 9.154
R3153 GND.n1291 GND.n1290 9.154
R3154 GND.n1066 GND.n1065 9.154
R3155 GND.n1292 GND.n1066 9.154
R3156 GND.n1295 GND.n1294 9.154
R3157 GND.n1294 GND.n1293 9.154
R3158 GND.n1063 GND.n1062 9.154
R3159 GND.n1062 GND.n1061 9.154
R3160 GND.n1300 GND.n1299 9.154
R3161 GND.n1301 GND.n1300 9.154
R3162 GND.n1060 GND.n1059 9.154
R3163 GND.n1302 GND.n1060 9.154
R3164 GND.n1305 GND.n1304 9.154
R3165 GND.n1304 GND.n1303 9.154
R3166 GND.n1057 GND.n1056 9.154
R3167 GND.n1056 GND.n1055 9.154
R3168 GND.n1311 GND.n1310 9.154
R3169 GND.n1312 GND.n1311 9.154
R3170 GND.n1309 GND.n1054 9.154
R3171 GND.n881 GND.n880 9.154
R3172 GND.n886 GND.n885 9.154
R3173 GND.n887 GND.n886 9.154
R3174 GND.n879 GND.n878 9.154
R3175 GND.n888 GND.n879 9.154
R3176 GND.n891 GND.n890 9.154
R3177 GND.n890 GND.n889 9.154
R3178 GND.n876 GND.n875 9.154
R3179 GND.n875 GND.n874 9.154
R3180 GND.n897 GND.n896 9.154
R3181 GND.n898 GND.n897 9.154
R3182 GND.n873 GND.n872 9.154
R3183 GND.n899 GND.n873 9.154
R3184 GND.n903 GND.n902 9.154
R3185 GND.n902 GND.n901 9.154
R3186 GND.n868 GND.n867 9.154
R3187 GND.n900 GND.n867 9.154
R3188 GND.n908 GND.n907 9.154
R3189 GND.n909 GND.n908 9.154
R3190 GND.n866 GND.n865 9.154
R3191 GND.n910 GND.n866 9.154
R3192 GND.n913 GND.n912 9.154
R3193 GND.n912 GND.n911 9.154
R3194 GND.n863 GND.n862 9.154
R3195 GND.n862 GND.n861 9.154
R3196 GND.n919 GND.n918 9.154
R3197 GND.n920 GND.n919 9.154
R3198 GND.n860 GND.n859 9.154
R3199 GND.n921 GND.n860 9.154
R3200 GND.n924 GND.n923 9.154
R3201 GND.n923 GND.n922 9.154
R3202 GND.n857 GND.n856 9.154
R3203 GND.n856 GND.n855 9.154
R3204 GND.n929 GND.n928 9.154
R3205 GND.n930 GND.n929 9.154
R3206 GND.n854 GND.n853 9.154
R3207 GND.n851 GND.n850 9.154
R3208 GND.n940 GND.n939 9.154
R3209 GND.n941 GND.n940 9.154
R3210 GND.n849 GND.n848 9.154
R3211 GND.n942 GND.n849 9.154
R3212 GND.n946 GND.n945 9.154
R3213 GND.n945 GND.n944 9.154
R3214 GND.n846 GND.n845 9.154
R3215 GND.n943 GND.n845 9.154
R3216 GND.n952 GND.n951 9.154
R3217 GND.n953 GND.n952 9.154
R3218 GND.n844 GND.n843 9.154
R3219 GND.n954 GND.n844 9.154
R3220 GND.n957 GND.n956 9.154
R3221 GND.n956 GND.n955 9.154
R3222 GND.n839 GND.n838 9.154
R3223 GND.n838 GND.n837 9.154
R3224 GND.n963 GND.n962 9.154
R3225 GND.n964 GND.n963 9.154
R3226 GND.n836 GND.n835 9.154
R3227 GND.n965 GND.n836 9.154
R3228 GND.n968 GND.n967 9.154
R3229 GND.n967 GND.n966 9.154
R3230 GND.n833 GND.n832 9.154
R3231 GND.n832 GND.n831 9.154
R3232 GND.n973 GND.n972 9.154
R3233 GND.n974 GND.n973 9.154
R3234 GND.n830 GND.n829 9.154
R3235 GND.n1052 GND.n1051 9.154
R3236 GND.n980 GND.n979 9.154
R3237 GND.n827 GND.n826 9.154
R3238 GND.n981 GND.n827 9.154
R3239 GND.n984 GND.n983 9.154
R3240 GND.n983 GND.n982 9.154
R3241 GND.n824 GND.n823 9.154
R3242 GND.n823 GND.n822 9.154
R3243 GND.n989 GND.n988 9.154
R3244 GND.n990 GND.n989 9.154
R3245 GND.n821 GND.n820 9.154
R3246 GND.n991 GND.n821 9.154
R3247 GND.n994 GND.n993 9.154
R3248 GND.n993 GND.n992 9.154
R3249 GND.n818 GND.n817 9.154
R3250 GND.n817 GND.n816 9.154
R3251 GND.n1000 GND.n999 9.154
R3252 GND.n1001 GND.n1000 9.154
R3253 GND.n815 GND.n814 9.154
R3254 GND.n1002 GND.n815 9.154
R3255 GND.n1005 GND.n1004 9.154
R3256 GND.n1004 GND.n1003 9.154
R3257 GND.n812 GND.n811 9.154
R3258 GND.n811 GND.n810 9.154
R3259 GND.n1013 GND.n1012 9.154
R3260 GND.n1014 GND.n1013 9.154
R3261 GND.n809 GND.n808 9.154
R3262 GND.n1015 GND.n809 9.154
R3263 GND.n1019 GND.n1018 9.154
R3264 GND.n1018 GND.n1017 9.154
R3265 GND.n807 GND.n806 9.154
R3266 GND.n1016 GND.n806 9.154
R3267 GND.n1025 GND.n1024 9.154
R3268 GND.n1026 GND.n1025 9.154
R3269 GND.n805 GND.n804 9.154
R3270 GND.n1027 GND.n805 9.154
R3271 GND.n1031 GND.n1030 9.154
R3272 GND.n1030 GND.n1029 9.154
R3273 GND.n802 GND.n801 9.154
R3274 GND.n1028 GND.n801 9.154
R3275 GND.n1036 GND.n1035 9.154
R3276 GND.n1037 GND.n1036 9.154
R3277 GND.n800 GND.n799 9.154
R3278 GND.n1038 GND.n800 9.154
R3279 GND.n1042 GND.n1041 9.154
R3280 GND.n1041 GND.n1040 9.154
R3281 GND.n797 GND.n796 9.154
R3282 GND.n1039 GND.n796 9.154
R3283 GND.n1048 GND.n1047 9.154
R3284 GND.n1049 GND.n1048 9.154
R3285 GND.n1046 GND.n795 9.154
R3286 GND.n1050 GND.n795 9.154
R3287 GND.n622 GND.n621 9.154
R3288 GND.n627 GND.n626 9.154
R3289 GND.n628 GND.n627 9.154
R3290 GND.n620 GND.n619 9.154
R3291 GND.n629 GND.n620 9.154
R3292 GND.n632 GND.n631 9.154
R3293 GND.n631 GND.n630 9.154
R3294 GND.n617 GND.n616 9.154
R3295 GND.n616 GND.n615 9.154
R3296 GND.n638 GND.n637 9.154
R3297 GND.n639 GND.n638 9.154
R3298 GND.n614 GND.n613 9.154
R3299 GND.n640 GND.n614 9.154
R3300 GND.n644 GND.n643 9.154
R3301 GND.n643 GND.n642 9.154
R3302 GND.n609 GND.n608 9.154
R3303 GND.n641 GND.n608 9.154
R3304 GND.n649 GND.n648 9.154
R3305 GND.n650 GND.n649 9.154
R3306 GND.n607 GND.n606 9.154
R3307 GND.n651 GND.n607 9.154
R3308 GND.n654 GND.n653 9.154
R3309 GND.n653 GND.n652 9.154
R3310 GND.n604 GND.n603 9.154
R3311 GND.n603 GND.n602 9.154
R3312 GND.n660 GND.n659 9.154
R3313 GND.n661 GND.n660 9.154
R3314 GND.n601 GND.n600 9.154
R3315 GND.n662 GND.n601 9.154
R3316 GND.n665 GND.n664 9.154
R3317 GND.n664 GND.n663 9.154
R3318 GND.n598 GND.n597 9.154
R3319 GND.n597 GND.n596 9.154
R3320 GND.n670 GND.n669 9.154
R3321 GND.n671 GND.n670 9.154
R3322 GND.n595 GND.n594 9.154
R3323 GND.n592 GND.n591 9.154
R3324 GND.n681 GND.n680 9.154
R3325 GND.n682 GND.n681 9.154
R3326 GND.n590 GND.n589 9.154
R3327 GND.n683 GND.n590 9.154
R3328 GND.n687 GND.n686 9.154
R3329 GND.n686 GND.n685 9.154
R3330 GND.n587 GND.n586 9.154
R3331 GND.n684 GND.n586 9.154
R3332 GND.n693 GND.n692 9.154
R3333 GND.n694 GND.n693 9.154
R3334 GND.n585 GND.n584 9.154
R3335 GND.n695 GND.n585 9.154
R3336 GND.n698 GND.n697 9.154
R3337 GND.n697 GND.n696 9.154
R3338 GND.n580 GND.n579 9.154
R3339 GND.n579 GND.n578 9.154
R3340 GND.n704 GND.n703 9.154
R3341 GND.n705 GND.n704 9.154
R3342 GND.n577 GND.n576 9.154
R3343 GND.n706 GND.n577 9.154
R3344 GND.n709 GND.n708 9.154
R3345 GND.n708 GND.n707 9.154
R3346 GND.n574 GND.n573 9.154
R3347 GND.n573 GND.n572 9.154
R3348 GND.n714 GND.n713 9.154
R3349 GND.n715 GND.n714 9.154
R3350 GND.n571 GND.n570 9.154
R3351 GND.n793 GND.n792 9.154
R3352 GND.n721 GND.n720 9.154
R3353 GND.n568 GND.n567 9.154
R3354 GND.n722 GND.n568 9.154
R3355 GND.n725 GND.n724 9.154
R3356 GND.n724 GND.n723 9.154
R3357 GND.n565 GND.n564 9.154
R3358 GND.n564 GND.n563 9.154
R3359 GND.n730 GND.n729 9.154
R3360 GND.n731 GND.n730 9.154
R3361 GND.n562 GND.n561 9.154
R3362 GND.n732 GND.n562 9.154
R3363 GND.n735 GND.n734 9.154
R3364 GND.n734 GND.n733 9.154
R3365 GND.n559 GND.n558 9.154
R3366 GND.n558 GND.n557 9.154
R3367 GND.n741 GND.n740 9.154
R3368 GND.n742 GND.n741 9.154
R3369 GND.n556 GND.n555 9.154
R3370 GND.n743 GND.n556 9.154
R3371 GND.n746 GND.n745 9.154
R3372 GND.n745 GND.n744 9.154
R3373 GND.n553 GND.n552 9.154
R3374 GND.n552 GND.n551 9.154
R3375 GND.n754 GND.n753 9.154
R3376 GND.n755 GND.n754 9.154
R3377 GND.n550 GND.n549 9.154
R3378 GND.n756 GND.n550 9.154
R3379 GND.n760 GND.n759 9.154
R3380 GND.n759 GND.n758 9.154
R3381 GND.n548 GND.n547 9.154
R3382 GND.n757 GND.n547 9.154
R3383 GND.n766 GND.n765 9.154
R3384 GND.n767 GND.n766 9.154
R3385 GND.n546 GND.n545 9.154
R3386 GND.n768 GND.n546 9.154
R3387 GND.n772 GND.n771 9.154
R3388 GND.n771 GND.n770 9.154
R3389 GND.n543 GND.n542 9.154
R3390 GND.n769 GND.n542 9.154
R3391 GND.n777 GND.n776 9.154
R3392 GND.n778 GND.n777 9.154
R3393 GND.n541 GND.n540 9.154
R3394 GND.n779 GND.n541 9.154
R3395 GND.n783 GND.n782 9.154
R3396 GND.n782 GND.n781 9.154
R3397 GND.n538 GND.n537 9.154
R3398 GND.n780 GND.n537 9.154
R3399 GND.n789 GND.n788 9.154
R3400 GND.n790 GND.n789 9.154
R3401 GND.n787 GND.n536 9.154
R3402 GND.n791 GND.n536 9.154
R3403 GND.n1660 GND.n1458 8.326
R3404 GND.n1532 GND.n1531 8.203
R3405 GND.n1667 GND.n1666 8.203
R3406 GND.n1763 GND.n1762 8.202
R3407 GND.n1659 GND.n1658 7.124
R3408 GND.n223 GND.n4 5.103
R3409 GND.n223 GND.n3 5.103
R3410 GND.n46 GND.n8 5.103
R3411 GND.n46 GND.n7 5.103
R3412 GND.n128 GND.n6 5.103
R3413 GND.n128 GND.n5 5.103
R3414 GND.n485 GND.n282 5.103
R3415 GND.n485 GND.n281 5.103
R3416 GND.n400 GND.n286 5.103
R3417 GND.n400 GND.n285 5.103
R3418 GND.n328 GND.n290 5.103
R3419 GND.n328 GND.n289 5.103
R3420 GND.n1829 GND.n1360 5.103
R3421 GND.n1830 GND.n1359 5.103
R3422 GND.n1703 GND.n1433 5.103
R3423 GND.n1715 GND.n1426 5.103
R3424 GND.n1588 GND.n1499 5.103
R3425 GND.n1599 GND.n1492 5.103
R3426 GND.n1285 GND.n1070 5.103
R3427 GND.n1230 GND.n1098 5.103
R3428 GND.n1176 GND.n1127 5.103
R3429 GND.n1010 GND.n1009 5.103
R3430 GND.n1010 GND.n1008 5.103
R3431 GND.n958 GND.n841 5.103
R3432 GND.n958 GND.n840 5.103
R3433 GND.n906 GND.n870 5.103
R3434 GND.n906 GND.n869 5.103
R3435 GND.n751 GND.n750 5.103
R3436 GND.n751 GND.n749 5.103
R3437 GND.n699 GND.n582 5.103
R3438 GND.n699 GND.n581 5.103
R3439 GND.n647 GND.n611 5.103
R3440 GND.n647 GND.n610 5.103
R3441 GND.n1545 GND.n1524 4.72
R3442 GND.n1549 GND.n1522 4.72
R3443 GND.n1555 GND.n1519 4.72
R3444 GND.n1559 GND.n1517 4.72
R3445 GND.n1565 GND.n1513 4.72
R3446 GND.n1570 GND.n1511 4.72
R3447 GND.n1576 GND.n1507 4.72
R3448 GND.n1580 GND.n1505 4.72
R3449 GND.n1586 GND.n1501 4.72
R3450 GND.n1590 GND.n1498 4.72
R3451 GND.n1596 GND.n1494 4.72
R3452 GND.n1600 GND.n1491 4.72
R3453 GND.n1606 GND.n1487 4.72
R3454 GND.n1610 GND.n1486 4.72
R3455 GND.n1616 GND.n1482 4.72
R3456 GND.n1621 GND.n1480 4.72
R3457 GND.n1627 GND.n1476 4.72
R3458 GND.n1631 GND.n1474 4.72
R3459 GND.n1638 GND.n1470 4.72
R3460 GND.n1642 GND.n1468 4.72
R3461 GND.n1649 GND.n1465 4.72
R3462 GND.n1656 GND.n1462 4.72
R3463 GND.n1652 GND.n1463 4.72
R3464 GND.n1661 GND.n1457 4.72
R3465 GND.n1538 GND.n1528 4.71
R3466 GND.n1534 GND.n1533 4.69
R3467 GND.n170 GND.n169 4.65
R3468 GND.n94 GND.n93 4.65
R3469 GND.n98 GND.n97 4.65
R3470 GND.n102 GND.n101 4.65
R3471 GND.n106 GND.n105 4.65
R3472 GND.n110 GND.n109 4.65
R3473 GND.n114 GND.n113 4.65
R3474 GND.n119 GND.n118 4.65
R3475 GND.n123 GND.n122 4.65
R3476 GND.n127 GND.n126 4.65
R3477 GND.n131 GND.n128 4.65
R3478 GND.n135 GND.n134 4.65
R3479 GND.n139 GND.n138 4.65
R3480 GND.n143 GND.n142 4.65
R3481 GND.n148 GND.n147 4.65
R3482 GND.n152 GND.n151 4.65
R3483 GND.n156 GND.n155 4.65
R3484 GND.n160 GND.n159 4.65
R3485 GND.n164 GND.n163 4.65
R3486 GND.n168 GND.n167 4.65
R3487 GND.n90 GND.n89 4.65
R3488 GND.n88 GND.n87 4.65
R3489 GND.n16 GND.n15 4.65
R3490 GND.n20 GND.n19 4.65
R3491 GND.n24 GND.n23 4.65
R3492 GND.n28 GND.n27 4.65
R3493 GND.n32 GND.n31 4.65
R3494 GND.n37 GND.n36 4.65
R3495 GND.n41 GND.n40 4.65
R3496 GND.n45 GND.n44 4.65
R3497 GND.n49 GND.n46 4.65
R3498 GND.n53 GND.n52 4.65
R3499 GND.n57 GND.n56 4.65
R3500 GND.n61 GND.n60 4.65
R3501 GND.n66 GND.n65 4.65
R3502 GND.n70 GND.n69 4.65
R3503 GND.n74 GND.n73 4.65
R3504 GND.n78 GND.n77 4.65
R3505 GND.n82 GND.n81 4.65
R3506 GND.n86 GND.n85 4.65
R3507 GND.n177 GND.n176 4.65
R3508 GND.n181 GND.n180 4.65
R3509 GND.n185 GND.n184 4.65
R3510 GND.n189 GND.n188 4.65
R3511 GND.n193 GND.n192 4.65
R3512 GND.n197 GND.n196 4.65
R3513 GND.n201 GND.n200 4.65
R3514 GND.n205 GND.n204 4.65
R3515 GND.n209 GND.n208 4.65
R3516 GND.n214 GND.n213 4.65
R3517 GND.n218 GND.n217 4.65
R3518 GND.n222 GND.n221 4.65
R3519 GND.n226 GND.n223 4.65
R3520 GND.n230 GND.n229 4.65
R3521 GND.n234 GND.n233 4.65
R3522 GND.n238 GND.n237 4.65
R3523 GND.n243 GND.n242 4.65
R3524 GND.n247 GND.n246 4.65
R3525 GND.n251 GND.n250 4.65
R3526 GND.n255 GND.n254 4.65
R3527 GND.n259 GND.n258 4.65
R3528 GND.n263 GND.n262 4.65
R3529 GND.n267 GND.n266 4.65
R3530 GND.n271 GND.n270 4.65
R3531 GND.n173 GND.n172 4.65
R3532 GND.n298 GND.n297 4.65
R3533 GND.n302 GND.n301 4.65
R3534 GND.n306 GND.n305 4.65
R3535 GND.n310 GND.n309 4.65
R3536 GND.n314 GND.n313 4.65
R3537 GND.n319 GND.n318 4.65
R3538 GND.n323 GND.n322 4.65
R3539 GND.n327 GND.n326 4.65
R3540 GND.n329 GND.n328 4.65
R3541 GND.n333 GND.n332 4.65
R3542 GND.n337 GND.n336 4.65
R3543 GND.n341 GND.n340 4.65
R3544 GND.n346 GND.n345 4.65
R3545 GND.n350 GND.n349 4.65
R3546 GND.n354 GND.n353 4.65
R3547 GND.n358 GND.n357 4.65
R3548 GND.n362 GND.n361 4.65
R3549 GND.n366 GND.n365 4.65
R3550 GND.n368 GND.n367 4.65
R3551 GND.n370 GND.n369 4.65
R3552 GND.n374 GND.n373 4.65
R3553 GND.n378 GND.n377 4.65
R3554 GND.n382 GND.n381 4.65
R3555 GND.n386 GND.n385 4.65
R3556 GND.n391 GND.n390 4.65
R3557 GND.n395 GND.n394 4.65
R3558 GND.n399 GND.n398 4.65
R3559 GND.n401 GND.n400 4.65
R3560 GND.n405 GND.n404 4.65
R3561 GND.n409 GND.n408 4.65
R3562 GND.n413 GND.n412 4.65
R3563 GND.n418 GND.n417 4.65
R3564 GND.n422 GND.n421 4.65
R3565 GND.n426 GND.n425 4.65
R3566 GND.n430 GND.n429 4.65
R3567 GND.n432 GND.n431 4.65
R3568 GND.n435 GND.n434 4.65
R3569 GND.n439 GND.n438 4.65
R3570 GND.n443 GND.n442 4.65
R3571 GND.n447 GND.n446 4.65
R3572 GND.n451 GND.n450 4.65
R3573 GND.n455 GND.n454 4.65
R3574 GND.n459 GND.n458 4.65
R3575 GND.n463 GND.n462 4.65
R3576 GND.n467 GND.n466 4.65
R3577 GND.n471 GND.n470 4.65
R3578 GND.n476 GND.n475 4.65
R3579 GND.n480 GND.n479 4.65
R3580 GND.n484 GND.n483 4.65
R3581 GND.n486 GND.n485 4.65
R3582 GND.n490 GND.n489 4.65
R3583 GND.n494 GND.n493 4.65
R3584 GND.n498 GND.n497 4.65
R3585 GND.n503 GND.n502 4.65
R3586 GND.n507 GND.n506 4.65
R3587 GND.n511 GND.n510 4.65
R3588 GND.n515 GND.n514 4.65
R3589 GND.n519 GND.n518 4.65
R3590 GND.n523 GND.n522 4.65
R3591 GND.n527 GND.n526 4.65
R3592 GND.n531 GND.n530 4.65
R3593 GND.n1758 GND.n1757 4.65
R3594 GND.n1670 GND.n1669 4.65
R3595 GND.n1663 GND.n1453 4.65
R3596 GND.n1749 GND.n1407 4.65
R3597 GND.n1402 GND.n1401 4.65
R3598 GND.n1538 GND.n1537 4.65
R3599 GND.n1487 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/GND 4.65
R3600 GND.n1654 GND.n1463 4.65
R3601 GND.n1457 GND.n1456 4.65
R3602 GND.n1535 GND.n1534 4.65
R3603 GND.n1536 GND.n1528 4.65
R3604 GND.n1546 GND.n1545 4.65
R3605 GND.n1549 GND.n1548 4.65
R3606 GND.n1556 GND.n1555 4.65
R3607 GND.n1559 GND.n1558 4.65
R3608 GND.n1566 GND.n1565 4.65
R3609 GND.n1570 GND.n1569 4.65
R3610 GND.n1577 GND.n1576 4.65
R3611 GND.n1580 GND.n1579 4.65
R3612 GND.n1587 GND.n1586 4.65
R3613 GND.n1590 GND.n1589 4.65
R3614 GND.n1597 GND.n1596 4.65
R3615 GND.n1600 GND.n1599 4.65
R3616 GND.n1607 GND.n1606 4.65
R3617 GND.n1610 GND.n1609 4.65
R3618 GND.n1617 GND.n1616 4.65
R3619 GND.n1621 GND.n1620 4.65
R3620 GND.n1628 GND.n1627 4.65
R3621 GND.n1631 GND.n1630 4.65
R3622 GND.n1639 GND.n1638 4.65
R3623 GND.n1642 GND.n1641 4.65
R3624 GND.n1650 GND.n1649 4.65
R3625 GND.n1524 GND.n1523 4.65
R3626 GND.n1547 GND.n1522 4.65
R3627 GND.n1519 GND.n1518 4.65
R3628 GND.n1557 GND.n1517 4.65
R3629 GND.n1513 GND.n1512 4.65
R3630 GND.n1567 GND.n1511 4.65
R3631 GND.n1507 GND.n1506 4.65
R3632 GND.n1578 GND.n1505 4.65
R3633 GND.n1501 GND.n1500 4.65
R3634 GND.n1588 GND.n1498 4.65
R3635 GND.n1494 GND.n1493 4.65
R3636 GND.n1598 GND.n1491 4.65
R3637 GND.n1608 GND.n1486 4.65
R3638 GND.n1482 GND.n1481 4.65
R3639 GND.n1618 GND.n1480 4.65
R3640 GND.n1476 GND.n1475 4.65
R3641 GND.n1629 GND.n1474 4.65
R3642 GND.n1470 GND.n1469 4.65
R3643 GND.n1640 GND.n1468 4.65
R3644 GND.n1465 GND.n1464 4.65
R3645 GND.n1651 GND.n1462 4.65
R3646 GND.n1656 GND.n1655 4.65
R3647 GND.n1653 GND.n1652 4.65
R3648 GND.n1662 GND.n1661 4.65
R3649 GND.n1665 GND.n1664 4.65
R3650 GND.n1668 GND.n1452 4.65
R3651 GND.n1680 GND.n1679 4.65
R3652 GND.n1684 GND.n1683 4.65
R3653 GND.n1691 GND.n1690 4.65
R3654 GND.n1695 GND.n1694 4.65
R3655 GND.n1702 GND.n1701 4.65
R3656 GND.n1705 GND.n1704 4.65
R3657 GND.n1713 GND.n1712 4.65
R3658 GND.n1716 GND.n1715 4.65
R3659 GND.n1723 GND.n1722 4.65
R3660 GND.n1727 GND.n1726 4.65
R3661 GND.n1734 GND.n1733 4.65
R3662 GND.n1738 GND.n1737 4.65
R3663 GND.n1745 GND.n1744 4.65
R3664 GND.n1751 GND.n1750 4.65
R3665 GND.n1748 GND.n1747 4.65
R3666 GND.n1673 GND.n1672 4.65
R3667 GND.n1671 GND.n1451 4.65
R3668 GND.n1447 GND.n1446 4.65
R3669 GND.n1681 GND.n1445 4.65
R3670 GND.n1441 GND.n1440 4.65
R3671 GND.n1692 GND.n1439 4.65
R3672 GND.n1435 GND.n1434 4.65
R3673 GND.n1703 GND.n1432 4.65
R3674 GND.n1428 GND.n1427 4.65
R3675 GND.n1714 GND.n1425 4.65
R3676 GND.n1421 GND.n1420 4.65
R3677 GND.n1725 GND.n1419 4.65
R3678 GND.n1415 GND.n1414 4.65
R3679 GND.n1735 GND.n1413 4.65
R3680 GND.n1409 GND.n1408 4.65
R3681 GND.n1746 GND.n1406 4.65
R3682 GND.n1766 GND.n1765 4.65
R3683 GND.n1769 GND.n1768 4.65
R3684 GND.n1776 GND.n1775 4.65
R3685 GND.n1779 GND.n1778 4.65
R3686 GND.n1786 GND.n1785 4.65
R3687 GND.n1789 GND.n1788 4.65
R3688 GND.n1796 GND.n1795 4.65
R3689 GND.n1799 GND.n1798 4.65
R3690 GND.n1806 GND.n1805 4.65
R3691 GND.n1811 GND.n1810 4.65
R3692 GND.n1818 GND.n1817 4.65
R3693 GND.n1821 GND.n1820 4.65
R3694 GND.n1828 GND.n1827 4.65
R3695 GND.n1831 GND.n1830 4.65
R3696 GND.n1838 GND.n1837 4.65
R3697 GND.n1841 GND.n1840 4.65
R3698 GND.n1848 GND.n1847 4.65
R3699 GND.n1853 GND.n1852 4.65
R3700 GND.n1860 GND.n1859 4.65
R3701 GND.n1863 GND.n1862 4.65
R3702 GND.n1870 GND.n1869 4.65
R3703 GND.n1873 GND.n1872 4.65
R3704 GND.n1880 GND.n1879 4.65
R3705 GND.n1883 GND.n1882 4.65
R3706 GND.n1890 GND.n1889 4.65
R3707 GND.n1893 GND.n1892 4.65
R3708 GND.n1759 GND.n1398 4.65
R3709 GND.n1761 GND.n1760 4.65
R3710 GND.n1764 GND.n1397 4.65
R3711 GND.n1767 GND.n1396 4.65
R3712 GND.n1392 GND.n1391 4.65
R3713 GND.n1777 GND.n1390 4.65
R3714 GND.n1386 GND.n1385 4.65
R3715 GND.n1787 GND.n1384 4.65
R3716 GND.n1380 GND.n1379 4.65
R3717 GND.n1797 GND.n1378 4.65
R3718 GND.n1374 GND.n1373 4.65
R3719 GND.n1807 GND.n1372 4.65
R3720 GND.n1368 GND.n1367 4.65
R3721 GND.n1819 GND.n1366 4.65
R3722 GND.n1362 GND.n1361 4.65
R3723 GND.n1829 GND.n1358 4.65
R3724 GND.n1354 GND.n1353 4.65
R3725 GND.n1839 GND.n1352 4.65
R3726 GND.n1348 GND.n1347 4.65
R3727 GND.n1850 GND.n1346 4.65
R3728 GND.n1342 GND.n1341 4.65
R3729 GND.n1861 GND.n1340 4.65
R3730 GND.n1336 GND.n1335 4.65
R3731 GND.n1871 GND.n1334 4.65
R3732 GND.n1330 GND.n1329 4.65
R3733 GND.n1881 GND.n1328 4.65
R3734 GND.n1324 GND.n1323 4.65
R3735 GND.n1891 GND.n1321 4.65
R3736 GND.n1146 GND.n1145 4.65
R3737 GND.n1139 GND.n1138 4.65
R3738 GND.n1154 GND.n1153 4.65
R3739 GND.n1155 GND.n1137 4.65
R3740 GND.n1157 GND.n1156 4.65
R3741 GND.n1134 GND.n1133 4.65
R3742 GND.n1165 GND.n1164 4.65
R3743 GND.n1167 GND.n1132 4.65
R3744 GND.n1169 GND.n1168 4.65
R3745 GND.n1129 GND.n1128 4.65
R3746 GND.n1176 GND.n1175 4.65
R3747 GND.n1177 GND.n1126 4.65
R3748 GND.n1180 GND.n1179 4.65
R3749 GND.n1178 GND.n1122 4.65
R3750 GND.n1187 GND.n1186 4.65
R3751 GND.n1188 GND.n1120 4.65
R3752 GND.n1190 GND.n1189 4.65
R3753 GND.n1116 GND.n1115 4.65
R3754 GND.n1197 GND.n1196 4.65
R3755 GND.n1198 GND.n1114 4.65
R3756 GND.n1200 GND.n1199 4.65
R3757 GND.n1110 GND.n1109 4.65
R3758 GND.n1205 GND.n1204 4.65
R3759 GND.n1208 GND.n1207 4.65
R3760 GND.n1209 GND.n1108 4.65
R3761 GND.n1211 GND.n1210 4.65
R3762 GND.n1105 GND.n1104 4.65
R3763 GND.n1219 GND.n1218 4.65
R3764 GND.n1221 GND.n1103 4.65
R3765 GND.n1223 GND.n1222 4.65
R3766 GND.n1100 GND.n1099 4.65
R3767 GND.n1230 GND.n1229 4.65
R3768 GND.n1231 GND.n1097 4.65
R3769 GND.n1234 GND.n1233 4.65
R3770 GND.n1232 GND.n1093 4.65
R3771 GND.n1241 GND.n1240 4.65
R3772 GND.n1242 GND.n1091 4.65
R3773 GND.n1244 GND.n1243 4.65
R3774 GND.n1087 GND.n1086 4.65
R3775 GND.n1249 GND.n1248 4.65
R3776 GND.n1252 GND.n1251 4.65
R3777 GND.n1253 GND.n1085 4.65
R3778 GND.n1255 GND.n1254 4.65
R3779 GND.n1082 GND.n1081 4.65
R3780 GND.n1263 GND.n1262 4.65
R3781 GND.n1264 GND.n1080 4.65
R3782 GND.n1266 GND.n1265 4.65
R3783 GND.n1077 GND.n1076 4.65
R3784 GND.n1274 GND.n1273 4.65
R3785 GND.n1276 GND.n1075 4.65
R3786 GND.n1278 GND.n1277 4.65
R3787 GND.n1072 GND.n1071 4.65
R3788 GND.n1285 GND.n1284 4.65
R3789 GND.n1286 GND.n1069 4.65
R3790 GND.n1289 GND.n1288 4.65
R3791 GND.n1287 GND.n1065 4.65
R3792 GND.n1296 GND.n1295 4.65
R3793 GND.n1297 GND.n1063 4.65
R3794 GND.n1299 GND.n1298 4.65
R3795 GND.n1059 GND.n1058 4.65
R3796 GND.n1306 GND.n1305 4.65
R3797 GND.n1307 GND.n1057 4.65
R3798 GND.n1310 GND.n1308 4.65
R3799 GND.n885 GND.n884 4.65
R3800 GND.n878 GND.n877 4.65
R3801 GND.n892 GND.n891 4.65
R3802 GND.n893 GND.n876 4.65
R3803 GND.n896 GND.n895 4.65
R3804 GND.n872 GND.n871 4.65
R3805 GND.n904 GND.n903 4.65
R3806 GND.n905 GND.n868 4.65
R3807 GND.n907 GND.n906 4.65
R3808 GND.n865 GND.n864 4.65
R3809 GND.n914 GND.n913 4.65
R3810 GND.n915 GND.n863 4.65
R3811 GND.n918 GND.n917 4.65
R3812 GND.n859 GND.n858 4.65
R3813 GND.n925 GND.n924 4.65
R3814 GND.n926 GND.n857 4.65
R3815 GND.n928 GND.n927 4.65
R3816 GND.n853 GND.n852 4.65
R3817 GND.n933 GND.n932 4.65
R3818 GND.n936 GND.n935 4.65
R3819 GND.n937 GND.n851 4.65
R3820 GND.n939 GND.n938 4.65
R3821 GND.n848 GND.n847 4.65
R3822 GND.n947 GND.n946 4.65
R3823 GND.n949 GND.n846 4.65
R3824 GND.n951 GND.n950 4.65
R3825 GND.n843 GND.n842 4.65
R3826 GND.n958 GND.n957 4.65
R3827 GND.n959 GND.n839 4.65
R3828 GND.n962 GND.n961 4.65
R3829 GND.n960 GND.n835 4.65
R3830 GND.n969 GND.n968 4.65
R3831 GND.n970 GND.n833 4.65
R3832 GND.n972 GND.n971 4.65
R3833 GND.n829 GND.n828 4.65
R3834 GND.n977 GND.n976 4.65
R3835 GND.n979 GND.n978 4.65
R3836 GND.n826 GND.n825 4.65
R3837 GND.n985 GND.n984 4.65
R3838 GND.n986 GND.n824 4.65
R3839 GND.n988 GND.n987 4.65
R3840 GND.n820 GND.n819 4.65
R3841 GND.n995 GND.n994 4.65
R3842 GND.n996 GND.n818 4.65
R3843 GND.n999 GND.n998 4.65
R3844 GND.n997 GND.n814 4.65
R3845 GND.n1006 GND.n1005 4.65
R3846 GND.n1007 GND.n812 4.65
R3847 GND.n1012 GND.n1011 4.65
R3848 GND.n1010 GND.n808 4.65
R3849 GND.n1020 GND.n1019 4.65
R3850 GND.n1021 GND.n807 4.65
R3851 GND.n1024 GND.n1023 4.65
R3852 GND.n804 GND.n803 4.65
R3853 GND.n1032 GND.n1031 4.65
R3854 GND.n1033 GND.n802 4.65
R3855 GND.n1035 GND.n1034 4.65
R3856 GND.n799 GND.n798 4.65
R3857 GND.n1043 GND.n1042 4.65
R3858 GND.n1044 GND.n797 4.65
R3859 GND.n1047 GND.n1045 4.65
R3860 GND.n626 GND.n625 4.65
R3861 GND.n619 GND.n618 4.65
R3862 GND.n633 GND.n632 4.65
R3863 GND.n634 GND.n617 4.65
R3864 GND.n637 GND.n636 4.65
R3865 GND.n613 GND.n612 4.65
R3866 GND.n645 GND.n644 4.65
R3867 GND.n646 GND.n609 4.65
R3868 GND.n648 GND.n647 4.65
R3869 GND.n606 GND.n605 4.65
R3870 GND.n655 GND.n654 4.65
R3871 GND.n656 GND.n604 4.65
R3872 GND.n659 GND.n658 4.65
R3873 GND.n600 GND.n599 4.65
R3874 GND.n666 GND.n665 4.65
R3875 GND.n667 GND.n598 4.65
R3876 GND.n669 GND.n668 4.65
R3877 GND.n594 GND.n593 4.65
R3878 GND.n674 GND.n673 4.65
R3879 GND.n677 GND.n676 4.65
R3880 GND.n678 GND.n592 4.65
R3881 GND.n680 GND.n679 4.65
R3882 GND.n589 GND.n588 4.65
R3883 GND.n688 GND.n687 4.65
R3884 GND.n690 GND.n587 4.65
R3885 GND.n692 GND.n691 4.65
R3886 GND.n584 GND.n583 4.65
R3887 GND.n699 GND.n698 4.65
R3888 GND.n700 GND.n580 4.65
R3889 GND.n703 GND.n702 4.65
R3890 GND.n701 GND.n576 4.65
R3891 GND.n710 GND.n709 4.65
R3892 GND.n711 GND.n574 4.65
R3893 GND.n713 GND.n712 4.65
R3894 GND.n570 GND.n569 4.65
R3895 GND.n718 GND.n717 4.65
R3896 GND.n720 GND.n719 4.65
R3897 GND.n567 GND.n566 4.65
R3898 GND.n726 GND.n725 4.65
R3899 GND.n727 GND.n565 4.65
R3900 GND.n729 GND.n728 4.65
R3901 GND.n561 GND.n560 4.65
R3902 GND.n736 GND.n735 4.65
R3903 GND.n737 GND.n559 4.65
R3904 GND.n740 GND.n739 4.65
R3905 GND.n738 GND.n555 4.65
R3906 GND.n747 GND.n746 4.65
R3907 GND.n748 GND.n553 4.65
R3908 GND.n753 GND.n752 4.65
R3909 GND.n751 GND.n549 4.65
R3910 GND.n761 GND.n760 4.65
R3911 GND.n762 GND.n548 4.65
R3912 GND.n765 GND.n764 4.65
R3913 GND.n545 GND.n544 4.65
R3914 GND.n773 GND.n772 4.65
R3915 GND.n774 GND.n543 4.65
R3916 GND.n776 GND.n775 4.65
R3917 GND.n540 GND.n539 4.65
R3918 GND.n784 GND.n783 4.65
R3919 GND.n785 GND.n538 4.65
R3920 GND.n788 GND.n786 4.65
R3921 GND.n1898 GND.n1316 4.467
R3922 EESPFAL_s1_0/GND GND.n1898 4.432
R3923 EESPFAL_s2_0/GND GND.n1315 4.379
R3924 EESPFAL_s0_0/GND GND.n1899 4.37
R3925 GND.n1764 GND.n1398 3.28
R3926 GND.n1765 GND.n1396 3.28
R3927 GND.n1769 GND.n1392 3.28
R3928 GND.n1775 GND.n1390 3.28
R3929 GND.n1779 GND.n1386 3.28
R3930 GND.n1785 GND.n1384 3.28
R3931 GND.n1789 GND.n1380 3.28
R3932 GND.n1795 GND.n1378 3.28
R3933 GND.n1799 GND.n1374 3.28
R3934 GND.n1805 GND.n1372 3.28
R3935 GND.n1811 GND.n1368 3.28
R3936 GND.n1817 GND.n1366 3.28
R3937 GND.n1821 GND.n1362 3.28
R3938 GND.n1827 GND.n1358 3.28
R3939 GND.n1831 GND.n1354 3.28
R3940 GND.n1837 GND.n1352 3.28
R3941 GND.n1841 GND.n1348 3.28
R3942 GND.n1847 GND.n1346 3.28
R3943 GND.n1853 GND.n1342 3.28
R3944 GND.n1859 GND.n1340 3.28
R3945 GND.n1863 GND.n1336 3.28
R3946 GND.n1869 GND.n1334 3.28
R3947 GND.n1873 GND.n1330 3.28
R3948 GND.n1879 GND.n1328 3.28
R3949 GND.n1883 GND.n1324 3.28
R3950 GND.n1889 GND.n1321 3.28
R3951 GND.n1893 GND.n1322 3.28
R3952 GND.n1665 GND.n1453 3.18
R3953 GND.n1668 GND.n1453 3.18
R3954 GND.n1669 GND.n1668 3.18
R3955 GND.n1669 GND.n1451 3.18
R3956 GND.n1673 GND.n1451 3.18
R3957 GND.n1673 GND.n1447 3.18
R3958 GND.n1679 GND.n1447 3.18
R3959 GND.n1679 GND.n1445 3.18
R3960 GND.n1684 GND.n1445 3.18
R3961 GND.n1684 GND.n1441 3.18
R3962 GND.n1690 GND.n1441 3.18
R3963 GND.n1690 GND.n1439 3.18
R3964 GND.n1695 GND.n1439 3.18
R3965 GND.n1695 GND.n1435 3.18
R3966 GND.n1701 GND.n1435 3.18
R3967 GND.n1701 GND.n1432 3.18
R3968 GND.n1705 GND.n1432 3.18
R3969 GND.n1705 GND.n1428 3.18
R3970 GND.n1712 GND.n1428 3.18
R3971 GND.n1712 GND.n1425 3.18
R3972 GND.n1716 GND.n1425 3.18
R3973 GND.n1716 GND.n1421 3.18
R3974 GND.n1722 GND.n1421 3.18
R3975 GND.n1722 GND.n1419 3.18
R3976 GND.n1727 GND.n1419 3.18
R3977 GND.n1727 GND.n1415 3.18
R3978 GND.n1733 GND.n1415 3.18
R3979 GND.n1733 GND.n1413 3.18
R3980 GND.n1738 GND.n1413 3.18
R3981 GND.n1738 GND.n1409 3.18
R3982 GND.n1744 GND.n1409 3.18
R3983 GND.n1744 GND.n1406 3.18
R3984 GND.n1751 GND.n1406 3.18
R3985 GND.n1751 GND.n1407 3.18
R3986 GND.n1747 GND.n1407 3.18
R3987 GND.n1747 GND.n1402 3.18
R3988 GND.n1757 GND.n1402 3.18
R3989 GND.n1761 GND.n1398 3.12
R3990 GND.n1765 GND.n1764 3.12
R3991 GND.n1769 GND.n1396 3.12
R3992 GND.n1775 GND.n1392 3.12
R3993 GND.n1779 GND.n1390 3.12
R3994 GND.n1785 GND.n1386 3.12
R3995 GND.n1789 GND.n1384 3.12
R3996 GND.n1795 GND.n1380 3.12
R3997 GND.n1799 GND.n1378 3.12
R3998 GND.n1805 GND.n1374 3.12
R3999 GND.n1811 GND.n1372 3.12
R4000 GND.n1817 GND.n1368 3.12
R4001 GND.n1821 GND.n1366 3.12
R4002 GND.n1827 GND.n1362 3.12
R4003 GND.n1831 GND.n1358 3.12
R4004 GND.n1837 GND.n1354 3.12
R4005 GND.n1841 GND.n1352 3.12
R4006 GND.n1847 GND.n1348 3.12
R4007 GND.n1853 GND.n1346 3.12
R4008 GND.n1859 GND.n1342 3.12
R4009 GND.n1863 GND.n1340 3.12
R4010 GND.n1869 GND.n1336 3.12
R4011 GND.n1873 GND.n1334 3.12
R4012 GND.n1879 GND.n1330 3.12
R4013 GND.n1883 GND.n1328 3.12
R4014 GND.n1889 GND.n1324 3.12
R4015 GND.n1893 GND.n1321 3.12
R4016 GND.n292 GND.n291 2.791
R4017 GND.n372 GND.n371 2.791
R4018 GND.n882 GND.n880 2.791
R4019 GND.n934 GND.n850 2.791
R4020 GND.n623 GND.n621 2.791
R4021 GND.n675 GND.n591 2.791
R4022 GND.n10 GND.n9 2.791
R4023 GND.n92 GND.n91 2.791
R4024 GND.n166 GND.n165 2.791
R4025 GND.n84 GND.n83 2.791
R4026 GND.n364 GND.n363 2.791
R4027 GND.n428 GND.n427 2.791
R4028 GND.n931 GND.n854 2.791
R4029 GND.n975 GND.n830 2.791
R4030 GND.n672 GND.n595 2.791
R4031 GND.n716 GND.n571 2.791
R4032 GND.n274 GND.n272 2.739
R4033 GND.n534 GND.n532 2.739
R4034 GND.n1314 GND.n1053 2.739
R4035 GND.n1052 GND.n794 2.739
R4036 GND.n793 GND.n535 2.739
R4037 GND.n294 GND.n293 2.682
R4038 GND.n1144 GND.n1142 2.682
R4039 GND.n883 GND.n881 2.682
R4040 GND.n624 GND.n622 2.682
R4041 GND.n12 GND.n11 2.682
R4042 GND.n272 GND.n2 2.682
R4043 GND.n532 GND.n278 2.682
R4044 GND.n1309 GND.n1053 2.682
R4045 GND.n1046 GND.n794 2.682
R4046 GND.n787 GND.n535 2.682
R4047 GND.n1658 GND.n1657 1.92
R4048 GND.n1897 GND.n1317 1.912
R4049 GND.n1322 GND.n1317 1.889
R4050 GND.n1143 GND.n1141 1.873
R4051 GND.n1206 GND.n1107 1.873
R4052 GND.n1313 GND.n1054 1.873
R4053 GND.n1203 GND.n1111 1.873
R4054 GND.n1247 GND.n1088 1.873
R4055 GND.n1250 GND.n1084 1.873
R4056 GND.n1538 GND.n1524 1.68
R4057 GND.n1545 GND.n1522 1.68
R4058 GND.n1549 GND.n1519 1.68
R4059 GND.n1555 GND.n1517 1.68
R4060 GND.n1559 GND.n1513 1.68
R4061 GND.n1565 GND.n1511 1.68
R4062 GND.n1570 GND.n1507 1.68
R4063 GND.n1576 GND.n1505 1.68
R4064 GND.n1580 GND.n1501 1.68
R4065 GND.n1586 GND.n1498 1.68
R4066 GND.n1590 GND.n1494 1.68
R4067 GND.n1596 GND.n1491 1.68
R4068 GND.n1600 GND.n1487 1.68
R4069 GND.n1606 GND.n1486 1.68
R4070 GND.n1610 GND.n1482 1.68
R4071 GND.n1616 GND.n1480 1.68
R4072 GND.n1621 GND.n1476 1.68
R4073 GND.n1627 GND.n1474 1.68
R4074 GND.n1631 GND.n1470 1.68
R4075 GND.n1638 GND.n1468 1.68
R4076 GND.n1642 GND.n1465 1.68
R4077 GND.n1649 GND.n1462 1.68
R4078 GND.n1656 GND.n1463 1.68
R4079 GND.n1652 GND.n1457 1.68
R4080 GND.n1534 GND.n1528 1.669
R4081 GND.n1533 GND.n1529 1.588
R4082 GND.n275 GND 1.565
R4083 GND.n1892 GND.n1317 1.417
R4084 GND.n298 GND.n294 1.096
R4085 GND.n1145 GND.n1144 1.096
R4086 GND.n884 GND.n883 1.096
R4087 GND.n625 GND.n624 1.096
R4088 GND.n16 GND.n12 1.095
R4089 GND.n272 GND.n271 1.095
R4090 GND.n532 GND.n531 1.095
R4091 GND.n1308 GND.n1053 1.095
R4092 GND.n1045 GND.n794 1.095
R4093 GND.n786 GND.n535 1.095
R4094 GND.n1535 GND.n1529 0.813
R4095 GND.n719 GND.n718 0.662
R4096 GND.n435 GND.n432 0.637
R4097 GND.n978 GND.n977 0.637
R4098 GND.n173 GND.n170 0.6
R4099 GND.n1252 GND.n1249 0.562
R4100 GND.n370 GND.n368 0.55
R4101 GND.n1208 GND.n1205 0.55
R4102 GND.n936 GND.n933 0.55
R4103 GND.n677 GND.n674 0.548
R4104 GND.n90 GND.n88 0.525
R4105 GND.n1660 GND.n1659 0.484
R4106 GND.n1531 GND.n1530 0.477
R4107 GND.n1666 GND.n1455 0.477
R4108 GND.n1762 GND.n1400 0.477
R4109 GND.n1896 GND.n1318 0.196
R4110 GND.n1760 GND.n1758 0.172
R4111 GND.n1664 GND.n1662 0.165
R4112 GND.n20 GND.n16 0.1
R4113 GND.n24 GND.n20 0.1
R4114 GND.n28 GND.n24 0.1
R4115 GND.n32 GND.n28 0.1
R4116 GND.n41 GND.n37 0.1
R4117 GND.n45 GND.n41 0.1
R4118 GND.n46 GND.n45 0.1
R4119 GND.n57 GND.n53 0.1
R4120 GND.n61 GND.n57 0.1
R4121 GND.n70 GND.n66 0.1
R4122 GND.n74 GND.n70 0.1
R4123 GND.n78 GND.n74 0.1
R4124 GND.n82 GND.n78 0.1
R4125 GND.n86 GND.n82 0.1
R4126 GND.n88 GND.n86 0.1
R4127 GND.n94 GND.n90 0.1
R4128 GND.n98 GND.n94 0.1
R4129 GND.n102 GND.n98 0.1
R4130 GND.n106 GND.n102 0.1
R4131 GND.n110 GND.n106 0.1
R4132 GND.n114 GND.n110 0.1
R4133 GND.n123 GND.n119 0.1
R4134 GND.n127 GND.n123 0.1
R4135 GND.n128 GND.n127 0.1
R4136 GND.n139 GND.n135 0.1
R4137 GND.n143 GND.n139 0.1
R4138 GND.n152 GND.n148 0.1
R4139 GND.n156 GND.n152 0.1
R4140 GND.n160 GND.n156 0.1
R4141 GND.n164 GND.n160 0.1
R4142 GND.n168 GND.n164 0.1
R4143 GND.n170 GND.n168 0.1
R4144 GND.n177 GND.n173 0.1
R4145 GND.n181 GND.n177 0.1
R4146 GND.n185 GND.n181 0.1
R4147 GND.n189 GND.n185 0.1
R4148 GND.n193 GND.n189 0.1
R4149 GND.n197 GND.n193 0.1
R4150 GND.n201 GND.n197 0.1
R4151 GND.n205 GND.n201 0.1
R4152 GND.n209 GND.n205 0.1
R4153 GND.n218 GND.n214 0.1
R4154 GND.n222 GND.n218 0.1
R4155 GND.n223 GND.n222 0.1
R4156 GND.n234 GND.n230 0.1
R4157 GND.n238 GND.n234 0.1
R4158 GND.n247 GND.n243 0.1
R4159 GND.n251 GND.n247 0.1
R4160 GND.n255 GND.n251 0.1
R4161 GND.n259 GND.n255 0.1
R4162 GND.n263 GND.n259 0.1
R4163 GND.n267 GND.n263 0.1
R4164 GND.n271 GND.n267 0.1
R4165 GND.n302 GND.n298 0.1
R4166 GND.n306 GND.n302 0.1
R4167 GND.n310 GND.n306 0.1
R4168 GND.n314 GND.n310 0.1
R4169 GND.n323 GND.n319 0.1
R4170 GND.n327 GND.n323 0.1
R4171 GND.n328 GND.n327 0.1
R4172 GND.n337 GND.n333 0.1
R4173 GND.n341 GND.n337 0.1
R4174 GND.n350 GND.n346 0.1
R4175 GND.n354 GND.n350 0.1
R4176 GND.n358 GND.n354 0.1
R4177 GND.n362 GND.n358 0.1
R4178 GND.n366 GND.n362 0.1
R4179 GND.n368 GND.n366 0.1
R4180 GND.n374 GND.n370 0.1
R4181 GND.n378 GND.n374 0.1
R4182 GND.n382 GND.n378 0.1
R4183 GND.n386 GND.n382 0.1
R4184 GND.n395 GND.n391 0.1
R4185 GND.n399 GND.n395 0.1
R4186 GND.n400 GND.n399 0.1
R4187 GND.n409 GND.n405 0.1
R4188 GND.n413 GND.n409 0.1
R4189 GND.n422 GND.n418 0.1
R4190 GND.n426 GND.n422 0.1
R4191 GND.n430 GND.n426 0.1
R4192 GND.n432 GND.n430 0.1
R4193 GND.n439 GND.n435 0.1
R4194 GND.n443 GND.n439 0.1
R4195 GND.n447 GND.n443 0.1
R4196 GND.n451 GND.n447 0.1
R4197 GND.n455 GND.n451 0.1
R4198 GND.n459 GND.n455 0.1
R4199 GND.n463 GND.n459 0.1
R4200 GND.n467 GND.n463 0.1
R4201 GND.n471 GND.n467 0.1
R4202 GND.n480 GND.n476 0.1
R4203 GND.n484 GND.n480 0.1
R4204 GND.n485 GND.n484 0.1
R4205 GND.n494 GND.n490 0.1
R4206 GND.n498 GND.n494 0.1
R4207 GND.n507 GND.n503 0.1
R4208 GND.n511 GND.n507 0.1
R4209 GND.n515 GND.n511 0.1
R4210 GND.n519 GND.n515 0.1
R4211 GND.n523 GND.n519 0.1
R4212 GND.n527 GND.n523 0.1
R4213 GND.n531 GND.n527 0.1
R4214 GND.n1145 GND.n1138 0.1
R4215 GND.n1154 GND.n1138 0.1
R4216 GND.n1155 GND.n1154 0.1
R4217 GND.n1156 GND.n1155 0.1
R4218 GND.n1156 GND.n1133 0.1
R4219 GND.n1165 GND.n1133 0.1
R4220 GND.n1168 GND.n1167 0.1
R4221 GND.n1168 GND.n1128 0.1
R4222 GND.n1176 GND.n1128 0.1
R4223 GND.n1179 GND.n1177 0.1
R4224 GND.n1179 GND.n1178 0.1
R4225 GND.n1188 GND.n1187 0.1
R4226 GND.n1189 GND.n1188 0.1
R4227 GND.n1189 GND.n1115 0.1
R4228 GND.n1197 GND.n1115 0.1
R4229 GND.n1198 GND.n1197 0.1
R4230 GND.n1199 GND.n1198 0.1
R4231 GND.n1199 GND.n1109 0.1
R4232 GND.n1205 GND.n1109 0.1
R4233 GND.n1209 GND.n1208 0.1
R4234 GND.n1210 GND.n1209 0.1
R4235 GND.n1210 GND.n1104 0.1
R4236 GND.n1219 GND.n1104 0.1
R4237 GND.n1222 GND.n1221 0.1
R4238 GND.n1222 GND.n1099 0.1
R4239 GND.n1230 GND.n1099 0.1
R4240 GND.n1233 GND.n1231 0.1
R4241 GND.n1233 GND.n1232 0.1
R4242 GND.n1242 GND.n1241 0.1
R4243 GND.n1243 GND.n1242 0.1
R4244 GND.n1243 GND.n1086 0.1
R4245 GND.n1249 GND.n1086 0.1
R4246 GND.n1253 GND.n1252 0.1
R4247 GND.n1254 GND.n1253 0.1
R4248 GND.n1254 GND.n1081 0.1
R4249 GND.n1263 GND.n1081 0.1
R4250 GND.n1264 GND.n1263 0.1
R4251 GND.n1265 GND.n1264 0.1
R4252 GND.n1265 GND.n1076 0.1
R4253 GND.n1274 GND.n1076 0.1
R4254 GND.n1277 GND.n1276 0.1
R4255 GND.n1277 GND.n1071 0.1
R4256 GND.n1285 GND.n1071 0.1
R4257 GND.n1288 GND.n1286 0.1
R4258 GND.n1288 GND.n1287 0.1
R4259 GND.n1297 GND.n1296 0.1
R4260 GND.n1298 GND.n1297 0.1
R4261 GND.n1298 GND.n1058 0.1
R4262 GND.n1306 GND.n1058 0.1
R4263 GND.n1307 GND.n1306 0.1
R4264 GND.n1308 GND.n1307 0.1
R4265 GND.n884 GND.n877 0.1
R4266 GND.n892 GND.n877 0.1
R4267 GND.n893 GND.n892 0.1
R4268 GND.n895 GND.n893 0.1
R4269 GND.n904 GND.n871 0.1
R4270 GND.n905 GND.n904 0.1
R4271 GND.n906 GND.n905 0.1
R4272 GND.n914 GND.n864 0.1
R4273 GND.n915 GND.n914 0.1
R4274 GND.n917 GND.n858 0.1
R4275 GND.n925 GND.n858 0.1
R4276 GND.n926 GND.n925 0.1
R4277 GND.n927 GND.n926 0.1
R4278 GND.n927 GND.n852 0.1
R4279 GND.n933 GND.n852 0.1
R4280 GND.n937 GND.n936 0.1
R4281 GND.n938 GND.n937 0.1
R4282 GND.n938 GND.n847 0.1
R4283 GND.n947 GND.n847 0.1
R4284 GND.n950 GND.n949 0.1
R4285 GND.n950 GND.n842 0.1
R4286 GND.n958 GND.n842 0.1
R4287 GND.n961 GND.n959 0.1
R4288 GND.n961 GND.n960 0.1
R4289 GND.n970 GND.n969 0.1
R4290 GND.n971 GND.n970 0.1
R4291 GND.n971 GND.n828 0.1
R4292 GND.n977 GND.n828 0.1
R4293 GND.n978 GND.n825 0.1
R4294 GND.n985 GND.n825 0.1
R4295 GND.n986 GND.n985 0.1
R4296 GND.n987 GND.n986 0.1
R4297 GND.n987 GND.n819 0.1
R4298 GND.n995 GND.n819 0.1
R4299 GND.n996 GND.n995 0.1
R4300 GND.n998 GND.n996 0.1
R4301 GND.n998 GND.n997 0.1
R4302 GND.n1007 GND.n1006 0.1
R4303 GND.n1011 GND.n1007 0.1
R4304 GND.n1011 GND.n1010 0.1
R4305 GND.n1021 GND.n1020 0.1
R4306 GND.n1023 GND.n1021 0.1
R4307 GND.n1032 GND.n803 0.1
R4308 GND.n1033 GND.n1032 0.1
R4309 GND.n1034 GND.n1033 0.1
R4310 GND.n1034 GND.n798 0.1
R4311 GND.n1043 GND.n798 0.1
R4312 GND.n1044 GND.n1043 0.1
R4313 GND.n1045 GND.n1044 0.1
R4314 GND.n625 GND.n618 0.1
R4315 GND.n633 GND.n618 0.1
R4316 GND.n634 GND.n633 0.1
R4317 GND.n636 GND.n634 0.1
R4318 GND.n645 GND.n612 0.1
R4319 GND.n646 GND.n645 0.1
R4320 GND.n647 GND.n646 0.1
R4321 GND.n655 GND.n605 0.1
R4322 GND.n656 GND.n655 0.1
R4323 GND.n658 GND.n599 0.1
R4324 GND.n666 GND.n599 0.1
R4325 GND.n667 GND.n666 0.1
R4326 GND.n668 GND.n667 0.1
R4327 GND.n668 GND.n593 0.1
R4328 GND.n674 GND.n593 0.1
R4329 GND.n678 GND.n677 0.1
R4330 GND.n679 GND.n678 0.1
R4331 GND.n679 GND.n588 0.1
R4332 GND.n688 GND.n588 0.1
R4333 GND.n691 GND.n690 0.1
R4334 GND.n691 GND.n583 0.1
R4335 GND.n699 GND.n583 0.1
R4336 GND.n702 GND.n700 0.1
R4337 GND.n702 GND.n701 0.1
R4338 GND.n711 GND.n710 0.1
R4339 GND.n712 GND.n711 0.1
R4340 GND.n712 GND.n569 0.1
R4341 GND.n718 GND.n569 0.1
R4342 GND.n719 GND.n566 0.1
R4343 GND.n726 GND.n566 0.1
R4344 GND.n727 GND.n726 0.1
R4345 GND.n728 GND.n727 0.1
R4346 GND.n728 GND.n560 0.1
R4347 GND.n736 GND.n560 0.1
R4348 GND.n737 GND.n736 0.1
R4349 GND.n739 GND.n737 0.1
R4350 GND.n739 GND.n738 0.1
R4351 GND.n748 GND.n747 0.1
R4352 GND.n752 GND.n748 0.1
R4353 GND.n752 GND.n751 0.1
R4354 GND.n762 GND.n761 0.1
R4355 GND.n764 GND.n762 0.1
R4356 GND.n773 GND.n544 0.1
R4357 GND.n774 GND.n773 0.1
R4358 GND.n775 GND.n774 0.1
R4359 GND.n775 GND.n539 0.1
R4360 GND.n784 GND.n539 0.1
R4361 GND.n785 GND.n784 0.1
R4362 GND.n786 GND.n785 0.1
R4363 GND.n37 GND.n33 0.075
R4364 GND.n53 GND 0.075
R4365 GND.n62 GND.n61 0.075
R4366 GND.n119 GND.n115 0.075
R4367 GND.n135 EESPFAL_s0_0/EESPFAL_NAND_v3_1/GND 0.075
R4368 GND.n144 GND.n143 0.075
R4369 GND.n214 GND.n210 0.075
R4370 GND.n230 EESPFAL_s0_0/EESPFAL_NAND_v3_2/GND 0.075
R4371 GND.n239 GND.n238 0.075
R4372 GND.n319 GND.n315 0.075
R4373 GND.n333 EESPFAL_s1_0/EESPFAL_NAND_v3_0/GND 0.075
R4374 GND.n342 GND.n341 0.075
R4375 GND.n391 GND.n387 0.075
R4376 GND.n405 EESPFAL_s1_0/EESPFAL_INV4_2/GND 0.075
R4377 GND.n414 GND.n413 0.075
R4378 GND.n476 GND.n472 0.075
R4379 GND.n490 EESPFAL_s1_0/EESPFAL_XOR_v3_0/GND 0.075
R4380 GND.n499 GND.n498 0.075
R4381 GND.n1167 GND.n1166 0.075
R4382 GND.n1177 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/GND 0.075
R4383 GND.n1178 GND.n1121 0.075
R4384 GND.n1221 GND.n1220 0.075
R4385 GND.n1231 EESPFAL_s3_0/EESPFAL_INV4_0/GND 0.075
R4386 GND.n1232 GND.n1092 0.075
R4387 GND.n1276 GND.n1275 0.075
R4388 GND.n1286 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/GND 0.075
R4389 GND.n1287 GND.n1064 0.075
R4390 GND.n894 GND.n871 0.075
R4391 EESPFAL_s3_0/EESPFAL_NAND_v3_0/GND GND.n864 0.075
R4392 GND.n916 GND.n915 0.075
R4393 GND.n949 GND.n948 0.075
R4394 GND.n959 EESPFAL_s3_0/EESPFAL_INV4_2/GND 0.075
R4395 GND.n960 GND.n834 0.075
R4396 GND.n1006 GND.n813 0.075
R4397 GND.n1020 EESPFAL_s3_0/EESPFAL_XOR_v3_0/GND 0.075
R4398 GND.n1023 GND.n1022 0.075
R4399 GND.n635 GND.n612 0.075
R4400 EESPFAL_s2_0/EESPFAL_NAND_v3_1/GND GND.n605 0.075
R4401 GND.n657 GND.n656 0.075
R4402 GND.n690 GND.n689 0.075
R4403 GND.n700 EESPFAL_s2_0/EESPFAL_INV4_1/GND 0.075
R4404 GND.n701 GND.n575 0.075
R4405 GND.n747 GND.n554 0.075
R4406 GND.n761 EESPFAL_s2_0/EESPFAL_XOR_v3_0/GND 0.075
R4407 GND.n764 GND.n763 0.075
R4408 GND.n1537 GND.n1536 0.04
R4409 GND.n1546 GND.n1523 0.04
R4410 GND.n1548 GND.n1547 0.04
R4411 GND.n1556 GND.n1518 0.04
R4412 GND.n1558 GND.n1557 0.04
R4413 GND.n1566 GND.n1512 0.04
R4414 GND.n1577 GND.n1506 0.04
R4415 GND.n1579 GND.n1578 0.04
R4416 GND.n1587 GND.n1500 0.04
R4417 GND.n1597 GND.n1493 0.04
R4418 GND.n1599 GND.n1598 0.04
R4419 GND.n1607 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/GND 0.04
R4420 GND.n1609 GND.n1608 0.04
R4421 GND.n1617 GND.n1481 0.04
R4422 GND.n1628 GND.n1475 0.04
R4423 GND.n1630 GND.n1629 0.04
R4424 GND.n1639 GND.n1469 0.04
R4425 GND.n1641 GND.n1640 0.04
R4426 GND.n1650 GND.n1464 0.04
R4427 GND.n1655 GND.n1651 0.04
R4428 GND.n1654 GND.n1653 0.04
R4429 GND.n1662 GND.n1456 0.04
R4430 GND.n1315 EESPFAL_s3_0/GND 0.035
R4431 EESPFAL_s0_0/GND GND.n275 0.035
R4432 GND.n1899 EESPFAL_s1_0/GND 0.035
R4433 GND.n1759 GND.n1397 0.028
R4434 GND.n1767 GND.n1766 0.028
R4435 GND.n1768 GND.n1391 0.028
R4436 GND.n1777 GND.n1776 0.028
R4437 GND.n1778 GND.n1385 0.028
R4438 GND.n1787 GND.n1786 0.028
R4439 GND.n1788 GND.n1379 0.028
R4440 GND.n1797 GND.n1796 0.028
R4441 GND.n1798 GND.n1373 0.028
R4442 GND.n1807 GND.n1806 0.028
R4443 GND.n1819 GND.n1818 0.028
R4444 GND.n1820 GND.n1361 0.028
R4445 GND.n1829 GND.n1828 0.028
R4446 GND.n1839 GND.n1838 0.028
R4447 GND.n1840 GND.n1347 0.028
R4448 GND.n1852 GND.n1341 0.028
R4449 GND.n1861 GND.n1860 0.028
R4450 GND.n1862 GND.n1335 0.028
R4451 GND.n1871 GND.n1870 0.028
R4452 GND.n1872 GND.n1329 0.028
R4453 GND.n1881 GND.n1880 0.028
R4454 GND.n1882 GND.n1323 0.028
R4455 GND.n1891 GND.n1890 0.028
R4456 GND.n1760 GND.n1759 0.027
R4457 GND.n1766 GND.n1397 0.027
R4458 GND.n1768 GND.n1767 0.027
R4459 GND.n1776 GND.n1391 0.027
R4460 GND.n1778 GND.n1777 0.027
R4461 GND.n1786 GND.n1385 0.027
R4462 GND.n1788 GND.n1787 0.027
R4463 GND.n1796 GND.n1379 0.027
R4464 GND.n1798 GND.n1797 0.027
R4465 GND.n1806 GND.n1373 0.027
R4466 GND.n1818 GND.n1367 0.027
R4467 GND.n1820 GND.n1819 0.027
R4468 GND.n1828 GND.n1361 0.027
R4469 GND.n1838 GND.n1353 0.027
R4470 GND.n1840 GND.n1839 0.027
R4471 GND.n1848 GND.n1347 0.027
R4472 GND.n1860 GND.n1341 0.027
R4473 GND.n1862 GND.n1861 0.027
R4474 GND.n1870 GND.n1335 0.027
R4475 GND.n1872 GND.n1871 0.027
R4476 GND.n1880 GND.n1329 0.027
R4477 GND.n1882 GND.n1881 0.027
R4478 GND.n1890 GND.n1323 0.027
R4479 GND.n1892 GND.n1891 0.027
R4480 GND.n1664 GND.n1663 0.027
R4481 GND.n1663 GND.n1452 0.027
R4482 GND.n1670 GND.n1452 0.027
R4483 GND.n1671 GND.n1670 0.027
R4484 GND.n1672 GND.n1671 0.027
R4485 GND.n1672 GND.n1446 0.027
R4486 GND.n1680 GND.n1446 0.027
R4487 GND.n1681 GND.n1680 0.027
R4488 GND.n1683 GND.n1440 0.027
R4489 GND.n1691 GND.n1440 0.027
R4490 GND.n1692 GND.n1691 0.027
R4491 GND.n1694 GND.n1692 0.027
R4492 GND.n1702 GND.n1434 0.027
R4493 GND.n1703 GND.n1702 0.027
R4494 GND.n1704 GND.n1427 0.027
R4495 GND.n1713 GND.n1427 0.027
R4496 GND.n1714 GND.n1713 0.027
R4497 GND.n1715 GND.n1714 0.027
R4498 GND.n1723 GND.n1420 0.027
R4499 GND.n1726 GND.n1725 0.027
R4500 GND.n1726 GND.n1414 0.027
R4501 GND.n1734 GND.n1414 0.027
R4502 GND.n1735 GND.n1734 0.027
R4503 GND.n1737 GND.n1408 0.027
R4504 GND.n1745 GND.n1408 0.027
R4505 GND.n1746 GND.n1745 0.027
R4506 GND.n1750 GND.n1746 0.027
R4507 GND.n1750 GND.n1749 0.027
R4508 GND.n1749 GND.n1748 0.027
R4509 GND.n1748 GND.n1401 0.027
R4510 GND.n1758 GND.n1401 0.027
R4511 GND.n1569 GND.n1568 0.027
R4512 GND.n1589 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/GND 0.027
R4513 GND.n1619 GND.n1618 0.027
R4514 GND.n1316 EESPFAL_s2_0/GND 0.026
R4515 GND.n33 GND.n32 0.025
R4516 GND.n46 GND 0.025
R4517 GND.n66 GND.n62 0.025
R4518 GND.n115 GND.n114 0.025
R4519 GND.n128 EESPFAL_s0_0/EESPFAL_NAND_v3_1/GND 0.025
R4520 GND.n148 GND.n144 0.025
R4521 GND.n210 GND.n209 0.025
R4522 GND.n223 EESPFAL_s0_0/EESPFAL_NAND_v3_2/GND 0.025
R4523 GND.n243 GND.n239 0.025
R4524 GND.n315 GND.n314 0.025
R4525 GND.n328 EESPFAL_s1_0/EESPFAL_NAND_v3_0/GND 0.025
R4526 GND.n346 GND.n342 0.025
R4527 GND.n387 GND.n386 0.025
R4528 GND.n400 EESPFAL_s1_0/EESPFAL_INV4_2/GND 0.025
R4529 GND.n418 GND.n414 0.025
R4530 GND.n472 GND.n471 0.025
R4531 GND.n485 EESPFAL_s1_0/EESPFAL_XOR_v3_0/GND 0.025
R4532 GND.n503 GND.n499 0.025
R4533 GND.n1166 GND.n1165 0.025
R4534 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/GND GND.n1176 0.025
R4535 GND.n1187 GND.n1121 0.025
R4536 GND.n1220 GND.n1219 0.025
R4537 EESPFAL_s3_0/EESPFAL_INV4_0/GND GND.n1230 0.025
R4538 GND.n1241 GND.n1092 0.025
R4539 GND.n1275 GND.n1274 0.025
R4540 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/GND GND.n1285 0.025
R4541 GND.n1296 GND.n1064 0.025
R4542 GND.n895 GND.n894 0.025
R4543 GND.n906 EESPFAL_s3_0/EESPFAL_NAND_v3_0/GND 0.025
R4544 GND.n917 GND.n916 0.025
R4545 GND.n948 GND.n947 0.025
R4546 EESPFAL_s3_0/EESPFAL_INV4_2/GND GND.n958 0.025
R4547 GND.n969 GND.n834 0.025
R4548 GND.n997 GND.n813 0.025
R4549 GND.n1010 EESPFAL_s3_0/EESPFAL_XOR_v3_0/GND 0.025
R4550 GND.n1022 GND.n803 0.025
R4551 GND.n636 GND.n635 0.025
R4552 GND.n647 EESPFAL_s2_0/EESPFAL_NAND_v3_1/GND 0.025
R4553 GND.n658 GND.n657 0.025
R4554 GND.n689 GND.n688 0.025
R4555 EESPFAL_s2_0/EESPFAL_INV4_1/GND GND.n699 0.025
R4556 GND.n710 GND.n575 0.025
R4557 GND.n738 GND.n554 0.025
R4558 GND.n751 EESPFAL_s2_0/EESPFAL_XOR_v3_0/GND 0.025
R4559 GND.n763 GND.n544 0.025
R4560 GND.n1809 GND.n1367 0.014
R4561 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/GND GND.n1353 0.014
R4562 GND.n1849 GND.n1848 0.014
R4563 GND.n1536 GND.n1535 0.014
R4564 GND.n1537 GND.n1523 0.014
R4565 GND.n1547 GND.n1546 0.014
R4566 GND.n1548 GND.n1518 0.014
R4567 GND.n1557 GND.n1556 0.014
R4568 GND.n1558 GND.n1512 0.014
R4569 GND.n1567 GND.n1566 0.014
R4570 GND.n1569 GND.n1506 0.014
R4571 GND.n1578 GND.n1577 0.014
R4572 GND.n1588 GND.n1587 0.014
R4573 GND.n1589 GND.n1493 0.014
R4574 GND.n1598 GND.n1597 0.014
R4575 GND.n1609 GND.n1481 0.014
R4576 GND.n1618 GND.n1617 0.014
R4577 GND.n1620 GND.n1475 0.014
R4578 GND.n1629 GND.n1628 0.014
R4579 GND.n1630 GND.n1469 0.014
R4580 GND.n1640 GND.n1639 0.014
R4581 GND.n1641 GND.n1464 0.014
R4582 GND.n1651 GND.n1650 0.014
R4583 GND.n1655 GND.n1654 0.014
R4584 GND.n1653 GND.n1456 0.014
R4585 GND.n1808 GND.n1807 0.013
R4586 GND.n1810 GND.n1808 0.013
R4587 GND.n1810 GND.n1809 0.013
R4588 EESPFAL_s2_0/EESPFAL_4in_NAND_0/GND GND.n1829 0.013
R4589 GND.n1830 EESPFAL_s2_0/EESPFAL_4in_NAND_0/GND 0.013
R4590 GND.n1830 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/GND 0.013
R4591 GND.n1850 GND.n1849 0.013
R4592 GND.n1851 GND.n1850 0.013
R4593 GND.n1852 GND.n1851 0.013
R4594 GND.n1682 GND.n1681 0.013
R4595 GND.n1683 GND.n1682 0.013
R4596 GND.n1694 GND.n1693 0.013
R4597 GND.n1693 GND.n1434 0.013
R4598 EESPFAL_s2_0/EESPFAL_INV4_2/GND GND.n1703 0.013
R4599 GND.n1704 EESPFAL_s2_0/EESPFAL_INV4_2/GND 0.013
R4600 GND.n1715 EESPFAL_s1_0/EESPFAL_INV4_0/GND 0.013
R4601 EESPFAL_s1_0/EESPFAL_INV4_0/GND GND.n1420 0.013
R4602 GND.n1724 GND.n1723 0.013
R4603 GND.n1725 GND.n1724 0.013
R4604 GND.n1736 GND.n1735 0.013
R4605 GND.n1737 GND.n1736 0.013
R4606 GND.n1568 GND.n1567 0.013
R4607 GND.n1579 GND.n1500 0.013
R4608 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/GND GND.n1588 0.013
R4609 GND.n1599 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/GND 0.013
R4610 GND.n1608 GND.n1607 0.013
R4611 GND.n1620 GND.n1619 0.013
R4612 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/A_bar 922.56
R4613 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t8 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t9 819.4
R4614 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t6 684.833
R4615 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t7 506.1
R4616 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t8 313.3
R4617 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t1 177.936
R4618 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n3 128.335
R4619 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n1 105.6
R4620 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t2 81.937
R4621 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n0 58.265
R4622 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n4 57.6
R4623 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n2 41.6
R4624 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t5 39.4
R4625 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t4 39.4
R4626 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t3 24
R4627 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t0 24
R4628 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n5 8.764
R4629 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n6 4.65
R4630 x1.n3 x1.t11 1176.57
R4631 x1.n2 x1.t1 1176.57
R4632 x1.n1 x1.t3 1176.57
R4633 x1.n3 x1.t5 1149.49
R4634 x1.n2 x1.t7 1149.49
R4635 x1.n1 x1.t8 1149.49
R4636 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B x1.t9 1106.75
R4637 x1 x1.t6 1026.78
R4638 EESPFAL_s3_0/EESPFAL_INV4_1/A x1.t0 778.1
R4639 EESPFAL_s0_0/EESPFAL_NAND_v3_2/B_bar x1.t4 527.366
R4640 EESPFAL_s2_0/EESPFAL_4in_NAND_0/B x1.t10 446.232
R4641 EESPFAL_s2_0/EESPFAL_INV4_1/A_bar x1.t2 392.5
R4642 x1.n0 EESPFAL_s0_0/EESPFAL_NAND_v3_2/B_bar 338.09
R4643 x1.n8 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B 290.41
R4644 x1.n6 EESPFAL_s2_0/EESPFAL_XOR_v3_1/A 254.89
R4645 x1.n7 EESPFAL_s2_0/EESPFAL_4in_NAND_0/B 254.89
R4646 x1.n4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/A 242.09
R4647 x1.n9 EESPFAL_s1_0/EESPFAL_XOR_v3_1/A 242.09
R4648 x1.n5 EESPFAL_s2_0/EESPFAL_INV4_1/A_bar 197.718
R4649 EESPFAL_s3_0/EESPFAL_XOR_v3_0/A x1.n3 128
R4650 EESPFAL_s2_0/EESPFAL_XOR_v3_1/A x1.n2 128
R4651 EESPFAL_s1_0/EESPFAL_XOR_v3_1/A x1.n1 128
R4652 EESPFAL_s3_0/x1 EESPFAL_s3_0/EESPFAL_INV4_1/A 44.476
R4653 EESPFAL_s0_0/x1 x1 23.476
R4654 x1.n8 x1.n7 3.546
R4655 EESPFAL_s1_0/x1 x1.n9 3.228
R4656 x1.n0 EESPFAL_s0_0/x1 2.51
R4657 x1.n6 x1.n5 2.168
R4658 EESPFAL_s1_0/x1 x1.n0 1.896
R4659 x1.n9 x1.n8 1.234
R4660 x1.n5 EESPFAL_s2_0/x1 1.153
R4661 EESPFAL_s2_0/x1 x1.n4 1.115
R4662 x1.n7 x1.n6 0.814
R4663 x1.n4 EESPFAL_s3_0/x1 0.084
R4664 CLK1.n277 CLK1.n276 407.048
R4665 CLK1.n232 CLK1.n223 407.048
R4666 CLK1.n1620 CLK1.n1619 407.048
R4667 CLK1.n1553 CLK1.n1552 407.048
R4668 CLK1.n1547 CLK1.n1546 407.048
R4669 CLK1.n1512 CLK1.n1503 407.048
R4670 CLK1.n1253 CLK1.n1252 407.048
R4671 CLK1.n1197 CLK1.n316 407.048
R4672 CLK1.n387 CLK1.n386 407.048
R4673 CLK1.n352 CLK1.n343 407.048
R4674 CLK1.n475 CLK1.n474 407.048
R4675 CLK1.n440 CLK1.n431 407.048
R4676 CLK1.n999 CLK1.n998 407.048
R4677 CLK1.n484 CLK1.n407 407.048
R4678 CLK1.n988 CLK1.n987 407.048
R4679 CLK1.n921 CLK1.n920 407.048
R4680 CLK1.n915 CLK1.n914 407.048
R4681 CLK1.n880 CLK1.n871 407.048
R4682 CLK1.n621 CLK1.n620 407.048
R4683 CLK1.n565 CLK1.n556 407.048
R4684 CLK1.n803 CLK1.n802 407.048
R4685 CLK1.n736 CLK1.n735 407.048
R4686 CLK1.n730 CLK1.n729 407.048
R4687 CLK1.n695 CLK1.n686 407.048
R4688 CLK1.n1435 CLK1.n1434 407.048
R4689 CLK1.n1368 CLK1.n1367 407.048
R4690 CLK1.n1362 CLK1.n1361 407.048
R4691 CLK1.n1327 CLK1.n1318 407.048
R4692 CLK1.n267 CLK1.n198 400
R4693 CLK1.n276 CLK1.n198 400
R4694 CLK1.n233 CLK1.n232 400
R4695 CLK1.n234 CLK1.n233 400
R4696 CLK1.n1607 CLK1.n1453 400
R4697 CLK1.n1608 CLK1.n1607 400
R4698 CLK1.n1609 CLK1.n1608 400
R4699 CLK1.n1609 CLK1.n1445 400
R4700 CLK1.n1619 CLK1.n1445 400
R4701 CLK1.n1553 CLK1.n1475 400
R4702 CLK1.n1562 CLK1.n1475 400
R4703 CLK1.n1563 CLK1.n1562 400
R4704 CLK1.n1564 CLK1.n1563 400
R4705 CLK1.n1564 CLK1.n1469 400
R4706 CLK1.n1242 CLK1.n1241 400
R4707 CLK1.n1243 CLK1.n1242 400
R4708 CLK1.n1243 CLK1.n285 400
R4709 CLK1.n1252 CLK1.n285 400
R4710 CLK1.n1198 CLK1.n1197 400
R4711 CLK1.n1199 CLK1.n1198 400
R4712 CLK1.n1199 CLK1.n310 400
R4713 CLK1.n1207 CLK1.n310 400
R4714 CLK1.n1010 CLK1.n506 400
R4715 CLK1.n1010 CLK1.n1009 400
R4716 CLK1.n1009 CLK1.n1008 400
R4717 CLK1.n1008 CLK1.n513 400
R4718 CLK1.n999 CLK1.n513 400
R4719 CLK1.n485 CLK1.n484 400
R4720 CLK1.n1050 CLK1.n485 400
R4721 CLK1.n1050 CLK1.n1049 400
R4722 CLK1.n1049 CLK1.n1048 400
R4723 CLK1.n1048 CLK1.n486 400
R4724 CLK1.n975 CLK1.n821 400
R4725 CLK1.n976 CLK1.n975 400
R4726 CLK1.n977 CLK1.n976 400
R4727 CLK1.n977 CLK1.n813 400
R4728 CLK1.n987 CLK1.n813 400
R4729 CLK1.n921 CLK1.n843 400
R4730 CLK1.n930 CLK1.n843 400
R4731 CLK1.n931 CLK1.n930 400
R4732 CLK1.n932 CLK1.n931 400
R4733 CLK1.n932 CLK1.n837 400
R4734 CLK1.n610 CLK1.n609 400
R4735 CLK1.n611 CLK1.n610 400
R4736 CLK1.n611 CLK1.n525 400
R4737 CLK1.n620 CLK1.n525 400
R4738 CLK1.n566 CLK1.n565 400
R4739 CLK1.n567 CLK1.n566 400
R4740 CLK1.n567 CLK1.n550 400
R4741 CLK1.n575 CLK1.n550 400
R4742 CLK1.n790 CLK1.n636 400
R4743 CLK1.n791 CLK1.n790 400
R4744 CLK1.n792 CLK1.n791 400
R4745 CLK1.n792 CLK1.n628 400
R4746 CLK1.n802 CLK1.n628 400
R4747 CLK1.n736 CLK1.n658 400
R4748 CLK1.n745 CLK1.n658 400
R4749 CLK1.n746 CLK1.n745 400
R4750 CLK1.n747 CLK1.n746 400
R4751 CLK1.n747 CLK1.n652 400
R4752 CLK1.n1422 CLK1.n1268 400
R4753 CLK1.n1423 CLK1.n1422 400
R4754 CLK1.n1424 CLK1.n1423 400
R4755 CLK1.n1424 CLK1.n1260 400
R4756 CLK1.n1434 CLK1.n1260 400
R4757 CLK1.n1368 CLK1.n1290 400
R4758 CLK1.n1377 CLK1.n1290 400
R4759 CLK1.n1378 CLK1.n1377 400
R4760 CLK1.n1379 CLK1.n1378 400
R4761 CLK1.n1379 CLK1.n1284 400
R4762 CLK1.n267 CLK1.n266 366.379
R4763 CLK1.n234 CLK1.n217 366.379
R4764 CLK1.n1599 CLK1.n1453 366.379
R4765 CLK1.n1573 CLK1.n1469 366.379
R4766 CLK1.n1546 CLK1.n1485 366.379
R4767 CLK1.n1513 CLK1.n1512 366.379
R4768 CLK1.n1241 CLK1.n292 366.379
R4769 CLK1.n1208 CLK1.n1207 366.379
R4770 CLK1.n386 CLK1.n325 366.379
R4771 CLK1.n353 CLK1.n352 366.379
R4772 CLK1.n474 CLK1.n413 366.379
R4773 CLK1.n441 CLK1.n440 366.379
R4774 CLK1.n1018 CLK1.n506 366.379
R4775 CLK1.n1040 CLK1.n486 366.379
R4776 CLK1.n967 CLK1.n821 366.379
R4777 CLK1.n941 CLK1.n837 366.379
R4778 CLK1.n914 CLK1.n853 366.379
R4779 CLK1.n881 CLK1.n880 366.379
R4780 CLK1.n609 CLK1.n532 366.379
R4781 CLK1.n576 CLK1.n575 366.379
R4782 CLK1.n782 CLK1.n636 366.379
R4783 CLK1.n756 CLK1.n652 366.379
R4784 CLK1.n729 CLK1.n668 366.379
R4785 CLK1.n696 CLK1.n695 366.379
R4786 CLK1.n1414 CLK1.n1268 366.379
R4787 CLK1.n1388 CLK1.n1284 366.379
R4788 CLK1.n1361 CLK1.n1300 366.379
R4789 CLK1.n1328 CLK1.n1327 366.379
R4790 CLK1.n1175 CLK1.n1174 240.502
R4791 CLK1.n1118 CLK1.n1117 240.501
R4792 CLK1.n1130 CLK1.n1103 236.76
R4793 CLK1.n1130 CLK1.n1129 236.76
R4794 CLK1.n1129 CLK1.n1128 236.76
R4795 CLK1.n1128 CLK1.n1104 236.76
R4796 CLK1.n1119 CLK1.n1104 236.76
R4797 CLK1.n1119 CLK1.n1118 236.76
R4798 CLK1.n1174 CLK1.n1173 236.76
R4799 CLK1.n1173 CLK1.n395 236.76
R4800 CLK1.n1164 CLK1.n395 236.76
R4801 CLK1.n1164 CLK1.n1163 236.76
R4802 CLK1.n1163 CLK1.n1162 236.76
R4803 CLK1.n1162 CLK1.n1069 236.76
R4804 CLK1.n1103 CLK1.n1095 215.793
R4805 CLK1.n1074 CLK1.n1069 215.793
R4806 CLK1.n243 CLK1.n217 131.034
R4807 CLK1.n244 CLK1.n243 131.034
R4808 CLK1.n246 CLK1.n245 131.034
R4809 CLK1.n256 CLK1.n255 131.034
R4810 CLK1.n265 CLK1.n205 131.034
R4811 CLK1.n266 CLK1.n265 131.034
R4812 CLK1.n1574 CLK1.n1573 131.034
R4813 CLK1.n1575 CLK1.n1574 131.034
R4814 CLK1.n1585 CLK1.n1463 131.034
R4815 CLK1.n1588 CLK1.n1587 131.034
R4816 CLK1.n1598 CLK1.n1597 131.034
R4817 CLK1.n1599 CLK1.n1598 131.034
R4818 CLK1.n1515 CLK1.n1513 131.034
R4819 CLK1.n1515 CLK1.n1514 131.034
R4820 CLK1.n1525 CLK1.n1524 131.034
R4821 CLK1.n1535 CLK1.n1491 131.034
R4822 CLK1.n1537 CLK1.n1536 131.034
R4823 CLK1.n1537 CLK1.n1485 131.034
R4824 CLK1.n1210 CLK1.n1208 131.034
R4825 CLK1.n1210 CLK1.n1209 131.034
R4826 CLK1.n1220 CLK1.n1219 131.034
R4827 CLK1.n1230 CLK1.n298 131.034
R4828 CLK1.n1232 CLK1.n1231 131.034
R4829 CLK1.n1232 CLK1.n292 131.034
R4830 CLK1.n355 CLK1.n353 131.034
R4831 CLK1.n355 CLK1.n354 131.034
R4832 CLK1.n365 CLK1.n364 131.034
R4833 CLK1.n375 CLK1.n331 131.034
R4834 CLK1.n377 CLK1.n376 131.034
R4835 CLK1.n377 CLK1.n325 131.034
R4836 CLK1.n443 CLK1.n441 131.034
R4837 CLK1.n443 CLK1.n442 131.034
R4838 CLK1.n453 CLK1.n452 131.034
R4839 CLK1.n463 CLK1.n419 131.034
R4840 CLK1.n465 CLK1.n464 131.034
R4841 CLK1.n465 CLK1.n413 131.034
R4842 CLK1.n1040 CLK1.n1039 131.034
R4843 CLK1.n1039 CLK1.n1038 131.034
R4844 CLK1.n1030 CLK1.n499 131.034
R4845 CLK1.n1028 CLK1.n500 131.034
R4846 CLK1.n1020 CLK1.n1019 131.034
R4847 CLK1.n1019 CLK1.n1018 131.034
R4848 CLK1.n942 CLK1.n941 131.034
R4849 CLK1.n943 CLK1.n942 131.034
R4850 CLK1.n953 CLK1.n831 131.034
R4851 CLK1.n956 CLK1.n955 131.034
R4852 CLK1.n966 CLK1.n965 131.034
R4853 CLK1.n967 CLK1.n966 131.034
R4854 CLK1.n883 CLK1.n881 131.034
R4855 CLK1.n883 CLK1.n882 131.034
R4856 CLK1.n893 CLK1.n892 131.034
R4857 CLK1.n903 CLK1.n859 131.034
R4858 CLK1.n905 CLK1.n904 131.034
R4859 CLK1.n905 CLK1.n853 131.034
R4860 CLK1.n578 CLK1.n576 131.034
R4861 CLK1.n578 CLK1.n577 131.034
R4862 CLK1.n588 CLK1.n587 131.034
R4863 CLK1.n598 CLK1.n538 131.034
R4864 CLK1.n600 CLK1.n599 131.034
R4865 CLK1.n600 CLK1.n532 131.034
R4866 CLK1.n757 CLK1.n756 131.034
R4867 CLK1.n758 CLK1.n757 131.034
R4868 CLK1.n768 CLK1.n646 131.034
R4869 CLK1.n771 CLK1.n770 131.034
R4870 CLK1.n781 CLK1.n780 131.034
R4871 CLK1.n782 CLK1.n781 131.034
R4872 CLK1.n698 CLK1.n696 131.034
R4873 CLK1.n698 CLK1.n697 131.034
R4874 CLK1.n708 CLK1.n707 131.034
R4875 CLK1.n718 CLK1.n674 131.034
R4876 CLK1.n720 CLK1.n719 131.034
R4877 CLK1.n720 CLK1.n668 131.034
R4878 CLK1.n1389 CLK1.n1388 131.034
R4879 CLK1.n1390 CLK1.n1389 131.034
R4880 CLK1.n1400 CLK1.n1278 131.034
R4881 CLK1.n1403 CLK1.n1402 131.034
R4882 CLK1.n1413 CLK1.n1412 131.034
R4883 CLK1.n1414 CLK1.n1413 131.034
R4884 CLK1.n1330 CLK1.n1328 131.034
R4885 CLK1.n1330 CLK1.n1329 131.034
R4886 CLK1.n1340 CLK1.n1339 131.034
R4887 CLK1.n1350 CLK1.n1306 131.034
R4888 CLK1.n1352 CLK1.n1351 131.034
R4889 CLK1.n1352 CLK1.n1300 131.034
R4890 CLK1.n254 CLK1.t166 122.844
R4891 CLK1.t16 CLK1.n254 122.844
R4892 CLK1.n1586 CLK1.t41 122.844
R4893 CLK1.t150 CLK1.n1586 122.844
R4894 CLK1.n1526 CLK1.t82 122.844
R4895 CLK1.n1526 CLK1.t0 122.844
R4896 CLK1.n1221 CLK1.t34 122.844
R4897 CLK1.n1221 CLK1.t135 122.844
R4898 CLK1.n366 CLK1.t145 122.844
R4899 CLK1.n366 CLK1.t102 122.844
R4900 CLK1.n454 CLK1.t121 122.844
R4901 CLK1.n454 CLK1.t8 122.844
R4902 CLK1.t123 CLK1.n1029 122.844
R4903 CLK1.n1029 CLK1.t141 122.844
R4904 CLK1.n954 CLK1.t112 122.844
R4905 CLK1.t38 CLK1.n954 122.844
R4906 CLK1.n894 CLK1.t72 122.844
R4907 CLK1.n894 CLK1.t127 122.844
R4908 CLK1.n589 CLK1.t158 122.844
R4909 CLK1.n589 CLK1.t156 122.844
R4910 CLK1.n769 CLK1.t152 122.844
R4911 CLK1.t179 CLK1.n769 122.844
R4912 CLK1.n709 CLK1.t78 122.844
R4913 CLK1.n709 CLK1.t43 122.844
R4914 CLK1.n1401 CLK1.t29 122.844
R4915 CLK1.t130 CLK1.n1401 122.844
R4916 CLK1.n1341 CLK1.t175 122.844
R4917 CLK1.n1341 CLK1.t14 122.844
R4918 CLK1.n246 CLK1.t164 106.465
R4919 CLK1.n256 CLK1.t18 106.465
R4920 CLK1.t177 CLK1.n1463 106.465
R4921 CLK1.n1587 CLK1.t51 106.465
R4922 CLK1.n1524 CLK1.t80 106.465
R4923 CLK1.t2 CLK1.n1535 106.465
R4924 CLK1.n1219 CLK1.t36 106.465
R4925 CLK1.t137 CLK1.n1230 106.465
R4926 CLK1.n364 CLK1.t143 106.465
R4927 CLK1.t104 CLK1.n375 106.465
R4928 CLK1.n452 CLK1.t119 106.465
R4929 CLK1.t10 CLK1.n463 106.465
R4930 CLK1.n499 CLK1.t193 106.465
R4931 CLK1.t47 CLK1.n500 106.465
R4932 CLK1.t20 CLK1.n831 106.465
R4933 CLK1.n955 CLK1.t184 106.465
R4934 CLK1.n892 CLK1.t74 106.465
R4935 CLK1.t125 CLK1.n903 106.465
R4936 CLK1.n587 CLK1.t160 106.465
R4937 CLK1.t154 CLK1.n598 106.465
R4938 CLK1.t92 CLK1.n646 106.465
R4939 CLK1.n770 CLK1.t139 106.465
R4940 CLK1.n707 CLK1.t76 106.465
R4941 CLK1.t45 CLK1.n718 106.465
R4942 CLK1.t69 CLK1.n1278 106.465
R4943 CLK1.n1402 CLK1.t132 106.465
R4944 CLK1.n1339 CLK1.t173 106.465
R4945 CLK1.t12 CLK1.n1350 106.465
R4946 CLK1.n231 CLK1.n224 96
R4947 CLK1.n231 CLK1.n222 96
R4948 CLK1.n235 CLK1.n222 96
R4949 CLK1.n235 CLK1.n218 96
R4950 CLK1.n242 CLK1.n218 96
R4951 CLK1.n242 CLK1.n216 96
R4952 CLK1.n247 CLK1.n216 96
R4953 CLK1.n247 CLK1.n211 96
R4954 CLK1.n253 CLK1.n211 96
R4955 CLK1.n253 CLK1.n210 96
R4956 CLK1.n257 CLK1.n210 96
R4957 CLK1.n257 CLK1.n206 96
R4958 CLK1.n264 CLK1.n206 96
R4959 CLK1.n264 CLK1.n204 96
R4960 CLK1.n268 CLK1.n204 96
R4961 CLK1.n268 CLK1.n199 96
R4962 CLK1.n275 CLK1.n199 96
R4963 CLK1.n275 CLK1.n197 96
R4964 CLK1.n1554 CLK1.n1481 96
R4965 CLK1.n1554 CLK1.n1476 96
R4966 CLK1.n1561 CLK1.n1476 96
R4967 CLK1.n1561 CLK1.n1474 96
R4968 CLK1.n1565 CLK1.n1474 96
R4969 CLK1.n1565 CLK1.n1470 96
R4970 CLK1.n1572 CLK1.n1470 96
R4971 CLK1.n1572 CLK1.n1468 96
R4972 CLK1.n1576 CLK1.n1468 96
R4973 CLK1.n1576 CLK1.n1464 96
R4974 CLK1.n1584 CLK1.n1464 96
R4975 CLK1.n1584 CLK1.n1462 96
R4976 CLK1.n1589 CLK1.n1462 96
R4977 CLK1.n1589 CLK1.n1459 96
R4978 CLK1.n1596 CLK1.n1459 96
R4979 CLK1.n1596 CLK1.n1458 96
R4980 CLK1.n1600 CLK1.n1458 96
R4981 CLK1.n1600 CLK1.n1454 96
R4982 CLK1.n1606 CLK1.n1454 96
R4983 CLK1.n1606 CLK1.n1452 96
R4984 CLK1.n1610 CLK1.n1452 96
R4985 CLK1.n1610 CLK1.n1446 96
R4986 CLK1.n1618 CLK1.n1446 96
R4987 CLK1.n1618 CLK1.n1444 96
R4988 CLK1.n1511 CLK1.n1504 96
R4989 CLK1.n1511 CLK1.n1502 96
R4990 CLK1.n1516 CLK1.n1502 96
R4991 CLK1.n1516 CLK1.n1498 96
R4992 CLK1.n1523 CLK1.n1498 96
R4993 CLK1.n1523 CLK1.n1497 96
R4994 CLK1.n1527 CLK1.n1497 96
R4995 CLK1.n1527 CLK1.n1492 96
R4996 CLK1.n1534 CLK1.n1492 96
R4997 CLK1.n1534 CLK1.n1490 96
R4998 CLK1.n1538 CLK1.n1490 96
R4999 CLK1.n1538 CLK1.n1486 96
R5000 CLK1.n1545 CLK1.n1486 96
R5001 CLK1.n1545 CLK1.n1484 96
R5002 CLK1.n1196 CLK1.n317 96
R5003 CLK1.n1196 CLK1.n315 96
R5004 CLK1.n1200 CLK1.n315 96
R5005 CLK1.n1200 CLK1.n311 96
R5006 CLK1.n1206 CLK1.n311 96
R5007 CLK1.n1206 CLK1.n309 96
R5008 CLK1.n1211 CLK1.n309 96
R5009 CLK1.n1211 CLK1.n305 96
R5010 CLK1.n1218 CLK1.n305 96
R5011 CLK1.n1218 CLK1.n304 96
R5012 CLK1.n1222 CLK1.n304 96
R5013 CLK1.n1222 CLK1.n299 96
R5014 CLK1.n1229 CLK1.n299 96
R5015 CLK1.n1229 CLK1.n297 96
R5016 CLK1.n1233 CLK1.n297 96
R5017 CLK1.n1233 CLK1.n293 96
R5018 CLK1.n1240 CLK1.n293 96
R5019 CLK1.n1240 CLK1.n291 96
R5020 CLK1.n1244 CLK1.n291 96
R5021 CLK1.n1244 CLK1.n286 96
R5022 CLK1.n1251 CLK1.n286 96
R5023 CLK1.n1251 CLK1.n284 96
R5024 CLK1.n351 CLK1.n344 96
R5025 CLK1.n351 CLK1.n342 96
R5026 CLK1.n356 CLK1.n342 96
R5027 CLK1.n356 CLK1.n338 96
R5028 CLK1.n363 CLK1.n338 96
R5029 CLK1.n363 CLK1.n337 96
R5030 CLK1.n367 CLK1.n337 96
R5031 CLK1.n367 CLK1.n332 96
R5032 CLK1.n374 CLK1.n332 96
R5033 CLK1.n374 CLK1.n330 96
R5034 CLK1.n378 CLK1.n330 96
R5035 CLK1.n378 CLK1.n326 96
R5036 CLK1.n385 CLK1.n326 96
R5037 CLK1.n385 CLK1.n324 96
R5038 CLK1.n439 CLK1.n432 96
R5039 CLK1.n439 CLK1.n430 96
R5040 CLK1.n444 CLK1.n430 96
R5041 CLK1.n444 CLK1.n426 96
R5042 CLK1.n451 CLK1.n426 96
R5043 CLK1.n451 CLK1.n425 96
R5044 CLK1.n455 CLK1.n425 96
R5045 CLK1.n455 CLK1.n420 96
R5046 CLK1.n462 CLK1.n420 96
R5047 CLK1.n462 CLK1.n418 96
R5048 CLK1.n466 CLK1.n418 96
R5049 CLK1.n466 CLK1.n414 96
R5050 CLK1.n473 CLK1.n414 96
R5051 CLK1.n473 CLK1.n412 96
R5052 CLK1.n483 CLK1.n408 96
R5053 CLK1.n483 CLK1.n405 96
R5054 CLK1.n1051 CLK1.n405 96
R5055 CLK1.n1051 CLK1.n406 96
R5056 CLK1.n1047 CLK1.n406 96
R5057 CLK1.n1047 CLK1.n487 96
R5058 CLK1.n1041 CLK1.n487 96
R5059 CLK1.n1041 CLK1.n491 96
R5060 CLK1.n1037 CLK1.n491 96
R5061 CLK1.n1037 CLK1.n492 96
R5062 CLK1.n1031 CLK1.n492 96
R5063 CLK1.n1031 CLK1.n498 96
R5064 CLK1.n1027 CLK1.n498 96
R5065 CLK1.n1027 CLK1.n501 96
R5066 CLK1.n1021 CLK1.n501 96
R5067 CLK1.n1021 CLK1.n505 96
R5068 CLK1.n1017 CLK1.n505 96
R5069 CLK1.n1017 CLK1.n507 96
R5070 CLK1.n1011 CLK1.n507 96
R5071 CLK1.n1011 CLK1.n512 96
R5072 CLK1.n1007 CLK1.n512 96
R5073 CLK1.n1007 CLK1.n514 96
R5074 CLK1.n1000 CLK1.n514 96
R5075 CLK1.n1000 CLK1.n519 96
R5076 CLK1.n922 CLK1.n849 96
R5077 CLK1.n922 CLK1.n844 96
R5078 CLK1.n929 CLK1.n844 96
R5079 CLK1.n929 CLK1.n842 96
R5080 CLK1.n933 CLK1.n842 96
R5081 CLK1.n933 CLK1.n838 96
R5082 CLK1.n940 CLK1.n838 96
R5083 CLK1.n940 CLK1.n836 96
R5084 CLK1.n944 CLK1.n836 96
R5085 CLK1.n944 CLK1.n832 96
R5086 CLK1.n952 CLK1.n832 96
R5087 CLK1.n952 CLK1.n830 96
R5088 CLK1.n957 CLK1.n830 96
R5089 CLK1.n957 CLK1.n827 96
R5090 CLK1.n964 CLK1.n827 96
R5091 CLK1.n964 CLK1.n826 96
R5092 CLK1.n968 CLK1.n826 96
R5093 CLK1.n968 CLK1.n822 96
R5094 CLK1.n974 CLK1.n822 96
R5095 CLK1.n974 CLK1.n820 96
R5096 CLK1.n978 CLK1.n820 96
R5097 CLK1.n978 CLK1.n814 96
R5098 CLK1.n986 CLK1.n814 96
R5099 CLK1.n986 CLK1.n812 96
R5100 CLK1.n879 CLK1.n872 96
R5101 CLK1.n879 CLK1.n870 96
R5102 CLK1.n884 CLK1.n870 96
R5103 CLK1.n884 CLK1.n866 96
R5104 CLK1.n891 CLK1.n866 96
R5105 CLK1.n891 CLK1.n865 96
R5106 CLK1.n895 CLK1.n865 96
R5107 CLK1.n895 CLK1.n860 96
R5108 CLK1.n902 CLK1.n860 96
R5109 CLK1.n902 CLK1.n858 96
R5110 CLK1.n906 CLK1.n858 96
R5111 CLK1.n906 CLK1.n854 96
R5112 CLK1.n913 CLK1.n854 96
R5113 CLK1.n913 CLK1.n852 96
R5114 CLK1.n564 CLK1.n557 96
R5115 CLK1.n564 CLK1.n555 96
R5116 CLK1.n568 CLK1.n555 96
R5117 CLK1.n568 CLK1.n551 96
R5118 CLK1.n574 CLK1.n551 96
R5119 CLK1.n574 CLK1.n549 96
R5120 CLK1.n579 CLK1.n549 96
R5121 CLK1.n579 CLK1.n545 96
R5122 CLK1.n586 CLK1.n545 96
R5123 CLK1.n586 CLK1.n544 96
R5124 CLK1.n590 CLK1.n544 96
R5125 CLK1.n590 CLK1.n539 96
R5126 CLK1.n597 CLK1.n539 96
R5127 CLK1.n597 CLK1.n537 96
R5128 CLK1.n601 CLK1.n537 96
R5129 CLK1.n601 CLK1.n533 96
R5130 CLK1.n608 CLK1.n533 96
R5131 CLK1.n608 CLK1.n531 96
R5132 CLK1.n612 CLK1.n531 96
R5133 CLK1.n612 CLK1.n526 96
R5134 CLK1.n619 CLK1.n526 96
R5135 CLK1.n619 CLK1.n524 96
R5136 CLK1.n737 CLK1.n664 96
R5137 CLK1.n737 CLK1.n659 96
R5138 CLK1.n744 CLK1.n659 96
R5139 CLK1.n744 CLK1.n657 96
R5140 CLK1.n748 CLK1.n657 96
R5141 CLK1.n748 CLK1.n653 96
R5142 CLK1.n755 CLK1.n653 96
R5143 CLK1.n755 CLK1.n651 96
R5144 CLK1.n759 CLK1.n651 96
R5145 CLK1.n759 CLK1.n647 96
R5146 CLK1.n767 CLK1.n647 96
R5147 CLK1.n767 CLK1.n645 96
R5148 CLK1.n772 CLK1.n645 96
R5149 CLK1.n772 CLK1.n642 96
R5150 CLK1.n779 CLK1.n642 96
R5151 CLK1.n779 CLK1.n641 96
R5152 CLK1.n783 CLK1.n641 96
R5153 CLK1.n783 CLK1.n637 96
R5154 CLK1.n789 CLK1.n637 96
R5155 CLK1.n789 CLK1.n635 96
R5156 CLK1.n793 CLK1.n635 96
R5157 CLK1.n793 CLK1.n629 96
R5158 CLK1.n801 CLK1.n629 96
R5159 CLK1.n801 CLK1.n627 96
R5160 CLK1.n694 CLK1.n687 96
R5161 CLK1.n694 CLK1.n685 96
R5162 CLK1.n699 CLK1.n685 96
R5163 CLK1.n699 CLK1.n681 96
R5164 CLK1.n706 CLK1.n681 96
R5165 CLK1.n706 CLK1.n680 96
R5166 CLK1.n710 CLK1.n680 96
R5167 CLK1.n710 CLK1.n675 96
R5168 CLK1.n717 CLK1.n675 96
R5169 CLK1.n717 CLK1.n673 96
R5170 CLK1.n721 CLK1.n673 96
R5171 CLK1.n721 CLK1.n669 96
R5172 CLK1.n728 CLK1.n669 96
R5173 CLK1.n728 CLK1.n667 96
R5174 CLK1.n1369 CLK1.n1296 96
R5175 CLK1.n1369 CLK1.n1291 96
R5176 CLK1.n1376 CLK1.n1291 96
R5177 CLK1.n1376 CLK1.n1289 96
R5178 CLK1.n1380 CLK1.n1289 96
R5179 CLK1.n1380 CLK1.n1285 96
R5180 CLK1.n1387 CLK1.n1285 96
R5181 CLK1.n1387 CLK1.n1283 96
R5182 CLK1.n1391 CLK1.n1283 96
R5183 CLK1.n1391 CLK1.n1279 96
R5184 CLK1.n1399 CLK1.n1279 96
R5185 CLK1.n1399 CLK1.n1277 96
R5186 CLK1.n1404 CLK1.n1277 96
R5187 CLK1.n1404 CLK1.n1274 96
R5188 CLK1.n1411 CLK1.n1274 96
R5189 CLK1.n1411 CLK1.n1273 96
R5190 CLK1.n1415 CLK1.n1273 96
R5191 CLK1.n1415 CLK1.n1269 96
R5192 CLK1.n1421 CLK1.n1269 96
R5193 CLK1.n1421 CLK1.n1267 96
R5194 CLK1.n1425 CLK1.n1267 96
R5195 CLK1.n1425 CLK1.n1261 96
R5196 CLK1.n1433 CLK1.n1261 96
R5197 CLK1.n1433 CLK1.n1259 96
R5198 CLK1.n1326 CLK1.n1319 96
R5199 CLK1.n1326 CLK1.n1317 96
R5200 CLK1.n1331 CLK1.n1317 96
R5201 CLK1.n1331 CLK1.n1313 96
R5202 CLK1.n1338 CLK1.n1313 96
R5203 CLK1.n1338 CLK1.n1312 96
R5204 CLK1.n1342 CLK1.n1312 96
R5205 CLK1.n1342 CLK1.n1307 96
R5206 CLK1.n1349 CLK1.n1307 96
R5207 CLK1.n1349 CLK1.n1305 96
R5208 CLK1.n1353 CLK1.n1305 96
R5209 CLK1.n1353 CLK1.n1301 96
R5210 CLK1.n1360 CLK1.n1301 96
R5211 CLK1.n1360 CLK1.n1299 96
R5212 CLK1.n226 CLK1.n223 85.261
R5213 CLK1.n1552 CLK1.n1551 85.261
R5214 CLK1.n1506 CLK1.n1503 85.261
R5215 CLK1.n1191 CLK1.n316 85.261
R5216 CLK1.n478 CLK1.n407 85.261
R5217 CLK1.n920 CLK1.n919 85.261
R5218 CLK1.n874 CLK1.n871 85.261
R5219 CLK1.n559 CLK1.n556 85.261
R5220 CLK1.n735 CLK1.n734 85.261
R5221 CLK1.n689 CLK1.n686 85.261
R5222 CLK1.n1367 CLK1.n1366 85.261
R5223 CLK1.n1321 CLK1.n1318 85.261
R5224 CLK1.n278 CLK1.n277 85.261
R5225 CLK1.n1621 CLK1.n1620 85.261
R5226 CLK1.n1548 CLK1.n1547 85.261
R5227 CLK1.n1254 CLK1.n1253 85.261
R5228 CLK1.n346 CLK1.n343 85.261
R5229 CLK1.n388 CLK1.n387 85.261
R5230 CLK1.n434 CLK1.n431 85.261
R5231 CLK1.n476 CLK1.n475 85.261
R5232 CLK1.n998 CLK1.n997 85.261
R5233 CLK1.n989 CLK1.n988 85.261
R5234 CLK1.n916 CLK1.n915 85.261
R5235 CLK1.n622 CLK1.n621 85.261
R5236 CLK1.n804 CLK1.n803 85.261
R5237 CLK1.n731 CLK1.n730 85.261
R5238 CLK1.n1436 CLK1.n1435 85.261
R5239 CLK1.n1363 CLK1.n1362 85.261
R5240 CLK1.n1075 CLK1.n1074 69.028
R5241 CLK1.n1076 CLK1.n1075 69.028
R5242 CLK1.n1085 CLK1.n1084 69.028
R5243 CLK1.n1092 CLK1.n1087 69.028
R5244 CLK1.n1094 CLK1.n1093 69.028
R5245 CLK1.n1095 CLK1.n1094 69.028
R5246 CLK1.n1086 CLK1.t86 64.713
R5247 CLK1.t98 CLK1.n1086 64.713
R5248 CLK1.n1084 CLK1.t84 56.085
R5249 CLK1.t96 CLK1.n1092 56.085
R5250 CLK1.n239 CLK1.t165 44.338
R5251 CLK1.n261 CLK1.t19 44.338
R5252 CLK1.n1079 CLK1.t181 44.338
R5253 CLK1.n1090 CLK1.t106 44.338
R5254 CLK1.n702 CLK1.t77 44.338
R5255 CLK1.n671 CLK1.t46 44.338
R5256 CLK1.n649 CLK1.t93 44.338
R5257 CLK1.n776 CLK1.t140 44.338
R5258 CLK1.n447 CLK1.t120 44.338
R5259 CLK1.n416 CLK1.t11 44.338
R5260 CLK1.n494 CLK1.t194 44.338
R5261 CLK1.n503 CLK1.t48 44.338
R5262 CLK1.n1334 CLK1.t174 44.338
R5263 CLK1.n1303 CLK1.t13 44.338
R5264 CLK1.n1281 CLK1.t70 44.338
R5265 CLK1.n1408 CLK1.t133 44.338
R5266 CLK1.n155 CLK1.t5 44.337
R5267 CLK1.n128 CLK1.t64 44.337
R5268 CLK1.n61 CLK1.t111 44.337
R5269 CLK1.n34 CLK1.t189 44.337
R5270 CLK1.n1593 CLK1.t52 44.337
R5271 CLK1.n1466 CLK1.t178 44.337
R5272 CLK1.n1488 CLK1.t3 44.337
R5273 CLK1.n1519 CLK1.t81 44.337
R5274 CLK1.n295 CLK1.t138 44.337
R5275 CLK1.n1214 CLK1.t37 44.337
R5276 CLK1.n328 CLK1.t105 44.337
R5277 CLK1.n359 CLK1.t144 44.337
R5278 CLK1.n1079 CLK1.t85 44.337
R5279 CLK1.n1090 CLK1.t97 44.337
R5280 CLK1.n961 CLK1.t185 44.337
R5281 CLK1.n834 CLK1.t21 44.337
R5282 CLK1.n856 CLK1.t126 44.337
R5283 CLK1.n887 CLK1.t75 44.337
R5284 CLK1.n535 CLK1.t155 44.337
R5285 CLK1.n582 CLK1.t161 44.337
R5286 CLK1.n1176 CLK1.n394 39.834
R5287 CLK1.n1172 CLK1.n394 39.834
R5288 CLK1.n1172 CLK1.n396 39.834
R5289 CLK1.n1165 CLK1.n396 39.834
R5290 CLK1.n1165 CLK1.n1068 39.834
R5291 CLK1.n1161 CLK1.n1068 39.834
R5292 CLK1.n1161 CLK1.n1070 39.834
R5293 CLK1.n1155 CLK1.n1070 39.834
R5294 CLK1.n1155 CLK1.n1154 39.834
R5295 CLK1.n1154 CLK1.n1153 39.834
R5296 CLK1.n1153 CLK1.n1077 39.834
R5297 CLK1.n1147 CLK1.n1077 39.834
R5298 CLK1.n1147 CLK1.n1146 39.834
R5299 CLK1.n1146 CLK1.n1145 39.834
R5300 CLK1.n1145 CLK1.n1088 39.834
R5301 CLK1.n1139 CLK1.n1088 39.834
R5302 CLK1.n1139 CLK1.n1138 39.834
R5303 CLK1.n1138 CLK1.n1137 39.834
R5304 CLK1.n1137 CLK1.n1096 39.834
R5305 CLK1.n1131 CLK1.n1096 39.834
R5306 CLK1.n1131 CLK1.n1102 39.834
R5307 CLK1.n1127 CLK1.n1102 39.834
R5308 CLK1.n1127 CLK1.n1105 39.834
R5309 CLK1.n1120 CLK1.n1105 39.834
R5310 CLK1.n1120 CLK1.n1112 39.834
R5311 CLK1.n1116 CLK1.n1112 39.834
R5312 CLK1.n3 CLK1.t89 39.4
R5313 CLK1.n3 CLK1.t26 39.4
R5314 CLK1.n7 CLK1.t191 39.4
R5315 CLK1.n7 CLK1.t109 39.4
R5316 CLK1.n213 CLK1.t167 39.4
R5317 CLK1.n213 CLK1.t17 39.4
R5318 CLK1.n1580 CLK1.t42 39.4
R5319 CLK1.n1580 CLK1.t151 39.4
R5320 CLK1.n1494 CLK1.t83 39.4
R5321 CLK1.n1494 CLK1.t1 39.4
R5322 CLK1.n301 CLK1.t35 39.4
R5323 CLK1.n301 CLK1.t136 39.4
R5324 CLK1.n1081 CLK1.t87 39.4
R5325 CLK1.n1081 CLK1.t99 39.4
R5326 CLK1.n1080 CLK1.t182 39.4
R5327 CLK1.n1080 CLK1.t107 39.4
R5328 CLK1.n334 CLK1.t146 39.4
R5329 CLK1.n334 CLK1.t103 39.4
R5330 CLK1.n495 CLK1.t124 39.4
R5331 CLK1.n495 CLK1.t142 39.4
R5332 CLK1.n422 CLK1.t122 39.4
R5333 CLK1.n422 CLK1.t9 39.4
R5334 CLK1.n948 CLK1.t113 39.4
R5335 CLK1.n948 CLK1.t39 39.4
R5336 CLK1.n862 CLK1.t73 39.4
R5337 CLK1.n862 CLK1.t128 39.4
R5338 CLK1.n541 CLK1.t159 39.4
R5339 CLK1.n541 CLK1.t157 39.4
R5340 CLK1.n763 CLK1.t153 39.4
R5341 CLK1.n763 CLK1.t180 39.4
R5342 CLK1.n677 CLK1.t79 39.4
R5343 CLK1.n677 CLK1.t44 39.4
R5344 CLK1.n1395 CLK1.t30 39.4
R5345 CLK1.n1395 CLK1.t131 39.4
R5346 CLK1.n1309 CLK1.t176 39.4
R5347 CLK1.n1309 CLK1.t15 39.4
R5348 CLK1.n1117 CLK1.n1114 39.262
R5349 CLK1.n1175 CLK1.n392 38.088
R5350 CLK1.n227 CLK1.t95 30.776
R5351 CLK1.n86 CLK1.t117 30.775
R5352 CLK1.n282 CLK1.t24 30.775
R5353 CLK1.n522 CLK1.t116 30.775
R5354 CLK1.n560 CLK1.t50 30.775
R5355 CLK1.n690 CLK1.t56 29.713
R5356 CLK1.n665 CLK1.t149 29.713
R5357 CLK1.n435 CLK1.t118 29.713
R5358 CLK1.n410 CLK1.t58 29.713
R5359 CLK1.n1322 CLK1.t147 29.713
R5360 CLK1.n1297 CLK1.t115 29.713
R5361 CLK1.n1482 CLK1.t171 29.712
R5362 CLK1.n1507 CLK1.t192 29.712
R5363 CLK1.n322 CLK1.t22 29.712
R5364 CLK1.n347 CLK1.t27 29.712
R5365 CLK1.n850 CLK1.t198 29.712
R5366 CLK1.n875 CLK1.t134 29.712
R5367 CLK1.n129 CLK1.t63 24.568
R5368 CLK1.n151 CLK1.t4 24.568
R5369 CLK1.n35 CLK1.t188 24.568
R5370 CLK1.n57 CLK1.t110 24.568
R5371 CLK1.t164 CLK1.n244 24.568
R5372 CLK1.t18 CLK1.n205 24.568
R5373 CLK1.n1575 CLK1.t177 24.568
R5374 CLK1.n1597 CLK1.t51 24.568
R5375 CLK1.n1514 CLK1.t80 24.568
R5376 CLK1.n1536 CLK1.t2 24.568
R5377 CLK1.n1209 CLK1.t36 24.568
R5378 CLK1.n1231 CLK1.t137 24.568
R5379 CLK1.n354 CLK1.t143 24.568
R5380 CLK1.n376 CLK1.t104 24.568
R5381 CLK1.n442 CLK1.t119 24.568
R5382 CLK1.n464 CLK1.t10 24.568
R5383 CLK1.n1038 CLK1.t193 24.568
R5384 CLK1.n1020 CLK1.t47 24.568
R5385 CLK1.n943 CLK1.t20 24.568
R5386 CLK1.n965 CLK1.t184 24.568
R5387 CLK1.n882 CLK1.t74 24.568
R5388 CLK1.n904 CLK1.t125 24.568
R5389 CLK1.n577 CLK1.t160 24.568
R5390 CLK1.n599 CLK1.t154 24.568
R5391 CLK1.n758 CLK1.t92 24.568
R5392 CLK1.n780 CLK1.t139 24.568
R5393 CLK1.n697 CLK1.t76 24.568
R5394 CLK1.n719 CLK1.t45 24.568
R5395 CLK1.n1390 CLK1.t69 24.568
R5396 CLK1.n1412 CLK1.t132 24.568
R5397 CLK1.n1329 CLK1.t173 24.568
R5398 CLK1.n1351 CLK1.t12 24.568
R5399 CLK1.n0 CLK1.t40 24
R5400 CLK1.n0 CLK1.t100 24
R5401 CLK1.n4 CLK1.t197 24
R5402 CLK1.n4 CLK1.t71 24
R5403 CLK1.n8 CLK1.t57 24
R5404 CLK1.n8 CLK1.t33 24
R5405 CLK1.n201 CLK1.t49 24
R5406 CLK1.n201 CLK1.t60 24
R5407 CLK1.n1449 CLK1.t168 24
R5408 CLK1.n1449 CLK1.t67 24
R5409 CLK1.n1478 CLK1.t91 24
R5410 CLK1.n1478 CLK1.t23 24
R5411 CLK1.n288 CLK1.t163 24
R5412 CLK1.n288 CLK1.t187 24
R5413 CLK1.n1182 CLK1.t170 24
R5414 CLK1.n1099 CLK1.t183 24
R5415 CLK1.n1099 CLK1.t6 24
R5416 CLK1.n1109 CLK1.t114 24
R5417 CLK1.n1109 CLK1.t28 24
R5418 CLK1.n1108 CLK1.t55 24
R5419 CLK1.n1108 CLK1.t31 24
R5420 CLK1.n1057 CLK1.t94 24
R5421 CLK1.n1057 CLK1.t162 24
R5422 CLK1.n817 CLK1.t54 24
R5423 CLK1.n817 CLK1.t148 24
R5424 CLK1.n846 CLK1.t186 24
R5425 CLK1.n846 CLK1.t61 24
R5426 CLK1.n528 CLK1.t66 24
R5427 CLK1.n528 CLK1.t196 24
R5428 CLK1.n661 CLK1.t90 24
R5429 CLK1.n661 CLK1.t195 24
R5430 CLK1.n632 CLK1.t65 24
R5431 CLK1.n632 CLK1.t68 24
R5432 CLK1.n516 CLK1.t129 24
R5433 CLK1.n516 CLK1.t169 24
R5434 CLK1.n1061 CLK1.t7 24
R5435 CLK1.n1061 CLK1.t59 24
R5436 CLK1.n1186 CLK1.t172 24
R5437 CLK1.n1293 CLK1.t32 24
R5438 CLK1.n1293 CLK1.t53 24
R5439 CLK1.n1264 CLK1.t62 24
R5440 CLK1.n1264 CLK1.t101 24
R5441 CLK1.t84 CLK1.n1076 12.942
R5442 CLK1.n1093 CLK1.t96 12.942
R5443 CLK1.n145 CLK1.n142 12.8
R5444 CLK1.n51 CLK1.n48 12.8
R5445 CLK1.n226 CLK1.n225 12.8
R5446 CLK1.n230 CLK1.n225 12.8
R5447 CLK1.n230 CLK1.n221 12.8
R5448 CLK1.n236 CLK1.n221 12.8
R5449 CLK1.n236 CLK1.n219 12.8
R5450 CLK1.n241 CLK1.n219 12.8
R5451 CLK1.n241 CLK1.n215 12.8
R5452 CLK1.n248 CLK1.n215 12.8
R5453 CLK1.n248 CLK1.n212 12.8
R5454 CLK1.n252 CLK1.n212 12.8
R5455 CLK1.n252 CLK1.n209 12.8
R5456 CLK1.n258 CLK1.n209 12.8
R5457 CLK1.n258 CLK1.n207 12.8
R5458 CLK1.n263 CLK1.n207 12.8
R5459 CLK1.n263 CLK1.n203 12.8
R5460 CLK1.n269 CLK1.n203 12.8
R5461 CLK1.n269 CLK1.n200 12.8
R5462 CLK1.n274 CLK1.n200 12.8
R5463 CLK1.n274 CLK1.n196 12.8
R5464 CLK1.n278 CLK1.n196 12.8
R5465 CLK1.n1551 CLK1.n1480 12.8
R5466 CLK1.n1555 CLK1.n1480 12.8
R5467 CLK1.n1555 CLK1.n1477 12.8
R5468 CLK1.n1560 CLK1.n1477 12.8
R5469 CLK1.n1560 CLK1.n1473 12.8
R5470 CLK1.n1566 CLK1.n1473 12.8
R5471 CLK1.n1566 CLK1.n1471 12.8
R5472 CLK1.n1571 CLK1.n1471 12.8
R5473 CLK1.n1571 CLK1.n1467 12.8
R5474 CLK1.n1577 CLK1.n1467 12.8
R5475 CLK1.n1577 CLK1.n1465 12.8
R5476 CLK1.n1583 CLK1.n1465 12.8
R5477 CLK1.n1583 CLK1.n1461 12.8
R5478 CLK1.n1590 CLK1.n1461 12.8
R5479 CLK1.n1590 CLK1.n1460 12.8
R5480 CLK1.n1595 CLK1.n1460 12.8
R5481 CLK1.n1595 CLK1.n1457 12.8
R5482 CLK1.n1601 CLK1.n1457 12.8
R5483 CLK1.n1601 CLK1.n1455 12.8
R5484 CLK1.n1605 CLK1.n1455 12.8
R5485 CLK1.n1605 CLK1.n1451 12.8
R5486 CLK1.n1611 CLK1.n1451 12.8
R5487 CLK1.n1611 CLK1.n1447 12.8
R5488 CLK1.n1617 CLK1.n1447 12.8
R5489 CLK1.n1617 CLK1.n1448 12.8
R5490 CLK1.n1506 CLK1.n1505 12.8
R5491 CLK1.n1510 CLK1.n1505 12.8
R5492 CLK1.n1510 CLK1.n1501 12.8
R5493 CLK1.n1517 CLK1.n1501 12.8
R5494 CLK1.n1517 CLK1.n1499 12.8
R5495 CLK1.n1522 CLK1.n1499 12.8
R5496 CLK1.n1522 CLK1.n1496 12.8
R5497 CLK1.n1528 CLK1.n1496 12.8
R5498 CLK1.n1528 CLK1.n1493 12.8
R5499 CLK1.n1533 CLK1.n1493 12.8
R5500 CLK1.n1533 CLK1.n1489 12.8
R5501 CLK1.n1539 CLK1.n1489 12.8
R5502 CLK1.n1539 CLK1.n1487 12.8
R5503 CLK1.n1544 CLK1.n1487 12.8
R5504 CLK1.n1544 CLK1.n1483 12.8
R5505 CLK1.n1548 CLK1.n1483 12.8
R5506 CLK1.n1191 CLK1.n318 12.8
R5507 CLK1.n1195 CLK1.n318 12.8
R5508 CLK1.n1195 CLK1.n314 12.8
R5509 CLK1.n1201 CLK1.n314 12.8
R5510 CLK1.n1201 CLK1.n312 12.8
R5511 CLK1.n1205 CLK1.n312 12.8
R5512 CLK1.n1205 CLK1.n308 12.8
R5513 CLK1.n1212 CLK1.n308 12.8
R5514 CLK1.n1212 CLK1.n306 12.8
R5515 CLK1.n1217 CLK1.n306 12.8
R5516 CLK1.n1217 CLK1.n303 12.8
R5517 CLK1.n1223 CLK1.n303 12.8
R5518 CLK1.n1223 CLK1.n300 12.8
R5519 CLK1.n1228 CLK1.n300 12.8
R5520 CLK1.n1228 CLK1.n296 12.8
R5521 CLK1.n1234 CLK1.n296 12.8
R5522 CLK1.n1234 CLK1.n294 12.8
R5523 CLK1.n1239 CLK1.n294 12.8
R5524 CLK1.n1239 CLK1.n290 12.8
R5525 CLK1.n1245 CLK1.n290 12.8
R5526 CLK1.n1245 CLK1.n287 12.8
R5527 CLK1.n1250 CLK1.n287 12.8
R5528 CLK1.n1250 CLK1.n283 12.8
R5529 CLK1.n1254 CLK1.n283 12.8
R5530 CLK1.n1181 CLK1.n321 12.8
R5531 CLK1.n346 CLK1.n345 12.8
R5532 CLK1.n350 CLK1.n345 12.8
R5533 CLK1.n350 CLK1.n341 12.8
R5534 CLK1.n357 CLK1.n341 12.8
R5535 CLK1.n357 CLK1.n339 12.8
R5536 CLK1.n362 CLK1.n339 12.8
R5537 CLK1.n362 CLK1.n336 12.8
R5538 CLK1.n368 CLK1.n336 12.8
R5539 CLK1.n368 CLK1.n333 12.8
R5540 CLK1.n373 CLK1.n333 12.8
R5541 CLK1.n373 CLK1.n329 12.8
R5542 CLK1.n379 CLK1.n329 12.8
R5543 CLK1.n379 CLK1.n327 12.8
R5544 CLK1.n384 CLK1.n327 12.8
R5545 CLK1.n384 CLK1.n323 12.8
R5546 CLK1.n388 CLK1.n323 12.8
R5547 CLK1.n1058 CLK1.n400 12.8
R5548 CLK1.n434 CLK1.n433 12.8
R5549 CLK1.n438 CLK1.n433 12.8
R5550 CLK1.n438 CLK1.n429 12.8
R5551 CLK1.n445 CLK1.n429 12.8
R5552 CLK1.n445 CLK1.n427 12.8
R5553 CLK1.n450 CLK1.n427 12.8
R5554 CLK1.n450 CLK1.n424 12.8
R5555 CLK1.n456 CLK1.n424 12.8
R5556 CLK1.n456 CLK1.n421 12.8
R5557 CLK1.n461 CLK1.n421 12.8
R5558 CLK1.n461 CLK1.n417 12.8
R5559 CLK1.n467 CLK1.n417 12.8
R5560 CLK1.n467 CLK1.n415 12.8
R5561 CLK1.n472 CLK1.n415 12.8
R5562 CLK1.n472 CLK1.n411 12.8
R5563 CLK1.n476 CLK1.n411 12.8
R5564 CLK1.n478 CLK1.n409 12.8
R5565 CLK1.n482 CLK1.n409 12.8
R5566 CLK1.n482 CLK1.n403 12.8
R5567 CLK1.n1052 CLK1.n403 12.8
R5568 CLK1.n1052 CLK1.n404 12.8
R5569 CLK1.n1046 CLK1.n404 12.8
R5570 CLK1.n1046 CLK1.n488 12.8
R5571 CLK1.n1042 CLK1.n488 12.8
R5572 CLK1.n1042 CLK1.n490 12.8
R5573 CLK1.n1036 CLK1.n490 12.8
R5574 CLK1.n1036 CLK1.n493 12.8
R5575 CLK1.n1032 CLK1.n493 12.8
R5576 CLK1.n1032 CLK1.n497 12.8
R5577 CLK1.n1026 CLK1.n497 12.8
R5578 CLK1.n1026 CLK1.n502 12.8
R5579 CLK1.n1022 CLK1.n502 12.8
R5580 CLK1.n1022 CLK1.n504 12.8
R5581 CLK1.n1016 CLK1.n504 12.8
R5582 CLK1.n1016 CLK1.n508 12.8
R5583 CLK1.n1012 CLK1.n508 12.8
R5584 CLK1.n1012 CLK1.n511 12.8
R5585 CLK1.n1006 CLK1.n511 12.8
R5586 CLK1.n1006 CLK1.n515 12.8
R5587 CLK1.n1001 CLK1.n515 12.8
R5588 CLK1.n1001 CLK1.n518 12.8
R5589 CLK1.n997 CLK1.n518 12.8
R5590 CLK1.n919 CLK1.n848 12.8
R5591 CLK1.n923 CLK1.n848 12.8
R5592 CLK1.n923 CLK1.n845 12.8
R5593 CLK1.n928 CLK1.n845 12.8
R5594 CLK1.n928 CLK1.n841 12.8
R5595 CLK1.n934 CLK1.n841 12.8
R5596 CLK1.n934 CLK1.n839 12.8
R5597 CLK1.n939 CLK1.n839 12.8
R5598 CLK1.n939 CLK1.n835 12.8
R5599 CLK1.n945 CLK1.n835 12.8
R5600 CLK1.n945 CLK1.n833 12.8
R5601 CLK1.n951 CLK1.n833 12.8
R5602 CLK1.n951 CLK1.n829 12.8
R5603 CLK1.n958 CLK1.n829 12.8
R5604 CLK1.n958 CLK1.n828 12.8
R5605 CLK1.n963 CLK1.n828 12.8
R5606 CLK1.n963 CLK1.n825 12.8
R5607 CLK1.n969 CLK1.n825 12.8
R5608 CLK1.n969 CLK1.n823 12.8
R5609 CLK1.n973 CLK1.n823 12.8
R5610 CLK1.n973 CLK1.n819 12.8
R5611 CLK1.n979 CLK1.n819 12.8
R5612 CLK1.n979 CLK1.n815 12.8
R5613 CLK1.n985 CLK1.n815 12.8
R5614 CLK1.n985 CLK1.n816 12.8
R5615 CLK1.n874 CLK1.n873 12.8
R5616 CLK1.n878 CLK1.n873 12.8
R5617 CLK1.n878 CLK1.n869 12.8
R5618 CLK1.n885 CLK1.n869 12.8
R5619 CLK1.n885 CLK1.n867 12.8
R5620 CLK1.n890 CLK1.n867 12.8
R5621 CLK1.n890 CLK1.n864 12.8
R5622 CLK1.n896 CLK1.n864 12.8
R5623 CLK1.n896 CLK1.n861 12.8
R5624 CLK1.n901 CLK1.n861 12.8
R5625 CLK1.n901 CLK1.n857 12.8
R5626 CLK1.n907 CLK1.n857 12.8
R5627 CLK1.n907 CLK1.n855 12.8
R5628 CLK1.n912 CLK1.n855 12.8
R5629 CLK1.n912 CLK1.n851 12.8
R5630 CLK1.n916 CLK1.n851 12.8
R5631 CLK1.n559 CLK1.n558 12.8
R5632 CLK1.n563 CLK1.n558 12.8
R5633 CLK1.n563 CLK1.n554 12.8
R5634 CLK1.n569 CLK1.n554 12.8
R5635 CLK1.n569 CLK1.n552 12.8
R5636 CLK1.n573 CLK1.n552 12.8
R5637 CLK1.n573 CLK1.n548 12.8
R5638 CLK1.n580 CLK1.n548 12.8
R5639 CLK1.n580 CLK1.n546 12.8
R5640 CLK1.n585 CLK1.n546 12.8
R5641 CLK1.n585 CLK1.n543 12.8
R5642 CLK1.n591 CLK1.n543 12.8
R5643 CLK1.n591 CLK1.n540 12.8
R5644 CLK1.n596 CLK1.n540 12.8
R5645 CLK1.n596 CLK1.n536 12.8
R5646 CLK1.n602 CLK1.n536 12.8
R5647 CLK1.n602 CLK1.n534 12.8
R5648 CLK1.n607 CLK1.n534 12.8
R5649 CLK1.n607 CLK1.n530 12.8
R5650 CLK1.n613 CLK1.n530 12.8
R5651 CLK1.n613 CLK1.n527 12.8
R5652 CLK1.n618 CLK1.n527 12.8
R5653 CLK1.n618 CLK1.n523 12.8
R5654 CLK1.n622 CLK1.n523 12.8
R5655 CLK1.n734 CLK1.n663 12.8
R5656 CLK1.n738 CLK1.n663 12.8
R5657 CLK1.n738 CLK1.n660 12.8
R5658 CLK1.n743 CLK1.n660 12.8
R5659 CLK1.n743 CLK1.n656 12.8
R5660 CLK1.n749 CLK1.n656 12.8
R5661 CLK1.n749 CLK1.n654 12.8
R5662 CLK1.n754 CLK1.n654 12.8
R5663 CLK1.n754 CLK1.n650 12.8
R5664 CLK1.n760 CLK1.n650 12.8
R5665 CLK1.n760 CLK1.n648 12.8
R5666 CLK1.n766 CLK1.n648 12.8
R5667 CLK1.n766 CLK1.n644 12.8
R5668 CLK1.n773 CLK1.n644 12.8
R5669 CLK1.n773 CLK1.n643 12.8
R5670 CLK1.n778 CLK1.n643 12.8
R5671 CLK1.n778 CLK1.n640 12.8
R5672 CLK1.n784 CLK1.n640 12.8
R5673 CLK1.n784 CLK1.n638 12.8
R5674 CLK1.n788 CLK1.n638 12.8
R5675 CLK1.n788 CLK1.n634 12.8
R5676 CLK1.n794 CLK1.n634 12.8
R5677 CLK1.n794 CLK1.n630 12.8
R5678 CLK1.n800 CLK1.n630 12.8
R5679 CLK1.n800 CLK1.n631 12.8
R5680 CLK1.n689 CLK1.n688 12.8
R5681 CLK1.n693 CLK1.n688 12.8
R5682 CLK1.n693 CLK1.n684 12.8
R5683 CLK1.n700 CLK1.n684 12.8
R5684 CLK1.n700 CLK1.n682 12.8
R5685 CLK1.n705 CLK1.n682 12.8
R5686 CLK1.n705 CLK1.n679 12.8
R5687 CLK1.n711 CLK1.n679 12.8
R5688 CLK1.n711 CLK1.n676 12.8
R5689 CLK1.n716 CLK1.n676 12.8
R5690 CLK1.n716 CLK1.n672 12.8
R5691 CLK1.n722 CLK1.n672 12.8
R5692 CLK1.n722 CLK1.n670 12.8
R5693 CLK1.n727 CLK1.n670 12.8
R5694 CLK1.n727 CLK1.n666 12.8
R5695 CLK1.n731 CLK1.n666 12.8
R5696 CLK1.n1063 CLK1.n398 12.8
R5697 CLK1.n1188 CLK1.n1187 12.8
R5698 CLK1.n1366 CLK1.n1295 12.8
R5699 CLK1.n1370 CLK1.n1295 12.8
R5700 CLK1.n1370 CLK1.n1292 12.8
R5701 CLK1.n1375 CLK1.n1292 12.8
R5702 CLK1.n1375 CLK1.n1288 12.8
R5703 CLK1.n1381 CLK1.n1288 12.8
R5704 CLK1.n1381 CLK1.n1286 12.8
R5705 CLK1.n1386 CLK1.n1286 12.8
R5706 CLK1.n1386 CLK1.n1282 12.8
R5707 CLK1.n1392 CLK1.n1282 12.8
R5708 CLK1.n1392 CLK1.n1280 12.8
R5709 CLK1.n1398 CLK1.n1280 12.8
R5710 CLK1.n1398 CLK1.n1276 12.8
R5711 CLK1.n1405 CLK1.n1276 12.8
R5712 CLK1.n1405 CLK1.n1275 12.8
R5713 CLK1.n1410 CLK1.n1275 12.8
R5714 CLK1.n1410 CLK1.n1272 12.8
R5715 CLK1.n1416 CLK1.n1272 12.8
R5716 CLK1.n1416 CLK1.n1270 12.8
R5717 CLK1.n1420 CLK1.n1270 12.8
R5718 CLK1.n1420 CLK1.n1266 12.8
R5719 CLK1.n1426 CLK1.n1266 12.8
R5720 CLK1.n1426 CLK1.n1262 12.8
R5721 CLK1.n1432 CLK1.n1262 12.8
R5722 CLK1.n1432 CLK1.n1263 12.8
R5723 CLK1.n1321 CLK1.n1320 12.8
R5724 CLK1.n1325 CLK1.n1320 12.8
R5725 CLK1.n1325 CLK1.n1316 12.8
R5726 CLK1.n1332 CLK1.n1316 12.8
R5727 CLK1.n1332 CLK1.n1314 12.8
R5728 CLK1.n1337 CLK1.n1314 12.8
R5729 CLK1.n1337 CLK1.n1311 12.8
R5730 CLK1.n1343 CLK1.n1311 12.8
R5731 CLK1.n1343 CLK1.n1308 12.8
R5732 CLK1.n1348 CLK1.n1308 12.8
R5733 CLK1.n1348 CLK1.n1304 12.8
R5734 CLK1.n1354 CLK1.n1304 12.8
R5735 CLK1.n1354 CLK1.n1302 12.8
R5736 CLK1.n1359 CLK1.n1302 12.8
R5737 CLK1.n1359 CLK1.n1298 12.8
R5738 CLK1.n1363 CLK1.n1298 12.8
R5739 CLK1.n1448 CLK1.n1443 11.36
R5740 CLK1.n816 CLK1.n811 11.36
R5741 CLK1.n631 CLK1.n626 11.36
R5742 CLK1.n1263 CLK1.n1258 11.36
R5743 CLK1.n1443 CLK1.n1442 9.3
R5744 CLK1.n811 CLK1.n810 9.3
R5745 CLK1.n626 CLK1.n625 9.3
R5746 CLK1.n1258 CLK1.n1257 9.3
R5747 CLK1.n11 CLK1.n10 8.855
R5748 CLK1.n15 CLK1.n14 8.855
R5749 CLK1.n14 CLK1.n13 8.855
R5750 CLK1.n20 CLK1.n19 8.855
R5751 CLK1.n19 CLK1.n18 8.855
R5752 CLK1.n24 CLK1.n23 8.855
R5753 CLK1.n23 CLK1.n22 8.855
R5754 CLK1.n28 CLK1.n27 8.855
R5755 CLK1.n27 CLK1.n26 8.855
R5756 CLK1.n32 CLK1.n31 8.855
R5757 CLK1.n31 CLK1.n30 8.855
R5758 CLK1.n37 CLK1.n36 8.855
R5759 CLK1.n36 CLK1.n35 8.855
R5760 CLK1.n41 CLK1.n40 8.855
R5761 CLK1.n40 CLK1.n39 8.855
R5762 CLK1.n45 CLK1.n44 8.855
R5763 CLK1.n44 CLK1.n43 8.855
R5764 CLK1.n48 CLK1.n6 8.855
R5765 CLK1.n6 CLK1.n5 8.855
R5766 CLK1.n51 CLK1.n50 8.855
R5767 CLK1.n50 CLK1.n49 8.855
R5768 CLK1.n55 CLK1.n54 8.855
R5769 CLK1.n54 CLK1.n53 8.855
R5770 CLK1.n59 CLK1.n58 8.855
R5771 CLK1.n58 CLK1.n57 8.855
R5772 CLK1.n64 CLK1.n63 8.855
R5773 CLK1.n63 CLK1.n62 8.855
R5774 CLK1.n68 CLK1.n67 8.855
R5775 CLK1.n67 CLK1.n66 8.855
R5776 CLK1.n72 CLK1.n71 8.855
R5777 CLK1.n71 CLK1.n70 8.855
R5778 CLK1.n76 CLK1.n75 8.855
R5779 CLK1.n75 CLK1.n74 8.855
R5780 CLK1.n80 CLK1.n79 8.855
R5781 CLK1.n79 CLK1.n78 8.855
R5782 CLK1.n84 CLK1.n83 8.855
R5783 CLK1.n93 CLK1.n92 8.855
R5784 CLK1.n97 CLK1.n96 8.855
R5785 CLK1.n96 CLK1.n95 8.855
R5786 CLK1.n101 CLK1.n100 8.855
R5787 CLK1.n100 CLK1.n99 8.855
R5788 CLK1.n106 CLK1.n105 8.855
R5789 CLK1.n105 CLK1.n104 8.855
R5790 CLK1.n110 CLK1.n109 8.855
R5791 CLK1.n109 CLK1.n108 8.855
R5792 CLK1.n114 CLK1.n113 8.855
R5793 CLK1.n113 CLK1.n112 8.855
R5794 CLK1.n118 CLK1.n117 8.855
R5795 CLK1.n117 CLK1.n116 8.855
R5796 CLK1.n122 CLK1.n121 8.855
R5797 CLK1.n121 CLK1.n120 8.855
R5798 CLK1.n126 CLK1.n125 8.855
R5799 CLK1.n125 CLK1.n124 8.855
R5800 CLK1.n131 CLK1.n130 8.855
R5801 CLK1.n130 CLK1.n129 8.855
R5802 CLK1.n135 CLK1.n134 8.855
R5803 CLK1.n134 CLK1.n133 8.855
R5804 CLK1.n139 CLK1.n138 8.855
R5805 CLK1.n138 CLK1.n137 8.855
R5806 CLK1.n142 CLK1.n2 8.855
R5807 CLK1.n2 CLK1.n1 8.855
R5808 CLK1.n145 CLK1.n144 8.855
R5809 CLK1.n144 CLK1.n143 8.855
R5810 CLK1.n149 CLK1.n148 8.855
R5811 CLK1.n148 CLK1.n147 8.855
R5812 CLK1.n153 CLK1.n152 8.855
R5813 CLK1.n152 CLK1.n151 8.855
R5814 CLK1.n158 CLK1.n157 8.855
R5815 CLK1.n157 CLK1.n156 8.855
R5816 CLK1.n162 CLK1.n161 8.855
R5817 CLK1.n161 CLK1.n160 8.855
R5818 CLK1.n166 CLK1.n165 8.855
R5819 CLK1.n165 CLK1.n164 8.855
R5820 CLK1.n170 CLK1.n169 8.855
R5821 CLK1.n169 CLK1.n168 8.855
R5822 CLK1.n174 CLK1.n173 8.855
R5823 CLK1.n173 CLK1.n172 8.855
R5824 CLK1.n178 CLK1.n177 8.855
R5825 CLK1.n177 CLK1.n176 8.855
R5826 CLK1.n183 CLK1.n182 8.855
R5827 CLK1.n182 CLK1.n181 8.855
R5828 CLK1.n187 CLK1.n186 8.855
R5829 CLK1.n186 CLK1.n185 8.855
R5830 CLK1.n191 CLK1.n190 8.855
R5831 CLK1.n225 CLK1.n224 8.855
R5832 CLK1.n231 CLK1.n230 8.855
R5833 CLK1.n232 CLK1.n231 8.855
R5834 CLK1.n222 CLK1.n221 8.855
R5835 CLK1.n233 CLK1.n222 8.855
R5836 CLK1.n236 CLK1.n235 8.855
R5837 CLK1.n235 CLK1.n234 8.855
R5838 CLK1.n219 CLK1.n218 8.855
R5839 CLK1.n218 CLK1.n217 8.855
R5840 CLK1.n242 CLK1.n241 8.855
R5841 CLK1.n243 CLK1.n242 8.855
R5842 CLK1.n216 CLK1.n215 8.855
R5843 CLK1.n244 CLK1.n216 8.855
R5844 CLK1.n248 CLK1.n247 8.855
R5845 CLK1.n247 CLK1.n246 8.855
R5846 CLK1.n212 CLK1.n211 8.855
R5847 CLK1.n245 CLK1.n211 8.855
R5848 CLK1.n253 CLK1.n252 8.855
R5849 CLK1.n254 CLK1.n253 8.855
R5850 CLK1.n210 CLK1.n209 8.855
R5851 CLK1.n255 CLK1.n210 8.855
R5852 CLK1.n258 CLK1.n257 8.855
R5853 CLK1.n257 CLK1.n256 8.855
R5854 CLK1.n207 CLK1.n206 8.855
R5855 CLK1.n206 CLK1.n205 8.855
R5856 CLK1.n264 CLK1.n263 8.855
R5857 CLK1.n265 CLK1.n264 8.855
R5858 CLK1.n204 CLK1.n203 8.855
R5859 CLK1.n266 CLK1.n204 8.855
R5860 CLK1.n269 CLK1.n268 8.855
R5861 CLK1.n268 CLK1.n267 8.855
R5862 CLK1.n200 CLK1.n199 8.855
R5863 CLK1.n199 CLK1.n198 8.855
R5864 CLK1.n275 CLK1.n274 8.855
R5865 CLK1.n276 CLK1.n275 8.855
R5866 CLK1.n197 CLK1.n196 8.855
R5867 CLK1.n1505 CLK1.n1504 8.855
R5868 CLK1.n1511 CLK1.n1510 8.855
R5869 CLK1.n1512 CLK1.n1511 8.855
R5870 CLK1.n1502 CLK1.n1501 8.855
R5871 CLK1.n1513 CLK1.n1502 8.855
R5872 CLK1.n1517 CLK1.n1516 8.855
R5873 CLK1.n1516 CLK1.n1515 8.855
R5874 CLK1.n1499 CLK1.n1498 8.855
R5875 CLK1.n1514 CLK1.n1498 8.855
R5876 CLK1.n1523 CLK1.n1522 8.855
R5877 CLK1.n1524 CLK1.n1523 8.855
R5878 CLK1.n1497 CLK1.n1496 8.855
R5879 CLK1.n1525 CLK1.n1497 8.855
R5880 CLK1.n1528 CLK1.n1527 8.855
R5881 CLK1.n1527 CLK1.n1526 8.855
R5882 CLK1.n1493 CLK1.n1492 8.855
R5883 CLK1.n1492 CLK1.n1491 8.855
R5884 CLK1.n1534 CLK1.n1533 8.855
R5885 CLK1.n1535 CLK1.n1534 8.855
R5886 CLK1.n1490 CLK1.n1489 8.855
R5887 CLK1.n1536 CLK1.n1490 8.855
R5888 CLK1.n1539 CLK1.n1538 8.855
R5889 CLK1.n1538 CLK1.n1537 8.855
R5890 CLK1.n1487 CLK1.n1486 8.855
R5891 CLK1.n1486 CLK1.n1485 8.855
R5892 CLK1.n1545 CLK1.n1544 8.855
R5893 CLK1.n1546 CLK1.n1545 8.855
R5894 CLK1.n1484 CLK1.n1483 8.855
R5895 CLK1.n1481 CLK1.n1480 8.855
R5896 CLK1.n1555 CLK1.n1554 8.855
R5897 CLK1.n1554 CLK1.n1553 8.855
R5898 CLK1.n1477 CLK1.n1476 8.855
R5899 CLK1.n1476 CLK1.n1475 8.855
R5900 CLK1.n1561 CLK1.n1560 8.855
R5901 CLK1.n1562 CLK1.n1561 8.855
R5902 CLK1.n1474 CLK1.n1473 8.855
R5903 CLK1.n1563 CLK1.n1474 8.855
R5904 CLK1.n1566 CLK1.n1565 8.855
R5905 CLK1.n1565 CLK1.n1564 8.855
R5906 CLK1.n1471 CLK1.n1470 8.855
R5907 CLK1.n1470 CLK1.n1469 8.855
R5908 CLK1.n1572 CLK1.n1571 8.855
R5909 CLK1.n1573 CLK1.n1572 8.855
R5910 CLK1.n1468 CLK1.n1467 8.855
R5911 CLK1.n1574 CLK1.n1468 8.855
R5912 CLK1.n1577 CLK1.n1576 8.855
R5913 CLK1.n1576 CLK1.n1575 8.855
R5914 CLK1.n1465 CLK1.n1464 8.855
R5915 CLK1.n1464 CLK1.n1463 8.855
R5916 CLK1.n1584 CLK1.n1583 8.855
R5917 CLK1.n1585 CLK1.n1584 8.855
R5918 CLK1.n1462 CLK1.n1461 8.855
R5919 CLK1.n1586 CLK1.n1462 8.855
R5920 CLK1.n1590 CLK1.n1589 8.855
R5921 CLK1.n1589 CLK1.n1588 8.855
R5922 CLK1.n1460 CLK1.n1459 8.855
R5923 CLK1.n1587 CLK1.n1459 8.855
R5924 CLK1.n1596 CLK1.n1595 8.855
R5925 CLK1.n1597 CLK1.n1596 8.855
R5926 CLK1.n1458 CLK1.n1457 8.855
R5927 CLK1.n1598 CLK1.n1458 8.855
R5928 CLK1.n1601 CLK1.n1600 8.855
R5929 CLK1.n1600 CLK1.n1599 8.855
R5930 CLK1.n1455 CLK1.n1454 8.855
R5931 CLK1.n1454 CLK1.n1453 8.855
R5932 CLK1.n1606 CLK1.n1605 8.855
R5933 CLK1.n1607 CLK1.n1606 8.855
R5934 CLK1.n1452 CLK1.n1451 8.855
R5935 CLK1.n1608 CLK1.n1452 8.855
R5936 CLK1.n1611 CLK1.n1610 8.855
R5937 CLK1.n1610 CLK1.n1609 8.855
R5938 CLK1.n1447 CLK1.n1446 8.855
R5939 CLK1.n1446 CLK1.n1445 8.855
R5940 CLK1.n1618 CLK1.n1617 8.855
R5941 CLK1.n1619 CLK1.n1618 8.855
R5942 CLK1.n1448 CLK1.n1444 8.855
R5943 CLK1.n1182 CLK1.n1181 8.855
R5944 CLK1.n345 CLK1.n344 8.855
R5945 CLK1.n351 CLK1.n350 8.855
R5946 CLK1.n352 CLK1.n351 8.855
R5947 CLK1.n342 CLK1.n341 8.855
R5948 CLK1.n353 CLK1.n342 8.855
R5949 CLK1.n357 CLK1.n356 8.855
R5950 CLK1.n356 CLK1.n355 8.855
R5951 CLK1.n339 CLK1.n338 8.855
R5952 CLK1.n354 CLK1.n338 8.855
R5953 CLK1.n363 CLK1.n362 8.855
R5954 CLK1.n364 CLK1.n363 8.855
R5955 CLK1.n337 CLK1.n336 8.855
R5956 CLK1.n365 CLK1.n337 8.855
R5957 CLK1.n368 CLK1.n367 8.855
R5958 CLK1.n367 CLK1.n366 8.855
R5959 CLK1.n333 CLK1.n332 8.855
R5960 CLK1.n332 CLK1.n331 8.855
R5961 CLK1.n374 CLK1.n373 8.855
R5962 CLK1.n375 CLK1.n374 8.855
R5963 CLK1.n330 CLK1.n329 8.855
R5964 CLK1.n376 CLK1.n330 8.855
R5965 CLK1.n379 CLK1.n378 8.855
R5966 CLK1.n378 CLK1.n377 8.855
R5967 CLK1.n327 CLK1.n326 8.855
R5968 CLK1.n326 CLK1.n325 8.855
R5969 CLK1.n385 CLK1.n384 8.855
R5970 CLK1.n386 CLK1.n385 8.855
R5971 CLK1.n324 CLK1.n323 8.855
R5972 CLK1.n1058 CLK1.n1057 8.855
R5973 CLK1.n433 CLK1.n432 8.855
R5974 CLK1.n519 CLK1.n518 8.855
R5975 CLK1.n873 CLK1.n872 8.855
R5976 CLK1.n879 CLK1.n878 8.855
R5977 CLK1.n880 CLK1.n879 8.855
R5978 CLK1.n870 CLK1.n869 8.855
R5979 CLK1.n881 CLK1.n870 8.855
R5980 CLK1.n885 CLK1.n884 8.855
R5981 CLK1.n884 CLK1.n883 8.855
R5982 CLK1.n867 CLK1.n866 8.855
R5983 CLK1.n882 CLK1.n866 8.855
R5984 CLK1.n891 CLK1.n890 8.855
R5985 CLK1.n892 CLK1.n891 8.855
R5986 CLK1.n865 CLK1.n864 8.855
R5987 CLK1.n893 CLK1.n865 8.855
R5988 CLK1.n896 CLK1.n895 8.855
R5989 CLK1.n895 CLK1.n894 8.855
R5990 CLK1.n861 CLK1.n860 8.855
R5991 CLK1.n860 CLK1.n859 8.855
R5992 CLK1.n902 CLK1.n901 8.855
R5993 CLK1.n903 CLK1.n902 8.855
R5994 CLK1.n858 CLK1.n857 8.855
R5995 CLK1.n904 CLK1.n858 8.855
R5996 CLK1.n907 CLK1.n906 8.855
R5997 CLK1.n906 CLK1.n905 8.855
R5998 CLK1.n855 CLK1.n854 8.855
R5999 CLK1.n854 CLK1.n853 8.855
R6000 CLK1.n913 CLK1.n912 8.855
R6001 CLK1.n914 CLK1.n913 8.855
R6002 CLK1.n852 CLK1.n851 8.855
R6003 CLK1.n849 CLK1.n848 8.855
R6004 CLK1.n923 CLK1.n922 8.855
R6005 CLK1.n922 CLK1.n921 8.855
R6006 CLK1.n845 CLK1.n844 8.855
R6007 CLK1.n844 CLK1.n843 8.855
R6008 CLK1.n929 CLK1.n928 8.855
R6009 CLK1.n930 CLK1.n929 8.855
R6010 CLK1.n842 CLK1.n841 8.855
R6011 CLK1.n931 CLK1.n842 8.855
R6012 CLK1.n934 CLK1.n933 8.855
R6013 CLK1.n933 CLK1.n932 8.855
R6014 CLK1.n839 CLK1.n838 8.855
R6015 CLK1.n838 CLK1.n837 8.855
R6016 CLK1.n940 CLK1.n939 8.855
R6017 CLK1.n941 CLK1.n940 8.855
R6018 CLK1.n836 CLK1.n835 8.855
R6019 CLK1.n942 CLK1.n836 8.855
R6020 CLK1.n945 CLK1.n944 8.855
R6021 CLK1.n944 CLK1.n943 8.855
R6022 CLK1.n833 CLK1.n832 8.855
R6023 CLK1.n832 CLK1.n831 8.855
R6024 CLK1.n952 CLK1.n951 8.855
R6025 CLK1.n953 CLK1.n952 8.855
R6026 CLK1.n830 CLK1.n829 8.855
R6027 CLK1.n954 CLK1.n830 8.855
R6028 CLK1.n958 CLK1.n957 8.855
R6029 CLK1.n957 CLK1.n956 8.855
R6030 CLK1.n828 CLK1.n827 8.855
R6031 CLK1.n955 CLK1.n827 8.855
R6032 CLK1.n964 CLK1.n963 8.855
R6033 CLK1.n965 CLK1.n964 8.855
R6034 CLK1.n826 CLK1.n825 8.855
R6035 CLK1.n966 CLK1.n826 8.855
R6036 CLK1.n969 CLK1.n968 8.855
R6037 CLK1.n968 CLK1.n967 8.855
R6038 CLK1.n823 CLK1.n822 8.855
R6039 CLK1.n822 CLK1.n821 8.855
R6040 CLK1.n974 CLK1.n973 8.855
R6041 CLK1.n975 CLK1.n974 8.855
R6042 CLK1.n820 CLK1.n819 8.855
R6043 CLK1.n976 CLK1.n820 8.855
R6044 CLK1.n979 CLK1.n978 8.855
R6045 CLK1.n978 CLK1.n977 8.855
R6046 CLK1.n815 CLK1.n814 8.855
R6047 CLK1.n814 CLK1.n813 8.855
R6048 CLK1.n986 CLK1.n985 8.855
R6049 CLK1.n987 CLK1.n986 8.855
R6050 CLK1.n816 CLK1.n812 8.855
R6051 CLK1.n558 CLK1.n557 8.855
R6052 CLK1.n564 CLK1.n563 8.855
R6053 CLK1.n565 CLK1.n564 8.855
R6054 CLK1.n555 CLK1.n554 8.855
R6055 CLK1.n566 CLK1.n555 8.855
R6056 CLK1.n569 CLK1.n568 8.855
R6057 CLK1.n568 CLK1.n567 8.855
R6058 CLK1.n552 CLK1.n551 8.855
R6059 CLK1.n551 CLK1.n550 8.855
R6060 CLK1.n574 CLK1.n573 8.855
R6061 CLK1.n575 CLK1.n574 8.855
R6062 CLK1.n549 CLK1.n548 8.855
R6063 CLK1.n576 CLK1.n549 8.855
R6064 CLK1.n580 CLK1.n579 8.855
R6065 CLK1.n579 CLK1.n578 8.855
R6066 CLK1.n546 CLK1.n545 8.855
R6067 CLK1.n577 CLK1.n545 8.855
R6068 CLK1.n586 CLK1.n585 8.855
R6069 CLK1.n587 CLK1.n586 8.855
R6070 CLK1.n544 CLK1.n543 8.855
R6071 CLK1.n588 CLK1.n544 8.855
R6072 CLK1.n591 CLK1.n590 8.855
R6073 CLK1.n590 CLK1.n589 8.855
R6074 CLK1.n540 CLK1.n539 8.855
R6075 CLK1.n539 CLK1.n538 8.855
R6076 CLK1.n597 CLK1.n596 8.855
R6077 CLK1.n598 CLK1.n597 8.855
R6078 CLK1.n537 CLK1.n536 8.855
R6079 CLK1.n599 CLK1.n537 8.855
R6080 CLK1.n602 CLK1.n601 8.855
R6081 CLK1.n601 CLK1.n600 8.855
R6082 CLK1.n534 CLK1.n533 8.855
R6083 CLK1.n533 CLK1.n532 8.855
R6084 CLK1.n608 CLK1.n607 8.855
R6085 CLK1.n609 CLK1.n608 8.855
R6086 CLK1.n531 CLK1.n530 8.855
R6087 CLK1.n610 CLK1.n531 8.855
R6088 CLK1.n613 CLK1.n612 8.855
R6089 CLK1.n612 CLK1.n611 8.855
R6090 CLK1.n527 CLK1.n526 8.855
R6091 CLK1.n526 CLK1.n525 8.855
R6092 CLK1.n619 CLK1.n618 8.855
R6093 CLK1.n620 CLK1.n619 8.855
R6094 CLK1.n524 CLK1.n523 8.855
R6095 CLK1.n688 CLK1.n687 8.855
R6096 CLK1.n694 CLK1.n693 8.855
R6097 CLK1.n695 CLK1.n694 8.855
R6098 CLK1.n685 CLK1.n684 8.855
R6099 CLK1.n696 CLK1.n685 8.855
R6100 CLK1.n700 CLK1.n699 8.855
R6101 CLK1.n699 CLK1.n698 8.855
R6102 CLK1.n682 CLK1.n681 8.855
R6103 CLK1.n697 CLK1.n681 8.855
R6104 CLK1.n706 CLK1.n705 8.855
R6105 CLK1.n707 CLK1.n706 8.855
R6106 CLK1.n680 CLK1.n679 8.855
R6107 CLK1.n708 CLK1.n680 8.855
R6108 CLK1.n711 CLK1.n710 8.855
R6109 CLK1.n710 CLK1.n709 8.855
R6110 CLK1.n676 CLK1.n675 8.855
R6111 CLK1.n675 CLK1.n674 8.855
R6112 CLK1.n717 CLK1.n716 8.855
R6113 CLK1.n718 CLK1.n717 8.855
R6114 CLK1.n673 CLK1.n672 8.855
R6115 CLK1.n719 CLK1.n673 8.855
R6116 CLK1.n722 CLK1.n721 8.855
R6117 CLK1.n721 CLK1.n720 8.855
R6118 CLK1.n670 CLK1.n669 8.855
R6119 CLK1.n669 CLK1.n668 8.855
R6120 CLK1.n728 CLK1.n727 8.855
R6121 CLK1.n729 CLK1.n728 8.855
R6122 CLK1.n667 CLK1.n666 8.855
R6123 CLK1.n664 CLK1.n663 8.855
R6124 CLK1.n738 CLK1.n737 8.855
R6125 CLK1.n737 CLK1.n736 8.855
R6126 CLK1.n660 CLK1.n659 8.855
R6127 CLK1.n659 CLK1.n658 8.855
R6128 CLK1.n744 CLK1.n743 8.855
R6129 CLK1.n745 CLK1.n744 8.855
R6130 CLK1.n657 CLK1.n656 8.855
R6131 CLK1.n746 CLK1.n657 8.855
R6132 CLK1.n749 CLK1.n748 8.855
R6133 CLK1.n748 CLK1.n747 8.855
R6134 CLK1.n654 CLK1.n653 8.855
R6135 CLK1.n653 CLK1.n652 8.855
R6136 CLK1.n755 CLK1.n754 8.855
R6137 CLK1.n756 CLK1.n755 8.855
R6138 CLK1.n651 CLK1.n650 8.855
R6139 CLK1.n757 CLK1.n651 8.855
R6140 CLK1.n760 CLK1.n759 8.855
R6141 CLK1.n759 CLK1.n758 8.855
R6142 CLK1.n648 CLK1.n647 8.855
R6143 CLK1.n647 CLK1.n646 8.855
R6144 CLK1.n767 CLK1.n766 8.855
R6145 CLK1.n768 CLK1.n767 8.855
R6146 CLK1.n645 CLK1.n644 8.855
R6147 CLK1.n769 CLK1.n645 8.855
R6148 CLK1.n773 CLK1.n772 8.855
R6149 CLK1.n772 CLK1.n771 8.855
R6150 CLK1.n643 CLK1.n642 8.855
R6151 CLK1.n770 CLK1.n642 8.855
R6152 CLK1.n779 CLK1.n778 8.855
R6153 CLK1.n780 CLK1.n779 8.855
R6154 CLK1.n641 CLK1.n640 8.855
R6155 CLK1.n781 CLK1.n641 8.855
R6156 CLK1.n784 CLK1.n783 8.855
R6157 CLK1.n783 CLK1.n782 8.855
R6158 CLK1.n638 CLK1.n637 8.855
R6159 CLK1.n637 CLK1.n636 8.855
R6160 CLK1.n789 CLK1.n788 8.855
R6161 CLK1.n790 CLK1.n789 8.855
R6162 CLK1.n635 CLK1.n634 8.855
R6163 CLK1.n791 CLK1.n635 8.855
R6164 CLK1.n794 CLK1.n793 8.855
R6165 CLK1.n793 CLK1.n792 8.855
R6166 CLK1.n630 CLK1.n629 8.855
R6167 CLK1.n629 CLK1.n628 8.855
R6168 CLK1.n801 CLK1.n800 8.855
R6169 CLK1.n802 CLK1.n801 8.855
R6170 CLK1.n631 CLK1.n627 8.855
R6171 CLK1.n439 CLK1.n438 8.855
R6172 CLK1.n440 CLK1.n439 8.855
R6173 CLK1.n430 CLK1.n429 8.855
R6174 CLK1.n441 CLK1.n430 8.855
R6175 CLK1.n445 CLK1.n444 8.855
R6176 CLK1.n444 CLK1.n443 8.855
R6177 CLK1.n427 CLK1.n426 8.855
R6178 CLK1.n442 CLK1.n426 8.855
R6179 CLK1.n451 CLK1.n450 8.855
R6180 CLK1.n452 CLK1.n451 8.855
R6181 CLK1.n425 CLK1.n424 8.855
R6182 CLK1.n453 CLK1.n425 8.855
R6183 CLK1.n456 CLK1.n455 8.855
R6184 CLK1.n455 CLK1.n454 8.855
R6185 CLK1.n421 CLK1.n420 8.855
R6186 CLK1.n420 CLK1.n419 8.855
R6187 CLK1.n462 CLK1.n461 8.855
R6188 CLK1.n463 CLK1.n462 8.855
R6189 CLK1.n418 CLK1.n417 8.855
R6190 CLK1.n464 CLK1.n418 8.855
R6191 CLK1.n467 CLK1.n466 8.855
R6192 CLK1.n466 CLK1.n465 8.855
R6193 CLK1.n415 CLK1.n414 8.855
R6194 CLK1.n414 CLK1.n413 8.855
R6195 CLK1.n473 CLK1.n472 8.855
R6196 CLK1.n474 CLK1.n473 8.855
R6197 CLK1.n412 CLK1.n411 8.855
R6198 CLK1.n409 CLK1.n408 8.855
R6199 CLK1.n483 CLK1.n482 8.855
R6200 CLK1.n484 CLK1.n483 8.855
R6201 CLK1.n405 CLK1.n403 8.855
R6202 CLK1.n485 CLK1.n405 8.855
R6203 CLK1.n1052 CLK1.n1051 8.855
R6204 CLK1.n1051 CLK1.n1050 8.855
R6205 CLK1.n406 CLK1.n404 8.855
R6206 CLK1.n1049 CLK1.n406 8.855
R6207 CLK1.n1047 CLK1.n1046 8.855
R6208 CLK1.n1048 CLK1.n1047 8.855
R6209 CLK1.n488 CLK1.n487 8.855
R6210 CLK1.n487 CLK1.n486 8.855
R6211 CLK1.n1042 CLK1.n1041 8.855
R6212 CLK1.n1041 CLK1.n1040 8.855
R6213 CLK1.n491 CLK1.n490 8.855
R6214 CLK1.n1039 CLK1.n491 8.855
R6215 CLK1.n1037 CLK1.n1036 8.855
R6216 CLK1.n1038 CLK1.n1037 8.855
R6217 CLK1.n493 CLK1.n492 8.855
R6218 CLK1.n499 CLK1.n492 8.855
R6219 CLK1.n1032 CLK1.n1031 8.855
R6220 CLK1.n1031 CLK1.n1030 8.855
R6221 CLK1.n498 CLK1.n497 8.855
R6222 CLK1.n1029 CLK1.n498 8.855
R6223 CLK1.n1027 CLK1.n1026 8.855
R6224 CLK1.n1028 CLK1.n1027 8.855
R6225 CLK1.n502 CLK1.n501 8.855
R6226 CLK1.n501 CLK1.n500 8.855
R6227 CLK1.n1022 CLK1.n1021 8.855
R6228 CLK1.n1021 CLK1.n1020 8.855
R6229 CLK1.n505 CLK1.n504 8.855
R6230 CLK1.n1019 CLK1.n505 8.855
R6231 CLK1.n1017 CLK1.n1016 8.855
R6232 CLK1.n1018 CLK1.n1017 8.855
R6233 CLK1.n508 CLK1.n507 8.855
R6234 CLK1.n507 CLK1.n506 8.855
R6235 CLK1.n1012 CLK1.n1011 8.855
R6236 CLK1.n1011 CLK1.n1010 8.855
R6237 CLK1.n512 CLK1.n511 8.855
R6238 CLK1.n1009 CLK1.n512 8.855
R6239 CLK1.n1007 CLK1.n1006 8.855
R6240 CLK1.n1008 CLK1.n1007 8.855
R6241 CLK1.n515 CLK1.n514 8.855
R6242 CLK1.n514 CLK1.n513 8.855
R6243 CLK1.n1001 CLK1.n1000 8.855
R6244 CLK1.n1000 CLK1.n999 8.855
R6245 CLK1.n1061 CLK1.n398 8.855
R6246 CLK1.n1187 CLK1.n1186 8.855
R6247 CLK1.n318 CLK1.n317 8.855
R6248 CLK1.n1196 CLK1.n1195 8.855
R6249 CLK1.n1197 CLK1.n1196 8.855
R6250 CLK1.n315 CLK1.n314 8.855
R6251 CLK1.n1198 CLK1.n315 8.855
R6252 CLK1.n1201 CLK1.n1200 8.855
R6253 CLK1.n1200 CLK1.n1199 8.855
R6254 CLK1.n312 CLK1.n311 8.855
R6255 CLK1.n311 CLK1.n310 8.855
R6256 CLK1.n1206 CLK1.n1205 8.855
R6257 CLK1.n1207 CLK1.n1206 8.855
R6258 CLK1.n309 CLK1.n308 8.855
R6259 CLK1.n1208 CLK1.n309 8.855
R6260 CLK1.n1212 CLK1.n1211 8.855
R6261 CLK1.n1211 CLK1.n1210 8.855
R6262 CLK1.n306 CLK1.n305 8.855
R6263 CLK1.n1209 CLK1.n305 8.855
R6264 CLK1.n1218 CLK1.n1217 8.855
R6265 CLK1.n1219 CLK1.n1218 8.855
R6266 CLK1.n304 CLK1.n303 8.855
R6267 CLK1.n1220 CLK1.n304 8.855
R6268 CLK1.n1223 CLK1.n1222 8.855
R6269 CLK1.n1222 CLK1.n1221 8.855
R6270 CLK1.n300 CLK1.n299 8.855
R6271 CLK1.n299 CLK1.n298 8.855
R6272 CLK1.n1229 CLK1.n1228 8.855
R6273 CLK1.n1230 CLK1.n1229 8.855
R6274 CLK1.n297 CLK1.n296 8.855
R6275 CLK1.n1231 CLK1.n297 8.855
R6276 CLK1.n1234 CLK1.n1233 8.855
R6277 CLK1.n1233 CLK1.n1232 8.855
R6278 CLK1.n294 CLK1.n293 8.855
R6279 CLK1.n293 CLK1.n292 8.855
R6280 CLK1.n1240 CLK1.n1239 8.855
R6281 CLK1.n1241 CLK1.n1240 8.855
R6282 CLK1.n291 CLK1.n290 8.855
R6283 CLK1.n1242 CLK1.n291 8.855
R6284 CLK1.n1245 CLK1.n1244 8.855
R6285 CLK1.n1244 CLK1.n1243 8.855
R6286 CLK1.n287 CLK1.n286 8.855
R6287 CLK1.n286 CLK1.n285 8.855
R6288 CLK1.n1251 CLK1.n1250 8.855
R6289 CLK1.n1252 CLK1.n1251 8.855
R6290 CLK1.n284 CLK1.n283 8.855
R6291 CLK1.n1320 CLK1.n1319 8.855
R6292 CLK1.n1326 CLK1.n1325 8.855
R6293 CLK1.n1327 CLK1.n1326 8.855
R6294 CLK1.n1317 CLK1.n1316 8.855
R6295 CLK1.n1328 CLK1.n1317 8.855
R6296 CLK1.n1332 CLK1.n1331 8.855
R6297 CLK1.n1331 CLK1.n1330 8.855
R6298 CLK1.n1314 CLK1.n1313 8.855
R6299 CLK1.n1329 CLK1.n1313 8.855
R6300 CLK1.n1338 CLK1.n1337 8.855
R6301 CLK1.n1339 CLK1.n1338 8.855
R6302 CLK1.n1312 CLK1.n1311 8.855
R6303 CLK1.n1340 CLK1.n1312 8.855
R6304 CLK1.n1343 CLK1.n1342 8.855
R6305 CLK1.n1342 CLK1.n1341 8.855
R6306 CLK1.n1308 CLK1.n1307 8.855
R6307 CLK1.n1307 CLK1.n1306 8.855
R6308 CLK1.n1349 CLK1.n1348 8.855
R6309 CLK1.n1350 CLK1.n1349 8.855
R6310 CLK1.n1305 CLK1.n1304 8.855
R6311 CLK1.n1351 CLK1.n1305 8.855
R6312 CLK1.n1354 CLK1.n1353 8.855
R6313 CLK1.n1353 CLK1.n1352 8.855
R6314 CLK1.n1302 CLK1.n1301 8.855
R6315 CLK1.n1301 CLK1.n1300 8.855
R6316 CLK1.n1360 CLK1.n1359 8.855
R6317 CLK1.n1361 CLK1.n1360 8.855
R6318 CLK1.n1299 CLK1.n1298 8.855
R6319 CLK1.n1296 CLK1.n1295 8.855
R6320 CLK1.n1370 CLK1.n1369 8.855
R6321 CLK1.n1369 CLK1.n1368 8.855
R6322 CLK1.n1292 CLK1.n1291 8.855
R6323 CLK1.n1291 CLK1.n1290 8.855
R6324 CLK1.n1376 CLK1.n1375 8.855
R6325 CLK1.n1377 CLK1.n1376 8.855
R6326 CLK1.n1289 CLK1.n1288 8.855
R6327 CLK1.n1378 CLK1.n1289 8.855
R6328 CLK1.n1381 CLK1.n1380 8.855
R6329 CLK1.n1380 CLK1.n1379 8.855
R6330 CLK1.n1286 CLK1.n1285 8.855
R6331 CLK1.n1285 CLK1.n1284 8.855
R6332 CLK1.n1387 CLK1.n1386 8.855
R6333 CLK1.n1388 CLK1.n1387 8.855
R6334 CLK1.n1283 CLK1.n1282 8.855
R6335 CLK1.n1389 CLK1.n1283 8.855
R6336 CLK1.n1392 CLK1.n1391 8.855
R6337 CLK1.n1391 CLK1.n1390 8.855
R6338 CLK1.n1280 CLK1.n1279 8.855
R6339 CLK1.n1279 CLK1.n1278 8.855
R6340 CLK1.n1399 CLK1.n1398 8.855
R6341 CLK1.n1400 CLK1.n1399 8.855
R6342 CLK1.n1277 CLK1.n1276 8.855
R6343 CLK1.n1401 CLK1.n1277 8.855
R6344 CLK1.n1405 CLK1.n1404 8.855
R6345 CLK1.n1404 CLK1.n1403 8.855
R6346 CLK1.n1275 CLK1.n1274 8.855
R6347 CLK1.n1402 CLK1.n1274 8.855
R6348 CLK1.n1411 CLK1.n1410 8.855
R6349 CLK1.n1412 CLK1.n1411 8.855
R6350 CLK1.n1273 CLK1.n1272 8.855
R6351 CLK1.n1413 CLK1.n1273 8.855
R6352 CLK1.n1416 CLK1.n1415 8.855
R6353 CLK1.n1415 CLK1.n1414 8.855
R6354 CLK1.n1270 CLK1.n1269 8.855
R6355 CLK1.n1269 CLK1.n1268 8.855
R6356 CLK1.n1421 CLK1.n1420 8.855
R6357 CLK1.n1422 CLK1.n1421 8.855
R6358 CLK1.n1267 CLK1.n1266 8.855
R6359 CLK1.n1423 CLK1.n1267 8.855
R6360 CLK1.n1426 CLK1.n1425 8.855
R6361 CLK1.n1425 CLK1.n1424 8.855
R6362 CLK1.n1262 CLK1.n1261 8.855
R6363 CLK1.n1261 CLK1.n1260 8.855
R6364 CLK1.n1433 CLK1.n1432 8.855
R6365 CLK1.n1434 CLK1.n1433 8.855
R6366 CLK1.n1263 CLK1.n1259 8.855
R6367 CLK1.n1056 CLK1.n1055 8.365
R6368 CLK1.n1190 CLK1.n319 8.365
R6369 CLK1.n137 CLK1.t88 8.189
R6370 CLK1.n143 CLK1.t25 8.189
R6371 CLK1.n43 CLK1.t190 8.189
R6372 CLK1.n49 CLK1.t108 8.189
R6373 CLK1.n245 CLK1.t166 8.189
R6374 CLK1.n255 CLK1.t16 8.189
R6375 CLK1.t41 CLK1.n1585 8.189
R6376 CLK1.n1588 CLK1.t150 8.189
R6377 CLK1.t82 CLK1.n1525 8.189
R6378 CLK1.t0 CLK1.n1491 8.189
R6379 CLK1.t34 CLK1.n1220 8.189
R6380 CLK1.t135 CLK1.n298 8.189
R6381 CLK1.t145 CLK1.n365 8.189
R6382 CLK1.t102 CLK1.n331 8.189
R6383 CLK1.t121 CLK1.n453 8.189
R6384 CLK1.t8 CLK1.n419 8.189
R6385 CLK1.n1030 CLK1.t123 8.189
R6386 CLK1.t141 CLK1.n1028 8.189
R6387 CLK1.t112 CLK1.n953 8.189
R6388 CLK1.n956 CLK1.t38 8.189
R6389 CLK1.t72 CLK1.n893 8.189
R6390 CLK1.t127 CLK1.n859 8.189
R6391 CLK1.t158 CLK1.n588 8.189
R6392 CLK1.t156 CLK1.n538 8.189
R6393 CLK1.t152 CLK1.n768 8.189
R6394 CLK1.n771 CLK1.t179 8.189
R6395 CLK1.t78 CLK1.n708 8.189
R6396 CLK1.t43 CLK1.n674 8.189
R6397 CLK1.t29 CLK1.n1400 8.189
R6398 CLK1.n1403 CLK1.t130 8.189
R6399 CLK1.t175 CLK1.n1340 8.189
R6400 CLK1.t14 CLK1.n1306 8.189
R6401 CLK1.n1100 CLK1.n1099 7.776
R6402 CLK1.n1110 CLK1.n1109 7.776
R6403 CLK1.n180 CLK1.n0 6.776
R6404 CLK1.n103 CLK1.n4 6.776
R6405 CLK1.n17 CLK1.n8 6.776
R6406 CLK1.n272 CLK1.n201 6.776
R6407 CLK1.n1613 CLK1.n1449 6.776
R6408 CLK1.n1558 CLK1.n1478 6.776
R6409 CLK1.n289 CLK1.n288 6.776
R6410 CLK1.n1124 CLK1.n1108 6.776
R6411 CLK1.n981 CLK1.n817 6.776
R6412 CLK1.n926 CLK1.n846 6.776
R6413 CLK1.n529 CLK1.n528 6.776
R6414 CLK1.n741 CLK1.n661 6.776
R6415 CLK1.n796 CLK1.n632 6.776
R6416 CLK1.n1004 CLK1.n516 6.776
R6417 CLK1.n1373 CLK1.n1293 6.776
R6418 CLK1.n1428 CLK1.n1264 6.776
R6419 CLK1.n1062 CLK1.n1060 6.754
R6420 CLK1.n1184 CLK1.n1183 6.754
R6421 CLK1.n141 CLK1.n3 4.938
R6422 CLK1.n47 CLK1.n7 4.938
R6423 CLK1.n251 CLK1.n213 4.938
R6424 CLK1.n1581 CLK1.n1580 4.938
R6425 CLK1.n1529 CLK1.n1494 4.938
R6426 CLK1.n1224 CLK1.n301 4.938
R6427 CLK1.n1082 CLK1.n1080 4.938
R6428 CLK1.n1082 CLK1.n1081 4.938
R6429 CLK1.n369 CLK1.n334 4.938
R6430 CLK1.n496 CLK1.n495 4.938
R6431 CLK1.n457 CLK1.n422 4.938
R6432 CLK1.n949 CLK1.n948 4.938
R6433 CLK1.n897 CLK1.n862 4.938
R6434 CLK1.n592 CLK1.n541 4.938
R6435 CLK1.n764 CLK1.n763 4.938
R6436 CLK1.n712 CLK1.n677 4.938
R6437 CLK1.n1396 CLK1.n1395 4.938
R6438 CLK1.n1344 CLK1.n1309 4.938
R6439 CLK1.n560 CLK1.n559 4.687
R6440 CLK1.n1192 CLK1.n1191 4.687
R6441 CLK1.n227 CLK1.n226 4.675
R6442 CLK1.n1507 CLK1.n1506 4.662
R6443 CLK1.n347 CLK1.n346 4.662
R6444 CLK1.n875 CLK1.n874 4.662
R6445 CLK1.n690 CLK1.n689 4.662
R6446 CLK1.n435 CLK1.n434 4.662
R6447 CLK1.n1322 CLK1.n1321 4.662
R6448 CLK1.n16 CLK1.n15 4.65
R6449 CLK1.n21 CLK1.n20 4.65
R6450 CLK1.n25 CLK1.n24 4.65
R6451 CLK1.n29 CLK1.n28 4.65
R6452 CLK1.n33 CLK1.n32 4.65
R6453 CLK1.n38 CLK1.n37 4.65
R6454 CLK1.n42 CLK1.n41 4.65
R6455 CLK1.n46 CLK1.n45 4.65
R6456 CLK1.n48 CLK1.n47 4.65
R6457 CLK1.n52 CLK1.n51 4.65
R6458 CLK1.n56 CLK1.n55 4.65
R6459 CLK1.n60 CLK1.n59 4.65
R6460 CLK1.n65 CLK1.n64 4.65
R6461 CLK1.n69 CLK1.n68 4.65
R6462 CLK1.n73 CLK1.n72 4.65
R6463 CLK1.n77 CLK1.n76 4.65
R6464 CLK1.n81 CLK1.n80 4.65
R6465 CLK1.n85 CLK1.n84 4.65
R6466 CLK1.n88 CLK1.n87 4.65
R6467 CLK1.n90 CLK1.n89 4.65
R6468 CLK1.n94 CLK1.n93 4.65
R6469 CLK1.n98 CLK1.n97 4.65
R6470 CLK1.n102 CLK1.n101 4.65
R6471 CLK1.n107 CLK1.n106 4.65
R6472 CLK1.n111 CLK1.n110 4.65
R6473 CLK1.n115 CLK1.n114 4.65
R6474 CLK1.n119 CLK1.n118 4.65
R6475 CLK1.n123 CLK1.n122 4.65
R6476 CLK1.n127 CLK1.n126 4.65
R6477 CLK1.n132 CLK1.n131 4.65
R6478 CLK1.n136 CLK1.n135 4.65
R6479 CLK1.n140 CLK1.n139 4.65
R6480 CLK1.n142 CLK1.n141 4.65
R6481 CLK1.n146 CLK1.n145 4.65
R6482 CLK1.n150 CLK1.n149 4.65
R6483 CLK1.n154 CLK1.n153 4.65
R6484 CLK1.n159 CLK1.n158 4.65
R6485 CLK1.n163 CLK1.n162 4.65
R6486 CLK1.n167 CLK1.n166 4.65
R6487 CLK1.n171 CLK1.n170 4.65
R6488 CLK1.n175 CLK1.n174 4.65
R6489 CLK1.n179 CLK1.n178 4.65
R6490 CLK1.n184 CLK1.n183 4.65
R6491 CLK1.n188 CLK1.n187 4.65
R6492 CLK1.n192 CLK1.n191 4.65
R6493 CLK1.n194 CLK1.n193 4.65
R6494 CLK1.n228 CLK1.n225 4.65
R6495 CLK1.n230 CLK1.n229 4.65
R6496 CLK1.n221 CLK1.n220 4.65
R6497 CLK1.n237 CLK1.n236 4.65
R6498 CLK1.n238 CLK1.n219 4.65
R6499 CLK1.n241 CLK1.n240 4.65
R6500 CLK1.n215 CLK1.n214 4.65
R6501 CLK1.n249 CLK1.n248 4.65
R6502 CLK1.n250 CLK1.n212 4.65
R6503 CLK1.n252 CLK1.n251 4.65
R6504 CLK1.n209 CLK1.n208 4.65
R6505 CLK1.n259 CLK1.n258 4.65
R6506 CLK1.n260 CLK1.n207 4.65
R6507 CLK1.n263 CLK1.n262 4.65
R6508 CLK1.n203 CLK1.n202 4.65
R6509 CLK1.n270 CLK1.n269 4.65
R6510 CLK1.n271 CLK1.n200 4.65
R6511 CLK1.n274 CLK1.n273 4.65
R6512 CLK1.n196 CLK1.n195 4.65
R6513 CLK1.n279 CLK1.n278 4.65
R6514 CLK1.n1508 CLK1.n1505 4.65
R6515 CLK1.n1510 CLK1.n1509 4.65
R6516 CLK1.n1501 CLK1.n1500 4.65
R6517 CLK1.n1518 CLK1.n1517 4.65
R6518 CLK1.n1520 CLK1.n1499 4.65
R6519 CLK1.n1522 CLK1.n1521 4.65
R6520 CLK1.n1496 CLK1.n1495 4.65
R6521 CLK1.n1529 CLK1.n1528 4.65
R6522 CLK1.n1530 CLK1.n1493 4.65
R6523 CLK1.n1533 CLK1.n1532 4.65
R6524 CLK1.n1531 CLK1.n1489 4.65
R6525 CLK1.n1540 CLK1.n1539 4.65
R6526 CLK1.n1541 CLK1.n1487 4.65
R6527 CLK1.n1544 CLK1.n1543 4.65
R6528 CLK1.n1542 CLK1.n1483 4.65
R6529 CLK1.n1549 CLK1.n1548 4.65
R6530 CLK1.n1551 CLK1.n1550 4.65
R6531 CLK1.n1480 CLK1.n1479 4.65
R6532 CLK1.n1556 CLK1.n1555 4.65
R6533 CLK1.n1557 CLK1.n1477 4.65
R6534 CLK1.n1560 CLK1.n1559 4.65
R6535 CLK1.n1473 CLK1.n1472 4.65
R6536 CLK1.n1567 CLK1.n1566 4.65
R6537 CLK1.n1568 CLK1.n1471 4.65
R6538 CLK1.n1571 CLK1.n1570 4.65
R6539 CLK1.n1569 CLK1.n1467 4.65
R6540 CLK1.n1578 CLK1.n1577 4.65
R6541 CLK1.n1579 CLK1.n1465 4.65
R6542 CLK1.n1583 CLK1.n1582 4.65
R6543 CLK1.n1581 CLK1.n1461 4.65
R6544 CLK1.n1591 CLK1.n1590 4.65
R6545 CLK1.n1592 CLK1.n1460 4.65
R6546 CLK1.n1595 CLK1.n1594 4.65
R6547 CLK1.n1457 CLK1.n1456 4.65
R6548 CLK1.n1602 CLK1.n1601 4.65
R6549 CLK1.n1603 CLK1.n1455 4.65
R6550 CLK1.n1605 CLK1.n1604 4.65
R6551 CLK1.n1451 CLK1.n1450 4.65
R6552 CLK1.n1612 CLK1.n1611 4.65
R6553 CLK1.n1614 CLK1.n1447 4.65
R6554 CLK1.n1617 CLK1.n1616 4.65
R6555 CLK1.n1615 CLK1.n1448 4.65
R6556 CLK1.n389 CLK1.n388 4.65
R6557 CLK1.n348 CLK1.n345 4.65
R6558 CLK1.n350 CLK1.n349 4.65
R6559 CLK1.n341 CLK1.n340 4.65
R6560 CLK1.n358 CLK1.n357 4.65
R6561 CLK1.n360 CLK1.n339 4.65
R6562 CLK1.n362 CLK1.n361 4.65
R6563 CLK1.n336 CLK1.n335 4.65
R6564 CLK1.n369 CLK1.n368 4.65
R6565 CLK1.n370 CLK1.n333 4.65
R6566 CLK1.n373 CLK1.n372 4.65
R6567 CLK1.n371 CLK1.n329 4.65
R6568 CLK1.n380 CLK1.n379 4.65
R6569 CLK1.n381 CLK1.n327 4.65
R6570 CLK1.n384 CLK1.n383 4.65
R6571 CLK1.n382 CLK1.n323 4.65
R6572 CLK1.n876 CLK1.n873 4.65
R6573 CLK1.n878 CLK1.n877 4.65
R6574 CLK1.n869 CLK1.n868 4.65
R6575 CLK1.n886 CLK1.n885 4.65
R6576 CLK1.n888 CLK1.n867 4.65
R6577 CLK1.n890 CLK1.n889 4.65
R6578 CLK1.n864 CLK1.n863 4.65
R6579 CLK1.n897 CLK1.n896 4.65
R6580 CLK1.n898 CLK1.n861 4.65
R6581 CLK1.n901 CLK1.n900 4.65
R6582 CLK1.n899 CLK1.n857 4.65
R6583 CLK1.n908 CLK1.n907 4.65
R6584 CLK1.n909 CLK1.n855 4.65
R6585 CLK1.n912 CLK1.n911 4.65
R6586 CLK1.n910 CLK1.n851 4.65
R6587 CLK1.n917 CLK1.n916 4.65
R6588 CLK1.n919 CLK1.n918 4.65
R6589 CLK1.n848 CLK1.n847 4.65
R6590 CLK1.n924 CLK1.n923 4.65
R6591 CLK1.n925 CLK1.n845 4.65
R6592 CLK1.n928 CLK1.n927 4.65
R6593 CLK1.n841 CLK1.n840 4.65
R6594 CLK1.n935 CLK1.n934 4.65
R6595 CLK1.n936 CLK1.n839 4.65
R6596 CLK1.n939 CLK1.n938 4.65
R6597 CLK1.n937 CLK1.n835 4.65
R6598 CLK1.n946 CLK1.n945 4.65
R6599 CLK1.n947 CLK1.n833 4.65
R6600 CLK1.n951 CLK1.n950 4.65
R6601 CLK1.n949 CLK1.n829 4.65
R6602 CLK1.n959 CLK1.n958 4.65
R6603 CLK1.n960 CLK1.n828 4.65
R6604 CLK1.n963 CLK1.n962 4.65
R6605 CLK1.n825 CLK1.n824 4.65
R6606 CLK1.n970 CLK1.n969 4.65
R6607 CLK1.n971 CLK1.n823 4.65
R6608 CLK1.n973 CLK1.n972 4.65
R6609 CLK1.n819 CLK1.n818 4.65
R6610 CLK1.n980 CLK1.n979 4.65
R6611 CLK1.n982 CLK1.n815 4.65
R6612 CLK1.n985 CLK1.n984 4.65
R6613 CLK1.n983 CLK1.n816 4.65
R6614 CLK1.n561 CLK1.n558 4.65
R6615 CLK1.n563 CLK1.n562 4.65
R6616 CLK1.n554 CLK1.n553 4.65
R6617 CLK1.n570 CLK1.n569 4.65
R6618 CLK1.n571 CLK1.n552 4.65
R6619 CLK1.n573 CLK1.n572 4.65
R6620 CLK1.n548 CLK1.n547 4.65
R6621 CLK1.n581 CLK1.n580 4.65
R6622 CLK1.n583 CLK1.n546 4.65
R6623 CLK1.n585 CLK1.n584 4.65
R6624 CLK1.n543 CLK1.n542 4.65
R6625 CLK1.n592 CLK1.n591 4.65
R6626 CLK1.n593 CLK1.n540 4.65
R6627 CLK1.n596 CLK1.n595 4.65
R6628 CLK1.n594 CLK1.n536 4.65
R6629 CLK1.n603 CLK1.n602 4.65
R6630 CLK1.n604 CLK1.n534 4.65
R6631 CLK1.n607 CLK1.n606 4.65
R6632 CLK1.n605 CLK1.n530 4.65
R6633 CLK1.n614 CLK1.n613 4.65
R6634 CLK1.n615 CLK1.n527 4.65
R6635 CLK1.n618 CLK1.n617 4.65
R6636 CLK1.n616 CLK1.n523 4.65
R6637 CLK1.n623 CLK1.n622 4.65
R6638 CLK1.n691 CLK1.n688 4.65
R6639 CLK1.n693 CLK1.n692 4.65
R6640 CLK1.n684 CLK1.n683 4.65
R6641 CLK1.n701 CLK1.n700 4.65
R6642 CLK1.n703 CLK1.n682 4.65
R6643 CLK1.n705 CLK1.n704 4.65
R6644 CLK1.n679 CLK1.n678 4.65
R6645 CLK1.n712 CLK1.n711 4.65
R6646 CLK1.n713 CLK1.n676 4.65
R6647 CLK1.n716 CLK1.n715 4.65
R6648 CLK1.n714 CLK1.n672 4.65
R6649 CLK1.n723 CLK1.n722 4.65
R6650 CLK1.n724 CLK1.n670 4.65
R6651 CLK1.n727 CLK1.n726 4.65
R6652 CLK1.n725 CLK1.n666 4.65
R6653 CLK1.n732 CLK1.n731 4.65
R6654 CLK1.n734 CLK1.n733 4.65
R6655 CLK1.n663 CLK1.n662 4.65
R6656 CLK1.n739 CLK1.n738 4.65
R6657 CLK1.n740 CLK1.n660 4.65
R6658 CLK1.n743 CLK1.n742 4.65
R6659 CLK1.n656 CLK1.n655 4.65
R6660 CLK1.n750 CLK1.n749 4.65
R6661 CLK1.n751 CLK1.n654 4.65
R6662 CLK1.n754 CLK1.n753 4.65
R6663 CLK1.n752 CLK1.n650 4.65
R6664 CLK1.n761 CLK1.n760 4.65
R6665 CLK1.n762 CLK1.n648 4.65
R6666 CLK1.n766 CLK1.n765 4.65
R6667 CLK1.n764 CLK1.n644 4.65
R6668 CLK1.n774 CLK1.n773 4.65
R6669 CLK1.n775 CLK1.n643 4.65
R6670 CLK1.n778 CLK1.n777 4.65
R6671 CLK1.n640 CLK1.n639 4.65
R6672 CLK1.n785 CLK1.n784 4.65
R6673 CLK1.n786 CLK1.n638 4.65
R6674 CLK1.n788 CLK1.n787 4.65
R6675 CLK1.n634 CLK1.n633 4.65
R6676 CLK1.n795 CLK1.n794 4.65
R6677 CLK1.n797 CLK1.n630 4.65
R6678 CLK1.n800 CLK1.n799 4.65
R6679 CLK1.n798 CLK1.n631 4.65
R6680 CLK1.n518 CLK1.n517 4.65
R6681 CLK1.n477 CLK1.n476 4.65
R6682 CLK1.n436 CLK1.n433 4.65
R6683 CLK1.n438 CLK1.n437 4.65
R6684 CLK1.n429 CLK1.n428 4.65
R6685 CLK1.n446 CLK1.n445 4.65
R6686 CLK1.n448 CLK1.n427 4.65
R6687 CLK1.n450 CLK1.n449 4.65
R6688 CLK1.n424 CLK1.n423 4.65
R6689 CLK1.n457 CLK1.n456 4.65
R6690 CLK1.n458 CLK1.n421 4.65
R6691 CLK1.n461 CLK1.n460 4.65
R6692 CLK1.n459 CLK1.n417 4.65
R6693 CLK1.n468 CLK1.n467 4.65
R6694 CLK1.n469 CLK1.n415 4.65
R6695 CLK1.n472 CLK1.n471 4.65
R6696 CLK1.n470 CLK1.n411 4.65
R6697 CLK1.n479 CLK1.n478 4.65
R6698 CLK1.n480 CLK1.n409 4.65
R6699 CLK1.n482 CLK1.n481 4.65
R6700 CLK1.n403 CLK1.n401 4.65
R6701 CLK1.n1053 CLK1.n1052 4.65
R6702 CLK1.n404 CLK1.n402 4.65
R6703 CLK1.n1046 CLK1.n1045 4.65
R6704 CLK1.n1044 CLK1.n488 4.65
R6705 CLK1.n1043 CLK1.n1042 4.65
R6706 CLK1.n490 CLK1.n489 4.65
R6707 CLK1.n1036 CLK1.n1035 4.65
R6708 CLK1.n1034 CLK1.n493 4.65
R6709 CLK1.n1033 CLK1.n1032 4.65
R6710 CLK1.n497 CLK1.n496 4.65
R6711 CLK1.n1026 CLK1.n1025 4.65
R6712 CLK1.n1024 CLK1.n502 4.65
R6713 CLK1.n1023 CLK1.n1022 4.65
R6714 CLK1.n509 CLK1.n504 4.65
R6715 CLK1.n1016 CLK1.n1015 4.65
R6716 CLK1.n1014 CLK1.n508 4.65
R6717 CLK1.n1013 CLK1.n1012 4.65
R6718 CLK1.n511 CLK1.n510 4.65
R6719 CLK1.n1006 CLK1.n1005 4.65
R6720 CLK1.n1003 CLK1.n515 4.65
R6721 CLK1.n1002 CLK1.n1001 4.65
R6722 CLK1.n400 CLK1.n399 4.65
R6723 CLK1.n1065 CLK1.n398 4.65
R6724 CLK1.n1064 CLK1.n1063 4.65
R6725 CLK1.n321 CLK1.n320 4.65
R6726 CLK1.n1181 CLK1.n1180 4.65
R6727 CLK1.n1189 CLK1.n1188 4.65
R6728 CLK1.n1193 CLK1.n318 4.65
R6729 CLK1.n1195 CLK1.n1194 4.65
R6730 CLK1.n314 CLK1.n313 4.65
R6731 CLK1.n1202 CLK1.n1201 4.65
R6732 CLK1.n1203 CLK1.n312 4.65
R6733 CLK1.n1205 CLK1.n1204 4.65
R6734 CLK1.n308 CLK1.n307 4.65
R6735 CLK1.n1213 CLK1.n1212 4.65
R6736 CLK1.n1215 CLK1.n306 4.65
R6737 CLK1.n1217 CLK1.n1216 4.65
R6738 CLK1.n303 CLK1.n302 4.65
R6739 CLK1.n1224 CLK1.n1223 4.65
R6740 CLK1.n1225 CLK1.n300 4.65
R6741 CLK1.n1228 CLK1.n1227 4.65
R6742 CLK1.n1226 CLK1.n296 4.65
R6743 CLK1.n1235 CLK1.n1234 4.65
R6744 CLK1.n1236 CLK1.n294 4.65
R6745 CLK1.n1239 CLK1.n1238 4.65
R6746 CLK1.n1237 CLK1.n290 4.65
R6747 CLK1.n1246 CLK1.n1245 4.65
R6748 CLK1.n1247 CLK1.n287 4.65
R6749 CLK1.n1250 CLK1.n1249 4.65
R6750 CLK1.n1248 CLK1.n283 4.65
R6751 CLK1.n1255 CLK1.n1254 4.65
R6752 CLK1.n1323 CLK1.n1320 4.65
R6753 CLK1.n1325 CLK1.n1324 4.65
R6754 CLK1.n1316 CLK1.n1315 4.65
R6755 CLK1.n1333 CLK1.n1332 4.65
R6756 CLK1.n1335 CLK1.n1314 4.65
R6757 CLK1.n1337 CLK1.n1336 4.65
R6758 CLK1.n1311 CLK1.n1310 4.65
R6759 CLK1.n1344 CLK1.n1343 4.65
R6760 CLK1.n1345 CLK1.n1308 4.65
R6761 CLK1.n1348 CLK1.n1347 4.65
R6762 CLK1.n1346 CLK1.n1304 4.65
R6763 CLK1.n1355 CLK1.n1354 4.65
R6764 CLK1.n1356 CLK1.n1302 4.65
R6765 CLK1.n1359 CLK1.n1358 4.65
R6766 CLK1.n1357 CLK1.n1298 4.65
R6767 CLK1.n1364 CLK1.n1363 4.65
R6768 CLK1.n1366 CLK1.n1365 4.65
R6769 CLK1.n1295 CLK1.n1294 4.65
R6770 CLK1.n1371 CLK1.n1370 4.65
R6771 CLK1.n1372 CLK1.n1292 4.65
R6772 CLK1.n1375 CLK1.n1374 4.65
R6773 CLK1.n1288 CLK1.n1287 4.65
R6774 CLK1.n1382 CLK1.n1381 4.65
R6775 CLK1.n1383 CLK1.n1286 4.65
R6776 CLK1.n1386 CLK1.n1385 4.65
R6777 CLK1.n1384 CLK1.n1282 4.65
R6778 CLK1.n1393 CLK1.n1392 4.65
R6779 CLK1.n1394 CLK1.n1280 4.65
R6780 CLK1.n1398 CLK1.n1397 4.65
R6781 CLK1.n1396 CLK1.n1276 4.65
R6782 CLK1.n1406 CLK1.n1405 4.65
R6783 CLK1.n1407 CLK1.n1275 4.65
R6784 CLK1.n1410 CLK1.n1409 4.65
R6785 CLK1.n1272 CLK1.n1271 4.65
R6786 CLK1.n1417 CLK1.n1416 4.65
R6787 CLK1.n1418 CLK1.n1270 4.65
R6788 CLK1.n1420 CLK1.n1419 4.65
R6789 CLK1.n1266 CLK1.n1265 4.65
R6790 CLK1.n1427 CLK1.n1426 4.65
R6791 CLK1.n1429 CLK1.n1262 4.65
R6792 CLK1.n1432 CLK1.n1431 4.65
R6793 CLK1.n1430 CLK1.n1263 4.65
R6794 CLK1.n1177 CLK1.n392 4.633
R6795 CLK1.n1177 CLK1.n393 4.633
R6796 CLK1.n1171 CLK1.n393 4.633
R6797 CLK1.n1171 CLK1.n397 4.633
R6798 CLK1.n1166 CLK1.n397 4.633
R6799 CLK1.n1166 CLK1.n1067 4.633
R6800 CLK1.n1160 CLK1.n1067 4.633
R6801 CLK1.n1160 CLK1.n1071 4.633
R6802 CLK1.n1156 CLK1.n1071 4.633
R6803 CLK1.n1156 CLK1.n1073 4.633
R6804 CLK1.n1152 CLK1.n1073 4.633
R6805 CLK1.n1152 CLK1.n1078 4.633
R6806 CLK1.n1148 CLK1.n1078 4.633
R6807 CLK1.n1148 CLK1.n1083 4.633
R6808 CLK1.n1144 CLK1.n1083 4.633
R6809 CLK1.n1144 CLK1.n1089 4.633
R6810 CLK1.n1140 CLK1.n1089 4.633
R6811 CLK1.n1140 CLK1.n1091 4.633
R6812 CLK1.n1136 CLK1.n1091 4.633
R6813 CLK1.n1136 CLK1.n1097 4.633
R6814 CLK1.n1132 CLK1.n1097 4.633
R6815 CLK1.n1132 CLK1.n1101 4.633
R6816 CLK1.n1126 CLK1.n1101 4.633
R6817 CLK1.n1126 CLK1.n1106 4.633
R6818 CLK1.n1121 CLK1.n1106 4.633
R6819 CLK1.n1121 CLK1.n1111 4.633
R6820 CLK1.n1115 CLK1.n1111 4.633
R6821 CLK1.n996 CLK1.n994 4.527
R6822 CLK1.n807 CLK1.n624 4.5
R6823 CLK1.n992 CLK1.n809 4.5
R6824 CLK1.n1439 CLK1.n1256 4.5
R6825 CLK1.n1624 CLK1.n1441 4.5
R6826 CLK1.n1177 CLK1.n1176 4.427
R6827 CLK1.n394 CLK1.n393 4.427
R6828 CLK1.n1174 CLK1.n394 4.427
R6829 CLK1.n1172 CLK1.n1171 4.427
R6830 CLK1.n1173 CLK1.n1172 4.427
R6831 CLK1.n397 CLK1.n396 4.427
R6832 CLK1.n396 CLK1.n395 4.427
R6833 CLK1.n1166 CLK1.n1165 4.427
R6834 CLK1.n1165 CLK1.n1164 4.427
R6835 CLK1.n1068 CLK1.n1067 4.427
R6836 CLK1.n1163 CLK1.n1068 4.427
R6837 CLK1.n1161 CLK1.n1160 4.427
R6838 CLK1.n1162 CLK1.n1161 4.427
R6839 CLK1.n1071 CLK1.n1070 4.427
R6840 CLK1.n1070 CLK1.n1069 4.427
R6841 CLK1.n1156 CLK1.n1155 4.427
R6842 CLK1.n1154 CLK1.n1073 4.427
R6843 CLK1.n1153 CLK1.n1152 4.427
R6844 CLK1.n1078 CLK1.n1077 4.427
R6845 CLK1.n1148 CLK1.n1147 4.427
R6846 CLK1.n1146 CLK1.n1083 4.427
R6847 CLK1.n1145 CLK1.n1144 4.427
R6848 CLK1.n1089 CLK1.n1088 4.427
R6849 CLK1.n1140 CLK1.n1139 4.427
R6850 CLK1.n1138 CLK1.n1091 4.427
R6851 CLK1.n1137 CLK1.n1136 4.427
R6852 CLK1.n1097 CLK1.n1096 4.427
R6853 CLK1.n1103 CLK1.n1096 4.427
R6854 CLK1.n1132 CLK1.n1131 4.427
R6855 CLK1.n1131 CLK1.n1130 4.427
R6856 CLK1.n1102 CLK1.n1101 4.427
R6857 CLK1.n1129 CLK1.n1102 4.427
R6858 CLK1.n1127 CLK1.n1126 4.427
R6859 CLK1.n1128 CLK1.n1127 4.427
R6860 CLK1.n1106 CLK1.n1105 4.427
R6861 CLK1.n1105 CLK1.n1104 4.427
R6862 CLK1.n1121 CLK1.n1120 4.427
R6863 CLK1.n1120 CLK1.n1119 4.427
R6864 CLK1.n1112 CLK1.n1111 4.427
R6865 CLK1.n1118 CLK1.n1112 4.427
R6866 CLK1.n1116 CLK1.n1115 4.427
R6867 CLK1.n1155 CLK1.n1074 4.427
R6868 CLK1.n1154 CLK1.n1075 4.427
R6869 CLK1.n1153 CLK1.n1076 4.427
R6870 CLK1.n1084 CLK1.n1077 4.427
R6871 CLK1.n1147 CLK1.n1085 4.427
R6872 CLK1.n1146 CLK1.n1086 4.427
R6873 CLK1.n1145 CLK1.n1087 4.427
R6874 CLK1.n1092 CLK1.n1088 4.427
R6875 CLK1.n1139 CLK1.n1093 4.427
R6876 CLK1.n1138 CLK1.n1094 4.427
R6877 CLK1.n1137 CLK1.n1095 4.427
R6878 CLK1.t86 CLK1.n1085 4.314
R6879 CLK1.n1087 CLK1.t98 4.314
R6880 CLK1.n1183 CLK1.n321 3.715
R6881 CLK1.n1056 CLK1.n400 3.715
R6882 CLK1.n1063 CLK1.n1062 3.715
R6883 CLK1.n1188 CLK1.n319 3.715
R6884 CLK1.n809 CLK1.n808 3.635
R6885 CLK1.n1441 CLK1.n1440 3.635
R6886 CLK1.n1185 CLK1.n1184 3.635
R6887 CLK1 CLK1.n1626 3.578
R6888 CLK1.n1622 CLK1.n1621 3.563
R6889 CLK1.n990 CLK1.n989 3.563
R6890 CLK1.n805 CLK1.n804 3.563
R6891 CLK1.n1437 CLK1.n1436 3.563
R6892 CLK1.n1180 CLK1.n1179 3.203
R6893 CLK1.n624 CLK1.n623 3.067
R6894 CLK1.n1256 CLK1.n1255 3.067
R6895 CLK1.n1059 CLK1.n1058 3.039
R6896 CLK1.n1187 CLK1.n1185 3.038
R6897 CLK1.n997 CLK1.n996 3.033
R6898 CLK1.n1060 CLK1.n1059 2.849
R6899 CLK1.n12 CLK1.n11 2.682
R6900 CLK1.n1626 CLK1.n279 2.625
R6901 CLK1.n1183 CLK1.n1182 2.57
R6902 CLK1.n1057 CLK1.n1056 2.57
R6903 CLK1.n1062 CLK1.n1061 2.57
R6904 CLK1.n1186 CLK1.n319 2.57
R6905 EESPFAL_s0_0/CLK1 CLK1.n194 2.35
R6906 CLK1.n1178 CLK1.n1177 2.325
R6907 CLK1.n393 CLK1.n391 2.325
R6908 CLK1.n1171 CLK1.n1170 2.325
R6909 CLK1.n1169 CLK1.n397 2.325
R6910 CLK1.n1167 CLK1.n1166 2.325
R6911 CLK1.n1067 CLK1.n1066 2.325
R6912 CLK1.n1160 CLK1.n1159 2.325
R6913 CLK1.n1158 CLK1.n1071 2.325
R6914 CLK1.n1157 CLK1.n1156 2.325
R6915 CLK1.n1073 CLK1.n1072 2.325
R6916 CLK1.n1152 CLK1.n1151 2.325
R6917 CLK1.n1150 CLK1.n1078 2.325
R6918 CLK1.n1149 CLK1.n1148 2.325
R6919 CLK1.n1083 CLK1.n1082 2.325
R6920 CLK1.n1144 CLK1.n1143 2.325
R6921 CLK1.n1142 CLK1.n1089 2.325
R6922 CLK1.n1141 CLK1.n1140 2.325
R6923 CLK1.n1098 CLK1.n1091 2.325
R6924 CLK1.n1136 CLK1.n1135 2.325
R6925 CLK1.n1134 CLK1.n1097 2.325
R6926 CLK1.n1133 CLK1.n1132 2.325
R6927 CLK1.n1107 CLK1.n1101 2.325
R6928 CLK1.n1126 CLK1.n1125 2.325
R6929 CLK1.n1123 CLK1.n1106 2.325
R6930 CLK1.n1122 CLK1.n1121 2.325
R6931 CLK1.n1113 CLK1.n1111 2.325
R6932 CLK1.n392 CLK1.n390 2.325
R6933 CLK1.n993 CLK1.n992 2.246
R6934 CLK1.n1625 CLK1.n1624 2.246
R6935 CLK1.n991 CLK1.n520 2.246
R6936 CLK1.n1623 CLK1.n280 2.246
R6937 CLK1.n808 CLK1.n807 2.245
R6938 CLK1.n1440 CLK1.n1439 2.245
R6939 CLK1.n806 CLK1.n521 2.245
R6940 CLK1.n1438 CLK1.n281 2.245
R6941 CLK1.n1055 CLK1.n1054 2.203
R6942 CLK1.n1168 CLK1.n1065 2.203
R6943 CLK1.n1192 CLK1.n1190 2.203
R6944 CLK1.n10 CLK1.n9 1.655
R6945 CLK1.n92 CLK1.n91 1.655
R6946 CLK1.n224 CLK1.n223 1.655
R6947 CLK1.n1504 CLK1.n1503 1.655
R6948 CLK1.n1552 CLK1.n1481 1.655
R6949 CLK1.n872 CLK1.n871 1.655
R6950 CLK1.n920 CLK1.n849 1.655
R6951 CLK1.n557 CLK1.n556 1.655
R6952 CLK1.n687 CLK1.n686 1.655
R6953 CLK1.n735 CLK1.n664 1.655
R6954 CLK1.n408 CLK1.n407 1.655
R6955 CLK1.n317 CLK1.n316 1.655
R6956 CLK1.n1319 CLK1.n1318 1.655
R6957 CLK1.n1367 CLK1.n1296 1.655
R6958 CLK1.n83 CLK1.n82 1.655
R6959 CLK1.n190 CLK1.n189 1.655
R6960 CLK1.n277 CLK1.n197 1.655
R6961 CLK1.n1547 CLK1.n1484 1.655
R6962 CLK1.n1620 CLK1.n1444 1.655
R6963 CLK1.n344 CLK1.n343 1.655
R6964 CLK1.n387 CLK1.n324 1.655
R6965 CLK1.n432 CLK1.n431 1.655
R6966 CLK1.n915 CLK1.n852 1.655
R6967 CLK1.n988 CLK1.n812 1.655
R6968 CLK1.n621 CLK1.n524 1.655
R6969 CLK1.n730 CLK1.n667 1.655
R6970 CLK1.n803 CLK1.n627 1.655
R6971 CLK1.n475 CLK1.n412 1.655
R6972 CLK1.n998 CLK1.n519 1.655
R6973 CLK1.n1253 CLK1.n284 1.655
R6974 CLK1.n1362 CLK1.n1299 1.655
R6975 CLK1.n1435 CLK1.n1259 1.655
R6976 CLK1.n1621 CLK1.n1443 1.44
R6977 CLK1.n989 CLK1.n811 1.44
R6978 CLK1.n804 CLK1.n626 1.44
R6979 CLK1.n1436 CLK1.n1258 1.44
R6980 CLK1.n1115 CLK1.n1114 1.156
R6981 CLK1.n16 CLK1.n12 1.096
R6982 CLK1.n995 EESPFAL_s2_0/CLK1 0.912
R6983 CLK1.n994 CLK1.n993 0.705
R6984 CLK1.n1626 CLK1.n1625 0.7
R6985 CLK1.n479 CLK1.n477 0.662
R6986 CLK1.n1550 CLK1.n1549 0.637
R6987 CLK1.n918 CLK1.n917 0.637
R6988 CLK1.n733 CLK1.n732 0.637
R6989 CLK1.n1365 CLK1.n1364 0.637
R6990 CLK1.n1114 CLK1.n1113 0.631
R6991 CLK1.n1176 CLK1.n1175 0.619
R6992 CLK1.n1117 CLK1.n1116 0.618
R6993 CLK1.n90 CLK1.n88 0.6
R6994 CLK1.n390 CLK1.n389 0.532
R6995 CLK1.n1055 CLK1.n399 0.125
R6996 CLK1.n1065 CLK1.n1064 0.125
R6997 CLK1.n1180 CLK1.n320 0.125
R6998 CLK1.n1190 CLK1.n1189 0.125
R6999 CLK1.n1064 CLK1.n1060 0.12
R7000 CLK1.n1189 CLK1.n1185 0.119
R7001 CLK1.n1059 CLK1.n399 0.119
R7002 CLK1.n1184 CLK1.n320 0.119
R7003 CLK1.n25 CLK1.n21 0.1
R7004 CLK1.n29 CLK1.n25 0.1
R7005 CLK1.n33 CLK1.n29 0.1
R7006 CLK1.n42 CLK1.n38 0.1
R7007 CLK1.n46 CLK1.n42 0.1
R7008 CLK1.n47 CLK1.n46 0.1
R7009 CLK1.n56 CLK1.n52 0.1
R7010 CLK1.n60 CLK1.n56 0.1
R7011 CLK1.n69 CLK1.n65 0.1
R7012 CLK1.n73 CLK1.n69 0.1
R7013 CLK1.n77 CLK1.n73 0.1
R7014 CLK1.n81 CLK1.n77 0.1
R7015 CLK1.n85 CLK1.n81 0.1
R7016 CLK1.n94 CLK1.n90 0.1
R7017 CLK1.n98 CLK1.n94 0.1
R7018 CLK1.n102 CLK1.n98 0.1
R7019 CLK1.n111 CLK1.n107 0.1
R7020 CLK1.n115 CLK1.n111 0.1
R7021 CLK1.n119 CLK1.n115 0.1
R7022 CLK1.n123 CLK1.n119 0.1
R7023 CLK1.n127 CLK1.n123 0.1
R7024 CLK1.n136 CLK1.n132 0.1
R7025 CLK1.n140 CLK1.n136 0.1
R7026 CLK1.n141 CLK1.n140 0.1
R7027 CLK1.n150 CLK1.n146 0.1
R7028 CLK1.n154 CLK1.n150 0.1
R7029 CLK1.n163 CLK1.n159 0.1
R7030 CLK1.n167 CLK1.n163 0.1
R7031 CLK1.n171 CLK1.n167 0.1
R7032 CLK1.n175 CLK1.n171 0.1
R7033 CLK1.n179 CLK1.n175 0.1
R7034 CLK1.n188 CLK1.n184 0.1
R7035 CLK1.n192 CLK1.n188 0.1
R7036 CLK1.n194 CLK1.n192 0.1
R7037 CLK1.n229 CLK1.n228 0.1
R7038 CLK1.n229 CLK1.n220 0.1
R7039 CLK1.n237 CLK1.n220 0.1
R7040 CLK1.n238 CLK1.n237 0.1
R7041 CLK1.n240 CLK1.n238 0.1
R7042 CLK1.n249 CLK1.n214 0.1
R7043 CLK1.n250 CLK1.n249 0.1
R7044 CLK1.n251 CLK1.n250 0.1
R7045 CLK1.n259 CLK1.n208 0.1
R7046 CLK1.n260 CLK1.n259 0.1
R7047 CLK1.n262 CLK1.n202 0.1
R7048 CLK1.n270 CLK1.n202 0.1
R7049 CLK1.n271 CLK1.n270 0.1
R7050 CLK1.n273 CLK1.n195 0.1
R7051 CLK1.n279 CLK1.n195 0.1
R7052 CLK1.n1509 CLK1.n1508 0.1
R7053 CLK1.n1509 CLK1.n1500 0.1
R7054 CLK1.n1518 CLK1.n1500 0.1
R7055 CLK1.n1521 CLK1.n1520 0.1
R7056 CLK1.n1521 CLK1.n1495 0.1
R7057 CLK1.n1529 CLK1.n1495 0.1
R7058 CLK1.n1532 CLK1.n1530 0.1
R7059 CLK1.n1532 CLK1.n1531 0.1
R7060 CLK1.n1541 CLK1.n1540 0.1
R7061 CLK1.n1543 CLK1.n1541 0.1
R7062 CLK1.n1543 CLK1.n1542 0.1
R7063 CLK1.n1550 CLK1.n1479 0.1
R7064 CLK1.n1556 CLK1.n1479 0.1
R7065 CLK1.n1557 CLK1.n1556 0.1
R7066 CLK1.n1559 CLK1.n1472 0.1
R7067 CLK1.n1567 CLK1.n1472 0.1
R7068 CLK1.n1568 CLK1.n1567 0.1
R7069 CLK1.n1570 CLK1.n1568 0.1
R7070 CLK1.n1570 CLK1.n1569 0.1
R7071 CLK1.n1579 CLK1.n1578 0.1
R7072 CLK1.n1582 CLK1.n1579 0.1
R7073 CLK1.n1582 CLK1.n1581 0.1
R7074 CLK1.n1592 CLK1.n1591 0.1
R7075 CLK1.n1594 CLK1.n1592 0.1
R7076 CLK1.n1602 CLK1.n1456 0.1
R7077 CLK1.n1603 CLK1.n1602 0.1
R7078 CLK1.n1604 CLK1.n1603 0.1
R7079 CLK1.n1604 CLK1.n1450 0.1
R7080 CLK1.n1612 CLK1.n1450 0.1
R7081 CLK1.n1616 CLK1.n1614 0.1
R7082 CLK1.n1616 CLK1.n1615 0.1
R7083 CLK1.n349 CLK1.n348 0.1
R7084 CLK1.n349 CLK1.n340 0.1
R7085 CLK1.n358 CLK1.n340 0.1
R7086 CLK1.n361 CLK1.n360 0.1
R7087 CLK1.n361 CLK1.n335 0.1
R7088 CLK1.n369 CLK1.n335 0.1
R7089 CLK1.n372 CLK1.n370 0.1
R7090 CLK1.n372 CLK1.n371 0.1
R7091 CLK1.n381 CLK1.n380 0.1
R7092 CLK1.n383 CLK1.n381 0.1
R7093 CLK1.n383 CLK1.n382 0.1
R7094 CLK1.n877 CLK1.n876 0.1
R7095 CLK1.n877 CLK1.n868 0.1
R7096 CLK1.n886 CLK1.n868 0.1
R7097 CLK1.n889 CLK1.n888 0.1
R7098 CLK1.n889 CLK1.n863 0.1
R7099 CLK1.n897 CLK1.n863 0.1
R7100 CLK1.n900 CLK1.n898 0.1
R7101 CLK1.n900 CLK1.n899 0.1
R7102 CLK1.n909 CLK1.n908 0.1
R7103 CLK1.n911 CLK1.n909 0.1
R7104 CLK1.n911 CLK1.n910 0.1
R7105 CLK1.n918 CLK1.n847 0.1
R7106 CLK1.n924 CLK1.n847 0.1
R7107 CLK1.n925 CLK1.n924 0.1
R7108 CLK1.n927 CLK1.n840 0.1
R7109 CLK1.n935 CLK1.n840 0.1
R7110 CLK1.n936 CLK1.n935 0.1
R7111 CLK1.n938 CLK1.n936 0.1
R7112 CLK1.n938 CLK1.n937 0.1
R7113 CLK1.n947 CLK1.n946 0.1
R7114 CLK1.n950 CLK1.n947 0.1
R7115 CLK1.n950 CLK1.n949 0.1
R7116 CLK1.n960 CLK1.n959 0.1
R7117 CLK1.n962 CLK1.n960 0.1
R7118 CLK1.n970 CLK1.n824 0.1
R7119 CLK1.n971 CLK1.n970 0.1
R7120 CLK1.n972 CLK1.n971 0.1
R7121 CLK1.n972 CLK1.n818 0.1
R7122 CLK1.n980 CLK1.n818 0.1
R7123 CLK1.n984 CLK1.n982 0.1
R7124 CLK1.n984 CLK1.n983 0.1
R7125 CLK1.n562 CLK1.n561 0.1
R7126 CLK1.n562 CLK1.n553 0.1
R7127 CLK1.n570 CLK1.n553 0.1
R7128 CLK1.n571 CLK1.n570 0.1
R7129 CLK1.n572 CLK1.n571 0.1
R7130 CLK1.n572 CLK1.n547 0.1
R7131 CLK1.n581 CLK1.n547 0.1
R7132 CLK1.n584 CLK1.n583 0.1
R7133 CLK1.n584 CLK1.n542 0.1
R7134 CLK1.n592 CLK1.n542 0.1
R7135 CLK1.n595 CLK1.n593 0.1
R7136 CLK1.n595 CLK1.n594 0.1
R7137 CLK1.n604 CLK1.n603 0.1
R7138 CLK1.n606 CLK1.n604 0.1
R7139 CLK1.n606 CLK1.n605 0.1
R7140 CLK1.n615 CLK1.n614 0.1
R7141 CLK1.n617 CLK1.n615 0.1
R7142 CLK1.n617 CLK1.n616 0.1
R7143 CLK1.n692 CLK1.n691 0.1
R7144 CLK1.n692 CLK1.n683 0.1
R7145 CLK1.n701 CLK1.n683 0.1
R7146 CLK1.n704 CLK1.n703 0.1
R7147 CLK1.n704 CLK1.n678 0.1
R7148 CLK1.n712 CLK1.n678 0.1
R7149 CLK1.n715 CLK1.n713 0.1
R7150 CLK1.n715 CLK1.n714 0.1
R7151 CLK1.n724 CLK1.n723 0.1
R7152 CLK1.n726 CLK1.n724 0.1
R7153 CLK1.n726 CLK1.n725 0.1
R7154 CLK1.n733 CLK1.n662 0.1
R7155 CLK1.n739 CLK1.n662 0.1
R7156 CLK1.n740 CLK1.n739 0.1
R7157 CLK1.n742 CLK1.n655 0.1
R7158 CLK1.n750 CLK1.n655 0.1
R7159 CLK1.n751 CLK1.n750 0.1
R7160 CLK1.n753 CLK1.n751 0.1
R7161 CLK1.n753 CLK1.n752 0.1
R7162 CLK1.n762 CLK1.n761 0.1
R7163 CLK1.n765 CLK1.n762 0.1
R7164 CLK1.n765 CLK1.n764 0.1
R7165 CLK1.n775 CLK1.n774 0.1
R7166 CLK1.n777 CLK1.n775 0.1
R7167 CLK1.n785 CLK1.n639 0.1
R7168 CLK1.n786 CLK1.n785 0.1
R7169 CLK1.n787 CLK1.n786 0.1
R7170 CLK1.n787 CLK1.n633 0.1
R7171 CLK1.n795 CLK1.n633 0.1
R7172 CLK1.n799 CLK1.n797 0.1
R7173 CLK1.n799 CLK1.n798 0.1
R7174 CLK1.n437 CLK1.n436 0.1
R7175 CLK1.n437 CLK1.n428 0.1
R7176 CLK1.n446 CLK1.n428 0.1
R7177 CLK1.n449 CLK1.n448 0.1
R7178 CLK1.n449 CLK1.n423 0.1
R7179 CLK1.n457 CLK1.n423 0.1
R7180 CLK1.n460 CLK1.n458 0.1
R7181 CLK1.n460 CLK1.n459 0.1
R7182 CLK1.n469 CLK1.n468 0.1
R7183 CLK1.n471 CLK1.n469 0.1
R7184 CLK1.n471 CLK1.n470 0.1
R7185 CLK1.n480 CLK1.n479 0.1
R7186 CLK1.n481 CLK1.n480 0.1
R7187 CLK1.n481 CLK1.n401 0.1
R7188 CLK1.n1053 CLK1.n402 0.1
R7189 CLK1.n1045 CLK1.n402 0.1
R7190 CLK1.n1045 CLK1.n1044 0.1
R7191 CLK1.n1044 CLK1.n1043 0.1
R7192 CLK1.n1043 CLK1.n489 0.1
R7193 CLK1.n1035 CLK1.n1034 0.1
R7194 CLK1.n1034 CLK1.n1033 0.1
R7195 CLK1.n1033 CLK1.n496 0.1
R7196 CLK1.n1025 CLK1.n1024 0.1
R7197 CLK1.n1024 CLK1.n1023 0.1
R7198 CLK1.n1015 CLK1.n509 0.1
R7199 CLK1.n1015 CLK1.n1014 0.1
R7200 CLK1.n1014 CLK1.n1013 0.1
R7201 CLK1.n1013 CLK1.n510 0.1
R7202 CLK1.n1005 CLK1.n510 0.1
R7203 CLK1.n1003 CLK1.n1002 0.1
R7204 CLK1.n1002 CLK1.n517 0.1
R7205 CLK1.n1194 CLK1.n1193 0.1
R7206 CLK1.n1194 CLK1.n313 0.1
R7207 CLK1.n1202 CLK1.n313 0.1
R7208 CLK1.n1203 CLK1.n1202 0.1
R7209 CLK1.n1204 CLK1.n1203 0.1
R7210 CLK1.n1204 CLK1.n307 0.1
R7211 CLK1.n1213 CLK1.n307 0.1
R7212 CLK1.n1216 CLK1.n1215 0.1
R7213 CLK1.n1216 CLK1.n302 0.1
R7214 CLK1.n1224 CLK1.n302 0.1
R7215 CLK1.n1227 CLK1.n1225 0.1
R7216 CLK1.n1227 CLK1.n1226 0.1
R7217 CLK1.n1236 CLK1.n1235 0.1
R7218 CLK1.n1238 CLK1.n1236 0.1
R7219 CLK1.n1238 CLK1.n1237 0.1
R7220 CLK1.n1247 CLK1.n1246 0.1
R7221 CLK1.n1249 CLK1.n1247 0.1
R7222 CLK1.n1249 CLK1.n1248 0.1
R7223 CLK1.n1324 CLK1.n1323 0.1
R7224 CLK1.n1324 CLK1.n1315 0.1
R7225 CLK1.n1333 CLK1.n1315 0.1
R7226 CLK1.n1336 CLK1.n1335 0.1
R7227 CLK1.n1336 CLK1.n1310 0.1
R7228 CLK1.n1344 CLK1.n1310 0.1
R7229 CLK1.n1347 CLK1.n1345 0.1
R7230 CLK1.n1347 CLK1.n1346 0.1
R7231 CLK1.n1356 CLK1.n1355 0.1
R7232 CLK1.n1358 CLK1.n1356 0.1
R7233 CLK1.n1358 CLK1.n1357 0.1
R7234 CLK1.n1365 CLK1.n1294 0.1
R7235 CLK1.n1371 CLK1.n1294 0.1
R7236 CLK1.n1372 CLK1.n1371 0.1
R7237 CLK1.n1374 CLK1.n1287 0.1
R7238 CLK1.n1382 CLK1.n1287 0.1
R7239 CLK1.n1383 CLK1.n1382 0.1
R7240 CLK1.n1385 CLK1.n1383 0.1
R7241 CLK1.n1385 CLK1.n1384 0.1
R7242 CLK1.n1394 CLK1.n1393 0.1
R7243 CLK1.n1397 CLK1.n1394 0.1
R7244 CLK1.n1397 CLK1.n1396 0.1
R7245 CLK1.n1407 CLK1.n1406 0.1
R7246 CLK1.n1409 CLK1.n1407 0.1
R7247 CLK1.n1417 CLK1.n1271 0.1
R7248 CLK1.n1418 CLK1.n1417 0.1
R7249 CLK1.n1419 CLK1.n1418 0.1
R7250 CLK1.n1419 CLK1.n1265 0.1
R7251 CLK1.n1427 CLK1.n1265 0.1
R7252 CLK1.n1431 CLK1.n1429 0.1
R7253 CLK1.n1431 CLK1.n1430 0.1
R7254 CLK1.n995 CLK1.n517 0.094
R7255 CLK1.n1615 CLK1.n1442 0.088
R7256 CLK1.n983 CLK1.n810 0.088
R7257 CLK1.n798 CLK1.n625 0.088
R7258 CLK1.n1430 CLK1.n1257 0.088
R7259 CLK1.n21 CLK1.n17 0.087
R7260 CLK1.n272 CLK1.n271 0.087
R7261 CLK1.n1508 CLK1.n1507 0.087
R7262 CLK1.n1542 CLK1.n1482 0.087
R7263 CLK1.n348 CLK1.n347 0.087
R7264 CLK1.n382 CLK1.n322 0.087
R7265 CLK1.n876 CLK1.n875 0.087
R7266 CLK1.n910 CLK1.n850 0.087
R7267 CLK1.n605 CLK1.n529 0.087
R7268 CLK1.n691 CLK1.n690 0.087
R7269 CLK1.n725 CLK1.n665 0.087
R7270 CLK1.n436 CLK1.n435 0.087
R7271 CLK1.n470 CLK1.n410 0.087
R7272 CLK1.n1237 CLK1.n289 0.087
R7273 CLK1.n1323 CLK1.n1322 0.087
R7274 CLK1.n1357 CLK1.n1297 0.087
R7275 EESPFAL_s0_0/CLK1 CLK1 0.084
R7276 CLK1.n38 CLK1.n34 0.075
R7277 CLK1.n52 CLK1 0.075
R7278 CLK1.n61 CLK1.n60 0.075
R7279 CLK1.n86 CLK1.n85 0.075
R7280 CLK1.n107 CLK1.n103 0.075
R7281 CLK1.n132 CLK1.n128 0.075
R7282 CLK1.n146 EESPFAL_s0_0/EESPFAL_XOR_v3_0/CLK 0.075
R7283 CLK1.n155 CLK1.n154 0.075
R7284 CLK1.n180 CLK1.n179 0.075
R7285 CLK1.n228 CLK1.n227 0.075
R7286 CLK1.n239 CLK1.n214 0.075
R7287 EESPFAL_s0_0/EESPFAL_NAND_v3_2/CLK CLK1.n208 0.075
R7288 CLK1.n261 CLK1.n260 0.075
R7289 CLK1.n1520 CLK1.n1519 0.075
R7290 CLK1.n1530 EESPFAL_s1_0/EESPFAL_INV4_2/CLK 0.075
R7291 CLK1.n1531 CLK1.n1488 0.075
R7292 CLK1.n1559 CLK1.n1558 0.075
R7293 CLK1.n1578 CLK1.n1466 0.075
R7294 CLK1.n1591 EESPFAL_s1_0/EESPFAL_XOR_v3_0/CLK 0.075
R7295 CLK1.n1594 CLK1.n1593 0.075
R7296 CLK1.n1613 CLK1.n1612 0.075
R7297 CLK1.n360 CLK1.n359 0.075
R7298 CLK1.n370 EESPFAL_s2_0/EESPFAL_INV4_0/CLK 0.075
R7299 CLK1.n371 CLK1.n328 0.075
R7300 CLK1.n888 CLK1.n887 0.075
R7301 CLK1.n898 EESPFAL_s3_0/EESPFAL_INV4_2/CLK 0.075
R7302 CLK1.n899 CLK1.n856 0.075
R7303 CLK1.n927 CLK1.n926 0.075
R7304 CLK1.n946 CLK1.n834 0.075
R7305 CLK1.n959 EESPFAL_s3_0/EESPFAL_XOR_v3_0/CLK 0.075
R7306 CLK1.n962 CLK1.n961 0.075
R7307 CLK1.n981 CLK1.n980 0.075
R7308 CLK1.n583 CLK1.n582 0.075
R7309 CLK1.n593 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/CLK 0.075
R7310 CLK1.n594 CLK1.n535 0.075
R7311 CLK1.n703 CLK1.n702 0.075
R7312 CLK1.n713 EESPFAL_s3_0/EESPFAL_INV4_1/CLK 0.075
R7313 CLK1.n714 CLK1.n671 0.075
R7314 CLK1.n742 CLK1.n741 0.075
R7315 CLK1.n761 CLK1.n649 0.075
R7316 CLK1.n774 EESPFAL_s3_0/EESPFAL_XOR_v3_1/CLK 0.075
R7317 CLK1.n777 CLK1.n776 0.075
R7318 CLK1.n796 CLK1.n795 0.075
R7319 CLK1.n448 CLK1.n447 0.075
R7320 CLK1.n458 EESPFAL_s2_0/EESPFAL_INV4_1/CLK 0.075
R7321 CLK1.n459 CLK1.n416 0.075
R7322 CLK1.n1054 CLK1.n1053 0.075
R7323 CLK1.n1035 CLK1.n494 0.075
R7324 CLK1.n1025 EESPFAL_s2_0/EESPFAL_XOR_v3_0/CLK 0.075
R7325 CLK1.n1023 CLK1.n503 0.075
R7326 CLK1.n1005 CLK1.n1004 0.075
R7327 CLK1.n1215 CLK1.n1214 0.075
R7328 CLK1.n1225 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/CLK 0.075
R7329 CLK1.n1226 CLK1.n295 0.075
R7330 CLK1.n1335 CLK1.n1334 0.075
R7331 CLK1.n1345 EESPFAL_s1_0/EESPFAL_INV4_1/CLK 0.075
R7332 CLK1.n1346 CLK1.n1303 0.075
R7333 CLK1.n1374 CLK1.n1373 0.075
R7334 CLK1.n1393 CLK1.n1281 0.075
R7335 CLK1.n1406 EESPFAL_s1_0/EESPFAL_XOR_v3_1/CLK 0.075
R7336 CLK1.n1409 CLK1.n1408 0.075
R7337 CLK1.n1428 CLK1.n1427 0.075
R7338 CLK1.n561 CLK1.n560 0.062
R7339 CLK1.n616 CLK1.n522 0.062
R7340 CLK1.n1193 CLK1.n1192 0.062
R7341 CLK1.n1248 CLK1.n282 0.062
R7342 CLK1.n1178 CLK1.n391 0.041
R7343 CLK1.n1170 CLK1.n391 0.041
R7344 CLK1.n1170 CLK1.n1169 0.041
R7345 CLK1.n1167 CLK1.n1066 0.041
R7346 CLK1.n1159 CLK1.n1066 0.041
R7347 CLK1.n1159 CLK1.n1158 0.041
R7348 CLK1.n1158 CLK1.n1157 0.041
R7349 CLK1.n1157 CLK1.n1072 0.041
R7350 CLK1.n1151 CLK1.n1150 0.041
R7351 CLK1.n1150 CLK1.n1149 0.041
R7352 CLK1.n1149 CLK1.n1082 0.041
R7353 CLK1.n1143 CLK1.n1142 0.041
R7354 CLK1.n1142 CLK1.n1141 0.041
R7355 CLK1.n1135 CLK1.n1098 0.041
R7356 CLK1.n1135 CLK1.n1134 0.041
R7357 CLK1.n1134 CLK1.n1133 0.041
R7358 CLK1.n1125 CLK1.n1107 0.041
R7359 CLK1.n1123 CLK1.n1122 0.041
R7360 CLK1.n623 CLK1.n522 0.037
R7361 CLK1.n1255 CLK1.n282 0.037
R7362 CLK1.n1133 CLK1.n1100 0.036
R7363 CLK1.n624 CLK1.n521 0.034
R7364 CLK1.n1256 CLK1.n281 0.034
R7365 CLK1.n809 EESPFAL_s3_0/CLK1 0.032
R7366 CLK1.n1441 EESPFAL_s1_0/CLK1 0.032
R7367 CLK1.n1168 CLK1.n1167 0.031
R7368 CLK1.n1151 CLK1.n1079 0.031
R7369 CLK1.n1143 EESPFAL_s2_0/EESPFAL_XOR_v3_1/CLK 0.031
R7370 CLK1.n1141 CLK1.n1090 0.031
R7371 CLK1.n1125 CLK1.n1124 0.031
R7372 CLK1.n34 CLK1.n33 0.025
R7373 CLK1.n47 CLK1 0.025
R7374 CLK1.n65 CLK1.n61 0.025
R7375 CLK1.n88 CLK1.n86 0.025
R7376 CLK1.n103 CLK1.n102 0.025
R7377 CLK1.n128 CLK1.n127 0.025
R7378 CLK1.n141 EESPFAL_s0_0/EESPFAL_XOR_v3_0/CLK 0.025
R7379 CLK1.n159 CLK1.n155 0.025
R7380 CLK1.n184 CLK1.n180 0.025
R7381 CLK1.n240 CLK1.n239 0.025
R7382 CLK1.n251 EESPFAL_s0_0/EESPFAL_NAND_v3_2/CLK 0.025
R7383 CLK1.n262 CLK1.n261 0.025
R7384 CLK1.n1519 CLK1.n1518 0.025
R7385 EESPFAL_s1_0/EESPFAL_INV4_2/CLK CLK1.n1529 0.025
R7386 CLK1.n1540 CLK1.n1488 0.025
R7387 CLK1.n1558 CLK1.n1557 0.025
R7388 CLK1.n1569 CLK1.n1466 0.025
R7389 CLK1.n1581 EESPFAL_s1_0/EESPFAL_XOR_v3_0/CLK 0.025
R7390 CLK1.n1593 CLK1.n1456 0.025
R7391 CLK1.n1614 CLK1.n1613 0.025
R7392 CLK1.n359 CLK1.n358 0.025
R7393 EESPFAL_s2_0/EESPFAL_INV4_0/CLK CLK1.n369 0.025
R7394 CLK1.n380 CLK1.n328 0.025
R7395 CLK1.n887 CLK1.n886 0.025
R7396 EESPFAL_s3_0/EESPFAL_INV4_2/CLK CLK1.n897 0.025
R7397 CLK1.n908 CLK1.n856 0.025
R7398 CLK1.n926 CLK1.n925 0.025
R7399 CLK1.n937 CLK1.n834 0.025
R7400 CLK1.n949 EESPFAL_s3_0/EESPFAL_XOR_v3_0/CLK 0.025
R7401 CLK1.n961 CLK1.n824 0.025
R7402 CLK1.n982 CLK1.n981 0.025
R7403 CLK1.n582 CLK1.n581 0.025
R7404 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/CLK CLK1.n592 0.025
R7405 CLK1.n603 CLK1.n535 0.025
R7406 CLK1.n702 CLK1.n701 0.025
R7407 EESPFAL_s3_0/EESPFAL_INV4_1/CLK CLK1.n712 0.025
R7408 CLK1.n723 CLK1.n671 0.025
R7409 CLK1.n741 CLK1.n740 0.025
R7410 CLK1.n752 CLK1.n649 0.025
R7411 CLK1.n764 EESPFAL_s3_0/EESPFAL_XOR_v3_1/CLK 0.025
R7412 CLK1.n776 CLK1.n639 0.025
R7413 CLK1.n797 CLK1.n796 0.025
R7414 CLK1.n447 CLK1.n446 0.025
R7415 EESPFAL_s2_0/EESPFAL_INV4_1/CLK CLK1.n457 0.025
R7416 CLK1.n468 CLK1.n416 0.025
R7417 CLK1.n1054 CLK1.n401 0.025
R7418 CLK1.n494 CLK1.n489 0.025
R7419 EESPFAL_s2_0/EESPFAL_XOR_v3_0/CLK CLK1.n496 0.025
R7420 CLK1.n509 CLK1.n503 0.025
R7421 CLK1.n1004 CLK1.n1003 0.025
R7422 CLK1.n1122 CLK1.n1110 0.025
R7423 CLK1.n1214 CLK1.n1213 0.025
R7424 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/CLK CLK1.n1224 0.025
R7425 CLK1.n1235 CLK1.n295 0.025
R7426 CLK1.n1334 CLK1.n1333 0.025
R7427 EESPFAL_s1_0/EESPFAL_INV4_1/CLK CLK1.n1344 0.025
R7428 CLK1.n1355 CLK1.n1303 0.025
R7429 CLK1.n1373 CLK1.n1372 0.025
R7430 CLK1.n1384 CLK1.n1281 0.025
R7431 CLK1.n1396 EESPFAL_s1_0/EESPFAL_XOR_v3_1/CLK 0.025
R7432 CLK1.n1408 CLK1.n1271 0.025
R7433 CLK1.n1429 CLK1.n1428 0.025
R7434 EESPFAL_s2_0/CLK1 CLK1.n994 0.02
R7435 CLK1.n1179 CLK1.n390 0.02
R7436 CLK1.n1179 CLK1.n1178 0.02
R7437 CLK1.n1622 CLK1.n1442 0.018
R7438 CLK1.n990 CLK1.n810 0.018
R7439 CLK1.n805 CLK1.n625 0.018
R7440 CLK1.n1437 CLK1.n1257 0.018
R7441 CLK1.n1625 CLK1.n280 0.016
R7442 CLK1.n993 CLK1.n520 0.016
R7443 CLK1.n808 CLK1.n521 0.016
R7444 CLK1.n1440 CLK1.n281 0.016
R7445 CLK1.n806 CLK1.n805 0.015
R7446 CLK1.n1438 CLK1.n1437 0.015
R7447 CLK1.n1113 CLK1.n1110 0.015
R7448 CLK1.n1623 CLK1.n1622 0.015
R7449 CLK1.n991 CLK1.n990 0.015
R7450 CLK1.n17 CLK1.n16 0.012
R7451 CLK1.n273 CLK1.n272 0.012
R7452 CLK1.n1549 CLK1.n1482 0.012
R7453 CLK1.n389 CLK1.n322 0.012
R7454 CLK1.n917 CLK1.n850 0.012
R7455 CLK1.n614 CLK1.n529 0.012
R7456 CLK1.n732 CLK1.n665 0.012
R7457 CLK1.n477 CLK1.n410 0.012
R7458 CLK1.n1246 CLK1.n289 0.012
R7459 CLK1.n1364 CLK1.n1297 0.012
R7460 CLK1.n807 CLK1.n806 0.011
R7461 CLK1.n1439 CLK1.n1438 0.011
R7462 CLK1.n992 CLK1.n991 0.01
R7463 CLK1.n1624 CLK1.n1623 0.01
R7464 CLK1.n1169 CLK1.n1168 0.01
R7465 CLK1.n1079 CLK1.n1072 0.01
R7466 EESPFAL_s2_0/EESPFAL_XOR_v3_1/CLK CLK1.n1082 0.01
R7467 CLK1.n1098 CLK1.n1090 0.01
R7468 CLK1.n1124 CLK1.n1123 0.01
R7469 CLK1.n996 CLK1.n995 0.006
R7470 CLK1.n1107 CLK1.n1100 0.005
R7471 EESPFAL_s3_0/CLK1 CLK1.n520 0.001
R7472 EESPFAL_s1_0/CLK1 CLK1.n280 0.001
R7473 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t8 819.4
R7474 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t9 736.033
R7475 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t6 514.133
R7476 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t7 305.266
R7477 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n5 192
R7478 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n0 166.734
R7479 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n4 105.6
R7480 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t3 97.937
R7481 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t2 97.937
R7482 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n1 76
R7483 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n3 73.939
R7484 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n2 57.6
R7485 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n6 56.157
R7486 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t5 39.4
R7487 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t0 39.4
R7488 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t4 24
R7489 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t1 24
R7490 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT 3.2
R7491 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t9 1074.82
R7492 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t8 819.4
R7493 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t7 506.1
R7494 EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 442.013
R7495 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t6 313.3
R7496 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t2 273.936
R7497 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n3 128.335
R7498 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n1 105.6
R7499 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t0 81.937
R7500 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n0 57.937
R7501 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n4 57.6
R7502 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n2 41.6
R7503 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t5 39.4
R7504 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t4 39.4
R7505 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t3 24
R7506 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t1 24
R7507 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n5 8.764
R7508 EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n6 4.65
R7509 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A x3_bar.t8 1271.5
R7510 x3_bar.n3 x3_bar.t11 1069.04
R7511 x3_bar.n3 x3_bar.t12 1015.9
R7512 x3_bar.n0 x3_bar.t4 810.772
R7513 x3_bar.n4 x3_bar.t6 810.772
R7514 x3_bar.n2 x3_bar.t10 810.772
R7515 EESPFAL_s3_0/EESPFAL_INV4_2/A x3_bar.t1 778.1
R7516 x3_bar.n0 x3_bar.t9 694.566
R7517 x3_bar.n4 x3_bar.t0 694.566
R7518 x3_bar.n2 x3_bar.t5 694.566
R7519 EESPFAL_s2_0/EESPFAL_4in_NAND_0/A x3_bar.t2 447.076
R7520 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C_bar x3_bar.t7 430.966
R7521 EESPFAL_s1_0/EESPFAL_INV4_2/A_bar x3_bar.t3 392.5
R7522 x3_bar.n11 EESPFAL_s1_0/EESPFAL_INV4_2/A_bar 179.64
R7523 x3_bar.n5 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C_bar 110.353
R7524 x3_bar.n9 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A 108.01
R7525 EESPFAL_s2_0/EESPFAL_XOR_v3_0/A_bar x3_bar.n3 89.6
R7526 x3_bar.n7 EESPFAL_s2_0/EESPFAL_XOR_v3_0/A_bar 72.49
R7527 x3_bar.n8 EESPFAL_s2_0/EESPFAL_4in_NAND_0/A 72.49
R7528 x3_bar.n1 x3_bar 59.69
R7529 x3_bar.n5 EESPFAL_s3_0/EESPFAL_XOR_v3_1/B_bar 59.69
R7530 x3_bar.n10 EESPFAL_s1_0/EESPFAL_XOR_v3_1/B_bar 59.69
R7531 x3_bar.n6 EESPFAL_s3_0/EESPFAL_INV4_2/A 40.836
R7532 x3_bar x3_bar.n0 25.6
R7533 EESPFAL_s3_0/EESPFAL_XOR_v3_1/B_bar x3_bar.n4 25.6
R7534 EESPFAL_s1_0/EESPFAL_XOR_v3_1/B_bar x3_bar.n2 25.6
R7535 EESPFAL_s1_0/x3_bar x3_bar.n1 4.084
R7536 x3_bar.n9 x3_bar.n8 3.984
R7537 x3_bar.n8 x3_bar.n7 3.717
R7538 EESPFAL_s3_0/x3_bar x3_bar.n5 2.634
R7539 x3_bar.n11 x3_bar.n10 1.69
R7540 x3_bar.n10 x3_bar.n9 1.578
R7541 EESPFAL_s2_0/x3_bar x3_bar.n6 1.206
R7542 EESPFAL_s1_0/x3_bar x3_bar.n11 0.912
R7543 x3_bar.n1 EESPFAL_s0_0/x3_bar 0.323
R7544 x3_bar.n6 EESPFAL_s3_0/x3_bar 0.181
R7545 x3_bar.n7 EESPFAL_s2_0/x3_bar 0.075
R7546 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t9 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t6 819.4
R7547 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t8 736.033
R7548 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t7 506.1
R7549 EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 367.829
R7550 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t9 313.3
R7551 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t0 273.937
R7552 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n0 128.334
R7553 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n2 105.6
R7554 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t1 81.937
R7555 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n1 57.937
R7556 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n4 57.6
R7557 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n3 41.6
R7558 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t5 39.4
R7559 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t2 39.4
R7560 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t3 24
R7561 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t4 24
R7562 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n5 8.764
R7563 EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n6 4.65
R7564 Dis2.n6 Dis2.n4 532.126
R7565 Dis2.n19 Dis2.t7 504.5
R7566 Dis2.n17 Dis2.t19 504.5
R7567 Dis2.n11 Dis2.t21 504.5
R7568 Dis2.n9 Dis2.t6 504.5
R7569 Dis2.n7 Dis2.t14 504.5
R7570 Dis2.n5 Dis2.t20 504.5
R7571 Dis2.n0 Dis2.t13 504.5
R7572 Dis2.n19 Dis2.t16 389.3
R7573 Dis2.n17 Dis2.t4 389.3
R7574 Dis2.n15 Dis2.t11 389.3
R7575 Dis2.n14 Dis2.t18 389.3
R7576 Dis2.n11 Dis2.t9 389.3
R7577 Dis2.n9 Dis2.t0 389.3
R7578 Dis2.n7 Dis2.t2 389.3
R7579 Dis2.n5 Dis2.t3 389.3
R7580 Dis2.n4 Dis2.t12 389.3
R7581 Dis2.n3 Dis2.t17 389.3
R7582 Dis2.n2 Dis2.t8 389.3
R7583 Dis2.n1 Dis2.t15 389.3
R7584 Dis2.n22 Dis2.t10 389.3
R7585 Dis2.n21 Dis2.t1 389.3
R7586 Dis2.n0 Dis2.t5 389.3
R7587 Dis2.n16 Dis2.n15 273.536
R7588 Dis2.n24 Dis2.n23 265.28
R7589 Dis2.n18 Dis2.n16 258.592
R7590 Dis2.n13 Dis2.n12 243.072
R7591 Dis2.n12 EESPFAL_s2_0/EESPFAL_NAND_v3_0/Dis 177.536
R7592 Dis2.n20 EESPFAL_s1_0/EESPFAL_NAND_v3_0/Dis 177.216
R7593 Dis2.n18 EESPFAL_s1_0/EESPFAL_NAND_v3_1/Dis 177.216
R7594 Dis2.n8 EESPFAL_s3_0/EESPFAL_NAND_v3_0/Dis 177.216
R7595 Dis2.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_1/Dis 177.216
R7596 Dis2.n10 EESPFAL_s2_0/EESPFAL_NAND_v3_1/Dis 176.896
R7597 Dis2.n13 Dis2.n2 165.061
R7598 Dis2.n24 Dis2 149.76
R7599 Dis2.n23 Dis2.n22 125.76
R7600 Dis2.n15 Dis2.n14 115.2
R7601 Dis2.n4 Dis2.n3 115.2
R7602 Dis2.n2 Dis2.n1 115.2
R7603 Dis2.n22 Dis2.n21 115.2
R7604 Dis2.n23 EESPFAL_s1_0/Dis2 9.259
R7605 Dis2 Dis2.n24 6.908
R7606 EESPFAL_s2_0/Dis2 EESPFAL_s3_0/Dis2 5.575
R7607 Dis2.n10 EESPFAL_s2_0/Dis2 3.357
R7608 EESPFAL_s1_0/Dis2 Dis2.n20 3.284
R7609 EESPFAL_s3_0/Dis2 Dis2.n8 3.284
R7610 EESPFAL_s1_0/EESPFAL_NAND_v3_0/Dis Dis2.n19 3.2
R7611 EESPFAL_s1_0/EESPFAL_NAND_v3_1/Dis Dis2.n17 3.2
R7612 Dis2.n14 EESPFAL_s1_0/EESPFAL_INV4_0/Dis 3.2
R7613 EESPFAL_s2_0/EESPFAL_NAND_v3_0/Dis Dis2.n11 3.2
R7614 EESPFAL_s2_0/EESPFAL_NAND_v3_1/Dis Dis2.n9 3.2
R7615 EESPFAL_s3_0/EESPFAL_NAND_v3_0/Dis Dis2.n7 3.2
R7616 EESPFAL_s3_0/EESPFAL_NAND_v3_1/Dis Dis2.n5 3.2
R7617 Dis2.n3 EESPFAL_s3_0/EESPFAL_INV4_0/Dis 3.2
R7618 Dis2.n1 EESPFAL_s2_0/EESPFAL_INV4_2/Dis 3.2
R7619 Dis2.n21 EESPFAL_s0_0/EESPFAL_NAND_v3_1/Dis 3.2
R7620 Dis2 Dis2.n0 3.2
R7621 Dis2.n16 Dis2.n13 2.039
R7622 Dis2.n12 Dis2.n10 0.627
R7623 Dis2.n8 Dis2.n6 0.623
R7624 Dis2.n20 Dis2.n18 0.623
R7625 EESPFAL_s0_0/Dis2 Dis2 0.162
R7626 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/A_bar 951.139
R7627 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t9 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t7 819.4
R7628 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t6 684.833
R7629 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n5 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t8 506.1
R7630 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n5 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t9 313.3
R7631 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n1 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t5 177.936
R7632 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n4 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n3 128.336
R7633 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n1 105.6
R7634 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n1 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t4 81.937
R7635 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n0 58.265
R7636 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n6 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n4 57.6
R7637 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n4 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n2 41.6
R7638 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n3 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t1 39.4
R7639 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n3 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t2 39.4
R7640 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n0 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t0 24
R7641 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n0 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t3 24
R7642 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n6 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n5 8.764
R7643 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n6 4.65
R7644 x0.n0 x0.t10 1176.57
R7645 x0.n0 x0.t6 1149.49
R7646 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B x0.t9 1106.75
R7647 x0.n3 x0.t8 800.452
R7648 x0.n2 x0.t0 800.452
R7649 x0.n1 x0.t5 800.452
R7650 x0.n3 x0.t4 787.997
R7651 x0.n2 x0.t1 787.997
R7652 x0.n1 x0.t3 787.997
R7653 EESPFAL_s2_0/EESPFAL_4in_NAND_0/C x0.t7 445.388
R7654 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C_bar x0.t2 430.966
R7655 x0.n4 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B 367.635
R7656 x0.n7 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C_bar 363.37
R7657 x0.n5 EESPFAL_s2_0/EESPFAL_XOR_v3_1/B 327.85
R7658 x0.n6 EESPFAL_s2_0/EESPFAL_4in_NAND_0/C 327.85
R7659 EESPFAL_s0_0/x0 x0 315.101
R7660 x0.n4 EESPFAL_s3_0/EESPFAL_XOR_v3_0/B 315.05
R7661 x0.n8 EESPFAL_s1_0/EESPFAL_XOR_v3_0/B 315.05
R7662 EESPFAL_s3_0/EESPFAL_XOR_v3_0/B x0.n3 169.6
R7663 EESPFAL_s2_0/EESPFAL_XOR_v3_1/B x0.n2 169.6
R7664 EESPFAL_s1_0/EESPFAL_XOR_v3_0/B x0.n1 169.6
R7665 x0 x0.n0 128
R7666 x0.n8 x0.n7 4.812
R7667 EESPFAL_s1_0/x0 EESPFAL_s0_0/x0 4.407
R7668 x0.n5 EESPFAL_s2_0/x0 2.976
R7669 x0.n7 x0.n6 2.781
R7670 x0.n6 x0.n5 1.346
R7671 EESPFAL_s2_0/x0 EESPFAL_s3_0/x0 1.2
R7672 EESPFAL_s1_0/x0 x0.n8 0.228
R7673 EESPFAL_s3_0/x0 x0.n4 0.228
R7674 s0.t8 s0.t6 819.4
R7675 s0.n2 s0.t8 514.133
R7676 s0.n2 s0.t7 305.266
R7677 s0.n3 s0.n1 166.734
R7678 s0.n4 s0.n3 99.2
R7679 s0.n5 s0.n4 99.2
R7680 s0.n4 s0.t5 97.937
R7681 s0.n5 s0.t4 91.537
R7682 s0 s0.n2 79.2
R7683 s0.n3 s0.n0 73.937
R7684 s0.n3 s0 54.4
R7685 s0.n1 s0.t3 39.4
R7686 s0.n1 s0.t1 39.4
R7687 s0.n0 s0.t2 24
R7688 s0.n0 s0.t0 24
R7689 s0 s0.n5 12.406
R7690 EESPFAL_s0_0/s0 s0 0.084
R7691 s0_bar.t7 s0_bar.t5 819.4
R7692 s0_bar.n4 s0_bar.t6 506.1
R7693 s0_bar.n4 s0_bar.t7 313.3
R7694 s0_bar.n1 s0_bar.t0 187.536
R7695 s0_bar.n3 s0_bar.n2 128.334
R7696 s0_bar.n1 s0_bar.n0 57.937
R7697 s0_bar.n5 s0_bar.n3 57.6
R7698 s0_bar.n3 s0_bar.n1 41.6
R7699 s0_bar.n2 s0_bar.t3 39.4
R7700 s0_bar.n2 s0_bar.t2 39.4
R7701 s0_bar.n0 s0_bar.t4 24
R7702 s0_bar.n0 s0_bar.t1 24
R7703 s0_bar.n5 s0_bar.n4 8.764
R7704 s0_bar s0_bar.n5 4.681
R7705 EESPFAL_s0_0/s0_bar s0_bar 0.081
R7706 CLK3.n414 CLK3.n413 407.048
R7707 CLK3.n37 CLK3.n28 407.048
R7708 CLK3.n345 CLK3.n344 407.048
R7709 CLK3.n400 CLK3.n399 407.048
R7710 CLK3.n270 CLK3.n269 407.048
R7711 CLK3.n324 CLK3.n323 407.048
R7712 CLK3.n199 CLK3.n198 407.048
R7713 CLK3.n254 CLK3.n253 407.048
R7714 CLK3.n72 CLK3.n3 400
R7715 CLK3.n413 CLK3.n3 400
R7716 CLK3.n38 CLK3.n37 400
R7717 CLK3.n39 CLK3.n38 400
R7718 CLK3.n346 CLK3.n345 400
R7719 CLK3.n346 CLK3.n108 400
R7720 CLK3.n354 CLK3.n108 400
R7721 CLK3.n355 CLK3.n354 400
R7722 CLK3.n389 CLK3.n388 400
R7723 CLK3.n389 CLK3.n83 400
R7724 CLK3.n398 CLK3.n83 400
R7725 CLK3.n399 CLK3.n398 400
R7726 CLK3.n281 CLK3.n280 400
R7727 CLK3.n280 CLK3.n147 400
R7728 CLK3.n271 CLK3.n147 400
R7729 CLK3.n271 CLK3.n270 400
R7730 CLK3.n323 CLK3.n322 400
R7731 CLK3.n322 CLK3.n122 400
R7732 CLK3.n314 CLK3.n122 400
R7733 CLK3.n314 CLK3.n313 400
R7734 CLK3.n200 CLK3.n199 400
R7735 CLK3.n200 CLK3.n187 400
R7736 CLK3.n208 CLK3.n187 400
R7737 CLK3.n209 CLK3.n208 400
R7738 CLK3.n243 CLK3.n242 400
R7739 CLK3.n243 CLK3.n162 400
R7740 CLK3.n252 CLK3.n162 400
R7741 CLK3.n253 CLK3.n252 400
R7742 CLK3.n72 CLK3.n71 366.379
R7743 CLK3.n39 CLK3.n22 366.379
R7744 CLK3.n356 CLK3.n355 366.379
R7745 CLK3.n388 CLK3.n387 366.379
R7746 CLK3.n282 CLK3.n281 366.379
R7747 CLK3.n313 CLK3.n312 366.379
R7748 CLK3.n210 CLK3.n209 366.379
R7749 CLK3.n242 CLK3.n241 366.379
R7750 CLK3.n48 CLK3.n22 131.034
R7751 CLK3.n49 CLK3.n48 131.034
R7752 CLK3.n51 CLK3.n50 131.034
R7753 CLK3.n61 CLK3.n60 131.034
R7754 CLK3.n70 CLK3.n10 131.034
R7755 CLK3.n71 CLK3.n70 131.034
R7756 CLK3.n356 CLK3.n102 131.034
R7757 CLK3.n365 CLK3.n102 131.034
R7758 CLK3.n368 CLK3.n366 131.034
R7759 CLK3.n377 CLK3.n376 131.034
R7760 CLK3.n378 CLK3.n90 131.034
R7761 CLK3.n387 CLK3.n90 131.034
R7762 CLK3.n312 CLK3.n128 131.034
R7763 CLK3.n303 CLK3.n128 131.034
R7764 CLK3.n302 CLK3.n301 131.034
R7765 CLK3.n293 CLK3.n292 131.034
R7766 CLK3.n291 CLK3.n141 131.034
R7767 CLK3.n282 CLK3.n141 131.034
R7768 CLK3.n210 CLK3.n181 131.034
R7769 CLK3.n219 CLK3.n181 131.034
R7770 CLK3.n222 CLK3.n220 131.034
R7771 CLK3.n231 CLK3.n230 131.034
R7772 CLK3.n232 CLK3.n169 131.034
R7773 CLK3.n241 CLK3.n169 131.034
R7774 CLK3.n59 CLK3.t24 122.844
R7775 CLK3.t18 CLK3.n59 122.844
R7776 CLK3.t43 CLK3.n367 122.844
R7777 CLK3.n367 CLK3.t32 122.844
R7778 CLK3.n140 CLK3.t36 122.844
R7779 CLK3.t16 CLK3.n140 122.844
R7780 CLK3.t45 CLK3.n221 122.844
R7781 CLK3.n221 CLK3.t30 122.844
R7782 CLK3.n51 CLK3.t26 106.465
R7783 CLK3.n61 CLK3.t20 106.465
R7784 CLK3.n366 CLK3.t41 106.465
R7785 CLK3.t34 CLK3.n377 106.465
R7786 CLK3.t12 CLK3.n302 106.465
R7787 CLK3.n292 CLK3.t2 106.465
R7788 CLK3.n220 CLK3.t5 106.465
R7789 CLK3.t7 CLK3.n231 106.465
R7790 CLK3.n36 CLK3.n29 96
R7791 CLK3.n36 CLK3.n27 96
R7792 CLK3.n40 CLK3.n27 96
R7793 CLK3.n40 CLK3.n23 96
R7794 CLK3.n47 CLK3.n23 96
R7795 CLK3.n47 CLK3.n21 96
R7796 CLK3.n52 CLK3.n21 96
R7797 CLK3.n52 CLK3.n16 96
R7798 CLK3.n58 CLK3.n16 96
R7799 CLK3.n58 CLK3.n15 96
R7800 CLK3.n62 CLK3.n15 96
R7801 CLK3.n62 CLK3.n11 96
R7802 CLK3.n69 CLK3.n11 96
R7803 CLK3.n69 CLK3.n9 96
R7804 CLK3.n73 CLK3.n9 96
R7805 CLK3.n73 CLK3.n4 96
R7806 CLK3.n412 CLK3.n4 96
R7807 CLK3.n412 CLK3.n2 96
R7808 CLK3.n343 CLK3.n113 96
R7809 CLK3.n347 CLK3.n113 96
R7810 CLK3.n347 CLK3.n109 96
R7811 CLK3.n353 CLK3.n109 96
R7812 CLK3.n353 CLK3.n107 96
R7813 CLK3.n357 CLK3.n107 96
R7814 CLK3.n357 CLK3.n103 96
R7815 CLK3.n364 CLK3.n103 96
R7816 CLK3.n364 CLK3.n101 96
R7817 CLK3.n369 CLK3.n101 96
R7818 CLK3.n369 CLK3.n96 96
R7819 CLK3.n375 CLK3.n96 96
R7820 CLK3.n375 CLK3.n95 96
R7821 CLK3.n379 CLK3.n95 96
R7822 CLK3.n379 CLK3.n91 96
R7823 CLK3.n386 CLK3.n91 96
R7824 CLK3.n386 CLK3.n89 96
R7825 CLK3.n390 CLK3.n89 96
R7826 CLK3.n390 CLK3.n84 96
R7827 CLK3.n397 CLK3.n84 96
R7828 CLK3.n397 CLK3.n82 96
R7829 CLK3.n401 CLK3.n82 96
R7830 CLK3.n325 CLK3.n121 96
R7831 CLK3.n321 CLK3.n121 96
R7832 CLK3.n321 CLK3.n123 96
R7833 CLK3.n315 CLK3.n123 96
R7834 CLK3.n315 CLK3.n127 96
R7835 CLK3.n311 CLK3.n127 96
R7836 CLK3.n311 CLK3.n129 96
R7837 CLK3.n304 CLK3.n129 96
R7838 CLK3.n304 CLK3.n133 96
R7839 CLK3.n300 CLK3.n133 96
R7840 CLK3.n300 CLK3.n134 96
R7841 CLK3.n294 CLK3.n134 96
R7842 CLK3.n294 CLK3.n139 96
R7843 CLK3.n290 CLK3.n139 96
R7844 CLK3.n290 CLK3.n142 96
R7845 CLK3.n283 CLK3.n142 96
R7846 CLK3.n283 CLK3.n146 96
R7847 CLK3.n279 CLK3.n146 96
R7848 CLK3.n279 CLK3.n148 96
R7849 CLK3.n272 CLK3.n148 96
R7850 CLK3.n272 CLK3.n153 96
R7851 CLK3.n268 CLK3.n153 96
R7852 CLK3.n197 CLK3.n192 96
R7853 CLK3.n201 CLK3.n192 96
R7854 CLK3.n201 CLK3.n188 96
R7855 CLK3.n207 CLK3.n188 96
R7856 CLK3.n207 CLK3.n186 96
R7857 CLK3.n211 CLK3.n186 96
R7858 CLK3.n211 CLK3.n182 96
R7859 CLK3.n218 CLK3.n182 96
R7860 CLK3.n218 CLK3.n180 96
R7861 CLK3.n223 CLK3.n180 96
R7862 CLK3.n223 CLK3.n175 96
R7863 CLK3.n229 CLK3.n175 96
R7864 CLK3.n229 CLK3.n174 96
R7865 CLK3.n233 CLK3.n174 96
R7866 CLK3.n233 CLK3.n170 96
R7867 CLK3.n240 CLK3.n170 96
R7868 CLK3.n240 CLK3.n168 96
R7869 CLK3.n244 CLK3.n168 96
R7870 CLK3.n244 CLK3.n163 96
R7871 CLK3.n251 CLK3.n163 96
R7872 CLK3.n251 CLK3.n161 96
R7873 CLK3.n255 CLK3.n161 96
R7874 CLK3.n31 CLK3.n28 85.261
R7875 CLK3.n400 CLK3.n79 85.261
R7876 CLK3.n324 CLK3.n118 85.261
R7877 CLK3.n254 CLK3.n158 85.261
R7878 CLK3.n415 CLK3.n414 85.261
R7879 CLK3.n344 CLK3.n114 85.261
R7880 CLK3.n269 CLK3.n154 85.261
R7881 CLK3.n198 CLK3.n193 85.261
R7882 CLK3.n307 CLK3.t13 44.338
R7883 CLK3.n287 CLK3.t3 44.338
R7884 CLK3.n44 CLK3.t27 44.338
R7885 CLK3.n66 CLK3.t21 44.338
R7886 CLK3.n382 CLK3.t35 44.337
R7887 CLK3.n361 CLK3.t42 44.337
R7888 CLK3.n236 CLK3.t8 44.337
R7889 CLK3.n215 CLK3.t6 44.337
R7890 CLK3.n407 CLK3.n406 44.163
R7891 CLK3.n18 CLK3.t25 39.4
R7892 CLK3.n18 CLK3.t19 39.4
R7893 CLK3.n98 CLK3.t44 39.4
R7894 CLK3.n98 CLK3.t33 39.4
R7895 CLK3.n136 CLK3.t37 39.4
R7896 CLK3.n136 CLK3.t17 39.4
R7897 CLK3.n177 CLK3.t46 39.4
R7898 CLK3.n177 CLK3.t31 39.4
R7899 CLK3.n264 CLK3.t0 30.776
R7900 CLK3.n32 CLK3.t23 30.776
R7901 CLK3.n404 CLK3.t1 30.775
R7902 CLK3.n258 CLK3.t39 30.775
R7903 CLK3.n194 CLK3.t14 30.775
R7904 CLK3.t26 CLK3.n49 24.568
R7905 CLK3.t20 CLK3.n10 24.568
R7906 CLK3.t41 CLK3.n365 24.568
R7907 CLK3.n378 CLK3.t34 24.568
R7908 CLK3.n303 CLK3.t12 24.568
R7909 CLK3.t2 CLK3.n291 24.568
R7910 CLK3.t5 CLK3.n219 24.568
R7911 CLK3.n232 CLK3.t7 24.568
R7912 CLK3.n86 CLK3.t15 24
R7913 CLK3.n86 CLK3.t11 24
R7914 CLK3.n331 CLK3.t38 24
R7915 CLK3.n165 CLK3.t40 24
R7916 CLK3.n165 CLK3.t9 24
R7917 CLK3.n150 CLK3.t22 24
R7918 CLK3.n150 CLK3.t29 24
R7919 CLK3.n335 CLK3.t4 24
R7920 CLK3.n6 CLK3.t28 24
R7921 CLK3.n6 CLK3.t10 24
R7922 CLK3.n31 CLK3.n30 12.8
R7923 CLK3.n35 CLK3.n30 12.8
R7924 CLK3.n35 CLK3.n26 12.8
R7925 CLK3.n41 CLK3.n26 12.8
R7926 CLK3.n41 CLK3.n24 12.8
R7927 CLK3.n46 CLK3.n24 12.8
R7928 CLK3.n46 CLK3.n20 12.8
R7929 CLK3.n53 CLK3.n20 12.8
R7930 CLK3.n53 CLK3.n17 12.8
R7931 CLK3.n57 CLK3.n17 12.8
R7932 CLK3.n57 CLK3.n14 12.8
R7933 CLK3.n63 CLK3.n14 12.8
R7934 CLK3.n63 CLK3.n12 12.8
R7935 CLK3.n68 CLK3.n12 12.8
R7936 CLK3.n68 CLK3.n8 12.8
R7937 CLK3.n74 CLK3.n8 12.8
R7938 CLK3.n74 CLK3.n5 12.8
R7939 CLK3.n411 CLK3.n5 12.8
R7940 CLK3.n411 CLK3.n1 12.8
R7941 CLK3.n415 CLK3.n1 12.8
R7942 CLK3.n342 CLK3.n114 12.8
R7943 CLK3.n342 CLK3.n112 12.8
R7944 CLK3.n348 CLK3.n112 12.8
R7945 CLK3.n348 CLK3.n110 12.8
R7946 CLK3.n352 CLK3.n110 12.8
R7947 CLK3.n352 CLK3.n106 12.8
R7948 CLK3.n358 CLK3.n106 12.8
R7949 CLK3.n358 CLK3.n104 12.8
R7950 CLK3.n363 CLK3.n104 12.8
R7951 CLK3.n363 CLK3.n100 12.8
R7952 CLK3.n370 CLK3.n100 12.8
R7953 CLK3.n370 CLK3.n97 12.8
R7954 CLK3.n374 CLK3.n97 12.8
R7955 CLK3.n374 CLK3.n94 12.8
R7956 CLK3.n380 CLK3.n94 12.8
R7957 CLK3.n380 CLK3.n92 12.8
R7958 CLK3.n385 CLK3.n92 12.8
R7959 CLK3.n385 CLK3.n88 12.8
R7960 CLK3.n391 CLK3.n88 12.8
R7961 CLK3.n391 CLK3.n85 12.8
R7962 CLK3.n396 CLK3.n85 12.8
R7963 CLK3.n396 CLK3.n81 12.8
R7964 CLK3.n402 CLK3.n81 12.8
R7965 CLK3.n402 CLK3.n79 12.8
R7966 CLK3.n330 CLK3.n117 12.8
R7967 CLK3.n326 CLK3.n118 12.8
R7968 CLK3.n326 CLK3.n120 12.8
R7969 CLK3.n320 CLK3.n120 12.8
R7970 CLK3.n320 CLK3.n124 12.8
R7971 CLK3.n316 CLK3.n124 12.8
R7972 CLK3.n316 CLK3.n126 12.8
R7973 CLK3.n310 CLK3.n126 12.8
R7974 CLK3.n310 CLK3.n130 12.8
R7975 CLK3.n305 CLK3.n130 12.8
R7976 CLK3.n305 CLK3.n132 12.8
R7977 CLK3.n299 CLK3.n132 12.8
R7978 CLK3.n299 CLK3.n135 12.8
R7979 CLK3.n295 CLK3.n135 12.8
R7980 CLK3.n295 CLK3.n138 12.8
R7981 CLK3.n289 CLK3.n138 12.8
R7982 CLK3.n289 CLK3.n143 12.8
R7983 CLK3.n284 CLK3.n143 12.8
R7984 CLK3.n284 CLK3.n145 12.8
R7985 CLK3.n278 CLK3.n145 12.8
R7986 CLK3.n278 CLK3.n149 12.8
R7987 CLK3.n273 CLK3.n149 12.8
R7988 CLK3.n273 CLK3.n152 12.8
R7989 CLK3.n196 CLK3.n193 12.8
R7990 CLK3.n196 CLK3.n191 12.8
R7991 CLK3.n202 CLK3.n191 12.8
R7992 CLK3.n202 CLK3.n189 12.8
R7993 CLK3.n206 CLK3.n189 12.8
R7994 CLK3.n206 CLK3.n185 12.8
R7995 CLK3.n212 CLK3.n185 12.8
R7996 CLK3.n212 CLK3.n183 12.8
R7997 CLK3.n217 CLK3.n183 12.8
R7998 CLK3.n217 CLK3.n179 12.8
R7999 CLK3.n224 CLK3.n179 12.8
R8000 CLK3.n224 CLK3.n176 12.8
R8001 CLK3.n228 CLK3.n176 12.8
R8002 CLK3.n228 CLK3.n173 12.8
R8003 CLK3.n234 CLK3.n173 12.8
R8004 CLK3.n234 CLK3.n171 12.8
R8005 CLK3.n239 CLK3.n171 12.8
R8006 CLK3.n239 CLK3.n167 12.8
R8007 CLK3.n245 CLK3.n167 12.8
R8008 CLK3.n245 CLK3.n164 12.8
R8009 CLK3.n250 CLK3.n164 12.8
R8010 CLK3.n250 CLK3.n160 12.8
R8011 CLK3.n256 CLK3.n160 12.8
R8012 CLK3.n256 CLK3.n158 12.8
R8013 CLK3.n337 CLK3.n336 12.8
R8014 CLK3.n155 CLK3.n152 12.32
R8015 CLK3.n156 CLK3.n154 10.56
R8016 CLK3 CLK3.n416 9.726
R8017 CLK3.n265 CLK3.n156 9.3
R8018 CLK3.n267 CLK3.n266 9.3
R8019 CLK3.n412 CLK3.n411 8.855
R8020 CLK3.n331 CLK3.n330 8.855
R8021 CLK3.n153 CLK3.n152 8.855
R8022 CLK3.n197 CLK3.n196 8.855
R8023 CLK3.n192 CLK3.n191 8.855
R8024 CLK3.n199 CLK3.n192 8.855
R8025 CLK3.n202 CLK3.n201 8.855
R8026 CLK3.n201 CLK3.n200 8.855
R8027 CLK3.n189 CLK3.n188 8.855
R8028 CLK3.n188 CLK3.n187 8.855
R8029 CLK3.n207 CLK3.n206 8.855
R8030 CLK3.n208 CLK3.n207 8.855
R8031 CLK3.n186 CLK3.n185 8.855
R8032 CLK3.n209 CLK3.n186 8.855
R8033 CLK3.n212 CLK3.n211 8.855
R8034 CLK3.n211 CLK3.n210 8.855
R8035 CLK3.n183 CLK3.n182 8.855
R8036 CLK3.n182 CLK3.n181 8.855
R8037 CLK3.n218 CLK3.n217 8.855
R8038 CLK3.n219 CLK3.n218 8.855
R8039 CLK3.n180 CLK3.n179 8.855
R8040 CLK3.n220 CLK3.n180 8.855
R8041 CLK3.n224 CLK3.n223 8.855
R8042 CLK3.n223 CLK3.n222 8.855
R8043 CLK3.n176 CLK3.n175 8.855
R8044 CLK3.n221 CLK3.n175 8.855
R8045 CLK3.n229 CLK3.n228 8.855
R8046 CLK3.n230 CLK3.n229 8.855
R8047 CLK3.n174 CLK3.n173 8.855
R8048 CLK3.n231 CLK3.n174 8.855
R8049 CLK3.n234 CLK3.n233 8.855
R8050 CLK3.n233 CLK3.n232 8.855
R8051 CLK3.n171 CLK3.n170 8.855
R8052 CLK3.n170 CLK3.n169 8.855
R8053 CLK3.n240 CLK3.n239 8.855
R8054 CLK3.n241 CLK3.n240 8.855
R8055 CLK3.n168 CLK3.n167 8.855
R8056 CLK3.n242 CLK3.n168 8.855
R8057 CLK3.n245 CLK3.n244 8.855
R8058 CLK3.n244 CLK3.n243 8.855
R8059 CLK3.n164 CLK3.n163 8.855
R8060 CLK3.n163 CLK3.n162 8.855
R8061 CLK3.n251 CLK3.n250 8.855
R8062 CLK3.n252 CLK3.n251 8.855
R8063 CLK3.n161 CLK3.n160 8.855
R8064 CLK3.n253 CLK3.n161 8.855
R8065 CLK3.n256 CLK3.n255 8.855
R8066 CLK3.n326 CLK3.n325 8.855
R8067 CLK3.n121 CLK3.n120 8.855
R8068 CLK3.n323 CLK3.n121 8.855
R8069 CLK3.n321 CLK3.n320 8.855
R8070 CLK3.n322 CLK3.n321 8.855
R8071 CLK3.n124 CLK3.n123 8.855
R8072 CLK3.n123 CLK3.n122 8.855
R8073 CLK3.n316 CLK3.n315 8.855
R8074 CLK3.n315 CLK3.n314 8.855
R8075 CLK3.n127 CLK3.n126 8.855
R8076 CLK3.n313 CLK3.n127 8.855
R8077 CLK3.n311 CLK3.n310 8.855
R8078 CLK3.n312 CLK3.n311 8.855
R8079 CLK3.n130 CLK3.n129 8.855
R8080 CLK3.n129 CLK3.n128 8.855
R8081 CLK3.n305 CLK3.n304 8.855
R8082 CLK3.n304 CLK3.n303 8.855
R8083 CLK3.n133 CLK3.n132 8.855
R8084 CLK3.n302 CLK3.n133 8.855
R8085 CLK3.n300 CLK3.n299 8.855
R8086 CLK3.n301 CLK3.n300 8.855
R8087 CLK3.n135 CLK3.n134 8.855
R8088 CLK3.n140 CLK3.n134 8.855
R8089 CLK3.n295 CLK3.n294 8.855
R8090 CLK3.n294 CLK3.n293 8.855
R8091 CLK3.n139 CLK3.n138 8.855
R8092 CLK3.n292 CLK3.n139 8.855
R8093 CLK3.n290 CLK3.n289 8.855
R8094 CLK3.n291 CLK3.n290 8.855
R8095 CLK3.n143 CLK3.n142 8.855
R8096 CLK3.n142 CLK3.n141 8.855
R8097 CLK3.n284 CLK3.n283 8.855
R8098 CLK3.n283 CLK3.n282 8.855
R8099 CLK3.n146 CLK3.n145 8.855
R8100 CLK3.n281 CLK3.n146 8.855
R8101 CLK3.n279 CLK3.n278 8.855
R8102 CLK3.n280 CLK3.n279 8.855
R8103 CLK3.n149 CLK3.n148 8.855
R8104 CLK3.n148 CLK3.n147 8.855
R8105 CLK3.n273 CLK3.n272 8.855
R8106 CLK3.n272 CLK3.n271 8.855
R8107 CLK3.n270 CLK3.n153 8.855
R8108 CLK3.n268 CLK3.n267 8.855
R8109 CLK3.n336 CLK3.n335 8.855
R8110 CLK3.n343 CLK3.n342 8.855
R8111 CLK3.n113 CLK3.n112 8.855
R8112 CLK3.n345 CLK3.n113 8.855
R8113 CLK3.n348 CLK3.n347 8.855
R8114 CLK3.n347 CLK3.n346 8.855
R8115 CLK3.n110 CLK3.n109 8.855
R8116 CLK3.n109 CLK3.n108 8.855
R8117 CLK3.n353 CLK3.n352 8.855
R8118 CLK3.n354 CLK3.n353 8.855
R8119 CLK3.n107 CLK3.n106 8.855
R8120 CLK3.n355 CLK3.n107 8.855
R8121 CLK3.n358 CLK3.n357 8.855
R8122 CLK3.n357 CLK3.n356 8.855
R8123 CLK3.n104 CLK3.n103 8.855
R8124 CLK3.n103 CLK3.n102 8.855
R8125 CLK3.n364 CLK3.n363 8.855
R8126 CLK3.n365 CLK3.n364 8.855
R8127 CLK3.n101 CLK3.n100 8.855
R8128 CLK3.n366 CLK3.n101 8.855
R8129 CLK3.n370 CLK3.n369 8.855
R8130 CLK3.n369 CLK3.n368 8.855
R8131 CLK3.n97 CLK3.n96 8.855
R8132 CLK3.n367 CLK3.n96 8.855
R8133 CLK3.n375 CLK3.n374 8.855
R8134 CLK3.n376 CLK3.n375 8.855
R8135 CLK3.n95 CLK3.n94 8.855
R8136 CLK3.n377 CLK3.n95 8.855
R8137 CLK3.n380 CLK3.n379 8.855
R8138 CLK3.n379 CLK3.n378 8.855
R8139 CLK3.n92 CLK3.n91 8.855
R8140 CLK3.n91 CLK3.n90 8.855
R8141 CLK3.n386 CLK3.n385 8.855
R8142 CLK3.n387 CLK3.n386 8.855
R8143 CLK3.n89 CLK3.n88 8.855
R8144 CLK3.n388 CLK3.n89 8.855
R8145 CLK3.n391 CLK3.n390 8.855
R8146 CLK3.n390 CLK3.n389 8.855
R8147 CLK3.n85 CLK3.n84 8.855
R8148 CLK3.n84 CLK3.n83 8.855
R8149 CLK3.n397 CLK3.n396 8.855
R8150 CLK3.n398 CLK3.n397 8.855
R8151 CLK3.n82 CLK3.n81 8.855
R8152 CLK3.n399 CLK3.n82 8.855
R8153 CLK3.n402 CLK3.n401 8.855
R8154 CLK3.n30 CLK3.n29 8.855
R8155 CLK3.n36 CLK3.n35 8.855
R8156 CLK3.n37 CLK3.n36 8.855
R8157 CLK3.n27 CLK3.n26 8.855
R8158 CLK3.n38 CLK3.n27 8.855
R8159 CLK3.n41 CLK3.n40 8.855
R8160 CLK3.n40 CLK3.n39 8.855
R8161 CLK3.n24 CLK3.n23 8.855
R8162 CLK3.n23 CLK3.n22 8.855
R8163 CLK3.n47 CLK3.n46 8.855
R8164 CLK3.n48 CLK3.n47 8.855
R8165 CLK3.n21 CLK3.n20 8.855
R8166 CLK3.n49 CLK3.n21 8.855
R8167 CLK3.n53 CLK3.n52 8.855
R8168 CLK3.n52 CLK3.n51 8.855
R8169 CLK3.n17 CLK3.n16 8.855
R8170 CLK3.n50 CLK3.n16 8.855
R8171 CLK3.n58 CLK3.n57 8.855
R8172 CLK3.n59 CLK3.n58 8.855
R8173 CLK3.n15 CLK3.n14 8.855
R8174 CLK3.n60 CLK3.n15 8.855
R8175 CLK3.n63 CLK3.n62 8.855
R8176 CLK3.n62 CLK3.n61 8.855
R8177 CLK3.n12 CLK3.n11 8.855
R8178 CLK3.n11 CLK3.n10 8.855
R8179 CLK3.n69 CLK3.n68 8.855
R8180 CLK3.n70 CLK3.n69 8.855
R8181 CLK3.n9 CLK3.n8 8.855
R8182 CLK3.n71 CLK3.n9 8.855
R8183 CLK3.n74 CLK3.n73 8.855
R8184 CLK3.n73 CLK3.n72 8.855
R8185 CLK3.n5 CLK3.n4 8.855
R8186 CLK3.n4 CLK3.n3 8.855
R8187 CLK3.n413 CLK3.n412 8.855
R8188 CLK3.n2 CLK3.n1 8.855
R8189 CLK3.n339 CLK3.n115 8.365
R8190 CLK3.n50 CLK3.t24 8.189
R8191 CLK3.n60 CLK3.t18 8.189
R8192 CLK3.n368 CLK3.t43 8.189
R8193 CLK3.n376 CLK3.t32 8.189
R8194 CLK3.n301 CLK3.t36 8.189
R8195 CLK3.n293 CLK3.t16 8.189
R8196 CLK3.n222 CLK3.t45 8.189
R8197 CLK3.n230 CLK3.t30 8.189
R8198 CLK3.n393 CLK3.n86 6.776
R8199 CLK3.n247 CLK3.n165 6.776
R8200 CLK3.n276 CLK3.n150 6.776
R8201 CLK3.n77 CLK3.n6 6.776
R8202 CLK3.n333 CLK3.n332 6.754
R8203 EESPFAL_s3_0/CLK3 CLK3.n259 5.161
R8204 CLK3.n406 CLK3.n405 4.966
R8205 CLK3.n56 CLK3.n18 4.938
R8206 CLK3.n372 CLK3.n98 4.938
R8207 CLK3.n297 CLK3.n136 4.938
R8208 CLK3.n226 CLK3.n177 4.938
R8209 CLK3.n194 CLK3.n193 4.687
R8210 CLK3.n328 CLK3.n118 4.687
R8211 CLK3.n264 CLK3.n154 4.687
R8212 CLK3.n340 CLK3.n114 4.687
R8213 CLK3.n32 CLK3.n31 4.675
R8214 CLK3.n196 CLK3.n195 4.65
R8215 CLK3.n191 CLK3.n190 4.65
R8216 CLK3.n203 CLK3.n202 4.65
R8217 CLK3.n204 CLK3.n189 4.65
R8218 CLK3.n206 CLK3.n205 4.65
R8219 CLK3.n185 CLK3.n184 4.65
R8220 CLK3.n213 CLK3.n212 4.65
R8221 CLK3.n214 CLK3.n183 4.65
R8222 CLK3.n217 CLK3.n216 4.65
R8223 CLK3.n179 CLK3.n178 4.65
R8224 CLK3.n225 CLK3.n224 4.65
R8225 CLK3.n226 CLK3.n176 4.65
R8226 CLK3.n228 CLK3.n227 4.65
R8227 CLK3.n173 CLK3.n172 4.65
R8228 CLK3.n235 CLK3.n234 4.65
R8229 CLK3.n237 CLK3.n171 4.65
R8230 CLK3.n239 CLK3.n238 4.65
R8231 CLK3.n167 CLK3.n166 4.65
R8232 CLK3.n246 CLK3.n245 4.65
R8233 CLK3.n248 CLK3.n164 4.65
R8234 CLK3.n250 CLK3.n249 4.65
R8235 CLK3.n160 CLK3.n159 4.65
R8236 CLK3.n257 CLK3.n256 4.65
R8237 CLK3.n152 CLK3.n151 4.65
R8238 CLK3.n327 CLK3.n326 4.65
R8239 CLK3.n120 CLK3.n119 4.65
R8240 CLK3.n320 CLK3.n319 4.65
R8241 CLK3.n318 CLK3.n124 4.65
R8242 CLK3.n317 CLK3.n316 4.65
R8243 CLK3.n126 CLK3.n125 4.65
R8244 CLK3.n310 CLK3.n309 4.65
R8245 CLK3.n308 CLK3.n130 4.65
R8246 CLK3.n306 CLK3.n305 4.65
R8247 CLK3.n132 CLK3.n131 4.65
R8248 CLK3.n299 CLK3.n298 4.65
R8249 CLK3.n297 CLK3.n135 4.65
R8250 CLK3.n296 CLK3.n295 4.65
R8251 CLK3.n138 CLK3.n137 4.65
R8252 CLK3.n289 CLK3.n288 4.65
R8253 CLK3.n286 CLK3.n143 4.65
R8254 CLK3.n285 CLK3.n284 4.65
R8255 CLK3.n145 CLK3.n144 4.65
R8256 CLK3.n278 CLK3.n277 4.65
R8257 CLK3.n275 CLK3.n149 4.65
R8258 CLK3.n274 CLK3.n273 4.65
R8259 CLK3.n117 CLK3.n116 4.65
R8260 CLK3.n330 CLK3.n329 4.65
R8261 CLK3.n338 CLK3.n337 4.65
R8262 CLK3.n342 CLK3.n341 4.65
R8263 CLK3.n112 CLK3.n111 4.65
R8264 CLK3.n349 CLK3.n348 4.65
R8265 CLK3.n350 CLK3.n110 4.65
R8266 CLK3.n352 CLK3.n351 4.65
R8267 CLK3.n106 CLK3.n105 4.65
R8268 CLK3.n359 CLK3.n358 4.65
R8269 CLK3.n360 CLK3.n104 4.65
R8270 CLK3.n363 CLK3.n362 4.65
R8271 CLK3.n100 CLK3.n99 4.65
R8272 CLK3.n371 CLK3.n370 4.65
R8273 CLK3.n372 CLK3.n97 4.65
R8274 CLK3.n374 CLK3.n373 4.65
R8275 CLK3.n94 CLK3.n93 4.65
R8276 CLK3.n381 CLK3.n380 4.65
R8277 CLK3.n383 CLK3.n92 4.65
R8278 CLK3.n385 CLK3.n384 4.65
R8279 CLK3.n88 CLK3.n87 4.65
R8280 CLK3.n392 CLK3.n391 4.65
R8281 CLK3.n394 CLK3.n85 4.65
R8282 CLK3.n396 CLK3.n395 4.65
R8283 CLK3.n81 CLK3.n80 4.65
R8284 CLK3.n403 CLK3.n402 4.65
R8285 CLK3.n411 CLK3.n410 4.65
R8286 CLK3.n33 CLK3.n30 4.65
R8287 CLK3.n35 CLK3.n34 4.65
R8288 CLK3.n26 CLK3.n25 4.65
R8289 CLK3.n42 CLK3.n41 4.65
R8290 CLK3.n43 CLK3.n24 4.65
R8291 CLK3.n46 CLK3.n45 4.65
R8292 CLK3.n20 CLK3.n19 4.65
R8293 CLK3.n54 CLK3.n53 4.65
R8294 CLK3.n55 CLK3.n17 4.65
R8295 CLK3.n57 CLK3.n56 4.65
R8296 CLK3.n14 CLK3.n13 4.65
R8297 CLK3.n64 CLK3.n63 4.65
R8298 CLK3.n65 CLK3.n12 4.65
R8299 CLK3.n68 CLK3.n67 4.65
R8300 CLK3.n8 CLK3.n7 4.65
R8301 CLK3.n75 CLK3.n74 4.65
R8302 CLK3.n76 CLK3.n5 4.65
R8303 CLK3.n416 CLK3.n415 4.65
R8304 CLK3.n262 CLK3.n261 4.5
R8305 CLK3.n263 CLK3.n262 4.5
R8306 CLK3.n263 CLK3.n155 4.5
R8307 CLK3.n408 CLK3.n0 4.5
R8308 CLK3.n409 CLK3.n408 4.5
R8309 CLK3.n260 EESPFAL_s2_0/CLK3 4.449
R8310 CLK3.n334 CLK3.n333 3.724
R8311 CLK3.n332 CLK3.n117 3.715
R8312 CLK3.n337 CLK3.n115 3.715
R8313 CLK3.n336 CLK3.n334 3.039
R8314 CLK3.n259 CLK3.n158 3.038
R8315 CLK3.n405 CLK3.n79 3.038
R8316 CLK3.n78 CLK3.n1 3.033
R8317 CLK3.n332 CLK3.n331 2.57
R8318 CLK3.n335 CLK3.n115 2.57
R8319 CLK3.n267 CLK3.n156 2.24
R8320 CLK3.n329 CLK3.n328 2.203
R8321 CLK3.n340 CLK3.n339 2.203
R8322 CLK3.n255 CLK3.n254 1.655
R8323 CLK3.n325 CLK3.n324 1.655
R8324 CLK3.n401 CLK3.n400 1.655
R8325 CLK3.n29 CLK3.n28 1.655
R8326 CLK3.n344 CLK3.n343 1.655
R8327 CLK3.n198 CLK3.n197 1.655
R8328 CLK3.n269 CLK3.n268 1.655
R8329 CLK3.n414 CLK3.n2 1.655
R8330 CLK3.n260 CLK3.n157 1.497
R8331 CLK3.n407 CLK3.n78 1.121
R8332 EESPFAL_s2_0/CLK3 EESPFAL_s3_0/CLK3 1.018
R8333 CLK3.n267 CLK3.n155 0.48
R8334 CLK3.n406 EESPFAL_s1_0/CLK3 0.195
R8335 CLK3.n329 CLK3.n116 0.125
R8336 CLK3.n339 CLK3.n338 0.125
R8337 CLK3.n333 CLK3.n116 0.119
R8338 CLK3.n338 CLK3.n334 0.119
R8339 CLK3.n195 CLK3.n190 0.1
R8340 CLK3.n203 CLK3.n190 0.1
R8341 CLK3.n204 CLK3.n203 0.1
R8342 CLK3.n205 CLK3.n204 0.1
R8343 CLK3.n205 CLK3.n184 0.1
R8344 CLK3.n213 CLK3.n184 0.1
R8345 CLK3.n214 CLK3.n213 0.1
R8346 CLK3.n216 CLK3.n178 0.1
R8347 CLK3.n225 CLK3.n178 0.1
R8348 CLK3.n226 CLK3.n225 0.1
R8349 CLK3.n227 CLK3.n172 0.1
R8350 CLK3.n235 CLK3.n172 0.1
R8351 CLK3.n238 CLK3.n237 0.1
R8352 CLK3.n238 CLK3.n166 0.1
R8353 CLK3.n246 CLK3.n166 0.1
R8354 CLK3.n249 CLK3.n248 0.1
R8355 CLK3.n249 CLK3.n159 0.1
R8356 CLK3.n257 CLK3.n159 0.1
R8357 CLK3.n327 CLK3.n119 0.1
R8358 CLK3.n319 CLK3.n119 0.1
R8359 CLK3.n319 CLK3.n318 0.1
R8360 CLK3.n318 CLK3.n317 0.1
R8361 CLK3.n317 CLK3.n125 0.1
R8362 CLK3.n309 CLK3.n125 0.1
R8363 CLK3.n309 CLK3.n308 0.1
R8364 CLK3.n306 CLK3.n131 0.1
R8365 CLK3.n298 CLK3.n131 0.1
R8366 CLK3.n298 CLK3.n297 0.1
R8367 CLK3.n296 CLK3.n137 0.1
R8368 CLK3.n288 CLK3.n137 0.1
R8369 CLK3.n286 CLK3.n285 0.1
R8370 CLK3.n285 CLK3.n144 0.1
R8371 CLK3.n277 CLK3.n144 0.1
R8372 CLK3.n275 CLK3.n274 0.1
R8373 CLK3.n274 CLK3.n151 0.1
R8374 CLK3.n341 CLK3.n111 0.1
R8375 CLK3.n349 CLK3.n111 0.1
R8376 CLK3.n350 CLK3.n349 0.1
R8377 CLK3.n351 CLK3.n350 0.1
R8378 CLK3.n351 CLK3.n105 0.1
R8379 CLK3.n359 CLK3.n105 0.1
R8380 CLK3.n360 CLK3.n359 0.1
R8381 CLK3.n362 CLK3.n99 0.1
R8382 CLK3.n371 CLK3.n99 0.1
R8383 CLK3.n372 CLK3.n371 0.1
R8384 CLK3.n373 CLK3.n93 0.1
R8385 CLK3.n381 CLK3.n93 0.1
R8386 CLK3.n384 CLK3.n383 0.1
R8387 CLK3.n384 CLK3.n87 0.1
R8388 CLK3.n392 CLK3.n87 0.1
R8389 CLK3.n395 CLK3.n394 0.1
R8390 CLK3.n395 CLK3.n80 0.1
R8391 CLK3.n403 CLK3.n80 0.1
R8392 CLK3.n34 CLK3.n33 0.1
R8393 CLK3.n34 CLK3.n25 0.1
R8394 CLK3.n42 CLK3.n25 0.1
R8395 CLK3.n43 CLK3.n42 0.1
R8396 CLK3.n45 CLK3.n43 0.1
R8397 CLK3.n54 CLK3.n19 0.1
R8398 CLK3.n55 CLK3.n54 0.1
R8399 CLK3.n56 CLK3.n55 0.1
R8400 CLK3.n64 CLK3.n13 0.1
R8401 CLK3.n65 CLK3.n64 0.1
R8402 CLK3.n67 CLK3.n7 0.1
R8403 CLK3.n75 CLK3.n7 0.1
R8404 CLK3.n76 CLK3.n75 0.1
R8405 EESPFAL_s0_0/CLK3 CLK3 0.1
R8406 CLK3.n247 CLK3.n246 0.087
R8407 CLK3.n277 CLK3.n276 0.087
R8408 CLK3.n393 CLK3.n392 0.087
R8409 CLK3.n77 CLK3.n76 0.087
R8410 CLK3.n216 CLK3.n215 0.075
R8411 CLK3.n227 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/CLK 0.075
R8412 CLK3.n236 CLK3.n235 0.075
R8413 CLK3.n307 CLK3.n306 0.075
R8414 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/CLK CLK3.n296 0.075
R8415 CLK3.n288 CLK3.n287 0.075
R8416 CLK3.n362 CLK3.n361 0.075
R8417 CLK3.n373 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/CLK 0.075
R8418 CLK3.n382 CLK3.n381 0.075
R8419 CLK3.n33 CLK3.n32 0.075
R8420 CLK3.n44 CLK3.n19 0.075
R8421 CLK3 CLK3.n13 0.075
R8422 CLK3.n66 CLK3.n65 0.075
R8423 CLK3.n410 CLK3.n409 0.073
R8424 CLK3.n416 CLK3.n0 0.072
R8425 CLK3.n261 CLK3.n151 0.063
R8426 CLK3.n195 CLK3.n194 0.062
R8427 CLK3.n258 CLK3.n257 0.062
R8428 CLK3.n328 CLK3.n327 0.062
R8429 CLK3.n341 CLK3.n340 0.062
R8430 CLK3.n404 CLK3.n403 0.062
R8431 CLK3.n265 CLK3.n264 0.045
R8432 CLK3.n259 CLK3.n258 0.034
R8433 CLK3.n405 CLK3.n404 0.034
R8434 CLK3.n78 CLK3.n0 0.027
R8435 CLK3.n409 CLK3.n78 0.026
R8436 CLK3.n215 CLK3.n214 0.025
R8437 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/CLK CLK3.n226 0.025
R8438 CLK3.n237 CLK3.n236 0.025
R8439 CLK3.n308 CLK3.n307 0.025
R8440 CLK3.n297 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/CLK 0.025
R8441 CLK3.n287 CLK3.n286 0.025
R8442 CLK3.n361 CLK3.n360 0.025
R8443 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/CLK CLK3.n372 0.025
R8444 CLK3.n383 CLK3.n382 0.025
R8445 CLK3.n45 CLK3.n44 0.025
R8446 CLK3.n56 CLK3 0.025
R8447 CLK3.n67 CLK3.n66 0.025
R8448 CLK3.n266 CLK3.n265 0.017
R8449 CLK3.n261 CLK3.n157 0.016
R8450 CLK3.n263 CLK3.n157 0.016
R8451 CLK3.n262 CLK3.n260 0.012
R8452 CLK3.n248 CLK3.n247 0.012
R8453 CLK3.n276 CLK3.n275 0.012
R8454 CLK3.n394 CLK3.n393 0.012
R8455 CLK3.n410 CLK3.n77 0.012
R8456 CLK3.n408 CLK3.n407 0.01
R8457 CLK3.n266 CLK3.n263 0.003
R8458 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t6 1074.82
R8459 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t7 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t8 819.4
R8460 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t7 514.133
R8461 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t9 305.266
R8462 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n6 260.333
R8463 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n5 192
R8464 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n3 166.736
R8465 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n5 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n4 105.6
R8466 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t0 97.937
R8467 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n5 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t1 97.937
R8468 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n1 76
R8469 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n0 73.937
R8470 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n2 57.6
R8471 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t4 39.4
R8472 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t3 39.4
R8473 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n0 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t5 24
R8474 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n0 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t2 24
R8475 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n2 EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT 3.2
R8476 x1_bar.n4 x1_bar.t2 1069.04
R8477 x1_bar.n3 x1_bar.t5 1069.04
R8478 x1_bar.n2 x1_bar.t7 1069.04
R8479 x1_bar.n4 x1_bar.t10 1015.9
R8480 x1_bar.n3 x1_bar.t6 1015.9
R8481 x1_bar.n2 x1_bar.t0 1015.9
R8482 EESPFAL_s2_0/EESPFAL_4in_NAND_0/B_bar x1_bar.t4 912.566
R8483 EESPFAL_s0_0/EESPFAL_NAND_v3_2/B x1_bar.t1 881.55
R8484 EESPFAL_s2_0/EESPFAL_INV4_1/A x1_bar.t9 778.1
R8485 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B_bar x1_bar.t3 604.112
R8486 x1_bar x1_bar.t8 479.166
R8487 EESPFAL_s3_0/EESPFAL_INV4_1/A_bar x1_bar.t11 392.5
R8488 x1_bar.n1 EESPFAL_s0_0/EESPFAL_NAND_v3_2/B 301.61
R8489 x1_bar.n9 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B_bar 253.93
R8490 x1_bar.n7 EESPFAL_s2_0/EESPFAL_XOR_v3_1/A_bar 218.41
R8491 x1_bar.n8 EESPFAL_s2_0/EESPFAL_4in_NAND_0/B_bar 218.41
R8492 x1_bar.n5 EESPFAL_s3_0/EESPFAL_XOR_v3_0/A_bar 205.61
R8493 x1_bar.n10 EESPFAL_s1_0/EESPFAL_XOR_v3_1/A_bar 205.61
R8494 EESPFAL_s3_0/x1_bar EESPFAL_s3_0/EESPFAL_INV4_1/A_bar 184.875
R8495 EESPFAL_s3_0/EESPFAL_XOR_v3_0/A_bar x1_bar.n4 89.6
R8496 EESPFAL_s2_0/EESPFAL_XOR_v3_1/A_bar x1_bar.n3 89.6
R8497 EESPFAL_s1_0/EESPFAL_XOR_v3_1/A_bar x1_bar.n2 89.6
R8498 x1_bar.n6 EESPFAL_s2_0/EESPFAL_INV4_1/A 41.24
R8499 x1_bar.n0 x1_bar 23.191
R8500 x1_bar.n7 EESPFAL_s2_0/x1_bar 3.048
R8501 EESPFAL_s1_0/x1_bar x1_bar.n10 2.945
R8502 x1_bar.n9 x1_bar.n8 2.5
R8503 x1_bar.n10 x1_bar.n9 1.843
R8504 x1_bar.n1 x1_bar.n0 1.654
R8505 EESPFAL_s1_0/x1_bar x1_bar.n1 1.648
R8506 x1_bar.n8 x1_bar.n7 1.617
R8507 x1_bar.n6 x1_bar.n5 1.276
R8508 x1_bar.n0 EESPFAL_s0_0/x1_bar 1.104
R8509 EESPFAL_s2_0/x1_bar x1_bar.n6 0.09
R8510 x1_bar.n5 EESPFAL_s3_0/x1_bar 0.023
R8511 s2_bar.t5 s2_bar.t6 819.4
R8512 s2_bar.n4 s2_bar.t7 506.1
R8513 s2_bar.n4 s2_bar.t5 313.3
R8514 s2_bar.n1 s2_bar.t1 181.136
R8515 s2_bar.n3 s2_bar.n2 128.334
R8516 s2_bar.n1 s2_bar.n0 57.937
R8517 s2_bar.n5 s2_bar.n3 57.6
R8518 s2_bar.n3 s2_bar.n1 41.6
R8519 s2_bar.n2 s2_bar.t3 39.4
R8520 s2_bar.n2 s2_bar.t4 39.4
R8521 s2_bar.n0 s2_bar.t0 24
R8522 s2_bar.n0 s2_bar.t2 24
R8523 s2_bar.n5 s2_bar.n4 8.764
R8524 s2_bar s2_bar.n5 4.681
R8525 EESPFAL_s2_0/s2_bar s2_bar 0.065
R8526 s2.t7 s2.t9 819.4
R8527 s2.n3 s2.t7 514.133
R8528 s2.n3 s2.t8 305.266
R8529 s2.n4 s2.n2 166.734
R8530 s2.n5 s2.n4 105.6
R8531 s2.n5 s2.t5 97.937
R8532 s2.n6 s2.n5 96
R8533 s2 s2.n6 83.731
R8534 s2 s2.n3 79.2
R8535 s2.n4 s2.n1 73.937
R8536 s2.n6 s2.n0 73.937
R8537 s2.n4 s2 54.4
R8538 s2.n2 s2.t3 39.4
R8539 s2.n2 s2.t2 39.4
R8540 s2.n1 s2.t1 24
R8541 s2.n1 s2.t4 24
R8542 s2.n0 s2.t6 24
R8543 s2.n0 s2.t0 24
R8544 EESPFAL_s2_0/s2 s2 0.081
R8545 s1.t9 s1.t7 819.4
R8546 s1.n3 s1.t9 514.133
R8547 s1.n3 s1.t8 305.266
R8548 s1.n4 s1.n1 166.734
R8549 s1.n5 s1.n4 105.6
R8550 s1.n5 s1.t3 97.937
R8551 s1.n6 s1.n5 96
R8552 s1 s1.n6 83.588
R8553 s1 s1.n3 79.2
R8554 s1.n4 s1.n2 73.937
R8555 s1.n6 s1.n0 73.937
R8556 s1.n4 s1 54.4
R8557 s1.n1 s1.t5 39.4
R8558 s1.n1 s1.t6 39.4
R8559 s1.n2 s1.t1 24
R8560 s1.n2 s1.t4 24
R8561 s1.n0 s1.t2 24
R8562 s1.n0 s1.t0 24
R8563 EESPFAL_s1_0/s1 s1 0.096
R8564 s1_bar.t6 s1_bar.t7 819.4
R8565 s1_bar.n4 s1_bar.t5 506.1
R8566 s1_bar.n4 s1_bar.t6 313.3
R8567 s1_bar.n2 s1_bar.t4 181.136
R8568 s1_bar.n3 s1_bar.n0 128.334
R8569 s1_bar.n2 s1_bar.n1 57.937
R8570 s1_bar.n5 s1_bar.n3 57.6
R8571 s1_bar.n3 s1_bar.n2 41.6
R8572 s1_bar.n0 s1_bar.t3 39.4
R8573 s1_bar.n0 s1_bar.t2 39.4
R8574 s1_bar.n1 s1_bar.t0 24
R8575 s1_bar.n1 s1_bar.t1 24
R8576 s1_bar.n5 s1_bar.n4 8.764
R8577 s1_bar s1_bar.n5 4.681
R8578 EESPFAL_s1_0/s1_bar s1_bar 0.103
R8579 x3.n4 x3.t7 1176.57
R8580 x3.n4 x3.t10 1149.49
R8581 EESPFAL_s2_0/EESPFAL_4in_NAND_0/A_bar x3.t3 1121.23
R8582 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C x3.t5 904.039
R8583 x3.n0 x3.t1 800.452
R8584 x3.n5 x3.t4 800.452
R8585 x3.n3 x3.t0 800.452
R8586 x3.n0 x3.t2 787.997
R8587 x3.n5 x3.t6 787.997
R8588 x3.n3 x3.t9 787.997
R8589 EESPFAL_s1_0/EESPFAL_INV4_2/A x3.t12 778.1
R8590 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A_bar x3.t11 696.166
R8591 EESPFAL_s3_0/EESPFAL_INV4_2/A_bar x3.t8 392.5
R8592 x3.n7 EESPFAL_s3_0/EESPFAL_INV4_2/A_bar 179.729
R8593 x3 x3.n0 169.6
R8594 EESPFAL_s3_0/EESPFAL_XOR_v3_1/B x3.n5 169.6
R8595 EESPFAL_s1_0/EESPFAL_XOR_v3_1/B x3.n3 169.6
R8596 x3.n6 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C 146.249
R8597 x3.n10 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A_bar 144.49
R8598 EESPFAL_s2_0/EESPFAL_XOR_v3_0/A x3.n4 128
R8599 x3.n8 EESPFAL_s2_0/EESPFAL_XOR_v3_0/A 108.97
R8600 x3.n9 EESPFAL_s2_0/EESPFAL_4in_NAND_0/A_bar 108.97
R8601 x3.n1 x3 96.17
R8602 x3.n6 EESPFAL_s3_0/EESPFAL_XOR_v3_1/B 96.17
R8603 x3.n11 EESPFAL_s1_0/EESPFAL_XOR_v3_1/B 96.17
R8604 x3.n2 EESPFAL_s1_0/EESPFAL_INV4_2/A 40.925
R8605 x3.n9 x3.n8 4.595
R8606 x3.n2 x3.n1 4.057
R8607 EESPFAL_s1_0/x3 x3.n11 2.854
R8608 x3.n10 x3.n9 2.74
R8609 x3.n11 x3.n10 1.915
R8610 x3.n7 x3.n6 1.878
R8611 EESPFAL_s2_0/x3 EESPFAL_s3_0/x3 1.196
R8612 EESPFAL_s3_0/x3 x3.n7 1.007
R8613 x3.n1 EESPFAL_s0_0/x3 0.262
R8614 EESPFAL_s1_0/x3 x3.n2 0.087
R8615 x3.n8 EESPFAL_s2_0/x3 0.042
R8616 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t9 1074.82
R8617 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t6 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t7 819.4
R8618 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t6 514.133
R8619 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t8 305.266
R8620 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n6 260.333
R8621 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n6 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n5 192
R8622 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n1 166.734
R8623 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n5 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n4 105.6
R8624 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n6 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t0 97.937
R8625 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n5 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t4 97.937
R8626 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n2 76
R8627 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n0 73.937
R8628 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n3 57.6
R8629 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t3 39.4
R8630 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t2 39.4
R8631 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n0 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t5 24
R8632 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n0 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t1 24
R8633 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n3 EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT 3.2
R8634 Dis3 Dis3.t4 392.5
R8635 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/Dis Dis3.t7 392.5
R8636 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/Dis Dis3.t1 392.5
R8637 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/Dis Dis3.t2 392.5
R8638 Dis3.n0 Dis3.t0 389.3
R8639 Dis3.n5 Dis3.t3 389.3
R8640 Dis3.n3 Dis3.t6 389.3
R8641 Dis3.n1 Dis3.t5 389.3
R8642 EESPFAL_s3_0/Dis3 Dis3.n1 297.172
R8643 Dis3.n6 Dis3.n5 285.061
R8644 Dis3.n4 Dis3.n3 284.736
R8645 Dis3.n0 Dis3 112
R8646 Dis3.n5 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/Dis 112
R8647 Dis3.n3 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/Dis 112
R8648 Dis3.n1 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/Dis 112
R8649 Dis3.n7 Dis3.n0 98.399
R8650 Dis3.n4 Dis3.n2 12.126
R8651 EESPFAL_s1_0/Dis3 Dis3.n6 12.061
R8652 Dis3.n7 EESPFAL_s1_0/Dis3 8.969
R8653 Dis3 Dis3.n7 4.678
R8654 EESPFAL_s2_0/Dis3 EESPFAL_s3_0/Dis3 1.73
R8655 Dis3.n6 Dis3.n4 1.496
R8656 EESPFAL_s0_0/Dis3 Dis3 0.106
R8657 Dis3.n2 EESPFAL_s2_0/Dis3 0.043
R8658 Dis3.n2 EESPFAL_s2_0/Dis3 0.031
R8659 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t9 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t6 819.4
R8660 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t7 736.033
R8661 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t9 514.133
R8662 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t8 305.266
R8663 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n5 192
R8664 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n0 166.734
R8665 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n4 105.6
R8666 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t2 97.937
R8667 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t5 97.937
R8668 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n1 76
R8669 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n3 73.939
R8670 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n2 57.6
R8671 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n6 56.157
R8672 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t0 39.4
R8673 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t3 39.4
R8674 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t4 24
R8675 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t1 24
R8676 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT 3.2
R8677 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t9 1074.82
R8678 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t8 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t6 819.4
R8679 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t7 506.1
R8680 EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 442.013
R8681 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t8 313.3
R8682 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t0 273.936
R8683 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n3 128.335
R8684 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n1 105.6
R8685 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t2 81.937
R8686 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n0 57.937
R8687 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n4 57.6
R8688 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n2 41.6
R8689 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t4 39.4
R8690 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t5 39.4
R8691 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t3 24
R8692 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t1 24
R8693 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n5 8.764
R8694 EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n6 4.65
R8695 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 819.4
R8696 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 506.1
R8697 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 313.3
R8698 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 305.997
R8699 EESPFAL_s3_0/EESPFAL_INV4_0/OUT EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 206.179
R8700 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 187.536
R8701 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 128.334
R8702 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 115.2
R8703 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 57.939
R8704 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 57.6
R8705 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 41.6
R8706 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 39.4
R8707 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 39.4
R8708 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 24
R8709 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 24
R8710 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 8.764
R8711 EESPFAL_s3_0/EESPFAL_INV4_0/OUT EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 4.65
R8712 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t5 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t6 819.4
R8713 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t8 775.706
R8714 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t5 514.133
R8715 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t7 305.266
R8716 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n4 166.735
R8717 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 163.511
R8718 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n2 102.4
R8719 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n1 88.255
R8720 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t4 81.937
R8721 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n6 76
R8722 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n5 57.6
R8723 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n0 51.537
R8724 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t3 39.4
R8725 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t2 39.4
R8726 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t0 24
R8727 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t1 24
R8728 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n3 6.4
R8729 EESPFAL_s3_0/EESPFAL_INV4_0/OUT_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n7 3.2
R8730 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t6 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t9 819.4
R8731 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t7 736.033
R8732 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t8 506.1
R8733 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t6 313.3
R8734 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t1 273.936
R8735 EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 266.318
R8736 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n3 128.336
R8737 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n1 105.6
R8738 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t0 81.937
R8739 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n0 57.937
R8740 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n4 57.6
R8741 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n2 41.6
R8742 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t4 39.4
R8743 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t3 39.4
R8744 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t2 24
R8745 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t5 24
R8746 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n5 8.764
R8747 EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n6 4.65
R8748 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/A_bar 922.56
R8749 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t8 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t9 819.4
R8750 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t7 684.833
R8751 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t6 506.1
R8752 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n5 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t8 313.3
R8753 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t4 177.936
R8754 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n3 128.335
R8755 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n1 105.6
R8756 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t5 81.937
R8757 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n0 58.265
R8758 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n4 57.6
R8759 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n2 41.6
R8760 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t2 39.4
R8761 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t1 39.4
R8762 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t0 24
R8763 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t3 24
R8764 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n5 8.764
R8765 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n6 4.65
R8766 x0_bar.n0 x0_bar.t9 1069.04
R8767 x0_bar.n0 x0_bar.t10 1015.9
R8768 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C x0_bar.t7 904.039
R8769 x0_bar.n4 x0_bar.t3 810.772
R8770 x0_bar.n3 x0_bar.t5 810.772
R8771 x0_bar.n2 x0_bar.t1 810.772
R8772 EESPFAL_s2_0/EESPFAL_4in_NAND_0/C_bar x0_bar.t4 703.9
R8773 x0_bar.n4 x0_bar.t0 694.566
R8774 x0_bar.n3 x0_bar.t2 694.566
R8775 x0_bar.n2 x0_bar.t6 694.566
R8776 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B_bar x0_bar.t8 604.112
R8777 x0_bar.n5 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B_bar 331.421
R8778 x0_bar.n8 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C 321.619
R8779 x0_bar.n6 EESPFAL_s2_0/EESPFAL_XOR_v3_1/B_bar 291.37
R8780 x0_bar.n7 EESPFAL_s2_0/EESPFAL_4in_NAND_0/C_bar 291.37
R8781 x0_bar.n1 x0_bar 278.57
R8782 x0_bar.n5 EESPFAL_s3_0/EESPFAL_XOR_v3_0/B_bar 278.57
R8783 x0_bar.n9 EESPFAL_s1_0/EESPFAL_XOR_v3_0/B_bar 278.57
R8784 x0_bar x0_bar.n0 89.6
R8785 EESPFAL_s3_0/EESPFAL_XOR_v3_0/B_bar x0_bar.n4 25.6
R8786 EESPFAL_s2_0/EESPFAL_XOR_v3_1/B_bar x0_bar.n3 25.6
R8787 EESPFAL_s1_0/EESPFAL_XOR_v3_0/B_bar x0_bar.n2 25.6
R8788 EESPFAL_s1_0/x0_bar x0_bar.n1 4.398
R8789 x0_bar.n9 x0_bar.n8 4.206
R8790 x0_bar.n6 EESPFAL_s2_0/x0_bar 2.695
R8791 x0_bar.n8 x0_bar.n7 2.604
R8792 x0_bar.n7 x0_bar.n6 2.126
R8793 EESPFAL_s2_0/x0_bar EESPFAL_s3_0/x0_bar 1.39
R8794 EESPFAL_s1_0/x0_bar x0_bar.n9 0.321
R8795 EESPFAL_s3_0/x0_bar x0_bar.n5 0.289
R8796 x0_bar.n1 EESPFAL_s0_0/x0_bar 0.009
R8797 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t8 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t9 819.4
R8798 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t6 736.033
R8799 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t8 514.133
R8800 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t7 305.266
R8801 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n5 192
R8802 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n1 166.734
R8803 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n6 160.887
R8804 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n4 105.6
R8805 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t0 97.937
R8806 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t1 97.937
R8807 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n2 76
R8808 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n0 73.937
R8809 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n3 57.6
R8810 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t5 39.4
R8811 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t3 39.4
R8812 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t4 24
R8813 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t2 24
R8814 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT 3.2
R8815 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n0 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t9 1071.3
R8816 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t7 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t8 819.4
R8817 EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 526.35
R8818 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n6 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t6 506.1
R8819 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n6 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t7 313.3
R8820 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t4 273.936
R8821 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n5 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n4 128.336
R8822 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n3 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n2 105.6
R8823 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t0 81.937
R8824 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n3 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n1 57.937
R8825 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n7 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n5 57.6
R8826 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n5 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n3 41.6
R8827 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t3 39.4
R8828 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n4 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t2 39.4
R8829 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n1 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t1 24
R8830 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n1 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t5 24
R8831 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n7 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n6 8.764
R8832 EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n7 4.65
R8833 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n0 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 3.52
R8834 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n0 2.607
R8835 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A x2_bar.t7 1271.5
R8836 x2_bar.n2 x2_bar.t11 1069.04
R8837 x2_bar.n5 x2_bar.t10 1069.04
R8838 x2_bar.n2 x2_bar.t4 1015.9
R8839 x2_bar.n5 x2_bar.t5 1015.9
R8840 x2_bar x2_bar.t0 833.352
R8841 x2_bar.n4 x2_bar.t1 810.772
R8842 EESPFAL_s2_0/EESPFAL_INV4_0/A x2_bar.t2 778.1
R8843 EESPFAL_s0_0/EESPFAL_NAND_v3_2/A_bar x2_bar.t6 736.033
R8844 x2_bar.n4 x2_bar.t8 694.566
R8845 EESPFAL_s2_0/EESPFAL_4in_NAND_0/D_bar x2_bar.t3 495.233
R8846 EESPFAL_s1_0/EESPFAL_INV4_1/A_bar x2_bar.t9 392.5
R8847 x2_bar.n1 EESPFAL_s0_0/EESPFAL_NAND_v3_2/A_bar 228.65
R8848 x2_bar.n10 EESPFAL_s1_0/EESPFAL_INV4_1/A_bar 182.7
R8849 x2_bar.n6 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A 182.235
R8850 x2_bar.n7 EESPFAL_s2_0/EESPFAL_XOR_v3_0/B_bar 145.45
R8851 x2_bar.n9 EESPFAL_s2_0/EESPFAL_4in_NAND_0/D_bar 145.45
R8852 x2_bar.n3 EESPFAL_s1_0/EESPFAL_XOR_v3_0/A_bar 132.65
R8853 x2_bar.n6 EESPFAL_s3_0/EESPFAL_XOR_v3_1/A_bar 132.65
R8854 EESPFAL_s1_0/EESPFAL_XOR_v3_0/A_bar x2_bar.n2 89.6
R8855 EESPFAL_s3_0/EESPFAL_XOR_v3_1/A_bar x2_bar.n5 89.6
R8856 x2_bar.n8 EESPFAL_s2_0/EESPFAL_INV4_0/A 41.057
R8857 EESPFAL_s2_0/EESPFAL_XOR_v3_0/B_bar x2_bar.n4 25.6
R8858 x2_bar.n0 x2_bar 22.325
R8859 x2_bar.n10 x2_bar.n9 4.913
R8860 EESPFAL_s3_0/x2_bar x2_bar.n6 2.946
R8861 x2_bar.n8 x2_bar.n7 2.782
R8862 x2_bar.n1 x2_bar.n0 2.568
R8863 EESPFAL_s1_0/x2_bar x2_bar.n10 1.998
R8864 x2_bar.n9 x2_bar.n8 1.843
R8865 x2_bar.n3 x2_bar.n1 1.79
R8866 EESPFAL_s2_0/x2_bar EESPFAL_s3_0/x2_bar 1.387
R8867 x2_bar.n7 EESPFAL_s2_0/x2_bar 0.415
R8868 x2_bar.n0 EESPFAL_s0_0/x2_bar 0.026
R8869 EESPFAL_s1_0/x2_bar x2_bar.n3 0.021
R8870 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t8 1074.82
R8871 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t6 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t7 819.4
R8872 EESPFAL_s0_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t10 736.033
R8873 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t6 514.133
R8874 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n2 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t9 305.266
R8875 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n5 192
R8876 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n0 166.734
R8877 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n4 105.6
R8878 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n6 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t0 97.939
R8879 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n5 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t2 97.937
R8880 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n7 76.565
R8881 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n2 76
R8882 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n1 73.937
R8883 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n3 57.6
R8884 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t1 39.4
R8885 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n0 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t3 39.4
R8886 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n7 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n6 25.6
R8887 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t5 24
R8888 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n1 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t4 24
R8889 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n7 EESPFAL_s0_0/EESPFAL_NAND_v3_1/A_bar 21.729
R8890 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n3 EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT 3.2
R8891 EESPFAL_s0_0/EESPFAL_NAND_v3_1/A EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t7 1074.82
R8892 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t6 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t8 819.4
R8893 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t9 736.033
R8894 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t10 506.1
R8895 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n6 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t6 313.3
R8896 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t1 273.936
R8897 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_s0_0/EESPFAL_NAND_v3_1/A 180.175
R8898 EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n0 161.141
R8899 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n4 128.335
R8900 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n2 105.6
R8901 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n2 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t0 81.937
R8902 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n7 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n5 64
R8903 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n3 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n1 57.937
R8904 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n5 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n3 41.6
R8905 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t5 39.4
R8906 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n4 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t4 39.4
R8907 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n0 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 24.135
R8908 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t3 24
R8909 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n1 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t2 24
R8910 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n7 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n6 8.764
R8911 EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n7 4.65
R8912 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t6 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t5 819.4
R8913 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t8 775.706
R8914 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t6 514.133
R8915 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t7 305.266
R8916 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n0 166.734
R8917 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 163.511
R8918 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n2 102.4
R8919 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n1 88.292
R8920 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t3 81.937
R8921 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n6 76
R8922 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n5 57.6
R8923 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n3 51.537
R8924 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t4 39.4
R8925 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t2 39.4
R8926 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t0 24
R8927 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t1 24
R8928 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n4 6.4
R8929 EESPFAL_s2_0/EESPFAL_INV4_2/OUT_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n7 3.2
R8930 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 819.4
R8931 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 506.1
R8932 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 313.3
R8933 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 305.997
R8934 EESPFAL_s2_0/EESPFAL_INV4_2/OUT EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 210.945
R8935 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 187.536
R8936 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 128.336
R8937 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 115.2
R8938 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 57.937
R8939 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 57.6
R8940 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 41.6
R8941 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 39.4
R8942 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 39.4
R8943 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 24
R8944 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 24
R8945 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 8.764
R8946 EESPFAL_s2_0/EESPFAL_INV4_2/OUT EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 4.65
R8947 s3.t7 s3.t8 819.4
R8948 s3.n3 s3.t7 514.133
R8949 s3.n3 s3.t9 305.266
R8950 s3.n4 s3.n1 166.734
R8951 s3.n5 s3.n4 105.6
R8952 s3.n5 s3.t4 97.937
R8953 s3.n6 s3.n5 96
R8954 s3 s3.n6 83.597
R8955 s3 s3.n3 79.2
R8956 s3.n4 s3.n2 73.937
R8957 s3.n6 s3.n0 73.937
R8958 s3.n4 s3 54.4
R8959 s3.n1 s3.t5 39.4
R8960 s3.n1 s3.t1 39.4
R8961 s3.n2 s3.t0 24
R8962 s3.n2 s3.t3 24
R8963 s3.n0 s3.t2 24
R8964 s3.n0 s3.t6 24
R8965 EESPFAL_s3_0/s3 s3 0.087
R8966 s3_bar.t7 s3_bar.t5 819.4
R8967 s3_bar.n4 s3_bar.t6 506.1
R8968 s3_bar.n4 s3_bar.t7 313.3
R8969 s3_bar.n2 s3_bar.t4 181.136
R8970 s3_bar.n3 s3_bar.n0 128.334
R8971 s3_bar.n2 s3_bar.n1 57.937
R8972 s3_bar.n5 s3_bar.n3 57.6
R8973 s3_bar.n3 s3_bar.n2 41.6
R8974 s3_bar.n0 s3_bar.t2 39.4
R8975 s3_bar.n0 s3_bar.t3 39.4
R8976 s3_bar.n1 s3_bar.t0 24
R8977 s3_bar.n1 s3_bar.t1 24
R8978 s3_bar.n5 s3_bar.n4 8.764
R8979 s3_bar s3_bar.n5 4.681
R8980 EESPFAL_s3_0/s3_bar s3_bar 0.09
R8981 x2.n5 x2.t10 1176.57
R8982 x2.n2 x2.t6 1176.57
R8983 x2.n5 x2.t11 1149.49
R8984 x2.n2 x2.t9 1149.49
R8985 EESPFAL_s0_0/EESPFAL_NAND_v3_2/A x2.t4 1074.82
R8986 x2.n4 x2.t3 800.452
R8987 x2.n4 x2.t5 787.997
R8988 EESPFAL_s1_0/EESPFAL_INV4_1/A x2.t1 778.1
R8989 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A_bar x2.t0 696.166
R8990 x2 x2.t2 687.833
R8991 EESPFAL_s2_0/EESPFAL_4in_NAND_0/D x2.t8 444.545
R8992 EESPFAL_s2_0/EESPFAL_INV4_0/A_bar x2.t7 392.5
R8993 x2.n1 EESPFAL_s0_0/EESPFAL_NAND_v3_2/A 265.13
R8994 x2.n6 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A_bar 219.021
R8995 x2.n8 EESPFAL_s2_0/EESPFAL_INV4_0/A_bar 196.579
R8996 x2.n7 EESPFAL_s2_0/EESPFAL_XOR_v3_0/B 181.93
R8997 x2.n9 EESPFAL_s2_0/EESPFAL_4in_NAND_0/D 181.93
R8998 EESPFAL_s2_0/EESPFAL_XOR_v3_0/B x2.n4 169.6
R8999 x2.n6 EESPFAL_s3_0/EESPFAL_XOR_v3_1/A 169.13
R9000 x2.n3 EESPFAL_s1_0/EESPFAL_XOR_v3_0/A 169.13
R9001 EESPFAL_s3_0/EESPFAL_XOR_v3_1/A x2.n5 128
R9002 EESPFAL_s1_0/EESPFAL_XOR_v3_0/A x2.n2 128
R9003 x2.n10 EESPFAL_s1_0/EESPFAL_INV4_1/A 41.1
R9004 x2.n0 x2 22.914
R9005 x2.n10 x2.n9 4.435
R9006 EESPFAL_s3_0/x2 x2.n6 3.203
R9007 EESPFAL_s1_0/x2 x2.n10 3.2
R9008 x2.n9 x2.n8 2.36
R9009 x2.n1 x2.n0 2.092
R9010 x2.n8 x2.n7 1.796
R9011 x2.n3 x2.n1 1.312
R9012 EESPFAL_s2_0/x2 EESPFAL_s3_0/x2 1.192
R9013 x2.n0 EESPFAL_s0_0/x2 0.956
R9014 x2.n7 EESPFAL_s2_0/x2 0.354
R9015 EESPFAL_s1_0/x2 x2.n3 0.051
C0 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_3070_n7750# 0.00fF
C1 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C2 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar s2 0.07fF
C3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.02fF
C4 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.07fF
C5 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.00fF
C6 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C7 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar Dis2 0.02fF
C8 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT Dis3 0.04fF
C9 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_6971_n4170# 0.00fF
C10 s1_bar EESPFAL_s1_0/EESPFAL_INV4_0/A 0.00fF
C11 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.02fF
C12 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.88fF
C13 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A Dis3 0.08fF
C14 a_2731_n4169# EESPFAL_s2_0/EESPFAL_INV4_2/A 0.00fF
C15 Dis2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.13fF
C16 a_2881_n4169# EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.01fF
C17 Dis2 a_7070_1471# 0.00fF
C18 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C19 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C20 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.02fF
C21 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C22 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.07fF
C23 Dis3 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar 0.00fF
C24 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 1.64fF
C25 s1 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C26 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C27 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.31fF
C28 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B CLK2 0.51fF
C29 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar Dis1 0.16fF
C30 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C Dis3 0.17fF
C31 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.10fF
C32 a_6821_n4170# CLK2 0.00fF
C33 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.11fF
C34 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C35 EESPFAL_s2_0/EESPFAL_INV4_2/A Dis1 0.12fF
C36 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.03fF
C37 s2 a_7190_n4930# 0.00fF
C38 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.56fF
C39 a_2770_n7070# EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C40 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B CLK2 0.42fF
C41 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C42 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.02fF
C43 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C44 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.02fF
C45 CLK1 CLK3 0.25fF
C46 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C47 Dis2 EESPFAL_s1_0/EESPFAL_INV4_0/A 0.05fF
C48 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.36fF
C49 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.08fF
C50 CLK2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.14fF
C51 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C52 a_7040_n4930# EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C53 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.09fF
C54 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C55 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.09fF
C56 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B a_2730_n2029# 0.00fF
C57 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.33fF
C58 s1 a_7190_n4930# 0.00fF
C59 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar a_2770_n7070# 0.00fF
C60 a_6800_n9890# CLK3 0.00fF
C61 CLK1 a_3030_n10570# 0.02fF
C62 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar s3 0.08fF
C63 a_2730_n9890# Dis1 0.00fF
C64 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B CLK3 0.01fF
C65 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.09fF
C66 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.09fF
C67 Dis1 a_1170_1471# 0.02fF
C68 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.09fF
C69 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar a_2730_791# 0.01fF
C70 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_2730_n10570# 0.01fF
C71 a_3030_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C72 a_2770_n7750# CLK1 0.02fF
C73 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.38fF
C74 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 1.00fF
C75 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C76 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C77 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar Dis2 0.01fF
C78 s0_bar CLK3 1.12fF
C79 s0 CLK2 0.18fF
C80 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C81 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.03fF
C82 Dis1 a_1170_n2029# 0.02fF
C83 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C84 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.75fF
C85 a_2920_n4929# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C86 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C CLK3 0.51fF
C87 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT a_6971_n12711# 0.00fF
C88 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar a_1470_n9890# 0.00fF
C89 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar a_3030_n2029# 0.00fF
C90 s2 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.00fF
C91 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.02fF
C92 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.04fF
C93 Dis3 a_6821_n12711# 0.00fF
C94 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar CLK3 0.34fF
C95 a_6821_n4170# s2 0.00fF
C96 Dis2 s3 0.02fF
C97 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.15fF
C98 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C99 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_1170_n1349# 0.01fF
C100 Dis1 a_2730_791# 0.00fF
C101 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar Dis2 0.01fF
C102 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.08fF
C103 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.04fF
C104 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A a_1470_n10570# 0.00fF
C105 a_1470_n9890# EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C106 s1_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.01fF
C107 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C108 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C109 CLK1 a_1170_n1349# 0.01fF
C110 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.02fF
C111 CLK2 a_6800_n1349# 0.02fF
C112 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.00fF
C113 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C114 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar Dis3 0.05fF
C115 s2 CLK2 0.12fF
C116 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar CLK1 0.04fF
C117 s2_bar CLK3 1.01fF
C118 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_1210_n7750# 0.00fF
C119 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar CLK1 1.26fF
C120 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.02fF
C121 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.01fF
C122 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.03fF
C123 Dis3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.02fF
C124 s1 a_6821_n4170# 0.00fF
C125 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C126 a_1210_n7070# Dis1 0.01fF
C127 a_7070_1471# Dis3 0.00fF
C128 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C129 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C130 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C131 s0_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.01fF
C132 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.01fF
C133 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C134 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C135 CLK3 a_5050_791# 0.00fF
C136 CLK3 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.32fF
C137 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B CLK1 0.83fF
C138 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar CLK2 0.04fF
C139 EESPFAL_s2_0/EESPFAL_INV4_2/A CLK2 0.66fF
C140 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B s3 0.00fF
C141 a_2731_n4169# CLK1 0.02fF
C142 s1 CLK2 0.11fF
C143 s1_bar CLK3 1.22fF
C144 a_2730_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C145 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.76fF
C146 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.06fF
C147 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.32fF
C148 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar s3 0.01fF
C149 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar CLK1 0.15fF
C150 Dis3 EESPFAL_s1_0/EESPFAL_INV4_0/A 0.00fF
C151 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.02fF
C152 Dis1 CLK1 11.99fF
C153 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C154 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C155 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.90fF
C156 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C157 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar 0.05fF
C158 CLK1 EESPFAL_s3_0/EESPFAL_INV4_0/A 1.05fF
C159 Dis2 CLK3 7.21fF
C160 a_3790_1471# CLK3 0.00fF
C161 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.02fF
C162 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B s0_bar 0.02fF
C163 Dis1 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.13fF
C164 Dis1 a_2730_1471# 0.00fF
C165 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.99fF
C166 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.12fF
C167 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_3030_n2029# 0.00fF
C168 a_3030_n1349# EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C169 s3 a_6971_n12711# 0.01fF
C170 a_5050_791# EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.00fF
C171 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_6800_n10570# 0.01fF
C172 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.10fF
C173 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT a_7040_n4930# 0.00fF
C174 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.06fF
C175 s2_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar 0.04fF
C176 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C177 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar 0.17fF
C178 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar CLK3 0.03fF
C179 a_2770_n4929# EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.00fF
C180 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar Dis3 0.02fF
C181 a_7190_n4930# EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C182 CLK3 a_6800_n2029# 0.00fF
C183 Dis1 a_2730_n2029# 0.00fF
C184 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar a_3070_n7070# 0.00fF
C185 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 2.14fF
C186 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A CLK3 0.03fF
C187 a_2920_n4929# CLK2 0.00fF
C188 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C Dis1 0.00fF
C189 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar a_3030_n9890# 0.01fF
C190 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C191 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.01fF
C192 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.34fF
C193 Dis3 s3 0.41fF
C194 EESPFAL_s2_0/EESPFAL_INV4_2/A s2 0.00fF
C195 CLK2 a_2730_791# 0.00fF
C196 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar Dis1 0.00fF
C197 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_7040_n4930# 0.00fF
C198 s1 s2 0.11fF
C199 CLK3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.09fF
C200 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_2730_n1349# 0.00fF
C201 s1_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar 0.00fF
C202 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar Dis3 0.00fF
C203 a_3030_n9890# EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C204 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A a_3030_n10570# 0.00fF
C205 CLK1 a_2730_n1349# 0.02fF
C206 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar s2_bar 1.69fF
C207 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B 1.76fF
C208 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.05fF
C209 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar CLK3 0.13fF
C210 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B a_5050_791# 0.00fF
C211 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C a_2731_n12710# 0.00fF
C212 a_6971_n4170# EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C213 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B a_3030_n10570# 0.00fF
C214 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_2770_n7750# 0.00fF
C215 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C a_7190_n4930# 0.00fF
C216 a_6859_n7070# CLK3 0.01fF
C217 a_2770_n7070# Dis1 0.01fF
C218 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C219 s1_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C220 Dis1 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C221 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B CLK1 1.04fF
C222 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B 0.00fF
C223 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.03fF
C224 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar Dis2 0.27fF
C225 Dis2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C226 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.04fF
C227 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.77fF
C228 CLK3 a_6971_n12711# 0.01fF
C229 s2_bar a_7190_n4930# 0.00fF
C230 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B CLK1 0.87fF
C231 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C232 EESPFAL_s3_0/EESPFAL_INV4_0/A EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.34fF
C233 CLK1 CLK2 4.79fF
C234 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.01fF
C235 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.07fF
C236 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_1510_n7070# 0.00fF
C237 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B a_3790_1471# 0.00fF
C238 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B Dis2 0.07fF
C239 CLK1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.87fF
C240 EESPFAL_s3_0/EESPFAL_INV4_0/A a_2881_n12710# 0.01fF
C241 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar 2.13fF
C242 s1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C243 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C244 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_1510_n7750# 0.00fF
C245 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 1.20fF
C246 s1_bar a_7190_n4930# 0.00fF
C247 CLK3 a_7070_791# 0.01fF
C248 a_6800_n9890# CLK2 0.02fF
C249 a_1170_n9890# CLK1 0.02fF
C250 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar a_3030_n1349# 0.00fF
C251 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_2881_n4169# 0.00fF
C252 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar s3_bar 1.83fF
C253 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar Dis2 0.24fF
C254 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B CLK2 0.37fF
C255 Dis3 CLK3 4.16fF
C256 Dis1 a_3790_1471# 0.00fF
C257 Dis1 Dis2 0.13fF
C258 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT a_6800_n10570# 0.01fF
C259 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C260 s0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.01fF
C261 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.01fF
C262 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C263 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.08fF
C264 Dis2 EESPFAL_s3_0/EESPFAL_INV4_0/A 0.04fF
C265 a_6821_n4170# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C266 EESPFAL_s2_0/EESPFAL_INV4_2/A a_2920_n4929# 0.01fF
C267 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B CLK3 0.04fF
C268 a_3070_n4929# EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.00fF
C269 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar Dis1 0.38fF
C270 s0_bar CLK2 0.29fF
C271 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C272 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.36fF
C273 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.07fF
C274 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar a_6859_n7070# 0.00fF
C275 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.01fF
C276 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C CLK2 1.11fF
C277 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A Dis1 0.33fF
C278 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.02fF
C279 a_7070_1471# EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.01fF
C280 s0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C281 s2_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.00fF
C282 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar CLK2 1.22fF
C283 a_6821_n4170# s2_bar 0.00fF
C284 Dis2 s3_bar 0.01fF
C285 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_6800_n1349# 0.01fF
C286 a_6859_n7750# Dis2 0.00fF
C287 Dis1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.09fF
C288 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B s0 0.00fF
C289 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 3.09fF
C290 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT a_7070_1471# 0.01fF
C291 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.05fF
C292 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C293 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.14fF
C294 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C a_6821_n12711# 0.00fF
C295 s2_bar CLK2 0.16fF
C296 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar Dis1 0.00fF
C297 CLK3 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.11fF
C298 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_INV4_0/A 0.01fF
C299 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.07fF
C300 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_INV4_0/A_bar 0.02fF
C301 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.05fF
C302 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar a_6859_n7070# 0.00fF
C303 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar a_6800_n1349# 0.00fF
C304 Dis1 a_1170_n10570# 0.02fF
C305 s1_bar a_6821_n4170# 0.00fF
C306 s2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C307 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.07fF
C308 s0_bar s0 1.62fF
C309 a_1470_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.00fF
C310 a_6859_n7750# EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.00fF
C311 CLK2 a_5050_791# 0.01fF
C312 CLK2 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.91fF
C313 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar Dis3 0.01fF
C314 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar CLK1 1.01fF
C315 EESPFAL_s2_0/EESPFAL_INV4_2/A CLK1 0.92fF
C316 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 1.45fF
C317 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C318 s1_bar CLK2 0.26fF
C319 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B s3_bar 0.01fF
C320 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar s0 0.10fF
C321 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.40fF
C322 CLK2 a_2881_n12710# 0.00fF
C323 a_6971_n4170# EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C324 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar s3_bar 0.05fF
C325 s1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C326 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.06fF
C327 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A a_1470_n2029# 0.00fF
C328 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B Dis3 0.14fF
C329 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_3070_n7070# 0.01fF
C330 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.02fF
C331 a_1510_n7070# EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C332 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B Dis2 0.05fF
C333 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C334 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_3070_n7750# 0.01fF
C335 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.02fF
C336 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C337 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.00fF
C338 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C339 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C340 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C s2 0.08fF
C341 a_2730_n9890# CLK1 0.02fF
C342 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B Dis2 0.05fF
C343 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_6971_n4170# 0.00fF
C344 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar Dis3 0.19fF
C345 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.01fF
C346 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_INV4_0/A 0.34fF
C347 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.78fF
C348 a_3790_1471# CLK2 0.00fF
C349 a_1170_1471# CLK1 0.01fF
C350 Dis1 Dis3 0.06fF
C351 Dis2 CLK2 5.28fF
C352 s0 a_5050_791# 0.00fF
C353 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.70fF
C354 Dis2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.03fF
C355 s3_bar a_6971_n12711# 0.00fF
C356 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar CLK3 0.03fF
C357 a_2881_n4169# EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C358 a_1170_n1349# EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C359 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C360 s2_bar s2 1.79fF
C361 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.04fF
C362 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_1170_n2029# 0.00fF
C363 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.02fF
C364 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.03fF
C365 Dis3 EESPFAL_s3_0/EESPFAL_INV4_0/A 0.00fF
C366 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.05fF
C367 s1 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C368 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar CLK2 0.18fF
C369 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B Dis1 0.09fF
C370 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.06fF
C371 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.03fF
C372 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 1.00fF
C373 CLK2 a_6800_n2029# 0.02fF
C374 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.38fF
C375 CLK1 a_1170_n2029# 0.01fF
C376 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.04fF
C377 a_7190_n4930# Dis3 0.00fF
C378 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A CLK2 0.79fF
C379 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT a_6821_n12711# 0.00fF
C380 a_2920_n4929# CLK1 0.02fF
C381 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.03fF
C382 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C383 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C384 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.41fF
C385 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.08fF
C386 CLK1 a_2730_791# 0.02fF
C387 EESPFAL_s2_0/EESPFAL_INV4_2/A s2_bar 0.00fF
C388 Dis3 s3_bar 0.28fF
C389 a_6859_n7750# Dis3 0.00fF
C390 CLK2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.50fF
C391 s1_bar s2 0.03fF
C392 s1 s2_bar 0.02fF
C393 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C394 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.15fF
C395 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C396 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A a_1170_n9890# 0.01fF
C397 Dis2 s0 0.02fF
C398 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C399 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.51fF
C400 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 1.27fF
C401 EESPFAL_s2_0/EESPFAL_INV4_2/A a_2770_n7070# 0.00fF
C402 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar CLK2 1.37fF
C403 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C s3 0.08fF
C404 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C405 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 1.64fF
C406 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C407 Dis1 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.38fF
C408 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.32fF
C409 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B a_2730_791# 0.01fF
C410 CLK3 a_6800_n10570# 0.00fF
C411 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_INV4_2/A_bar 0.00fF
C412 Dis1 a_2730_n10570# 0.00fF
C413 a_1210_n7070# CLK1 0.01fF
C414 s1_bar s1 2.12fF
C415 a_6859_n7070# CLK2 0.02fF
C416 a_3030_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.01fF
C417 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.66fF
C418 Dis2 a_6800_n1349# 0.00fF
C419 a_2881_n4169# EESPFAL_s2_0/EESPFAL_INV4_2/A_bar 0.00fF
C420 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.31fF
C421 a_7040_n4930# CLK3 0.02fF
C422 s2 Dis2 0.01fF
C423 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C424 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C425 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar CLK3 0.38fF
C426 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.03fF
C427 CLK2 a_6971_n12711# 0.00fF
C428 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C429 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 1.69fF
C430 a_2920_n4929# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C431 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.09fF
C432 a_1510_n7750# Dis1 0.02fF
C433 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT CLK3 0.69fF
C434 s2 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C435 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C436 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A a_3030_n2029# 0.01fF
C437 a_3070_n7070# EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C438 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B Dis3 0.06fF
C439 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.06fF
C440 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_1170_n1349# 0.00fF
C441 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.07fF
C442 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar Dis2 0.02fF
C443 a_6821_n4170# Dis3 0.00fF
C444 EESPFAL_s2_0/EESPFAL_INV4_2/A Dis2 0.04fF
C445 s1 Dis2 0.02fF
C446 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.01fF
C447 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 1.45fF
C448 s1_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C449 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C450 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C451 CLK2 a_7070_791# 0.00fF
C452 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C453 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.05fF
C454 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B Dis3 0.05fF
C455 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B CLK3 0.81fF
C456 a_7190_n4930# EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C457 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar a_1470_n10570# 0.01fF
C458 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B CLK1 0.97fF
C459 Dis3 CLK2 1.25fF
C460 a_2730_1471# CLK1 0.02fF
C461 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.04fF
C462 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.03fF
C463 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C464 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.03fF
C465 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C466 Dis3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.04fF
C467 a_3030_n9890# EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.00fF
C468 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C469 EESPFAL_s1_0/EESPFAL_INV4_0/A EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.74fF
C470 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar Dis1 0.16fF
C471 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.02fF
C472 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.01fF
C473 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C474 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C475 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.01fF
C476 a_2730_n1349# EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C477 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_2730_n2029# 0.00fF
C478 s0_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C479 CLK3 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.50fF
C480 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B CLK2 0.47fF
C481 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar CLK3 0.33fF
C482 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar s3 0.00fF
C483 a_2730_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.00fF
C484 CLK1 a_2730_n2029# 0.02fF
C485 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.03fF
C486 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.29fF
C487 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.01fF
C488 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT s3 0.05fF
C489 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C CLK1 0.10fF
C490 s0 a_7070_791# 0.00fF
C491 s0_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.03fF
C492 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar CLK1 0.02fF
C493 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar s3 0.02fF
C494 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C495 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C496 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.09fF
C497 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B s0_bar 0.00fF
C498 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A a_2730_n9890# 0.00fF
C499 Dis3 s0 0.20fF
C500 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C501 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C502 CLK2 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.85fF
C503 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.07fF
C504 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.10fF
C505 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.01fF
C506 a_5050_791# EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.00fF
C507 a_2770_n7070# CLK1 0.02fF
C508 s2_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C509 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar a_2730_n10570# 0.00fF
C510 a_7070_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.01fF
C511 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar 0.69fF
C512 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.80fF
C513 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar a_7040_n4930# 0.00fF
C514 CLK1 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.16fF
C515 CLK1 a_5050_791# 0.00fF
C516 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A CLK3 0.21fF
C517 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT 0.07fF
C518 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.02fF
C519 a_2770_n4929# EESPFAL_s1_0/EESPFAL_INV4_0/A 0.00fF
C520 s2 Dis3 0.42fF
C521 a_7190_n4930# EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C522 Dis1 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.02fF
C523 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar s0_bar 0.05fF
C524 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 1.23fF
C525 CLK1 a_2881_n12710# 0.02fF
C526 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar CLK3 0.03fF
C527 a_3070_n7750# Dis1 0.00fF
C528 s1_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.05fF
C529 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_s1_0/EESPFAL_INV4_0/A 0.06fF
C530 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 2.86fF
C531 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar 0.00fF
C532 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_2730_n1349# 0.01fF
C533 CLK3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C534 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar Dis3 0.04fF
C535 EESPFAL_s2_0/EESPFAL_INV4_2/A Dis3 0.00fF
C536 s0 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C537 s1 Dis3 0.43fF
C538 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar a_3030_n10570# 0.00fF
C539 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C s2_bar 0.11fF
C540 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar a_3030_1471# 0.00fF
C541 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_1210_n7070# 0.01fF
C542 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B 0.10fF
C543 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.48fF
C544 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C545 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT CLK3 1.16fF
C546 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar a_2731_n12710# 0.00fF
C547 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B Dis1 0.00fF
C548 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar a_3030_n9890# 0.00fF
C549 a_3790_1471# CLK1 0.02fF
C550 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar a_3030_n10570# 0.00fF
C551 Dis2 CLK1 0.32fF
C552 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s1_0/EESPFAL_INV4_0/A 0.00fF
C553 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_2770_n7750# 0.00fF
C554 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_1210_n7750# 0.01fF
C555 s0_bar a_5050_791# 0.00fF
C556 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.50fF
C557 Dis1 a_1470_n1349# 0.01fF
C558 CLK3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.38fF
C559 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar CLK2 0.13fF
C560 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_2731_n4169# 0.00fF
C561 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_6800_n2029# 0.00fF
C562 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.32fF
C563 s1_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C564 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar CLK1 1.98fF
C565 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C566 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C567 a_6800_n9890# Dis2 0.00fF
C568 Dis1 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C569 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_INV4_0/A_bar 0.01fF
C570 a_3790_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.00fF
C571 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar Dis1 0.00fF
C572 Dis2 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.04fF
C573 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.04fF
C574 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B a_7190_n4930# 0.00fF
C575 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.10fF
C576 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar a_2770_n4929# 0.00fF
C577 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A CLK1 1.93fF
C578 EESPFAL_s3_0/EESPFAL_INV4_0/A EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.07fF
C579 a_6971_n4170# CLK3 0.02fF
C580 a_6821_n4170# EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C581 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B a_6859_n7750# 0.00fF
C582 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar a_6800_n2029# 0.00fF
C583 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.07fF
C584 a_6800_n1349# EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C585 s1_bar s2_bar 0.02fF
C586 CLK1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.83fF
C587 s2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C588 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A a_6800_n9890# 0.01fF
C589 s1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C590 Dis2 s0_bar 0.01fF
C591 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.97fF
C592 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B a_3030_n1349# 0.00fF
C593 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar CLK1 0.05fF
C594 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_7190_n4930# 0.00fF
C595 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C s3_bar 0.12fF
C596 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C Dis2 0.39fF
C597 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar Dis2 0.24fF
C598 CLK2 a_6800_n10570# 0.02fF
C599 CLK1 a_1170_n10570# 0.01fF
C600 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar a_2881_n12710# 0.00fF
C601 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar a_6800_n9890# 0.00fF
C602 s1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.02fF
C603 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.02fF
C604 s0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C605 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C606 a_7040_n4930# CLK2 0.00fF
C607 a_3070_n4929# EESPFAL_s1_0/EESPFAL_INV4_0/A 0.00fF
C608 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A CLK3 0.03fF
C609 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A Dis1 0.29fF
C610 s2_bar Dis2 0.01fF
C611 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar CLK2 1.22fF
C612 a_1170_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C613 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.21fF
C614 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.98fF
C615 s2 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C616 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar Dis1 0.29fF
C617 a_7070_1471# EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.00fF
C618 s0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C619 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.08fF
C620 s2_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C621 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT CLK2 0.78fF
C622 Dis2 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.23fF
C623 Dis2 a_5050_791# 0.02fF
C624 a_6821_n4170# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B 0.00fF
C625 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_6821_n12711# 0.00fF
C626 Dis1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.32fF
C627 s1_bar Dis2 0.01fF
C628 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.08fF
C629 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar a_1170_n2029# 0.01fF
C630 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.12fF
C631 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.10fF
C632 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_2770_n7070# 0.00fF
C633 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.02fF
C634 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C635 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B CLK2 0.93fF
C636 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT Dis1 0.00fF
C637 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.00fF
C638 Dis3 CLK1 0.78fF
C639 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_INV4_0/A 0.01fF
C640 CLK3 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.04fF
C641 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.21fF
C642 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_6859_n7750# 0.00fF
C643 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_2770_n7750# 0.00fF
C644 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar a_2730_791# 0.01fF
C645 Dis1 a_3030_n1349# 0.00fF
C646 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C a_6859_n7070# 0.00fF
C647 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT a_6800_n1349# 0.01fF
C648 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_6821_n4170# 0.00fF
C649 Dis1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C650 s2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C651 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.07fF
C652 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar s0 0.69fF
C653 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_INV4_0/A 0.01fF
C654 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C655 CLK2 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 1.06fF
C656 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B CLK1 0.90fF
C657 a_2731_n4169# EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.01fF
C658 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C659 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar s3_bar 0.00fF
C660 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C661 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar CLK2 0.94fF
C662 Dis3 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.00fF
C663 Dis2 a_3790_1471# 0.00fF
C664 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT s0 0.06fF
C665 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.77fF
C666 a_6971_n4170# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C667 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar a_3070_n4929# 0.00fF
C668 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT s3_bar 0.07fF
C669 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C670 a_2881_n4169# CLK2 0.00fF
C671 s1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.04fF
C672 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B a_6800_n9890# 0.00fF
C673 s2 a_7040_n4930# 0.00fF
C674 s0_bar a_7070_791# 0.00fF
C675 Dis1 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.29fF
C676 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.05fF
C677 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C678 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar Dis2 0.02fF
C679 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar s3_bar 0.05fF
C680 Dis3 s0_bar 0.17fF
C681 Dis2 a_6800_n2029# 0.00fF
C682 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.07fF
C683 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C684 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C685 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C686 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT a_6800_n1349# 0.00fF
C687 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar a_7070_791# 0.00fF
C688 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A Dis2 0.02fF
C689 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C Dis3 0.19fF
C690 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_INV4_0/A 0.07fF
C691 CLK1 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 1.57fF
C692 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 1.68fF
C693 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 1.02fF
C694 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar Dis3 0.12fF
C695 s1 a_7040_n4930# 0.00fF
C696 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar a_6971_n12711# 0.00fF
C697 CLK1 a_2730_n10570# 0.02fF
C698 a_1470_n9890# Dis1 0.01fF
C699 Dis2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.06fF
C700 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar a_3070_n7750# 0.00fF
C701 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B s2 0.05fF
C702 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.02fF
C703 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.01fF
C704 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C705 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C706 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.01fF
C707 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C708 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar Dis2 0.33fF
C709 s2_bar Dis3 0.30fF
C710 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A CLK2 0.82fF
C711 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_1470_n10570# 0.00fF
C712 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A Dis1 0.34fF
C713 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 1.26fF
C714 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.26fF
C715 a_2730_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C716 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C717 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.31fF
C718 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar CLK2 0.10fF
C719 a_1510_n7750# CLK1 0.02fF
C720 a_6859_n7070# Dis2 0.00fF
C721 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C722 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C723 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.00fF
C724 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 1.05fF
C725 Dis3 a_5050_791# 0.00fF
C726 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 1.02fF
C727 Dis3 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.18fF
C728 a_2770_n4929# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C729 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar s2 0.00fF
C730 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B 0.00fF
C731 s1 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B 0.01fF
C732 CLK2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.09fF
C733 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C734 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A s3 0.02fF
C735 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT a_6821_n12711# 0.00fF
C736 s1_bar Dis3 0.29fF
C737 s0_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C738 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.06fF
C739 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar a_1170_n9890# 0.00fF
C740 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.07fF
C741 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.29fF
C742 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar a_2730_n2029# 0.00fF
C743 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.05fF
C744 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT CLK2 1.07fF
C745 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar s3 0.00fF
C746 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.02fF
C747 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A a_1170_n10570# 0.00fF
C748 a_1170_n9890# EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C749 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.02fF
C750 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C751 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.06fF
C752 Dis1 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.32fF
C753 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_6859_n7750# 0.01fF
C754 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.28fF
C755 CLK2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 1.23fF
C756 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_INV4_2/A 0.01fF
C757 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar s1 0.07fF
C758 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar CLK1 0.87fF
C759 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.09fF
C760 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar CLK3 0.21fF
C761 a_2881_n4169# EESPFAL_s2_0/EESPFAL_INV4_2/A 0.00fF
C762 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 3.15fF
C763 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C764 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C765 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B CLK3 0.43fF
C766 Dis2 Dis3 3.18fF
C767 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar a_2730_791# 0.00fF
C768 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 1.28fF
C769 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C770 a_6971_n4170# CLK2 0.00fF
C771 CLK2 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.08fF
C772 a_1470_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C773 s2 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.01fF
C774 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar a_5050_791# 0.01fF
C775 a_3070_n7070# EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C776 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar CLK3 0.02fF
C777 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar Dis3 0.03fF
C778 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.05fF
C779 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.04fF
C780 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.56fF
C781 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar a_6971_n12711# 0.00fF
C782 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B Dis2 0.05fF
C783 s2_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.01fF
C784 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.01fF
C785 s1_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C786 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.01fF
C787 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C788 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C789 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A Dis3 0.09fF
C790 a_7190_n4930# EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C791 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT CLK3 1.33fF
C792 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C793 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B a_3030_n2029# 0.00fF
C794 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.04fF
C795 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C796 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C797 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar a_3070_n7070# 0.00fF
C798 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.07fF
C799 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A CLK3 0.22fF
C800 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.87fF
C801 Dis3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.06fF
C802 a_3030_n9890# Dis1 0.00fF
C803 s1_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C804 Dis1 a_1470_1471# 0.01fF
C805 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.02fF
C806 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C807 s0_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C808 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.01fF
C809 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C810 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C811 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.03fF
C812 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_2730_n2029# 0.00fF
C813 a_2730_n1349# EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C814 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar Dis3 0.01fF
C815 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A CLK2 0.79fF
C816 s3 a_6821_n12711# 0.01fF
C817 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_3030_n10570# 0.01fF
C818 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C CLK3 0.50fF
C819 Dis2 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.11fF
C820 a_3790_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C821 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar CLK1 0.19fF
C822 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C823 s2_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C824 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.06fF
C825 a_3070_n7750# CLK1 0.02fF
C826 a_6859_n7070# Dis3 0.00fF
C827 a_7040_n4930# EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C828 s0_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.02fF
C829 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C830 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.68fF
C831 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C832 Dis1 a_1470_n2029# 0.01fF
C833 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT CLK1 0.00fF
C834 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar a_2770_n7070# 0.00fF
C835 a_3070_n4929# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C836 a_2770_n4929# CLK2 0.00fF
C837 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT s3 0.06fF
C838 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C839 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar a_2730_n9890# 0.01fF
C840 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.00fF
C841 a_6821_n4170# EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C842 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.14fF
C843 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.31fF
C844 Dis3 a_6971_n12711# 0.00fF
C845 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.02fF
C846 a_6971_n4170# s2 0.00fF
C847 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.17fF
C848 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_1470_n1349# 0.01fF
C849 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B CLK1 0.01fF
C850 a_2730_n9890# EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C851 CLK2 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.83fF
C852 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A a_2730_n10570# 0.00fF
C853 CLK1 a_1470_n1349# 0.02fF
C854 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.95fF
C855 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.00fF
C856 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.02fF
C857 a_5050_791# EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C858 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C859 a_6821_n4170# EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C860 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar s0_bar 0.15fF
C861 s2_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C862 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_1510_n7750# 0.00fF
C863 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar a_6800_n2029# 0.00fF
C864 Dis3 a_7070_791# 0.00fF
C865 CLK1 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.11fF
C866 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C a_7040_n4930# 0.00fF
C867 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.02fF
C868 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar 0.08fF
C869 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar 0.74fF
C870 s1 a_6971_n4170# 0.00fF
C871 s1 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.00fF
C872 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar Dis1 0.00fF
C873 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C874 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.01fF
C875 a_1510_n7070# Dis1 0.02fF
C876 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar CLK1 0.17fF
C877 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.26fF
C878 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT s0_bar 0.12fF
C879 Dis1 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.01fF
C880 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.94fF
C881 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar Dis2 0.02fF
C882 a_2881_n4169# CLK1 0.02fF
C883 a_3030_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C884 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.02fF
C885 s1_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.07fF
C886 CLK3 a_6821_n12711# 0.01fF
C887 s2_bar a_7040_n4930# 0.00fF
C888 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar 0.72fF
C889 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar Dis1 0.15fF
C890 Dis1 a_2731_n12710# 0.00fF
C891 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B Dis3 0.06fF
C892 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar 0.00fF
C893 a_6800_n10570# EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C894 s0 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.01fF
C895 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar a_7190_n4930# 0.00fF
C896 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B a_3030_1471# 0.00fF
C897 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.34fF
C898 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_1210_n7070# 0.00fF
C899 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C900 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B 1.45fF
C901 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C902 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar CLK3 0.03fF
C903 EESPFAL_s3_0/EESPFAL_INV4_0/A a_2731_n12710# 0.01fF
C904 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT Dis1 0.00fF
C905 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B a_3030_n9890# 0.00fF
C906 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar a_6859_n7750# 0.00fF
C907 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C908 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar a_5050_791# 0.00fF
C909 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_1210_n7750# 0.00fF
C910 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.03fF
C911 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C912 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C913 s1_bar a_7040_n4930# 0.00fF
C914 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar a_2730_n1349# 0.00fF
C915 CLK3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.76fF
C916 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A Dis1 0.28fF
C917 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_2731_n4169# 0.00fF
C918 a_7070_1471# CLK3 0.00fF
C919 Dis1 a_3030_1471# 0.00fF
C920 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B s2_bar 0.10fF
C921 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.16fF
C922 a_6800_n1349# EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.00fF
C923 Dis1 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar 0.27fF
C924 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C925 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A CLK1 1.47fF
C926 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C927 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_INV4_0/A 0.06fF
C928 Dis3 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.04fF
C929 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C Dis1 0.00fF
C930 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.08fF
C931 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT a_7190_n4930# 0.00fF
C932 Dis2 a_6800_n10570# 0.00fF
C933 EESPFAL_s2_0/EESPFAL_INV4_2/A a_2770_n4929# 0.01fF
C934 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar CLK1 1.34fF
C935 EESPFAL_s3_0/EESPFAL_INV4_0/A EESPFAL_s3_0/EESPFAL_INV4_0/A_bar 0.73fF
C936 a_2920_n4929# EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.00fF
C937 CLK3 EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C938 Dis1 a_3030_n2029# 0.00fF
C939 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT a_6859_n7750# 0.01fF
C940 a_6800_n1349# EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C941 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT a_6800_n2029# 0.01fF
C942 s1_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B 0.00fF
C943 CLK1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 1.67fF
C944 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar s2_bar 0.01fF
C945 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A s3_bar 0.03fF
C946 a_3070_n4929# CLK2 0.00fF
C947 s2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C948 a_3790_1471# EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.00fF
C949 s1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.02fF
C950 Dis2 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.30fF
C951 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.01fF
C952 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.16fF
C953 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_7190_n4930# 0.00fF
C954 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT CLK1 0.01fF
C955 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_3030_n1349# 0.00fF
C956 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 2.13fF
C957 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A a_6800_n10570# 0.00fF
C958 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.02fF
C959 CLK1 a_3030_n1349# 0.02fF
C960 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT Dis2 0.11fF
C961 CLK1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C962 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C a_2881_n12710# 0.00fF
C963 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar s1_bar 1.83fF
C964 s1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.06fF
C965 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT a_6800_n9890# 0.01fF
C966 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C967 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_3070_n7750# 0.00fF
C968 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.03fF
C969 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar CLK3 0.01fF
C970 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar CLK2 1.32fF
C971 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B Dis2 0.10fF
C972 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar a_6800_n10570# 0.00fF
C973 a_3070_n7070# Dis1 0.00fF
C974 a_6800_n9890# EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C975 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B CLK2 0.67fF
C976 a_1170_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.00fF
C977 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B a_3030_n1349# 0.00fF
C978 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.03fF
C979 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar Dis3 0.04fF
C980 CLK1 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 1.44fF
C981 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.03fF
C982 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.02fF
C983 s2_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.02fF
C984 CLK3 s3 1.06fF
C985 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar CLK2 0.06fF
C986 CLK2 a_2731_n12710# 0.00fF
C987 Dis2 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.41fF
C988 a_6821_n4170# EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C989 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar Dis2 0.25fF
C990 a_6971_n4170# EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C991 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C992 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C993 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C994 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.08fF
C995 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_2770_n7070# 0.01fF
C996 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A a_1170_n2029# 0.00fF
C997 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.02fF
C998 a_1210_n7070# EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C999 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar Dis1 0.17fF
C1000 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT CLK2 1.03fF
C1001 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.00fF
C1002 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar a_2770_n7750# 0.01fF
C1003 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A a_2730_791# 0.00fF
C1004 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A CLK2 0.95fF
C1005 a_1470_n9890# CLK1 0.02fF
C1006 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_6821_n4170# 0.00fF
C1007 Dis1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1008 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_6800_n2029# 0.00fF
C1009 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B s0 0.09fF
C1010 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.04fF
C1011 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.03fF
C1012 CLK2 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar 0.08fF
C1013 s3_bar a_6821_n12711# 0.00fF
C1014 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A CLK1 1.87fF
C1015 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C1016 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C1017 a_2731_n4169# EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C1018 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C CLK2 1.08fF
C1019 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_INV4_0/A 0.00fF
C1020 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.05fF
C1021 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar s0 0.01fF
C1022 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B a_6859_n7070# 0.01fF
C1023 a_6971_n4170# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1024 EESPFAL_s2_0/EESPFAL_INV4_2/A a_3070_n4929# 0.01fF
C1025 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C1026 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C1027 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.10fF
C1028 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_6800_n9890# 0.00fF
C1029 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B a_6800_n1349# 0.00fF
C1030 Dis1 EESPFAL_s1_0/EESPFAL_INV4_0/A 0.11fF
C1031 s2 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.01fF
C1032 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1033 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar a_7070_791# 0.02fF
C1034 a_7040_n4930# Dis3 0.00fF
C1035 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A Dis2 0.03fF
C1036 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.22fF
C1037 a_2770_n4929# CLK1 0.02fF
C1038 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT s3_bar 0.11fF
C1039 Dis3 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.47fF
C1040 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.01fF
C1041 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C1042 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.02fF
C1043 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C1044 a_6971_n4170# s2_bar 0.00fF
C1045 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT a_7070_791# 0.01fF
C1046 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar Dis2 0.02fF
C1047 CLK1 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 1.24fF
C1048 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 1.18fF
C1049 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 1.44fF
C1050 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B a_3070_n7070# 0.00fF
C1051 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT Dis3 0.08fF
C1052 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.09fF
C1053 Dis2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.04fF
C1054 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C a_6971_n12711# 0.00fF
C1055 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B a_3070_n7750# 0.00fF
C1056 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1057 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.03fF
C1058 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT s2 0.04fF
C1059 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.02fF
C1060 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1061 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.01fF
C1062 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1063 Dis1 a_1470_n10570# 0.01fF
C1064 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT Dis2 0.16fF
C1065 s1_bar a_6971_n4170# 0.00fF
C1066 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B Dis3 0.03fF
C1067 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar Dis1 0.31fF
C1068 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.32fF
C1069 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 3.15fF
C1070 a_2730_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.01fF
C1071 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C1072 Dis2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.31fF
C1073 a_2731_n4169# EESPFAL_s2_0/EESPFAL_INV4_2/A_bar 0.00fF
C1074 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.02fF
C1075 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.00fF
C1076 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.02fF
C1077 CLK2 a_6821_n12711# 0.00fF
C1078 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.09fF
C1079 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.09fF
C1080 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C1081 Dis3 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.18fF
C1082 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C1083 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C1084 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C s2 0.01fF
C1085 s1 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1086 a_1210_n7750# Dis1 0.01fF
C1087 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.04fF
C1088 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.56fF
C1089 s0_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.01fF
C1090 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar Dis1 0.39fF
C1091 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.05fF
C1092 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar Dis3 0.18fF
C1093 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.14fF
C1094 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.36fF
C1095 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.08fF
C1096 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A a_2730_n2029# 0.01fF
C1097 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_6859_n7070# 0.01fF
C1098 a_2770_n7070# EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C1099 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar CLK2 0.05fF
C1100 EESPFAL_s3_0/EESPFAL_INV4_0/A s3 0.00fF
C1101 Dis2 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.01fF
C1102 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.02fF
C1103 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1104 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 0.03fF
C1105 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.02fF
C1106 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1107 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.04fF
C1108 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.10fF
C1109 a_3030_n9890# CLK1 0.02fF
C1110 CLK2 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.94fF
C1111 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_INV4_2/A 0.01fF
C1112 a_7040_n4930# EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1113 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C s1 0.08fF
C1114 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.87fF
C1115 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.16fF
C1116 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar a_1170_n10570# 0.01fF
C1117 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C1118 a_7070_1471# CLK2 0.01fF
C1119 a_1470_1471# CLK1 0.02fF
C1120 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar CLK3 0.60fF
C1121 s3_bar s3 2.14fF
C1122 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1123 a_2730_n9890# EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.00fF
C1124 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 1.02fF
C1125 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.16fF
C1126 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_1470_n2029# 0.00fF
C1127 a_1470_n1349# EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1128 CLK2 EESPFAL_s1_0/EESPFAL_INV4_0/A 0.74fF
C1129 CLK1 a_1470_n2029# 0.02fF
C1130 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A a_5050_791# 0.00fF
C1131 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B CLK3 0.05fF
C1132 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.03fF
C1133 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A Dis3 0.01fF
C1134 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1135 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT a_6971_n12711# 0.00fF
C1136 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1137 a_3070_n4929# CLK1 0.02fF
C1138 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A Dis2 0.01fF
C1139 s2_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1140 s1_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.03fF
C1141 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1142 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.01fF
C1143 CLK1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 1.03fF
C1144 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar Dis3 0.08fF
C1145 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar CLK3 0.33fF
C1146 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar a_6971_n12711# 0.00fF
C1147 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A a_1470_n9890# 0.01fF
C1148 a_7070_1471# s0 0.00fF
C1149 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar a_3030_n2029# 0.00fF
C1150 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar 0.01fF
C1151 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.02fF
C1152 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.00fF
C1153 Dis1 CLK3 0.01fF
C1154 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.09fF
C1155 Dis3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar 0.08fF
C1156 EESPFAL_s2_0/EESPFAL_INV4_2/A a_3070_n7070# 0.00fF
C1157 s1_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.11fF
C1158 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.22fF
C1159 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1160 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/B 0.00fF
C1161 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.16fF
C1162 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1163 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/A 0.02fF
C1164 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C1165 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT Dis3 0.03fF
C1166 CLK3 EESPFAL_s3_0/EESPFAL_INV4_0/A 0.01fF
C1167 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar CLK1 0.05fF
C1168 Dis1 a_3030_n10570# 0.00fF
C1169 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar CLK2 0.09fF
C1170 a_1510_n7070# CLK1 0.01fF
C1171 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B CLK1 0.11fF
C1172 a_3790_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.01fF
C1173 Dis2 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.05fF
C1174 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.04fF
C1175 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.00fF
C1176 Dis3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar 0.01fF
C1177 a_7190_n4930# CLK3 0.02fF
C1178 a_7040_n4930# EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1179 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C1180 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar 0.01fF
C1181 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.02fF
C1182 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1183 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar CLK1 0.79fF
C1184 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C1185 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1186 CLK3 s3_bar 1.19fF
C1187 CLK2 s3 0.11fF
C1188 CLK1 a_2731_n12710# 0.02fF
C1189 a_3070_n4929# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1190 a_6859_n7750# CLK3 0.00fF
C1191 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar s3 0.00fF
C1192 a_2770_n7750# Dis1 0.01fF
C1193 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar CLK2 0.20fF
C1194 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.08fF
C1195 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.13fF
C1196 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A a_6800_n2029# 0.01fF
C1197 a_6859_n7070# EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C1198 Dis1 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.10fF
C1199 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_1470_n1349# 0.00fF
C1200 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1201 a_6971_n4170# Dis3 0.00fF
C1202 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT CLK1 0.01fF
C1203 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar a_2730_n10570# 0.00fF
C1204 Dis3 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.00fF
C1205 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.02fF
C1206 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar a_2730_1471# 0.00fF
C1207 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A CLK1 1.43fF
C1208 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.00fF
C1209 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B s0_bar 0.90fF
C1210 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1211 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar a_2730_n9890# 0.00fF
C1212 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar a_2730_n10570# 0.00fF
C1213 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT a_6800_n2029# 0.01fF
C1214 a_3030_1471# CLK1 0.01fF
C1215 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar 0.22fF
C1216 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.10fF
C1217 Dis1 a_1170_n1349# 0.02fF
C1218 CLK1 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar 1.42fF
C1219 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C1220 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar Dis1 0.00fF
C1221 s1 EESPFAL_s1_0/EESPFAL_INV4_0/A 0.00fF
C1222 a_6800_n9890# EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.00fF
C1223 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C CLK1 0.12fF
C1224 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar s0_bar 0.00fF
C1225 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar 0.08fF
C1226 Dis1 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar 0.30fF
C1227 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.01fF
C1228 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar a_3030_n1349# 0.00fF
C1229 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.47fF
C1230 a_3030_n1349# EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 0.00fF
C1231 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A a_3030_n2029# 0.00fF
C1232 CLK1 a_3030_n2029# 0.02fF
C1233 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar 0.10fF
C1234 a_3030_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_1/B 0.00fF
C1235 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.01fF
C1236 s2_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar 0.10fF
C1237 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B a_7040_n4930# 0.01fF
C1238 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B CLK3 0.08fF
C1239 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar 0.09fF
C1240 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B Dis1 0.08fF
C1241 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A Dis3 0.03fF
C1242 a_6800_n10570# EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1243 a_6821_n4170# CLK3 0.02fF
C1244 a_2731_n4169# Dis1 0.00fF
C1245 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar a_7190_n4930# 0.00fF
C1246 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.10fF
C1247 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar 0.08fF
C1248 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B CLK3 0.02fF
C1249 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar Dis1 0.00fF
C1250 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A a_3030_n9890# 0.00fF
C1251 CLK2 CLK3 5.57fF
C1252 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C1253 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s1_0/EESPFAL_INV4_0/A_bar 0.02fF
C1254 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar a_6859_n7750# 0.00fF
C1255 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.42fF
C1256 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.96fF
C1257 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B a_5050_791# 0.01fF
C1258 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_7040_n4930# 0.00fF
C1259 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar s2 0.00fF
C1260 CLK3 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.03fF
C1261 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A a_7070_791# 0.00fF
C1262 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT s2_bar 0.07fF
C1263 Dis2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.02fF
C1264 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C 0.01fF
C1265 Dis1 EESPFAL_s3_0/EESPFAL_INV4_0/A 0.11fF
C1266 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar a_5050_791# 0.00fF
C1267 a_3070_n7070# CLK1 0.02fF
C1268 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar a_2731_n12710# 0.00fF
C1269 a_6971_n4170# EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C1270 Dis3 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A 0.13fF
C1271 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar a_3030_n10570# 0.00fF
C1272 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.08fF
C1273 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar a_7190_n4930# 0.00fF
C1274 EESPFAL_s2_0/EESPFAL_INV4_2/A EESPFAL_s2_0/EESPFAL_INV4_2/A_bar 0.97fF
C1275 a_2920_n4929# EESPFAL_s1_0/EESPFAL_INV4_0/A 0.00fF
C1276 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B 0.00fF
C1277 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C s2_bar 0.00fF
C1278 s1_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1279 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar Dis2 0.28fF
C1280 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.03fF
C1281 s0 CLK3 0.87fF
C1282 Dis2 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.24fF
C1283 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.02fF
C1284 CLK2 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.48fF
C1285 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar a_3030_n1349# 0.01fF
C1286 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar CLK1 1.17fF
C1287 EESPFAL_s3_0/EESPFAL_INV4_0/A s3_bar 0.00fF
C1288 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C1289 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1290 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.16fF
C1291 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar Dis2 0.06fF
C1292 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_1510_n7070# 0.01fF
C1293 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar a_3790_1471# 0.00fF
C1294 CLK1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C1295 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar a_2881_n12710# 0.00fF
C1296 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C s1_bar 0.12fF
C1297 s1 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.00fF
C1298 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A a_3070_n7750# 0.00fF
C1299 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.02fF
C1300 CLK3 a_6800_n1349# 0.00fF
C1301 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A a_1510_n7750# 0.01fF
C1302 Dis1 a_2730_n1349# 0.00fF
C1303 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar a_2881_n4169# 0.00fF
C1304 s2 CLK3 1.10fF
C1305 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar CLK2 1.22fF
C1306 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT a_6800_n10570# 0.01fF
C1307 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT Dis2 0.11fF
C1308 a_6800_n9890# EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT 0.00fF
C1309 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar CLK2 0.03fF
C1310 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 1.57fF
C1311 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar 3.23fF
C1312 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A Dis2 0.04fF
C1313 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar a_6800_n10570# 0.00fF
C1314 CLK1 EESPFAL_s1_0/EESPFAL_INV4_0/A 1.07fF
C1315 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C1316 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B EESPFAL_s2_0/EESPFAL_NAND_v3_0/A 0.06fF
C1317 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar EESPFAL_s2_0/EESPFAL_NAND_v3_0/B 0.01fF
C1318 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1319 s0 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B 0.00fF
C1320 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B CLK2 0.44fF
C1321 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar a_2920_n4929# 0.00fF
C1322 a_6821_n4170# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C1323 Dis2 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar 0.01fF
C1324 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar CLK3 0.02fF
C1325 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B Dis1 0.09fF
C1326 EESPFAL_s2_0/EESPFAL_INV4_2/A CLK3 0.01fF
C1327 a_2731_n4169# CLK2 0.00fF
C1328 s1 CLK3 1.07fF
C1329 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C Dis2 0.43fF
C1330 a_6971_n4170# EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT 0.00fF
C1331 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_0/A 0.01fF
C1332 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/B 0.49fF
C1333 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT 0.01fF
C1334 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.07fF
C1335 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar a_6859_n7070# 0.00fF
C1336 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/A 0.00fF
C1337 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar CLK2 0.95fF
C1338 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B Dis1 0.10fF
C1339 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.02fF
C1340 a_7070_1471# s0_bar 0.00fF
C1341 Dis1 CLK2 0.10fF
C1342 Dis1 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar 0.16fF
C1343 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A EESPFAL_s3_0/EESPFAL_NAND_v3_1/B 1.06fF
C1344 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C a_6800_n2029# 0.00fF
C1345 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar 0.66fF
C1346 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar 0.01fF
C1347 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar a_7070_1471# 0.01fF
C1348 Dis3 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar 0.05fF
C1349 CLK2 EESPFAL_s3_0/EESPFAL_INV4_0/A 0.72fF
C1350 CLK1 a_1470_n10570# 0.02fF
C1351 a_1170_n9890# Dis1 0.03fF
C1352 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar a_6821_n12711# 0.00fF
C1353 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar CLK1 1.49fF
C1354 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar EESPFAL_s3_0/EESPFAL_NAND_v3_1/A 0.01fF
C1355 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.00fF
C1356 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar EESPFAL_s3_0/EESPFAL_INV4_0/A 0.01fF
C1357 CLK3 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar 0.03fF
C1358 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B s0 0.02fF
C1359 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar a_2770_n7750# 0.00fF
C1360 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT a_6859_n7070# 0.01fF
C1361 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C EESPFAL_s1_0/EESPFAL_INV4_0/A 0.01fF
C1362 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A a_1170_n10570# 0.00fF
C1363 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.10fF
C1364 a_1470_1471# EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar 0.01fF
C1365 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B a_7070_791# 0.00fF
C1366 s2 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar 0.02fF
C1367 CLK2 s3_bar 0.26fF
C1368 a_1210_n7750# CLK1 0.01fF
C1369 a_6859_n7750# CLK2 0.02fF
C1370 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar Dis3 0.01fF
C1371 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar s3_bar 0.00fF
C1372 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar 0.08fF
C1373 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C 0.04fF
C1374 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar CLK1 1.84fF
C1375 Dis3 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B 0.06fF
C1376 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar 0.00fF
C1377 a_6971_n4170# EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B 0.00fF
C1378 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar EESPFAL_s1_0/EESPFAL_NAND_v3_1/A 0.02fF
C1379 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar a_1470_n2029# 0.01fF
C1380 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar a_3070_n7070# 0.00fF
C1381 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar 0.00fF
C1382 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar EESPFAL_s2_0/EESPFAL_NAND_v3_1/B 0.15fF
C1383 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar Dis3 0.01fF
C1384 s1 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar 0.00fF
C1385 a_6971_n12711# GND 0.02fF
C1386 a_6821_n12711# GND 0.02fF
C1387 a_2881_n12710# GND 0.02fF
C1388 a_2731_n12710# GND 0.02fF
C1389 s3 GND 1.76fF
C1390 s3_bar GND 1.70fF
C1391 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar GND 1.26fF $ **FLOATING
C1392 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C GND 1.22fF $ **FLOATING
C1393 EESPFAL_s3_0/EESPFAL_INV4_0/A_bar GND 1.23fF
C1394 EESPFAL_s3_0/EESPFAL_INV4_0/A GND 1.36fF
C1395 a_6800_n10570# GND 0.02fF
C1396 a_3030_n10570# GND 0.01fF
C1397 a_2730_n10570# GND 0.01fF
C1398 a_1470_n10570# GND 0.01fF
C1399 a_1170_n10570# GND 0.01fF
C1400 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT_bar GND 1.49fF
C1401 EESPFAL_s3_0/EESPFAL_NAND_v3_1/OUT GND 1.14fF
C1402 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B_bar GND 1.09fF
C1403 EESPFAL_s3_0/EESPFAL_NAND_v3_1/B GND 1.28fF
C1404 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar GND 2.14fF $ **FLOATING
C1405 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A GND 2.42fF $ **FLOATING
C1406 a_6800_n9890# GND 0.02fF
C1407 a_3030_n9890# GND 0.01fF
C1408 a_2730_n9890# GND 0.01fF
C1409 a_1470_n9890# GND 0.01fF
C1410 a_1170_n9890# GND 0.01fF
C1411 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar GND 2.53fF $ **FLOATING
C1412 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT GND 1.73fF
C1413 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B_bar GND 1.10fF
C1414 EESPFAL_s3_0/EESPFAL_NAND_v3_0/B GND 1.34fF
C1415 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A GND 2.68fF $ **FLOATING
C1416 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar GND 1.89fF $ **FLOATING
C1417 a_6859_n7750# GND 0.02fF
C1418 a_3070_n7750# GND 0.01fF
C1419 a_2770_n7750# GND 0.01fF
C1420 a_1510_n7750# GND 0.02fF
C1421 a_1210_n7750# GND 0.01fF
C1422 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B_bar GND 1.14fF
C1423 EESPFAL_s2_0/EESPFAL_NAND_v3_1/B GND 1.34fF
C1424 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A GND 2.10fF $ **FLOATING
C1425 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar GND 1.65fF $ **FLOATING
C1426 a_6859_n7070# GND 0.02fF
C1427 a_3070_n7070# GND 0.01fF
C1428 a_2770_n7070# GND 0.01fF
C1429 a_1510_n7070# GND 0.02fF
C1430 a_1210_n7070# GND 0.01fF
C1431 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B_bar GND 1.09fF
C1432 EESPFAL_s2_0/EESPFAL_NAND_v3_0/B GND 1.24fF
C1433 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A_bar GND 1.57fF
C1434 EESPFAL_s2_0/EESPFAL_NAND_v3_0/A GND 1.41fF
C1435 a_7190_n4930# GND 0.02fF
C1436 a_7040_n4930# GND 0.02fF
C1437 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar GND 2.57fF $ **FLOATING
C1438 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B_bar GND 1.54fF
C1439 s2 GND 0.99fF
C1440 s2_bar GND 0.96fF
C1441 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/B GND 1.14fF
C1442 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT GND 1.69fF
C1443 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar GND 1.28fF $ **FLOATING
C1444 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C GND 1.25fF $ **FLOATING
C1445 a_3070_n4929# GND 0.02fF
C1446 a_2920_n4929# GND 0.02fF
C1447 a_2770_n4929# GND 0.02fF
C1448 EESPFAL_s2_0/EESPFAL_INV4_2/A_bar GND 1.71fF
C1449 EESPFAL_s2_0/EESPFAL_INV4_2/A GND 1.69fF
C1450 a_6971_n4170# GND 0.02fF
C1451 a_6821_n4170# GND 0.02fF
C1452 a_2881_n4169# GND 0.02fF
C1453 a_2731_n4169# GND 0.02fF
C1454 s1 GND 1.52fF
C1455 s1_bar GND 1.69fF
C1456 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar GND 1.28fF $ **FLOATING
C1457 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C GND 1.25fF $ **FLOATING
C1458 EESPFAL_s1_0/EESPFAL_INV4_0/A_bar GND 1.33fF
C1459 EESPFAL_s1_0/EESPFAL_INV4_0/A GND 1.35fF
C1460 a_6800_n2029# GND 0.02fF
C1461 a_3030_n2029# GND 0.01fF
C1462 a_2730_n2029# GND 0.01fF
C1463 a_1470_n2029# GND 0.01fF
C1464 a_1170_n2029# GND 0.01fF
C1465 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT_bar GND 1.50fF
C1466 EESPFAL_s1_0/EESPFAL_NAND_v3_1/OUT GND 1.14fF
C1467 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B GND 1.21fF
C1468 EESPFAL_s1_0/EESPFAL_NAND_v3_1/B_bar GND 1.11fF
C1469 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar GND 2.41fF $ **FLOATING
C1470 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A GND 2.46fF $ **FLOATING
C1471 a_6800_n1349# GND 0.02fF
C1472 a_3030_n1349# GND 0.01fF
C1473 a_2730_n1349# GND 0.01fF
C1474 a_1470_n1349# GND 0.01fF
C1475 a_1170_n1349# GND 0.01fF
C1476 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar GND 2.53fF $ **FLOATING
C1477 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT GND 1.74fF
C1478 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B_bar GND 1.10fF
C1479 EESPFAL_s1_0/EESPFAL_NAND_v3_0/B GND 1.33fF
C1480 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A GND 2.64fF $ **FLOATING
C1481 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar GND 1.90fF $ **FLOATING
C1482 a_7070_791# GND 0.01fF
C1483 a_5050_791# GND 0.01fF
C1484 a_2730_791# GND 0.02fF
C1485 s0 GND 0.86fF
C1486 s0_bar GND 0.79fF
C1487 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B_bar GND 1.44fF
C1488 EESPFAL_s0_0/EESPFAL_NOR_v3_0/B GND 1.10fF
C1489 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B_bar GND 1.32fF
C1490 EESPFAL_s0_0/EESPFAL_NAND_v3_1/B GND 1.29fF
C1491 Dis3 GND 9.86fF
C1492 a_7070_1471# GND 0.02fF
C1493 a_3790_1471# GND 0.02fF
C1494 a_3030_1471# GND 0.01fF
C1495 a_2730_1471# GND 0.01fF
C1496 a_1470_1471# GND 0.01fF
C1497 a_1170_1471# GND 0.01fF
C1498 Dis2 GND 17.94fF
C1499 Dis1 GND 30.27fF
C1500 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT_bar GND 1.73fF
C1501 EESPFAL_s0_0/EESPFAL_NAND_v3_0/OUT GND 1.61fF
C1502 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B_bar GND 1.17fF
C1503 EESPFAL_s0_0/EESPFAL_NAND_v3_0/B GND 1.33fF
C1504 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar GND 2.51fF $ **FLOATING
C1505 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A GND 3.06fF $ **FLOATING
C1506 CLK3 GND 14.75fF
C1507 CLK2 GND 34.13fF
C1508 CLK1 GND 61.59fF
C1509 EESPFAL_s0_0/x2 GND 0.52fF $ **FLOATING
C1510 x2.t2 GND 0.21fF
C1511 x2.n0 GND 4.69fF $ **FLOATING
C1512 x2.t4 GND 0.42fF
C1513 EESPFAL_s0_0/EESPFAL_NAND_v3_2/A GND 1.99fF $ **FLOATING
C1514 x2.n1 GND 1.90fF $ **FLOATING
C1515 x2.t9 GND 0.29fF
C1516 x2.t6 GND 0.26fF
C1517 x2.n2 GND 2.25fF $ **FLOATING
C1518 EESPFAL_s1_0/EESPFAL_XOR_v3_0/A GND 0.33fF $ **FLOATING
C1519 x2.n3 GND 0.88fF $ **FLOATING
C1520 x2.t1 GND 0.20fF
C1521 EESPFAL_s1_0/EESPFAL_INV4_1/A GND 1.05fF $ **FLOATING
C1522 x2.t8 GND 0.30fF
C1523 EESPFAL_s2_0/EESPFAL_4in_NAND_0/D GND 2.28fF $ **FLOATING
C1524 x2.t7 GND 0.15fF
C1525 EESPFAL_s2_0/EESPFAL_INV4_0/A_bar GND 0.53fF $ **FLOATING
C1526 x2.t3 GND 0.20fF
C1527 x2.t5 GND 0.19fF
C1528 x2.n4 GND 2.35fF $ **FLOATING
C1529 EESPFAL_s2_0/EESPFAL_XOR_v3_0/B GND 0.39fF $ **FLOATING
C1530 x2.t11 GND 0.29fF
C1531 x2.t10 GND 0.26fF
C1532 x2.n5 GND 2.25fF $ **FLOATING
C1533 EESPFAL_s3_0/EESPFAL_XOR_v3_1/A GND 0.33fF $ **FLOATING
C1534 x2.t0 GND 0.25fF
C1535 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A_bar GND 0.76fF $ **FLOATING
C1536 x2.n6 GND 4.56fF $ **FLOATING
C1537 EESPFAL_s3_0/x2 GND 1.96fF $ **FLOATING
C1538 EESPFAL_s2_0/x2 GND 0.69fF $ **FLOATING
C1539 x2.n7 GND 1.24fF $ **FLOATING
C1540 x2.n8 GND 5.70fF $ **FLOATING
C1541 x2.n9 GND 3.32fF $ **FLOATING
C1542 x2.n10 GND 8.07fF $ **FLOATING
C1543 EESPFAL_s1_0/x2 GND 1.45fF $ **FLOATING
C1544 s3_bar.t2 GND 0.05fF
C1545 s3_bar.t3 GND 0.05fF
C1546 s3_bar.n0 GND 0.12fF $ **FLOATING
C1547 s3_bar.t0 GND 0.05fF
C1548 s3_bar.t1 GND 0.05fF
C1549 s3_bar.n1 GND 0.14fF $ **FLOATING
C1550 s3_bar.t4 GND 0.27fF
C1551 s3_bar.n2 GND 0.19fF $ **FLOATING
C1552 s3_bar.n3 GND 0.13fF $ **FLOATING
C1553 s3_bar.t5 GND 0.06fF
C1554 s3_bar.t7 GND 0.06fF
C1555 s3_bar.t6 GND 0.04fF
C1556 s3_bar.n4 GND 0.07fF $ **FLOATING
C1557 s3_bar.n5 GND 0.05fF $ **FLOATING
C1558 EESPFAL_s3_0/s3_bar GND 0.01fF $ **FLOATING
C1559 s3.t2 GND 0.04fF
C1560 s3.t6 GND 0.04fF
C1561 s3.n0 GND 0.15fF $ **FLOATING
C1562 s3.t4 GND 0.19fF
C1563 s3.t5 GND 0.04fF
C1564 s3.t1 GND 0.04fF
C1565 s3.n1 GND 0.14fF $ **FLOATING
C1566 s3.t0 GND 0.04fF
C1567 s3.t3 GND 0.04fF
C1568 s3.n2 GND 0.15fF $ **FLOATING
C1569 s3.t8 GND 0.06fF
C1570 s3.t7 GND 0.06fF
C1571 s3.t9 GND 0.03fF
C1572 s3.n3 GND 0.06fF $ **FLOATING
C1573 s3.n4 GND 0.20fF $ **FLOATING
C1574 s3.n5 GND 0.17fF $ **FLOATING
C1575 s3.n6 GND 0.14fF $ **FLOATING
C1576 EESPFAL_s3_0/s3 GND 0.01fF $ **FLOATING
C1577 EESPFAL_s2_0/EESPFAL_INV4_2/OUT GND 0.23fF $ **FLOATING
C1578 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 GND 0.03fF
C1579 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 GND 0.63fF $ **FLOATING
C1580 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 GND 0.04fF
C1581 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 GND 0.04fF
C1582 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 GND 0.13fF $ **FLOATING
C1583 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 GND 0.25fF
C1584 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 GND 0.17fF $ **FLOATING
C1585 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 GND 0.04fF
C1586 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 GND 0.04fF
C1587 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 GND 0.11fF $ **FLOATING
C1588 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 GND 0.12fF $ **FLOATING
C1589 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 GND 0.04fF
C1590 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 GND 0.06fF
C1591 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 GND 0.05fF
C1592 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 GND 0.06fF $ **FLOATING
C1593 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 GND 0.04fF $ **FLOATING
C1594 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t4 GND 0.04fF
C1595 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t2 GND 0.04fF
C1596 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n0 GND 0.13fF $ **FLOATING
C1597 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t3 GND 0.17fF
C1598 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t8 GND 0.05fF
C1599 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n1 GND 0.78fF $ **FLOATING
C1600 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n2 GND 0.18fF $ **FLOATING
C1601 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t0 GND 0.04fF
C1602 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t1 GND 0.04fF
C1603 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n3 GND 0.12fF $ **FLOATING
C1604 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n4 GND 0.11fF $ **FLOATING
C1605 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n5 GND 0.11fF $ **FLOATING
C1606 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t7 GND 0.03fF
C1607 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t5 GND 0.06fF
C1608 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.t6 GND 0.06fF
C1609 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n6 GND 0.06fF $ **FLOATING
C1610 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/C.n7 GND 0.03fF $ **FLOATING
C1611 EESPFAL_s2_0/EESPFAL_INV4_2/OUT_bar GND 0.01fF $ **FLOATING
C1612 EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT_bar GND 0.12fF $ **FLOATING
C1613 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t9 GND 0.04fF
C1614 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t7 GND 0.07fF
C1615 EESPFAL_s0_0/EESPFAL_NAND_v3_1/A GND 0.34fF $ **FLOATING
C1616 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n0 GND 0.63fF $ **FLOATING
C1617 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t3 GND 0.03fF
C1618 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t2 GND 0.03fF
C1619 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n1 GND 0.08fF $ **FLOATING
C1620 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t0 GND 0.11fF
C1621 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t1 GND 0.18fF
C1622 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n2 GND 0.16fF $ **FLOATING
C1623 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n3 GND 0.07fF $ **FLOATING
C1624 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t5 GND 0.03fF
C1625 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t4 GND 0.03fF
C1626 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n4 GND 0.07fF $ **FLOATING
C1627 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n5 GND 0.08fF $ **FLOATING
C1628 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t8 GND 0.04fF
C1629 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t6 GND 0.03fF
C1630 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.t10 GND 0.03fF
C1631 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n6 GND 0.04fF $ **FLOATING
C1632 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A_bar.n7 GND 0.01fF $ **FLOATING
C1633 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t8 GND 0.08fF
C1634 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t10 GND 0.04fF
C1635 EESPFAL_s0_0/EESPFAL_NAND_v3_1/A_bar GND 0.16fF $ **FLOATING
C1636 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t2 GND 0.12fF
C1637 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t1 GND 0.03fF
C1638 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t3 GND 0.03fF
C1639 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n0 GND 0.09fF $ **FLOATING
C1640 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t5 GND 0.03fF
C1641 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t4 GND 0.03fF
C1642 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n1 GND 0.10fF $ **FLOATING
C1643 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t7 GND 0.04fF
C1644 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t6 GND 0.04fF
C1645 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t9 GND 0.02fF
C1646 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n2 GND 0.04fF $ **FLOATING
C1647 EESPFAL_s0_0/EESPFAL_XOR_v3_0/OUT GND 0.01fF $ **FLOATING
C1648 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n3 GND 0.02fF $ **FLOATING
C1649 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n4 GND 0.13fF $ **FLOATING
C1650 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n5 GND 0.13fF $ **FLOATING
C1651 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.t0 GND 0.12fF
C1652 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n6 GND 0.11fF $ **FLOATING
C1653 EESPFAL_s0_0/EESPFAL_NAND_v3_0/A.n7 GND 0.36fF $ **FLOATING
C1654 EESPFAL_s0_0/x2_bar GND 0.21fF $ **FLOATING
C1655 x2_bar.t0 GND 0.43fF
C1656 x2_bar.n0 GND 4.46fF $ **FLOATING
C1657 x2_bar.t6 GND 0.23fF
C1658 EESPFAL_s0_0/EESPFAL_NAND_v3_2/A_bar GND 0.68fF $ **FLOATING
C1659 x2_bar.n1 GND 2.39fF $ **FLOATING
C1660 x2_bar.t11 GND 0.44fF
C1661 x2_bar.t4 GND 0.25fF
C1662 x2_bar.n2 GND 2.34fF $ **FLOATING
C1663 EESPFAL_s1_0/EESPFAL_XOR_v3_0/A_bar GND 0.26fF $ **FLOATING
C1664 x2_bar.n3 GND 1.09fF $ **FLOATING
C1665 x2_bar.t9 GND 0.15fF
C1666 EESPFAL_s1_0/EESPFAL_INV4_1/A_bar GND 0.54fF $ **FLOATING
C1667 x2_bar.t3 GND 0.18fF
C1668 EESPFAL_s2_0/EESPFAL_4in_NAND_0/D_bar GND 0.46fF $ **FLOATING
C1669 x2_bar.t2 GND 0.21fF
C1670 EESPFAL_s2_0/EESPFAL_INV4_0/A GND 1.09fF $ **FLOATING
C1671 x2_bar.t1 GND 0.57fF
C1672 x2_bar.t8 GND 0.20fF
C1673 x2_bar.n4 GND 1.89fF $ **FLOATING
C1674 EESPFAL_s2_0/EESPFAL_XOR_v3_0/B_bar GND 0.20fF $ **FLOATING
C1675 x2_bar.t10 GND 0.44fF
C1676 x2_bar.t5 GND 0.25fF
C1677 x2_bar.n5 GND 2.34fF $ **FLOATING
C1678 EESPFAL_s3_0/EESPFAL_XOR_v3_1/A_bar GND 0.26fF $ **FLOATING
C1679 x2_bar.t7 GND 0.49fF
C1680 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/A GND 2.23fF $ **FLOATING
C1681 x2_bar.n6 GND 4.71fF $ **FLOATING
C1682 EESPFAL_s3_0/x2_bar GND 2.03fF $ **FLOATING
C1683 EESPFAL_s2_0/x2_bar GND 0.84fF $ **FLOATING
C1684 x2_bar.n7 GND 1.75fF $ **FLOATING
C1685 x2_bar.n8 GND 6.98fF $ **FLOATING
C1686 x2_bar.n9 GND 3.41fF $ **FLOATING
C1687 x2_bar.n10 GND 7.07fF $ **FLOATING
C1688 EESPFAL_s1_0/x2_bar GND 0.94fF $ **FLOATING
C1689 EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT_bar GND 0.35fF $ **FLOATING
C1690 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t9 GND 0.11fF
C1691 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n0 GND 0.43fF $ **FLOATING
C1692 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t1 GND 0.04fF
C1693 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t5 GND 0.04fF
C1694 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n1 GND 0.12fF $ **FLOATING
C1695 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t0 GND 0.15fF
C1696 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t4 GND 0.27fF
C1697 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n2 GND 0.23fF $ **FLOATING
C1698 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n3 GND 0.10fF $ **FLOATING
C1699 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t3 GND 0.04fF
C1700 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t2 GND 0.04fF
C1701 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n4 GND 0.10fF $ **FLOATING
C1702 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n5 GND 0.11fF $ **FLOATING
C1703 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t6 GND 0.04fF
C1704 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t8 GND 0.05fF
C1705 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.t7 GND 0.05fF
C1706 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n6 GND 0.06fF $ **FLOATING
C1707 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A.n7 GND 0.04fF $ **FLOATING
C1708 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t6 GND 0.07fF
C1709 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t1 GND 0.21fF
C1710 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t4 GND 0.05fF
C1711 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t2 GND 0.05fF
C1712 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n0 GND 0.17fF $ **FLOATING
C1713 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t5 GND 0.05fF
C1714 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t3 GND 0.05fF
C1715 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n1 GND 0.15fF $ **FLOATING
C1716 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t7 GND 0.04fF
C1717 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t9 GND 0.07fF
C1718 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t8 GND 0.07fF
C1719 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n2 GND 0.07fF $ **FLOATING
C1720 EESPFAL_s2_0/EESPFAL_XOR_v3_0/OUT GND 0.01fF $ **FLOATING
C1721 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n3 GND 0.04fF $ **FLOATING
C1722 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n4 GND 0.22fF $ **FLOATING
C1723 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n5 GND 0.22fF $ **FLOATING
C1724 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.t0 GND 0.21fF
C1725 EESPFAL_s2_0/EESPFAL_NAND_v3_1/A_bar.n6 GND 0.76fF $ **FLOATING
C1726 EESPFAL_s0_0/x0_bar GND 0.21fF $ **FLOATING
C1727 x0_bar.t9 GND 0.46fF
C1728 x0_bar.t10 GND 0.26fF
C1729 x0_bar.n0 GND 2.48fF $ **FLOATING
C1730 x0_bar.n1 GND 2.62fF $ **FLOATING
C1731 x0_bar.t1 GND 0.60fF
C1732 x0_bar.t6 GND 0.21fF
C1733 x0_bar.n2 GND 2.01fF $ **FLOATING
C1734 EESPFAL_s1_0/EESPFAL_XOR_v3_0/B_bar GND 0.38fF $ **FLOATING
C1735 x0_bar.t7 GND 0.54fF
C1736 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C GND 2.16fF $ **FLOATING
C1737 x0_bar.t4 GND 0.24fF
C1738 EESPFAL_s2_0/EESPFAL_4in_NAND_0/C_bar GND 0.79fF $ **FLOATING
C1739 x0_bar.t5 GND 0.60fF
C1740 x0_bar.t2 GND 0.21fF
C1741 x0_bar.n3 GND 2.01fF $ **FLOATING
C1742 EESPFAL_s2_0/EESPFAL_XOR_v3_1/B_bar GND 0.39fF $ **FLOATING
C1743 x0_bar.t3 GND 0.60fF
C1744 x0_bar.t0 GND 0.21fF
C1745 x0_bar.n4 GND 2.01fF $ **FLOATING
C1746 EESPFAL_s3_0/EESPFAL_XOR_v3_0/B_bar GND 0.38fF $ **FLOATING
C1747 x0_bar.t8 GND 0.23fF
C1748 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B_bar GND 0.87fF $ **FLOATING
C1749 x0_bar.n5 GND 6.64fF $ **FLOATING
C1750 EESPFAL_s3_0/x0_bar GND 0.83fF $ **FLOATING
C1751 EESPFAL_s2_0/x0_bar GND 2.03fF $ **FLOATING
C1752 x0_bar.n6 GND 2.84fF $ **FLOATING
C1753 x0_bar.n7 GND 2.79fF $ **FLOATING
C1754 x0_bar.n8 GND 3.87fF $ **FLOATING
C1755 x0_bar.n9 GND 2.68fF $ **FLOATING
C1756 EESPFAL_s1_0/x0_bar GND 2.34fF $ **FLOATING
C1757 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t7 GND 0.04fF
C1758 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/A_bar GND 0.53fF $ **FLOATING
C1759 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t0 GND 0.04fF
C1760 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t3 GND 0.04fF
C1761 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n0 GND 0.11fF $ **FLOATING
C1762 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t5 GND 0.13fF
C1763 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t4 GND 0.20fF
C1764 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n1 GND 0.19fF $ **FLOATING
C1765 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n2 GND 0.09fF $ **FLOATING
C1766 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t2 GND 0.04fF
C1767 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t1 GND 0.04fF
C1768 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n3 GND 0.09fF $ **FLOATING
C1769 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n4 GND 0.10fF $ **FLOATING
C1770 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t9 GND 0.05fF
C1771 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t8 GND 0.04fF
C1772 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.t6 GND 0.03fF
C1773 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n5 GND 0.05fF $ **FLOATING
C1774 EESPFAL_s1_0/EESPFAL_NAND_v3_0/OUT_bar.n6 GND 0.04fF $ **FLOATING
C1775 EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT_bar GND 0.32fF $ **FLOATING
C1776 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t7 GND 0.07fF
C1777 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t2 GND 0.05fF
C1778 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t5 GND 0.05fF
C1779 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n0 GND 0.16fF $ **FLOATING
C1780 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t0 GND 0.20fF
C1781 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t1 GND 0.34fF
C1782 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n1 GND 0.30fF $ **FLOATING
C1783 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n2 GND 0.13fF $ **FLOATING
C1784 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t4 GND 0.05fF
C1785 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t3 GND 0.05fF
C1786 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n3 GND 0.13fF $ **FLOATING
C1787 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n4 GND 0.14fF $ **FLOATING
C1788 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t8 GND 0.05fF
C1789 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t9 GND 0.07fF
C1790 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.t6 GND 0.06fF
C1791 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n5 GND 0.07fF $ **FLOATING
C1792 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A_bar.n6 GND 0.05fF $ **FLOATING
C1793 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t0 GND 0.04fF
C1794 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t1 GND 0.04fF
C1795 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n0 GND 0.12fF $ **FLOATING
C1796 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t4 GND 0.16fF
C1797 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t8 GND 0.05fF
C1798 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n1 GND 0.77fF $ **FLOATING
C1799 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n2 GND 0.18fF $ **FLOATING
C1800 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n3 GND 0.11fF $ **FLOATING
C1801 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t3 GND 0.04fF
C1802 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t2 GND 0.04fF
C1803 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n4 GND 0.13fF $ **FLOATING
C1804 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n5 GND 0.11fF $ **FLOATING
C1805 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t6 GND 0.06fF
C1806 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t5 GND 0.06fF
C1807 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.t7 GND 0.03fF
C1808 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n6 GND 0.06fF $ **FLOATING
C1809 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C.n7 GND 0.03fF $ **FLOATING
C1810 EESPFAL_s3_0/EESPFAL_INV4_0/OUT_bar GND 0.01fF $ **FLOATING
C1811 EESPFAL_s3_0/EESPFAL_INV4_0/OUT GND 0.23fF $ **FLOATING
C1812 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 GND 0.03fF
C1813 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 GND 0.63fF $ **FLOATING
C1814 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 GND 0.04fF
C1815 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 GND 0.04fF
C1816 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 GND 0.11fF $ **FLOATING
C1817 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 GND 0.25fF
C1818 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 GND 0.04fF
C1819 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 GND 0.04fF
C1820 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 GND 0.13fF $ **FLOATING
C1821 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 GND 0.17fF $ **FLOATING
C1822 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 GND 0.12fF $ **FLOATING
C1823 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 GND 0.06fF
C1824 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 GND 0.05fF
C1825 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 GND 0.04fF
C1826 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 GND 0.06fF $ **FLOATING
C1827 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 GND 0.04fF $ **FLOATING
C1828 EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT_bar GND 0.30fF $ **FLOATING
C1829 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t9 GND 0.12fF
C1830 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t3 GND 0.04fF
C1831 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t1 GND 0.04fF
C1832 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n0 GND 0.13fF $ **FLOATING
C1833 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t2 GND 0.17fF
C1834 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t0 GND 0.29fF
C1835 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n1 GND 0.26fF $ **FLOATING
C1836 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n2 GND 0.11fF $ **FLOATING
C1837 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t4 GND 0.04fF
C1838 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t5 GND 0.04fF
C1839 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n3 GND 0.11fF $ **FLOATING
C1840 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n4 GND 0.12fF $ **FLOATING
C1841 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t6 GND 0.06fF
C1842 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t8 GND 0.05fF
C1843 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.t7 GND 0.04fF
C1844 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n5 GND 0.06fF $ **FLOATING
C1845 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A.n6 GND 0.04fF $ **FLOATING
C1846 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t7 GND 0.08fF
C1847 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t5 GND 0.24fF
C1848 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t2 GND 0.24fF
C1849 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t0 GND 0.05fF
C1850 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t3 GND 0.05fF
C1851 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n0 GND 0.17fF $ **FLOATING
C1852 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t6 GND 0.07fF
C1853 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t9 GND 0.08fF
C1854 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t8 GND 0.04fF
C1855 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n1 GND 0.08fF $ **FLOATING
C1856 EESPFAL_s3_0/EESPFAL_XOR_v3_0/OUT GND 0.01fF $ **FLOATING
C1857 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n2 GND 0.04fF $ **FLOATING
C1858 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t4 GND 0.05fF
C1859 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.t1 GND 0.05fF
C1860 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n3 GND 0.18fF $ **FLOATING
C1861 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n4 GND 0.24fF $ **FLOATING
C1862 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n5 GND 0.24fF $ **FLOATING
C1863 EESPFAL_s3_0/EESPFAL_NAND_v3_0/A_bar.n6 GND 0.52fF $ **FLOATING
C1864 Dis3.t4 GND 0.14fF
C1865 Dis3.t0 GND 0.15fF
C1866 Dis3.n0 GND 0.44fF $ **FLOATING
C1867 Dis3.t2 GND 0.14fF
C1868 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/Dis GND -0.17fF $ **FLOATING
C1869 Dis3.t5 GND 0.15fF
C1870 Dis3.n1 GND 0.72fF $ **FLOATING
C1871 EESPFAL_s3_0/Dis3 GND 3.46fF $ **FLOATING
C1872 EESPFAL_s2_0/Dis3 GND 0.20fF $ **FLOATING
C1873 Dis3.n2 GND 1.38fF $ **FLOATING
C1874 Dis3.t1 GND 0.14fF
C1875 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/Dis GND -0.17fF $ **FLOATING
C1876 Dis3.t6 GND 0.15fF
C1877 Dis3.n3 GND 0.64fF $ **FLOATING
C1878 Dis3.n4 GND 2.12fF $ **FLOATING
C1879 Dis3.t7 GND 0.14fF
C1880 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/Dis GND -0.17fF $ **FLOATING
C1881 Dis3.t3 GND 0.15fF
C1882 Dis3.n5 GND 0.64fF $ **FLOATING
C1883 Dis3.n6 GND 2.14fF $ **FLOATING
C1884 EESPFAL_s1_0/Dis3 GND 2.12fF $ **FLOATING
C1885 Dis3.n7 GND 1.74fF $ **FLOATING
C1886 EESPFAL_s0_0/Dis3 GND 0.03fF $ **FLOATING
C1887 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t9 GND 0.13fF
C1888 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t4 GND 0.21fF
C1889 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t5 GND 0.05fF
C1890 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t1 GND 0.05fF
C1891 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n0 GND 0.16fF $ **FLOATING
C1892 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t3 GND 0.05fF
C1893 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t2 GND 0.05fF
C1894 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n1 GND 0.15fF $ **FLOATING
C1895 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t8 GND 0.04fF
C1896 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t7 GND 0.06fF
C1897 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t6 GND 0.07fF
C1898 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n2 GND 0.07fF $ **FLOATING
C1899 EESPFAL_s1_0/EESPFAL_XOR_v3_1/OUT GND 0.01fF $ **FLOATING
C1900 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n3 GND 0.04fF $ **FLOATING
C1901 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n4 GND 0.22fF $ **FLOATING
C1902 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n5 GND 0.22fF $ **FLOATING
C1903 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.t0 GND 0.21fF
C1904 EESPFAL_s1_0/EESPFAL_NAND_v3_1/A.n6 GND 0.31fF $ **FLOATING
C1905 EESPFAL_s0_0/x3 GND 0.23fF $ **FLOATING
C1906 x3.t2 GND 0.20fF
C1907 x3.t1 GND 0.21fF
C1908 x3.n0 GND 2.43fF $ **FLOATING
C1909 x3.n1 GND 2.19fF $ **FLOATING
C1910 x3.t12 GND 0.21fF
C1911 EESPFAL_s1_0/EESPFAL_INV4_2/A GND 1.05fF $ **FLOATING
C1912 x3.n2 GND 6.53fF $ **FLOATING
C1913 x3.t0 GND 0.21fF
C1914 x3.t9 GND 0.20fF
C1915 x3.n3 GND 2.43fF $ **FLOATING
C1916 EESPFAL_s1_0/EESPFAL_XOR_v3_1/B GND 0.31fF $ **FLOATING
C1917 x3.t11 GND 0.26fF
C1918 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A_bar GND 0.69fF $ **FLOATING
C1919 x3.t3 GND 0.31fF
C1920 EESPFAL_s2_0/EESPFAL_4in_NAND_0/A_bar GND 0.77fF $ **FLOATING
C1921 x3.t10 GND 0.31fF
C1922 x3.t7 GND 0.27fF
C1923 x3.n4 GND 2.34fF $ **FLOATING
C1924 EESPFAL_s2_0/EESPFAL_XOR_v3_0/A GND 0.27fF $ **FLOATING
C1925 x3.t8 GND 0.15fF
C1926 EESPFAL_s3_0/EESPFAL_INV4_2/A_bar GND 0.53fF $ **FLOATING
C1927 x3.t4 GND 0.21fF
C1928 x3.t6 GND 0.20fF
C1929 x3.n5 GND 2.43fF $ **FLOATING
C1930 EESPFAL_s3_0/EESPFAL_XOR_v3_1/B GND 0.31fF $ **FLOATING
C1931 x3.t5 GND 0.50fF
C1932 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C GND 1.83fF $ **FLOATING
C1933 x3.n6 GND 4.21fF $ **FLOATING
C1934 x3.n7 GND 5.01fF $ **FLOATING
C1935 EESPFAL_s3_0/x3 GND 1.02fF $ **FLOATING
C1936 EESPFAL_s2_0/x3 GND 0.57fF $ **FLOATING
C1937 x3.n8 GND 2.35fF $ **FLOATING
C1938 x3.n9 GND 3.60fF $ **FLOATING
C1939 x3.n10 GND 2.40fF $ **FLOATING
C1940 x3.n11 GND 2.40fF $ **FLOATING
C1941 EESPFAL_s1_0/x3 GND 1.36fF $ **FLOATING
C1942 EESPFAL_s1_0/s1_bar GND 0.01fF $ **FLOATING
C1943 s1_bar.t3 GND 0.05fF
C1944 s1_bar.t2 GND 0.05fF
C1945 s1_bar.n0 GND 0.12fF $ **FLOATING
C1946 s1_bar.t0 GND 0.05fF
C1947 s1_bar.t1 GND 0.05fF
C1948 s1_bar.n1 GND 0.14fF $ **FLOATING
C1949 s1_bar.t4 GND 0.27fF
C1950 s1_bar.n2 GND 0.19fF $ **FLOATING
C1951 s1_bar.n3 GND 0.13fF $ **FLOATING
C1952 s1_bar.t7 GND 0.06fF
C1953 s1_bar.t6 GND 0.06fF
C1954 s1_bar.t5 GND 0.04fF
C1955 s1_bar.n4 GND 0.07fF $ **FLOATING
C1956 s1_bar.n5 GND 0.05fF $ **FLOATING
C1957 EESPFAL_s1_0/s1 GND 0.01fF $ **FLOATING
C1958 s1.t2 GND 0.04fF
C1959 s1.t0 GND 0.04fF
C1960 s1.n0 GND 0.15fF $ **FLOATING
C1961 s1.t3 GND 0.19fF
C1962 s1.t5 GND 0.04fF
C1963 s1.t6 GND 0.04fF
C1964 s1.n1 GND 0.14fF $ **FLOATING
C1965 s1.t1 GND 0.04fF
C1966 s1.t4 GND 0.04fF
C1967 s1.n2 GND 0.15fF $ **FLOATING
C1968 s1.t7 GND 0.06fF
C1969 s1.t9 GND 0.06fF
C1970 s1.t8 GND 0.03fF
C1971 s1.n3 GND 0.06fF $ **FLOATING
C1972 s1.n4 GND 0.19fF $ **FLOATING
C1973 s1.n5 GND 0.16fF $ **FLOATING
C1974 s1.n6 GND 0.13fF $ **FLOATING
C1975 EESPFAL_s0_0/x1_bar GND 0.71fF $ **FLOATING
C1976 x1_bar.t8 GND 0.17fF
C1977 x1_bar.n0 GND 4.89fF $ **FLOATING
C1978 x1_bar.t1 GND 0.43fF
C1979 EESPFAL_s0_0/EESPFAL_NAND_v3_2/B GND 1.95fF $ **FLOATING
C1980 x1_bar.n1 GND 1.98fF $ **FLOATING
C1981 x1_bar.t7 GND 0.44fF
C1982 x1_bar.t0 GND 0.25fF
C1983 x1_bar.n2 GND 2.34fF $ **FLOATING
C1984 EESPFAL_s1_0/EESPFAL_XOR_v3_1/A_bar GND 0.34fF $ **FLOATING
C1985 x1_bar.t3 GND 0.22fF
C1986 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B_bar GND 0.69fF $ **FLOATING
C1987 x1_bar.t4 GND 0.27fF
C1988 EESPFAL_s2_0/EESPFAL_4in_NAND_0/B_bar GND 0.78fF $ **FLOATING
C1989 x1_bar.t5 GND 0.44fF
C1990 x1_bar.t6 GND 0.25fF
C1991 x1_bar.n3 GND 2.34fF $ **FLOATING
C1992 EESPFAL_s2_0/EESPFAL_XOR_v3_1/A_bar GND 0.36fF $ **FLOATING
C1993 x1_bar.t9 GND 0.21fF
C1994 EESPFAL_s2_0/EESPFAL_INV4_1/A GND 1.12fF $ **FLOATING
C1995 x1_bar.t2 GND 0.44fF
C1996 x1_bar.t10 GND 0.25fF
C1997 x1_bar.n4 GND 2.34fF $ **FLOATING
C1998 EESPFAL_s3_0/EESPFAL_XOR_v3_0/A_bar GND 0.34fF $ **FLOATING
C1999 x1_bar.t11 GND 0.15fF
C2000 EESPFAL_s3_0/EESPFAL_INV4_1/A_bar GND 0.64fF $ **FLOATING
C2001 EESPFAL_s3_0/x1_bar GND 9.57fF $ **FLOATING
C2002 x1_bar.n5 GND 0.93fF $ **FLOATING
C2003 x1_bar.n6 GND 5.68fF $ **FLOATING
C2004 EESPFAL_s2_0/x1_bar GND 1.47fF $ **FLOATING
C2005 x1_bar.n7 GND 2.52fF $ **FLOATING
C2006 x1_bar.n8 GND 2.26fF $ **FLOATING
C2007 x1_bar.n9 GND 2.41fF $ **FLOATING
C2008 x1_bar.n10 GND 2.56fF $ **FLOATING
C2009 EESPFAL_s1_0/x1_bar GND 2.15fF $ **FLOATING
C2010 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t6 GND 0.12fF
C2011 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t0 GND 0.20fF
C2012 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t1 GND 0.20fF
C2013 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t5 GND 0.05fF
C2014 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t2 GND 0.05fF
C2015 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n0 GND 0.16fF $ **FLOATING
C2016 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t9 GND 0.03fF
C2017 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t8 GND 0.06fF
C2018 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t7 GND 0.07fF
C2019 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n1 GND 0.07fF $ **FLOATING
C2020 EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT GND 0.01fF $ **FLOATING
C2021 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n2 GND 0.03fF $ **FLOATING
C2022 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t4 GND 0.05fF
C2023 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.t3 GND 0.05fF
C2024 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n3 GND 0.14fF $ **FLOATING
C2025 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n4 GND 0.21fF $ **FLOATING
C2026 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n5 GND 0.21fF $ **FLOATING
C2027 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A.n6 GND 0.30fF $ **FLOATING
C2028 CLK3.n0 GND 0.02fF $ **FLOATING
C2029 CLK3.n1 GND 0.02fF $ **FLOATING
C2030 CLK3.n2 GND 0.03fF $ **FLOATING
C2031 CLK3.n3 GND 0.06fF $ **FLOATING
C2032 CLK3.n4 GND 0.03fF $ **FLOATING
C2033 CLK3.n5 GND 0.02fF $ **FLOATING
C2034 CLK3.t28 GND 0.03fF
C2035 CLK3.t10 GND 0.03fF
C2036 CLK3.n6 GND 0.16fF $ **FLOATING
C2037 CLK3.n7 GND 0.03fF $ **FLOATING
C2038 CLK3.n8 GND 0.02fF $ **FLOATING
C2039 CLK3.n9 GND 0.03fF $ **FLOATING
C2040 CLK3.n10 GND 0.11fF $ **FLOATING
C2041 CLK3.n11 GND 0.03fF $ **FLOATING
C2042 CLK3.n12 GND 0.02fF $ **FLOATING
C2043 CLK3.t21 GND 0.05fF
C2044 CLK3.n13 GND 0.03fF $ **FLOATING
C2045 CLK3.n14 GND 0.02fF $ **FLOATING
C2046 CLK3.n15 GND 0.03fF $ **FLOATING
C2047 CLK3.t24 GND 0.09fF
C2048 CLK3.n16 GND 0.03fF $ **FLOATING
C2049 CLK3.n17 GND 0.02fF $ **FLOATING
C2050 CLK3.t25 GND 0.03fF
C2051 CLK3.t19 GND 0.03fF
C2052 CLK3.n18 GND 0.10fF $ **FLOATING
C2053 CLK3.n19 GND 0.03fF $ **FLOATING
C2054 CLK3.n20 GND 0.02fF $ **FLOATING
C2055 CLK3.n21 GND 0.03fF $ **FLOATING
C2056 CLK3.n22 GND 0.14fF $ **FLOATING
C2057 CLK3.n23 GND 0.03fF $ **FLOATING
C2058 CLK3.n24 GND 0.02fF $ **FLOATING
C2059 CLK3.n25 GND 0.03fF $ **FLOATING
C2060 CLK3.n26 GND 0.02fF $ **FLOATING
C2061 CLK3.n27 GND 0.03fF $ **FLOATING
C2062 CLK3.n28 GND 0.07fF $ **FLOATING
C2063 CLK3.n29 GND 0.03fF $ **FLOATING
C2064 CLK3.n30 GND 0.02fF $ **FLOATING
C2065 CLK3.t23 GND 0.08fF
C2066 CLK3.n31 GND 0.13fF $ **FLOATING
C2067 CLK3.n32 GND 0.36fF $ **FLOATING
C2068 CLK3.n33 GND 0.03fF $ **FLOATING
C2069 CLK3.n34 GND 0.03fF $ **FLOATING
C2070 CLK3.n35 GND 0.02fF $ **FLOATING
C2071 CLK3.n36 GND 0.03fF $ **FLOATING
C2072 CLK3.n37 GND 0.06fF $ **FLOATING
C2073 CLK3.n38 GND 0.06fF $ **FLOATING
C2074 CLK3.n39 GND 0.06fF $ **FLOATING
C2075 CLK3.n40 GND 0.03fF $ **FLOATING
C2076 CLK3.n41 GND 0.02fF $ **FLOATING
C2077 CLK3.n42 GND 0.03fF $ **FLOATING
C2078 CLK3.n43 GND 0.03fF $ **FLOATING
C2079 CLK3.t27 GND 0.05fF
C2080 CLK3.n44 GND 0.30fF $ **FLOATING
C2081 CLK3.n45 GND 0.02fF $ **FLOATING
C2082 CLK3.n46 GND 0.02fF $ **FLOATING
C2083 CLK3.n47 GND 0.03fF $ **FLOATING
C2084 CLK3.n48 GND 0.18fF $ **FLOATING
C2085 CLK3.n49 GND 0.11fF $ **FLOATING
C2086 CLK3.t26 GND 0.09fF
C2087 CLK3.n50 GND 0.10fF $ **FLOATING
C2088 CLK3.n51 GND 0.16fF $ **FLOATING
C2089 CLK3.n52 GND 0.03fF $ **FLOATING
C2090 CLK3.n53 GND 0.02fF $ **FLOATING
C2091 CLK3.n54 GND 0.03fF $ **FLOATING
C2092 CLK3.n55 GND 0.03fF $ **FLOATING
C2093 CLK3.n56 GND 0.18fF $ **FLOATING
C2094 CLK3.n57 GND 0.02fF $ **FLOATING
C2095 CLK3.n58 GND 0.03fF $ **FLOATING
C2096 CLK3.n59 GND 0.17fF $ **FLOATING
C2097 CLK3.t18 GND 0.09fF
C2098 CLK3.n60 GND 0.10fF $ **FLOATING
C2099 CLK3.t20 GND 0.09fF
C2100 CLK3.n61 GND 0.16fF $ **FLOATING
C2101 CLK3.n62 GND 0.03fF $ **FLOATING
C2102 CLK3.n63 GND 0.02fF $ **FLOATING
C2103 CLK3.n64 GND 0.03fF $ **FLOATING
C2104 CLK3.n65 GND 0.03fF $ **FLOATING
C2105 CLK3.n66 GND 0.30fF $ **FLOATING
C2106 CLK3.n67 GND 0.02fF $ **FLOATING
C2107 CLK3.n68 GND 0.02fF $ **FLOATING
C2108 CLK3.n69 GND 0.03fF $ **FLOATING
C2109 CLK3.n70 GND 0.18fF $ **FLOATING
C2110 CLK3.n71 GND 0.14fF $ **FLOATING
C2111 CLK3.n72 GND 0.06fF $ **FLOATING
C2112 CLK3.n73 GND 0.03fF $ **FLOATING
C2113 CLK3.n74 GND 0.02fF $ **FLOATING
C2114 CLK3.n75 GND 0.03fF $ **FLOATING
C2115 CLK3.n76 GND 0.03fF $ **FLOATING
C2116 CLK3.n77 GND 0.19fF $ **FLOATING
C2117 CLK3.n78 GND 0.01fF $ **FLOATING
C2118 CLK3.n79 GND 0.13fF $ **FLOATING
C2119 CLK3.t1 GND 0.08fF
C2120 CLK3.n80 GND 0.03fF $ **FLOATING
C2121 CLK3.n81 GND 0.02fF $ **FLOATING
C2122 CLK3.n82 GND 0.03fF $ **FLOATING
C2123 CLK3.n83 GND 0.06fF $ **FLOATING
C2124 CLK3.n84 GND 0.03fF $ **FLOATING
C2125 CLK3.n85 GND 0.02fF $ **FLOATING
C2126 CLK3.t15 GND 0.03fF
C2127 CLK3.t11 GND 0.03fF
C2128 CLK3.n86 GND 0.16fF $ **FLOATING
C2129 CLK3.n87 GND 0.03fF $ **FLOATING
C2130 CLK3.n88 GND 0.02fF $ **FLOATING
C2131 CLK3.n89 GND 0.03fF $ **FLOATING
C2132 CLK3.n90 GND 0.18fF $ **FLOATING
C2133 CLK3.n91 GND 0.03fF $ **FLOATING
C2134 CLK3.n92 GND 0.02fF $ **FLOATING
C2135 CLK3.t35 GND 0.05fF
C2136 CLK3.n93 GND 0.03fF $ **FLOATING
C2137 CLK3.n94 GND 0.02fF $ **FLOATING
C2138 CLK3.n95 GND 0.03fF $ **FLOATING
C2139 CLK3.t32 GND 0.09fF
C2140 CLK3.n96 GND 0.03fF $ **FLOATING
C2141 CLK3.n97 GND 0.02fF $ **FLOATING
C2142 CLK3.t44 GND 0.03fF
C2143 CLK3.t33 GND 0.03fF
C2144 CLK3.n98 GND 0.10fF $ **FLOATING
C2145 CLK3.n99 GND 0.03fF $ **FLOATING
C2146 CLK3.n100 GND 0.02fF $ **FLOATING
C2147 CLK3.n101 GND 0.03fF $ **FLOATING
C2148 CLK3.n102 GND 0.18fF $ **FLOATING
C2149 CLK3.n103 GND 0.03fF $ **FLOATING
C2150 CLK3.n104 GND 0.02fF $ **FLOATING
C2151 CLK3.t42 GND 0.05fF
C2152 CLK3.n105 GND 0.03fF $ **FLOATING
C2153 CLK3.n106 GND 0.02fF $ **FLOATING
C2154 CLK3.n107 GND 0.03fF $ **FLOATING
C2155 CLK3.n108 GND 0.06fF $ **FLOATING
C2156 CLK3.n109 GND 0.03fF $ **FLOATING
C2157 CLK3.n110 GND 0.02fF $ **FLOATING
C2158 CLK3.n111 GND 0.03fF $ **FLOATING
C2159 CLK3.n112 GND 0.02fF $ **FLOATING
C2160 CLK3.n113 GND 0.03fF $ **FLOATING
C2161 CLK3.n114 GND 0.13fF $ **FLOATING
C2162 CLK3.n115 GND 0.02fF $ **FLOATING
C2163 CLK3.n116 GND 0.02fF $ **FLOATING
C2164 CLK3.n117 GND 0.02fF $ **FLOATING
C2165 CLK3.t38 GND 0.03fF
C2166 CLK3.n118 GND 0.13fF $ **FLOATING
C2167 CLK3.n119 GND 0.03fF $ **FLOATING
C2168 CLK3.n120 GND 0.02fF $ **FLOATING
C2169 CLK3.n121 GND 0.03fF $ **FLOATING
C2170 CLK3.n122 GND 0.06fF $ **FLOATING
C2171 CLK3.n123 GND 0.03fF $ **FLOATING
C2172 CLK3.n124 GND 0.02fF $ **FLOATING
C2173 CLK3.n125 GND 0.03fF $ **FLOATING
C2174 CLK3.n126 GND 0.02fF $ **FLOATING
C2175 CLK3.n127 GND 0.03fF $ **FLOATING
C2176 CLK3.n128 GND 0.18fF $ **FLOATING
C2177 CLK3.n129 GND 0.03fF $ **FLOATING
C2178 CLK3.n130 GND 0.02fF $ **FLOATING
C2179 CLK3.t13 GND 0.05fF
C2180 CLK3.n131 GND 0.03fF $ **FLOATING
C2181 CLK3.n132 GND 0.02fF $ **FLOATING
C2182 CLK3.n133 GND 0.03fF $ **FLOATING
C2183 CLK3.t36 GND 0.09fF
C2184 CLK3.n134 GND 0.03fF $ **FLOATING
C2185 CLK3.n135 GND 0.02fF $ **FLOATING
C2186 CLK3.t37 GND 0.03fF
C2187 CLK3.t17 GND 0.03fF
C2188 CLK3.n136 GND 0.10fF $ **FLOATING
C2189 CLK3.n137 GND 0.03fF $ **FLOATING
C2190 CLK3.n138 GND 0.02fF $ **FLOATING
C2191 CLK3.n139 GND 0.03fF $ **FLOATING
C2192 CLK3.n140 GND 0.17fF $ **FLOATING
C2193 CLK3.t16 GND 0.09fF
C2194 CLK3.n141 GND 0.18fF $ **FLOATING
C2195 CLK3.n142 GND 0.03fF $ **FLOATING
C2196 CLK3.n143 GND 0.02fF $ **FLOATING
C2197 CLK3.t3 GND 0.05fF
C2198 CLK3.n144 GND 0.03fF $ **FLOATING
C2199 CLK3.n145 GND 0.02fF $ **FLOATING
C2200 CLK3.n146 GND 0.03fF $ **FLOATING
C2201 CLK3.n147 GND 0.06fF $ **FLOATING
C2202 CLK3.n148 GND 0.03fF $ **FLOATING
C2203 CLK3.n149 GND 0.02fF $ **FLOATING
C2204 CLK3.t22 GND 0.03fF
C2205 CLK3.t29 GND 0.03fF
C2206 CLK3.n150 GND 0.16fF $ **FLOATING
C2207 CLK3.n151 GND 0.03fF $ **FLOATING
C2208 CLK3.n152 GND 0.02fF $ **FLOATING
C2209 CLK3.n153 GND 0.03fF $ **FLOATING
C2210 CLK3.n154 GND 0.13fF $ **FLOATING
C2211 CLK3.n155 GND 0.01fF $ **FLOATING
C2212 CLK3.n156 GND 0.01fF $ **FLOATING
C2213 CLK3.n157 GND 0.01fF $ **FLOATING
C2214 CLK3.n158 GND 0.13fF $ **FLOATING
C2215 CLK3.t39 GND 0.08fF
C2216 CLK3.n159 GND 0.03fF $ **FLOATING
C2217 CLK3.n160 GND 0.02fF $ **FLOATING
C2218 CLK3.n161 GND 0.03fF $ **FLOATING
C2219 CLK3.n162 GND 0.06fF $ **FLOATING
C2220 CLK3.n163 GND 0.03fF $ **FLOATING
C2221 CLK3.n164 GND 0.02fF $ **FLOATING
C2222 CLK3.t40 GND 0.03fF
C2223 CLK3.t9 GND 0.03fF
C2224 CLK3.n165 GND 0.16fF $ **FLOATING
C2225 CLK3.n166 GND 0.03fF $ **FLOATING
C2226 CLK3.n167 GND 0.02fF $ **FLOATING
C2227 CLK3.n168 GND 0.03fF $ **FLOATING
C2228 CLK3.n169 GND 0.18fF $ **FLOATING
C2229 CLK3.n170 GND 0.03fF $ **FLOATING
C2230 CLK3.n171 GND 0.02fF $ **FLOATING
C2231 CLK3.t8 GND 0.05fF
C2232 CLK3.n172 GND 0.03fF $ **FLOATING
C2233 CLK3.n173 GND 0.02fF $ **FLOATING
C2234 CLK3.n174 GND 0.03fF $ **FLOATING
C2235 CLK3.t30 GND 0.09fF
C2236 CLK3.n175 GND 0.03fF $ **FLOATING
C2237 CLK3.n176 GND 0.02fF $ **FLOATING
C2238 CLK3.t46 GND 0.03fF
C2239 CLK3.t31 GND 0.03fF
C2240 CLK3.n177 GND 0.10fF $ **FLOATING
C2241 CLK3.n178 GND 0.03fF $ **FLOATING
C2242 CLK3.n179 GND 0.02fF $ **FLOATING
C2243 CLK3.n180 GND 0.03fF $ **FLOATING
C2244 CLK3.n181 GND 0.18fF $ **FLOATING
C2245 CLK3.n182 GND 0.03fF $ **FLOATING
C2246 CLK3.n183 GND 0.02fF $ **FLOATING
C2247 CLK3.t6 GND 0.05fF
C2248 CLK3.n184 GND 0.03fF $ **FLOATING
C2249 CLK3.n185 GND 0.02fF $ **FLOATING
C2250 CLK3.n186 GND 0.03fF $ **FLOATING
C2251 CLK3.n187 GND 0.06fF $ **FLOATING
C2252 CLK3.n188 GND 0.03fF $ **FLOATING
C2253 CLK3.n189 GND 0.02fF $ **FLOATING
C2254 CLK3.n190 GND 0.03fF $ **FLOATING
C2255 CLK3.n191 GND 0.02fF $ **FLOATING
C2256 CLK3.n192 GND 0.03fF $ **FLOATING
C2257 CLK3.n193 GND 0.13fF $ **FLOATING
C2258 CLK3.t14 GND 0.08fF
C2259 CLK3.n194 GND 0.36fF $ **FLOATING
C2260 CLK3.n195 GND 0.03fF $ **FLOATING
C2261 CLK3.n196 GND 0.02fF $ **FLOATING
C2262 CLK3.n197 GND 0.03fF $ **FLOATING
C2263 CLK3.n198 GND 0.07fF $ **FLOATING
C2264 CLK3.n199 GND 0.06fF $ **FLOATING
C2265 CLK3.n200 GND 0.06fF $ **FLOATING
C2266 CLK3.n201 GND 0.03fF $ **FLOATING
C2267 CLK3.n202 GND 0.02fF $ **FLOATING
C2268 CLK3.n203 GND 0.03fF $ **FLOATING
C2269 CLK3.n204 GND 0.03fF $ **FLOATING
C2270 CLK3.n205 GND 0.03fF $ **FLOATING
C2271 CLK3.n206 GND 0.02fF $ **FLOATING
C2272 CLK3.n207 GND 0.03fF $ **FLOATING
C2273 CLK3.n208 GND 0.06fF $ **FLOATING
C2274 CLK3.n209 GND 0.06fF $ **FLOATING
C2275 CLK3.n210 GND 0.14fF $ **FLOATING
C2276 CLK3.n211 GND 0.03fF $ **FLOATING
C2277 CLK3.n212 GND 0.02fF $ **FLOATING
C2278 CLK3.n213 GND 0.03fF $ **FLOATING
C2279 CLK3.n214 GND 0.02fF $ **FLOATING
C2280 CLK3.n215 GND 0.30fF $ **FLOATING
C2281 CLK3.n216 GND 0.03fF $ **FLOATING
C2282 CLK3.n217 GND 0.02fF $ **FLOATING
C2283 CLK3.n218 GND 0.03fF $ **FLOATING
C2284 CLK3.n219 GND 0.11fF $ **FLOATING
C2285 CLK3.t5 GND 0.09fF
C2286 CLK3.n220 GND 0.16fF $ **FLOATING
C2287 CLK3.n221 GND 0.17fF $ **FLOATING
C2288 CLK3.t45 GND 0.09fF
C2289 CLK3.n222 GND 0.10fF $ **FLOATING
C2290 CLK3.n223 GND 0.03fF $ **FLOATING
C2291 CLK3.n224 GND 0.02fF $ **FLOATING
C2292 CLK3.n225 GND 0.03fF $ **FLOATING
C2293 CLK3.n226 GND 0.18fF $ **FLOATING
C2294 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/CLK GND 0.02fF $ **FLOATING
C2295 CLK3.n227 GND 0.03fF $ **FLOATING
C2296 CLK3.n228 GND 0.02fF $ **FLOATING
C2297 CLK3.n229 GND 0.03fF $ **FLOATING
C2298 CLK3.n230 GND 0.10fF $ **FLOATING
C2299 CLK3.n231 GND 0.16fF $ **FLOATING
C2300 CLK3.t7 GND 0.09fF
C2301 CLK3.n232 GND 0.11fF $ **FLOATING
C2302 CLK3.n233 GND 0.03fF $ **FLOATING
C2303 CLK3.n234 GND 0.02fF $ **FLOATING
C2304 CLK3.n235 GND 0.03fF $ **FLOATING
C2305 CLK3.n236 GND 0.30fF $ **FLOATING
C2306 CLK3.n237 GND 0.02fF $ **FLOATING
C2307 CLK3.n238 GND 0.03fF $ **FLOATING
C2308 CLK3.n239 GND 0.02fF $ **FLOATING
C2309 CLK3.n240 GND 0.03fF $ **FLOATING
C2310 CLK3.n241 GND 0.14fF $ **FLOATING
C2311 CLK3.n242 GND 0.06fF $ **FLOATING
C2312 CLK3.n243 GND 0.06fF $ **FLOATING
C2313 CLK3.n244 GND 0.03fF $ **FLOATING
C2314 CLK3.n245 GND 0.02fF $ **FLOATING
C2315 CLK3.n246 GND 0.03fF $ **FLOATING
C2316 CLK3.n247 GND 0.19fF $ **FLOATING
C2317 CLK3.n248 GND 0.02fF $ **FLOATING
C2318 CLK3.n249 GND 0.03fF $ **FLOATING
C2319 CLK3.n250 GND 0.02fF $ **FLOATING
C2320 CLK3.n251 GND 0.03fF $ **FLOATING
C2321 CLK3.n252 GND 0.06fF $ **FLOATING
C2322 CLK3.n253 GND 0.06fF $ **FLOATING
C2323 CLK3.n254 GND 0.07fF $ **FLOATING
C2324 CLK3.n255 GND 0.03fF $ **FLOATING
C2325 CLK3.n256 GND 0.02fF $ **FLOATING
C2326 CLK3.n257 GND 0.03fF $ **FLOATING
C2327 CLK3.n258 GND 0.34fF $ **FLOATING
C2328 CLK3.n259 GND 0.41fF $ **FLOATING
C2329 EESPFAL_s3_0/CLK3 GND 0.61fF $ **FLOATING
C2330 EESPFAL_s2_0/CLK3 GND 0.55fF $ **FLOATING
C2331 CLK3.n260 GND 0.44fF $ **FLOATING
C2332 CLK3.n261 GND 0.01fF $ **FLOATING
C2333 CLK3.n262 GND 0.02fF $ **FLOATING
C2334 CLK3.n263 GND 0.00fF $ **FLOATING
C2335 CLK3.t0 GND 0.08fF
C2336 CLK3.n264 GND 0.36fF $ **FLOATING
C2337 CLK3.n265 GND 0.01fF $ **FLOATING
C2338 CLK3.n266 GND 0.00fF $ **FLOATING
C2339 CLK3.n267 GND 0.00fF $ **FLOATING
C2340 CLK3.n268 GND 0.03fF $ **FLOATING
C2341 CLK3.n269 GND 0.07fF $ **FLOATING
C2342 CLK3.n270 GND 0.06fF $ **FLOATING
C2343 CLK3.n271 GND 0.06fF $ **FLOATING
C2344 CLK3.n272 GND 0.03fF $ **FLOATING
C2345 CLK3.n273 GND 0.02fF $ **FLOATING
C2346 CLK3.n274 GND 0.03fF $ **FLOATING
C2347 CLK3.n275 GND 0.02fF $ **FLOATING
C2348 CLK3.n276 GND 0.19fF $ **FLOATING
C2349 CLK3.n277 GND 0.03fF $ **FLOATING
C2350 CLK3.n278 GND 0.02fF $ **FLOATING
C2351 CLK3.n279 GND 0.03fF $ **FLOATING
C2352 CLK3.n280 GND 0.06fF $ **FLOATING
C2353 CLK3.n281 GND 0.06fF $ **FLOATING
C2354 CLK3.n282 GND 0.14fF $ **FLOATING
C2355 CLK3.n283 GND 0.03fF $ **FLOATING
C2356 CLK3.n284 GND 0.02fF $ **FLOATING
C2357 CLK3.n285 GND 0.03fF $ **FLOATING
C2358 CLK3.n286 GND 0.02fF $ **FLOATING
C2359 CLK3.n287 GND 0.30fF $ **FLOATING
C2360 CLK3.n288 GND 0.03fF $ **FLOATING
C2361 CLK3.n289 GND 0.02fF $ **FLOATING
C2362 CLK3.n290 GND 0.03fF $ **FLOATING
C2363 CLK3.n291 GND 0.11fF $ **FLOATING
C2364 CLK3.t2 GND 0.09fF
C2365 CLK3.n292 GND 0.16fF $ **FLOATING
C2366 CLK3.n293 GND 0.10fF $ **FLOATING
C2367 CLK3.n294 GND 0.03fF $ **FLOATING
C2368 CLK3.n295 GND 0.02fF $ **FLOATING
C2369 CLK3.n296 GND 0.03fF $ **FLOATING
C2370 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/CLK GND 0.02fF $ **FLOATING
C2371 CLK3.n297 GND 0.18fF $ **FLOATING
C2372 CLK3.n298 GND 0.03fF $ **FLOATING
C2373 CLK3.n299 GND 0.02fF $ **FLOATING
C2374 CLK3.n300 GND 0.03fF $ **FLOATING
C2375 CLK3.n301 GND 0.10fF $ **FLOATING
C2376 CLK3.n302 GND 0.16fF $ **FLOATING
C2377 CLK3.t12 GND 0.09fF
C2378 CLK3.n303 GND 0.11fF $ **FLOATING
C2379 CLK3.n304 GND 0.03fF $ **FLOATING
C2380 CLK3.n305 GND 0.02fF $ **FLOATING
C2381 CLK3.n306 GND 0.03fF $ **FLOATING
C2382 CLK3.n307 GND 0.30fF $ **FLOATING
C2383 CLK3.n308 GND 0.02fF $ **FLOATING
C2384 CLK3.n309 GND 0.03fF $ **FLOATING
C2385 CLK3.n310 GND 0.02fF $ **FLOATING
C2386 CLK3.n311 GND 0.03fF $ **FLOATING
C2387 CLK3.n312 GND 0.14fF $ **FLOATING
C2388 CLK3.n313 GND 0.06fF $ **FLOATING
C2389 CLK3.n314 GND 0.06fF $ **FLOATING
C2390 CLK3.n315 GND 0.03fF $ **FLOATING
C2391 CLK3.n316 GND 0.02fF $ **FLOATING
C2392 CLK3.n317 GND 0.03fF $ **FLOATING
C2393 CLK3.n318 GND 0.03fF $ **FLOATING
C2394 CLK3.n319 GND 0.03fF $ **FLOATING
C2395 CLK3.n320 GND 0.02fF $ **FLOATING
C2396 CLK3.n321 GND 0.03fF $ **FLOATING
C2397 CLK3.n322 GND 0.06fF $ **FLOATING
C2398 CLK3.n323 GND 0.06fF $ **FLOATING
C2399 CLK3.n324 GND 0.07fF $ **FLOATING
C2400 CLK3.n325 GND 0.03fF $ **FLOATING
C2401 CLK3.n326 GND 0.02fF $ **FLOATING
C2402 CLK3.n327 GND 0.03fF $ **FLOATING
C2403 CLK3.n328 GND 0.09fF $ **FLOATING
C2404 CLK3.n329 GND 0.08fF $ **FLOATING
C2405 CLK3.n330 GND 0.03fF $ **FLOATING
C2406 CLK3.n331 GND 0.10fF $ **FLOATING
C2407 CLK3.n332 GND 0.01fF $ **FLOATING
C2408 CLK3.n333 GND 0.12fF $ **FLOATING
C2409 CLK3.n334 GND 0.10fF $ **FLOATING
C2410 CLK3.t4 GND 0.03fF
C2411 CLK3.n335 GND 0.10fF $ **FLOATING
C2412 CLK3.n336 GND 0.02fF $ **FLOATING
C2413 CLK3.n337 GND 0.02fF $ **FLOATING
C2414 CLK3.n338 GND 0.02fF $ **FLOATING
C2415 CLK3.n339 GND 0.09fF $ **FLOATING
C2416 CLK3.n340 GND 0.09fF $ **FLOATING
C2417 CLK3.n341 GND 0.03fF $ **FLOATING
C2418 CLK3.n342 GND 0.02fF $ **FLOATING
C2419 CLK3.n343 GND 0.03fF $ **FLOATING
C2420 CLK3.n344 GND 0.07fF $ **FLOATING
C2421 CLK3.n345 GND 0.06fF $ **FLOATING
C2422 CLK3.n346 GND 0.06fF $ **FLOATING
C2423 CLK3.n347 GND 0.03fF $ **FLOATING
C2424 CLK3.n348 GND 0.02fF $ **FLOATING
C2425 CLK3.n349 GND 0.03fF $ **FLOATING
C2426 CLK3.n350 GND 0.03fF $ **FLOATING
C2427 CLK3.n351 GND 0.03fF $ **FLOATING
C2428 CLK3.n352 GND 0.02fF $ **FLOATING
C2429 CLK3.n353 GND 0.03fF $ **FLOATING
C2430 CLK3.n354 GND 0.06fF $ **FLOATING
C2431 CLK3.n355 GND 0.06fF $ **FLOATING
C2432 CLK3.n356 GND 0.14fF $ **FLOATING
C2433 CLK3.n357 GND 0.03fF $ **FLOATING
C2434 CLK3.n358 GND 0.02fF $ **FLOATING
C2435 CLK3.n359 GND 0.03fF $ **FLOATING
C2436 CLK3.n360 GND 0.02fF $ **FLOATING
C2437 CLK3.n361 GND 0.30fF $ **FLOATING
C2438 CLK3.n362 GND 0.03fF $ **FLOATING
C2439 CLK3.n363 GND 0.02fF $ **FLOATING
C2440 CLK3.n364 GND 0.03fF $ **FLOATING
C2441 CLK3.n365 GND 0.11fF $ **FLOATING
C2442 CLK3.t41 GND 0.09fF
C2443 CLK3.n366 GND 0.16fF $ **FLOATING
C2444 CLK3.n367 GND 0.17fF $ **FLOATING
C2445 CLK3.t43 GND 0.09fF
C2446 CLK3.n368 GND 0.10fF $ **FLOATING
C2447 CLK3.n369 GND 0.03fF $ **FLOATING
C2448 CLK3.n370 GND 0.02fF $ **FLOATING
C2449 CLK3.n371 GND 0.03fF $ **FLOATING
C2450 CLK3.n372 GND 0.18fF $ **FLOATING
C2451 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/CLK GND 0.02fF $ **FLOATING
C2452 CLK3.n373 GND 0.03fF $ **FLOATING
C2453 CLK3.n374 GND 0.02fF $ **FLOATING
C2454 CLK3.n375 GND 0.03fF $ **FLOATING
C2455 CLK3.n376 GND 0.10fF $ **FLOATING
C2456 CLK3.n377 GND 0.16fF $ **FLOATING
C2457 CLK3.t34 GND 0.09fF
C2458 CLK3.n378 GND 0.11fF $ **FLOATING
C2459 CLK3.n379 GND 0.03fF $ **FLOATING
C2460 CLK3.n380 GND 0.02fF $ **FLOATING
C2461 CLK3.n381 GND 0.03fF $ **FLOATING
C2462 CLK3.n382 GND 0.30fF $ **FLOATING
C2463 CLK3.n383 GND 0.02fF $ **FLOATING
C2464 CLK3.n384 GND 0.03fF $ **FLOATING
C2465 CLK3.n385 GND 0.02fF $ **FLOATING
C2466 CLK3.n386 GND 0.03fF $ **FLOATING
C2467 CLK3.n387 GND 0.14fF $ **FLOATING
C2468 CLK3.n388 GND 0.06fF $ **FLOATING
C2469 CLK3.n389 GND 0.06fF $ **FLOATING
C2470 CLK3.n390 GND 0.03fF $ **FLOATING
C2471 CLK3.n391 GND 0.02fF $ **FLOATING
C2472 CLK3.n392 GND 0.03fF $ **FLOATING
C2473 CLK3.n393 GND 0.19fF $ **FLOATING
C2474 CLK3.n394 GND 0.02fF $ **FLOATING
C2475 CLK3.n395 GND 0.03fF $ **FLOATING
C2476 CLK3.n396 GND 0.02fF $ **FLOATING
C2477 CLK3.n397 GND 0.03fF $ **FLOATING
C2478 CLK3.n398 GND 0.06fF $ **FLOATING
C2479 CLK3.n399 GND 0.06fF $ **FLOATING
C2480 CLK3.n400 GND 0.07fF $ **FLOATING
C2481 CLK3.n401 GND 0.03fF $ **FLOATING
C2482 CLK3.n402 GND 0.02fF $ **FLOATING
C2483 CLK3.n403 GND 0.03fF $ **FLOATING
C2484 CLK3.n404 GND 0.34fF $ **FLOATING
C2485 CLK3.n405 GND 0.39fF $ **FLOATING
C2486 EESPFAL_s1_0/CLK3 GND 0.03fF $ **FLOATING
C2487 CLK3.n406 GND 0.58fF $ **FLOATING
C2488 CLK3.n407 GND 0.34fF $ **FLOATING
C2489 CLK3.n408 GND 0.02fF $ **FLOATING
C2490 CLK3.n409 GND 0.02fF $ **FLOATING
C2491 CLK3.n410 GND 0.01fF $ **FLOATING
C2492 CLK3.n411 GND 0.02fF $ **FLOATING
C2493 CLK3.n412 GND 0.03fF $ **FLOATING
C2494 CLK3.n413 GND 0.06fF $ **FLOATING
C2495 CLK3.n414 GND 0.07fF $ **FLOATING
C2496 CLK3.n415 GND 0.13fF $ **FLOATING
C2497 CLK3.n416 GND 0.25fF $ **FLOATING
C2498 EESPFAL_s0_0/CLK3 GND 0.01fF $ **FLOATING
C2499 x0.t6 GND 0.29fF
C2500 x0.t10 GND 0.25fF
C2501 x0.n0 GND 2.19fF $ **FLOATING
C2502 EESPFAL_s0_0/x0 GND 2.43fF $ **FLOATING
C2503 x0.t5 GND 0.20fF
C2504 x0.t3 GND 0.19fF
C2505 x0.n1 GND 2.28fF $ **FLOATING
C2506 EESPFAL_s1_0/EESPFAL_XOR_v3_0/B GND 0.52fF $ **FLOATING
C2507 x0.t2 GND 0.16fF
C2508 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/C_bar GND 0.64fF $ **FLOATING
C2509 x0.t7 GND 0.31fF
C2510 EESPFAL_s2_0/EESPFAL_4in_NAND_0/C GND 2.53fF $ **FLOATING
C2511 x0.t0 GND 0.20fF
C2512 x0.t1 GND 0.19fF
C2513 x0.n2 GND 2.28fF $ **FLOATING
C2514 EESPFAL_s2_0/EESPFAL_XOR_v3_1/B GND 0.53fF $ **FLOATING
C2515 x0.t8 GND 0.20fF
C2516 x0.t4 GND 0.19fF
C2517 x0.n3 GND 2.28fF $ **FLOATING
C2518 EESPFAL_s3_0/EESPFAL_XOR_v3_0/B GND 0.52fF $ **FLOATING
C2519 x0.t9 GND 0.48fF
C2520 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/B GND 2.10fF $ **FLOATING
C2521 x0.n4 GND 6.00fF $ **FLOATING
C2522 EESPFAL_s3_0/x0 GND 0.62fF $ **FLOATING
C2523 EESPFAL_s2_0/x0 GND 1.81fF $ **FLOATING
C2524 x0.n5 GND 2.31fF $ **FLOATING
C2525 x0.n6 GND 2.22fF $ **FLOATING
C2526 x0.n7 GND 3.77fF $ **FLOATING
C2527 x0.n8 GND 2.61fF $ **FLOATING
C2528 EESPFAL_s1_0/x0 GND 2.01fF $ **FLOATING
C2529 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t6 GND 0.04fF
C2530 EESPFAL_s2_0/EESPFAL_3in_NOR_v2_0/A_bar GND 0.53fF $ **FLOATING
C2531 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t0 GND 0.04fF
C2532 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t3 GND 0.04fF
C2533 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n0 GND 0.11fF $ **FLOATING
C2534 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t4 GND 0.14fF
C2535 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t5 GND 0.20fF
C2536 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n1 GND 0.19fF $ **FLOATING
C2537 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n2 GND 0.09fF $ **FLOATING
C2538 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t1 GND 0.04fF
C2539 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t2 GND 0.04fF
C2540 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n3 GND 0.09fF $ **FLOATING
C2541 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n4 GND 0.10fF $ **FLOATING
C2542 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t8 GND 0.03fF
C2543 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t7 GND 0.05fF
C2544 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.t9 GND 0.04fF
C2545 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n5 GND 0.05fF $ **FLOATING
C2546 EESPFAL_s2_0/EESPFAL_NAND_v3_1/OUT_bar.n6 GND 0.04fF $ **FLOATING
C2547 Dis2.t13 GND 0.24fF
C2548 Dis2.t5 GND 0.15fF
C2549 Dis2.n0 GND 0.61fF $ **FLOATING
C2550 Dis2.t8 GND 0.15fF
C2551 Dis2.t15 GND 0.15fF
C2552 EESPFAL_s2_0/EESPFAL_INV4_2/Dis GND -0.29fF $ **FLOATING
C2553 Dis2.n1 GND 0.32fF $ **FLOATING
C2554 Dis2.n2 GND 0.55fF $ **FLOATING
C2555 Dis2.t12 GND 0.15fF
C2556 Dis2.t17 GND 0.15fF
C2557 EESPFAL_s3_0/EESPFAL_INV4_0/Dis GND -0.29fF $ **FLOATING
C2558 Dis2.n3 GND 0.32fF $ **FLOATING
C2559 Dis2.n4 GND 1.49fF $ **FLOATING
C2560 Dis2.t20 GND 0.24fF
C2561 Dis2.t3 GND 0.15fF
C2562 Dis2.n5 GND 0.61fF $ **FLOATING
C2563 EESPFAL_s3_0/EESPFAL_NAND_v3_1/Dis GND 0.25fF $ **FLOATING
C2564 Dis2.n6 GND 2.97fF $ **FLOATING
C2565 Dis2.t14 GND 0.24fF
C2566 Dis2.t2 GND 0.15fF
C2567 Dis2.n7 GND 0.61fF $ **FLOATING
C2568 EESPFAL_s3_0/EESPFAL_NAND_v3_0/Dis GND 0.25fF $ **FLOATING
C2569 Dis2.n8 GND 0.96fF $ **FLOATING
C2570 EESPFAL_s3_0/Dis2 GND 0.75fF $ **FLOATING
C2571 EESPFAL_s2_0/Dis2 GND 0.76fF $ **FLOATING
C2572 Dis2.t6 GND 0.24fF
C2573 Dis2.t0 GND 0.15fF
C2574 Dis2.n9 GND 0.61fF $ **FLOATING
C2575 EESPFAL_s2_0/EESPFAL_NAND_v3_1/Dis GND 0.24fF $ **FLOATING
C2576 Dis2.n10 GND 0.97fF $ **FLOATING
C2577 Dis2.t21 GND 0.24fF
C2578 Dis2.t9 GND 0.15fF
C2579 Dis2.n11 GND 0.61fF $ **FLOATING
C2580 EESPFAL_s2_0/EESPFAL_NAND_v3_0/Dis GND 0.25fF $ **FLOATING
C2581 Dis2.n12 GND 2.09fF $ **FLOATING
C2582 Dis2.n13 GND 1.96fF $ **FLOATING
C2583 Dis2.t11 GND 0.15fF
C2584 Dis2.t18 GND 0.15fF
C2585 EESPFAL_s1_0/EESPFAL_INV4_0/Dis GND -0.29fF $ **FLOATING
C2586 Dis2.n14 GND 0.32fF $ **FLOATING
C2587 Dis2.n15 GND 0.68fF $ **FLOATING
C2588 Dis2.n16 GND 1.90fF $ **FLOATING
C2589 Dis2.t19 GND 0.24fF
C2590 Dis2.t4 GND 0.15fF
C2591 Dis2.n17 GND 0.61fF $ **FLOATING
C2592 EESPFAL_s1_0/EESPFAL_NAND_v3_1/Dis GND 0.25fF $ **FLOATING
C2593 Dis2.n18 GND 2.11fF $ **FLOATING
C2594 Dis2.t7 GND 0.24fF
C2595 Dis2.t16 GND 0.15fF
C2596 Dis2.n19 GND 0.61fF $ **FLOATING
C2597 EESPFAL_s1_0/EESPFAL_NAND_v3_0/Dis GND 0.25fF $ **FLOATING
C2598 Dis2.n20 GND 0.96fF $ **FLOATING
C2599 EESPFAL_s1_0/Dis2 GND 1.40fF $ **FLOATING
C2600 Dis2.t10 GND 0.15fF
C2601 Dis2.t1 GND 0.15fF
C2602 EESPFAL_s0_0/EESPFAL_NAND_v3_1/Dis GND -0.40fF $ **FLOATING
C2603 Dis2.n21 GND 0.32fF $ **FLOATING
C2604 Dis2.n22 GND 0.50fF $ **FLOATING
C2605 Dis2.n23 GND 1.09fF $ **FLOATING
C2606 Dis2.n24 GND 0.87fF $ **FLOATING
C2607 EESPFAL_s0_0/Dis2 GND 0.04fF $ **FLOATING
C2608 EESPFAL_s3_0/EESPFAL_XOR_v3_1/OUT_bar GND 0.50fF $ **FLOATING
C2609 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t8 GND 0.07fF
C2610 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t5 GND 0.05fF
C2611 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t2 GND 0.05fF
C2612 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n0 GND 0.13fF $ **FLOATING
C2613 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t3 GND 0.05fF
C2614 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t4 GND 0.05fF
C2615 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n1 GND 0.15fF $ **FLOATING
C2616 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t1 GND 0.19fF
C2617 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t0 GND 0.33fF
C2618 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n2 GND 0.29fF $ **FLOATING
C2619 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n3 GND 0.12fF $ **FLOATING
C2620 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n4 GND 0.14fF $ **FLOATING
C2621 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t7 GND 0.05fF
C2622 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t6 GND 0.06fF
C2623 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.t9 GND 0.06fF
C2624 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n5 GND 0.07fF $ **FLOATING
C2625 EESPFAL_s3_0/EESPFAL_NAND_v3_1/A_bar.n6 GND 0.05fF $ **FLOATING
C2626 EESPFAL_s0_0/x3_bar GND 0.32fF $ **FLOATING
C2627 x3_bar.t4 GND 0.53fF
C2628 x3_bar.t9 GND 0.18fF
C2629 x3_bar.n0 GND 1.78fF $ **FLOATING
C2630 x3_bar.n1 GND 2.08fF $ **FLOATING
C2631 x3_bar.t3 GND 0.14fF
C2632 EESPFAL_s1_0/EESPFAL_INV4_2/A_bar GND 0.50fF $ **FLOATING
C2633 x3_bar.t10 GND 0.53fF
C2634 x3_bar.t5 GND 0.18fF
C2635 x3_bar.n2 GND 1.78fF $ **FLOATING
C2636 EESPFAL_s1_0/EESPFAL_XOR_v3_1/B_bar GND 0.11fF $ **FLOATING
C2637 x3_bar.t8 GND 0.46fF
C2638 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/A GND 2.00fF $ **FLOATING
C2639 x3_bar.t2 GND 0.34fF
C2640 EESPFAL_s2_0/EESPFAL_4in_NAND_0/A GND 2.64fF $ **FLOATING
C2641 x3_bar.t11 GND 0.41fF
C2642 x3_bar.t12 GND 0.23fF
C2643 x3_bar.n3 GND 2.20fF $ **FLOATING
C2644 EESPFAL_s2_0/EESPFAL_XOR_v3_0/A_bar GND 0.18fF $ **FLOATING
C2645 x3_bar.t1 GND 0.20fF
C2646 EESPFAL_s3_0/EESPFAL_INV4_2/A GND 0.98fF $ **FLOATING
C2647 x3_bar.t6 GND 0.53fF
C2648 x3_bar.t0 GND 0.18fF
C2649 x3_bar.n4 GND 1.78fF $ **FLOATING
C2650 EESPFAL_s3_0/EESPFAL_XOR_v3_1/B_bar GND 0.11fF $ **FLOATING
C2651 x3_bar.t7 GND 0.16fF
C2652 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/C_bar GND 0.43fF $ **FLOATING
C2653 x3_bar.n5 GND 4.37fF $ **FLOATING
C2654 EESPFAL_s3_0/x3_bar GND 1.24fF $ **FLOATING
C2655 x3_bar.n6 GND 4.89fF $ **FLOATING
C2656 EESPFAL_s2_0/x3_bar GND 0.56fF $ **FLOATING
C2657 x3_bar.n7 GND 1.82fF $ **FLOATING
C2658 x3_bar.n8 GND 3.54fF $ **FLOATING
C2659 x3_bar.n9 GND 2.64fF $ **FLOATING
C2660 x3_bar.n10 GND 1.58fF $ **FLOATING
C2661 x3_bar.n11 GND 4.52fF $ **FLOATING
C2662 EESPFAL_s1_0/x3_bar GND 2.20fF $ **FLOATING
C2663 EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT_bar GND 0.30fF $ **FLOATING
C2664 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t9 GND 0.12fF
C2665 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t3 GND 0.04fF
C2666 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t1 GND 0.04fF
C2667 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n0 GND 0.13fF $ **FLOATING
C2668 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t0 GND 0.17fF
C2669 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t2 GND 0.29fF
C2670 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n1 GND 0.26fF $ **FLOATING
C2671 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n2 GND 0.11fF $ **FLOATING
C2672 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t5 GND 0.04fF
C2673 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t4 GND 0.04fF
C2674 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n3 GND 0.11fF $ **FLOATING
C2675 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n4 GND 0.12fF $ **FLOATING
C2676 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t8 GND 0.06fF
C2677 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t6 GND 0.05fF
C2678 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.t7 GND 0.04fF
C2679 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n5 GND 0.06fF $ **FLOATING
C2680 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A.n6 GND 0.04fF $ **FLOATING
C2681 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t9 GND 0.08fF
C2682 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t2 GND 0.24fF
C2683 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t3 GND 0.24fF
C2684 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t5 GND 0.05fF
C2685 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t0 GND 0.05fF
C2686 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n0 GND 0.17fF $ **FLOATING
C2687 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t8 GND 0.07fF
C2688 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t6 GND 0.08fF
C2689 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t7 GND 0.04fF
C2690 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n1 GND 0.08fF $ **FLOATING
C2691 EESPFAL_s1_0/EESPFAL_XOR_v3_0/OUT GND 0.01fF $ **FLOATING
C2692 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n2 GND 0.04fF $ **FLOATING
C2693 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t4 GND 0.05fF
C2694 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.t1 GND 0.05fF
C2695 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n3 GND 0.18fF $ **FLOATING
C2696 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n4 GND 0.24fF $ **FLOATING
C2697 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n5 GND 0.24fF $ **FLOATING
C2698 EESPFAL_s1_0/EESPFAL_NAND_v3_0/A_bar.n6 GND 0.52fF $ **FLOATING
C2699 CLK1.t40 GND 0.03fF
C2700 CLK1.t100 GND 0.03fF
C2701 CLK1.n0 GND 0.15fF $ **FLOATING
C2702 CLK1.t5 GND 0.05fF
C2703 EESPFAL_s0_0/EESPFAL_XOR_v3_0/CLK GND 0.02fF $ **FLOATING
C2704 CLK1.n1 GND 0.17fF $ **FLOATING
C2705 CLK1.n2 GND 0.03fF $ **FLOATING
C2706 CLK1.t89 GND 0.03fF
C2707 CLK1.t26 GND 0.03fF
C2708 CLK1.n3 GND 0.10fF $ **FLOATING
C2709 CLK1.t64 GND 0.05fF
C2710 CLK1.t197 GND 0.03fF
C2711 CLK1.t71 GND 0.03fF
C2712 CLK1.n4 GND 0.15fF $ **FLOATING
C2713 CLK1.t117 GND 0.08fF
C2714 CLK1.t111 GND 0.05fF
C2715 CLK1.n5 GND 0.17fF $ **FLOATING
C2716 CLK1.n6 GND 0.03fF $ **FLOATING
C2717 CLK1.t191 GND 0.03fF
C2718 CLK1.t109 GND 0.03fF
C2719 CLK1.n7 GND 0.10fF $ **FLOATING
C2720 CLK1.t189 GND 0.05fF
C2721 CLK1.t57 GND 0.03fF
C2722 CLK1.t33 GND 0.03fF
C2723 CLK1.n8 GND 0.15fF $ **FLOATING
C2724 CLK1.n9 GND 0.08fF $ **FLOATING
C2725 CLK1.n10 GND 0.03fF $ **FLOATING
C2726 CLK1.n11 GND 0.02fF $ **FLOATING
C2727 CLK1.n12 GND 0.13fF $ **FLOATING
C2728 CLK1.n13 GND 0.06fF $ **FLOATING
C2729 CLK1.n14 GND 0.03fF $ **FLOATING
C2730 CLK1.n15 GND 0.02fF $ **FLOATING
C2731 CLK1.n16 GND 0.07fF $ **FLOATING
C2732 CLK1.n17 GND 0.19fF $ **FLOATING
C2733 CLK1.n18 GND 0.06fF $ **FLOATING
C2734 CLK1.n19 GND 0.03fF $ **FLOATING
C2735 CLK1.n20 GND 0.02fF $ **FLOATING
C2736 CLK1.n21 GND 0.03fF $ **FLOATING
C2737 CLK1.n22 GND 0.06fF $ **FLOATING
C2738 CLK1.n23 GND 0.03fF $ **FLOATING
C2739 CLK1.n24 GND 0.02fF $ **FLOATING
C2740 CLK1.n25 GND 0.03fF $ **FLOATING
C2741 CLK1.n26 GND 0.14fF $ **FLOATING
C2742 CLK1.n27 GND 0.03fF $ **FLOATING
C2743 CLK1.n28 GND 0.02fF $ **FLOATING
C2744 CLK1.n29 GND 0.03fF $ **FLOATING
C2745 CLK1.n30 GND 0.18fF $ **FLOATING
C2746 CLK1.n31 GND 0.03fF $ **FLOATING
C2747 CLK1.n32 GND 0.02fF $ **FLOATING
C2748 CLK1.n33 GND 0.02fF $ **FLOATING
C2749 CLK1.n34 GND 0.29fF $ **FLOATING
C2750 CLK1.t188 GND 0.09fF
C2751 CLK1.n35 GND 0.11fF $ **FLOATING
C2752 CLK1.n36 GND 0.03fF $ **FLOATING
C2753 CLK1.n37 GND 0.02fF $ **FLOATING
C2754 CLK1.n38 GND 0.03fF $ **FLOATING
C2755 CLK1.n39 GND 0.16fF $ **FLOATING
C2756 CLK1.n40 GND 0.03fF $ **FLOATING
C2757 CLK1.n41 GND 0.02fF $ **FLOATING
C2758 CLK1.n42 GND 0.03fF $ **FLOATING
C2759 CLK1.t190 GND 0.09fF
C2760 CLK1.n43 GND 0.09fF $ **FLOATING
C2761 CLK1.n44 GND 0.03fF $ **FLOATING
C2762 CLK1.n45 GND 0.02fF $ **FLOATING
C2763 CLK1.n46 GND 0.03fF $ **FLOATING
C2764 CLK1.n47 GND 0.17fF $ **FLOATING
C2765 CLK1.n48 GND 0.02fF $ **FLOATING
C2766 CLK1.t108 GND 0.09fF
C2767 CLK1.n49 GND 0.09fF $ **FLOATING
C2768 CLK1.n50 GND 0.03fF $ **FLOATING
C2769 CLK1.n51 GND 0.02fF $ **FLOATING
C2770 CLK1.n52 GND 0.03fF $ **FLOATING
C2771 CLK1.n53 GND 0.16fF $ **FLOATING
C2772 CLK1.n54 GND 0.03fF $ **FLOATING
C2773 CLK1.n55 GND 0.02fF $ **FLOATING
C2774 CLK1.n56 GND 0.03fF $ **FLOATING
C2775 CLK1.t110 GND 0.09fF
C2776 CLK1.n57 GND 0.11fF $ **FLOATING
C2777 CLK1.n58 GND 0.03fF $ **FLOATING
C2778 CLK1.n59 GND 0.02fF $ **FLOATING
C2779 CLK1.n60 GND 0.03fF $ **FLOATING
C2780 CLK1.n61 GND 0.29fF $ **FLOATING
C2781 CLK1.n62 GND 0.18fF $ **FLOATING
C2782 CLK1.n63 GND 0.03fF $ **FLOATING
C2783 CLK1.n64 GND 0.02fF $ **FLOATING
C2784 CLK1.n65 GND 0.02fF $ **FLOATING
C2785 CLK1.n66 GND 0.14fF $ **FLOATING
C2786 CLK1.n67 GND 0.03fF $ **FLOATING
C2787 CLK1.n68 GND 0.02fF $ **FLOATING
C2788 CLK1.n69 GND 0.03fF $ **FLOATING
C2789 CLK1.n70 GND 0.06fF $ **FLOATING
C2790 CLK1.n71 GND 0.03fF $ **FLOATING
C2791 CLK1.n72 GND 0.02fF $ **FLOATING
C2792 CLK1.n73 GND 0.03fF $ **FLOATING
C2793 CLK1.n74 GND 0.06fF $ **FLOATING
C2794 CLK1.n75 GND 0.03fF $ **FLOATING
C2795 CLK1.n76 GND 0.02fF $ **FLOATING
C2796 CLK1.n77 GND 0.03fF $ **FLOATING
C2797 CLK1.n78 GND 0.06fF $ **FLOATING
C2798 CLK1.n79 GND 0.03fF $ **FLOATING
C2799 CLK1.n80 GND 0.02fF $ **FLOATING
C2800 CLK1.n81 GND 0.03fF $ **FLOATING
C2801 CLK1.n82 GND 0.07fF $ **FLOATING
C2802 CLK1.n83 GND 0.03fF $ **FLOATING
C2803 CLK1.n84 GND 0.02fF $ **FLOATING
C2804 CLK1.n85 GND 0.03fF $ **FLOATING
C2805 CLK1.n86 GND 0.34fF $ **FLOATING
C2806 CLK1.n87 GND 0.13fF $ **FLOATING
C2807 CLK1.n88 GND 0.10fF $ **FLOATING
C2808 CLK1.n89 GND 0.21fF $ **FLOATING
C2809 CLK1.n90 GND 0.11fF $ **FLOATING
C2810 CLK1.n91 GND 0.08fF $ **FLOATING
C2811 CLK1.n92 GND 0.03fF $ **FLOATING
C2812 CLK1.n93 GND 0.02fF $ **FLOATING
C2813 CLK1.n94 GND 0.03fF $ **FLOATING
C2814 CLK1.n95 GND 0.06fF $ **FLOATING
C2815 CLK1.n96 GND 0.03fF $ **FLOATING
C2816 CLK1.n97 GND 0.02fF $ **FLOATING
C2817 CLK1.n98 GND 0.03fF $ **FLOATING
C2818 CLK1.n99 GND 0.06fF $ **FLOATING
C2819 CLK1.n100 GND 0.03fF $ **FLOATING
C2820 CLK1.n101 GND 0.02fF $ **FLOATING
C2821 CLK1.n102 GND 0.02fF $ **FLOATING
C2822 CLK1.n103 GND 0.19fF $ **FLOATING
C2823 CLK1.n104 GND 0.06fF $ **FLOATING
C2824 CLK1.n105 GND 0.03fF $ **FLOATING
C2825 CLK1.n106 GND 0.02fF $ **FLOATING
C2826 CLK1.n107 GND 0.03fF $ **FLOATING
C2827 CLK1.n108 GND 0.06fF $ **FLOATING
C2828 CLK1.n109 GND 0.03fF $ **FLOATING
C2829 CLK1.n110 GND 0.02fF $ **FLOATING
C2830 CLK1.n111 GND 0.03fF $ **FLOATING
C2831 CLK1.n112 GND 0.06fF $ **FLOATING
C2832 CLK1.n113 GND 0.03fF $ **FLOATING
C2833 CLK1.n114 GND 0.02fF $ **FLOATING
C2834 CLK1.n115 GND 0.03fF $ **FLOATING
C2835 CLK1.n116 GND 0.06fF $ **FLOATING
C2836 CLK1.n117 GND 0.03fF $ **FLOATING
C2837 CLK1.n118 GND 0.02fF $ **FLOATING
C2838 CLK1.n119 GND 0.03fF $ **FLOATING
C2839 CLK1.n120 GND 0.14fF $ **FLOATING
C2840 CLK1.n121 GND 0.03fF $ **FLOATING
C2841 CLK1.n122 GND 0.02fF $ **FLOATING
C2842 CLK1.n123 GND 0.03fF $ **FLOATING
C2843 CLK1.n124 GND 0.18fF $ **FLOATING
C2844 CLK1.n125 GND 0.03fF $ **FLOATING
C2845 CLK1.n126 GND 0.02fF $ **FLOATING
C2846 CLK1.n127 GND 0.02fF $ **FLOATING
C2847 CLK1.n128 GND 0.29fF $ **FLOATING
C2848 CLK1.t63 GND 0.09fF
C2849 CLK1.n129 GND 0.11fF $ **FLOATING
C2850 CLK1.n130 GND 0.03fF $ **FLOATING
C2851 CLK1.n131 GND 0.02fF $ **FLOATING
C2852 CLK1.n132 GND 0.03fF $ **FLOATING
C2853 CLK1.n133 GND 0.16fF $ **FLOATING
C2854 CLK1.n134 GND 0.03fF $ **FLOATING
C2855 CLK1.n135 GND 0.02fF $ **FLOATING
C2856 CLK1.n136 GND 0.03fF $ **FLOATING
C2857 CLK1.t88 GND 0.09fF
C2858 CLK1.n137 GND 0.09fF $ **FLOATING
C2859 CLK1.n138 GND 0.03fF $ **FLOATING
C2860 CLK1.n139 GND 0.02fF $ **FLOATING
C2861 CLK1.n140 GND 0.03fF $ **FLOATING
C2862 CLK1.n141 GND 0.17fF $ **FLOATING
C2863 CLK1.n142 GND 0.02fF $ **FLOATING
C2864 CLK1.t25 GND 0.09fF
C2865 CLK1.n143 GND 0.09fF $ **FLOATING
C2866 CLK1.n144 GND 0.03fF $ **FLOATING
C2867 CLK1.n145 GND 0.02fF $ **FLOATING
C2868 CLK1.n146 GND 0.03fF $ **FLOATING
C2869 CLK1.n147 GND 0.16fF $ **FLOATING
C2870 CLK1.n148 GND 0.03fF $ **FLOATING
C2871 CLK1.n149 GND 0.02fF $ **FLOATING
C2872 CLK1.n150 GND 0.03fF $ **FLOATING
C2873 CLK1.t4 GND 0.09fF
C2874 CLK1.n151 GND 0.11fF $ **FLOATING
C2875 CLK1.n152 GND 0.03fF $ **FLOATING
C2876 CLK1.n153 GND 0.02fF $ **FLOATING
C2877 CLK1.n154 GND 0.03fF $ **FLOATING
C2878 CLK1.n155 GND 0.29fF $ **FLOATING
C2879 CLK1.n156 GND 0.18fF $ **FLOATING
C2880 CLK1.n157 GND 0.03fF $ **FLOATING
C2881 CLK1.n158 GND 0.02fF $ **FLOATING
C2882 CLK1.n159 GND 0.02fF $ **FLOATING
C2883 CLK1.n160 GND 0.14fF $ **FLOATING
C2884 CLK1.n161 GND 0.03fF $ **FLOATING
C2885 CLK1.n162 GND 0.02fF $ **FLOATING
C2886 CLK1.n163 GND 0.03fF $ **FLOATING
C2887 CLK1.n164 GND 0.06fF $ **FLOATING
C2888 CLK1.n165 GND 0.03fF $ **FLOATING
C2889 CLK1.n166 GND 0.02fF $ **FLOATING
C2890 CLK1.n167 GND 0.03fF $ **FLOATING
C2891 CLK1.n168 GND 0.06fF $ **FLOATING
C2892 CLK1.n169 GND 0.03fF $ **FLOATING
C2893 CLK1.n170 GND 0.02fF $ **FLOATING
C2894 CLK1.n171 GND 0.03fF $ **FLOATING
C2895 CLK1.n172 GND 0.06fF $ **FLOATING
C2896 CLK1.n173 GND 0.03fF $ **FLOATING
C2897 CLK1.n174 GND 0.02fF $ **FLOATING
C2898 CLK1.n175 GND 0.03fF $ **FLOATING
C2899 CLK1.n176 GND 0.06fF $ **FLOATING
C2900 CLK1.n177 GND 0.03fF $ **FLOATING
C2901 CLK1.n178 GND 0.02fF $ **FLOATING
C2902 CLK1.n179 GND 0.03fF $ **FLOATING
C2903 CLK1.n180 GND 0.19fF $ **FLOATING
C2904 CLK1.n181 GND 0.06fF $ **FLOATING
C2905 CLK1.n182 GND 0.03fF $ **FLOATING
C2906 CLK1.n183 GND 0.02fF $ **FLOATING
C2907 CLK1.n184 GND 0.02fF $ **FLOATING
C2908 CLK1.n185 GND 0.06fF $ **FLOATING
C2909 CLK1.n186 GND 0.03fF $ **FLOATING
C2910 CLK1.n187 GND 0.02fF $ **FLOATING
C2911 CLK1.n188 GND 0.03fF $ **FLOATING
C2912 CLK1.n189 GND 0.08fF $ **FLOATING
C2913 CLK1.n190 GND 0.03fF $ **FLOATING
C2914 CLK1.n191 GND 0.02fF $ **FLOATING
C2915 CLK1.n192 GND 0.03fF $ **FLOATING
C2916 CLK1.n193 GND 0.21fF $ **FLOATING
C2917 CLK1.n194 GND 0.05fF $ **FLOATING
C2918 CLK1.n195 GND 0.03fF $ **FLOATING
C2919 CLK1.n196 GND 0.02fF $ **FLOATING
C2920 CLK1.n197 GND 0.03fF $ **FLOATING
C2921 CLK1.n198 GND 0.06fF $ **FLOATING
C2922 CLK1.n199 GND 0.03fF $ **FLOATING
C2923 CLK1.n200 GND 0.02fF $ **FLOATING
C2924 CLK1.t49 GND 0.03fF
C2925 CLK1.t60 GND 0.03fF
C2926 CLK1.n201 GND 0.15fF $ **FLOATING
C2927 CLK1.n202 GND 0.03fF $ **FLOATING
C2928 CLK1.n203 GND 0.02fF $ **FLOATING
C2929 CLK1.n204 GND 0.03fF $ **FLOATING
C2930 CLK1.n205 GND 0.11fF $ **FLOATING
C2931 CLK1.n206 GND 0.03fF $ **FLOATING
C2932 CLK1.n207 GND 0.02fF $ **FLOATING
C2933 CLK1.t19 GND 0.05fF
C2934 CLK1.n208 GND 0.03fF $ **FLOATING
C2935 CLK1.n209 GND 0.02fF $ **FLOATING
C2936 CLK1.n210 GND 0.03fF $ **FLOATING
C2937 CLK1.t166 GND 0.09fF
C2938 CLK1.n211 GND 0.03fF $ **FLOATING
C2939 CLK1.n212 GND 0.02fF $ **FLOATING
C2940 CLK1.t167 GND 0.03fF
C2941 CLK1.t17 GND 0.03fF
C2942 CLK1.n213 GND 0.10fF $ **FLOATING
C2943 CLK1.n214 GND 0.03fF $ **FLOATING
C2944 CLK1.n215 GND 0.02fF $ **FLOATING
C2945 CLK1.n216 GND 0.03fF $ **FLOATING
C2946 CLK1.n217 GND 0.14fF $ **FLOATING
C2947 CLK1.n218 GND 0.03fF $ **FLOATING
C2948 CLK1.n219 GND 0.02fF $ **FLOATING
C2949 CLK1.n220 GND 0.03fF $ **FLOATING
C2950 CLK1.n221 GND 0.02fF $ **FLOATING
C2951 CLK1.n222 GND 0.03fF $ **FLOATING
C2952 CLK1.n223 GND 0.07fF $ **FLOATING
C2953 CLK1.n224 GND 0.03fF $ **FLOATING
C2954 CLK1.n225 GND 0.02fF $ **FLOATING
C2955 CLK1.t95 GND 0.08fF
C2956 CLK1.n226 GND 0.13fF $ **FLOATING
C2957 CLK1.n227 GND 0.35fF $ **FLOATING
C2958 CLK1.n228 GND 0.03fF $ **FLOATING
C2959 CLK1.n229 GND 0.03fF $ **FLOATING
C2960 CLK1.n230 GND 0.02fF $ **FLOATING
C2961 CLK1.n231 GND 0.03fF $ **FLOATING
C2962 CLK1.n232 GND 0.06fF $ **FLOATING
C2963 CLK1.n233 GND 0.06fF $ **FLOATING
C2964 CLK1.n234 GND 0.06fF $ **FLOATING
C2965 CLK1.n235 GND 0.03fF $ **FLOATING
C2966 CLK1.n236 GND 0.02fF $ **FLOATING
C2967 CLK1.n237 GND 0.03fF $ **FLOATING
C2968 CLK1.n238 GND 0.03fF $ **FLOATING
C2969 CLK1.t165 GND 0.05fF
C2970 CLK1.n239 GND 0.29fF $ **FLOATING
C2971 CLK1.n240 GND 0.02fF $ **FLOATING
C2972 CLK1.n241 GND 0.02fF $ **FLOATING
C2973 CLK1.n242 GND 0.03fF $ **FLOATING
C2974 CLK1.n243 GND 0.18fF $ **FLOATING
C2975 CLK1.n244 GND 0.11fF $ **FLOATING
C2976 CLK1.t164 GND 0.09fF
C2977 CLK1.n245 GND 0.09fF $ **FLOATING
C2978 CLK1.n246 GND 0.16fF $ **FLOATING
C2979 CLK1.n247 GND 0.03fF $ **FLOATING
C2980 CLK1.n248 GND 0.02fF $ **FLOATING
C2981 CLK1.n249 GND 0.03fF $ **FLOATING
C2982 CLK1.n250 GND 0.03fF $ **FLOATING
C2983 EESPFAL_s0_0/EESPFAL_NAND_v3_2/CLK GND 0.02fF $ **FLOATING
C2984 CLK1.n251 GND 0.17fF $ **FLOATING
C2985 CLK1.n252 GND 0.02fF $ **FLOATING
C2986 CLK1.n253 GND 0.03fF $ **FLOATING
C2987 CLK1.n254 GND 0.17fF $ **FLOATING
C2988 CLK1.t16 GND 0.09fF
C2989 CLK1.n255 GND 0.09fF $ **FLOATING
C2990 CLK1.t18 GND 0.09fF
C2991 CLK1.n256 GND 0.16fF $ **FLOATING
C2992 CLK1.n257 GND 0.03fF $ **FLOATING
C2993 CLK1.n258 GND 0.02fF $ **FLOATING
C2994 CLK1.n259 GND 0.03fF $ **FLOATING
C2995 CLK1.n260 GND 0.03fF $ **FLOATING
C2996 CLK1.n261 GND 0.29fF $ **FLOATING
C2997 CLK1.n262 GND 0.02fF $ **FLOATING
C2998 CLK1.n263 GND 0.02fF $ **FLOATING
C2999 CLK1.n264 GND 0.03fF $ **FLOATING
C3000 CLK1.n265 GND 0.18fF $ **FLOATING
C3001 CLK1.n266 GND 0.14fF $ **FLOATING
C3002 CLK1.n267 GND 0.06fF $ **FLOATING
C3003 CLK1.n268 GND 0.03fF $ **FLOATING
C3004 CLK1.n269 GND 0.02fF $ **FLOATING
C3005 CLK1.n270 GND 0.03fF $ **FLOATING
C3006 CLK1.n271 GND 0.03fF $ **FLOATING
C3007 CLK1.n272 GND 0.19fF $ **FLOATING
C3008 CLK1.n273 GND 0.02fF $ **FLOATING
C3009 CLK1.n274 GND 0.02fF $ **FLOATING
C3010 CLK1.n275 GND 0.03fF $ **FLOATING
C3011 CLK1.n276 GND 0.06fF $ **FLOATING
C3012 CLK1.n277 GND 0.07fF $ **FLOATING
C3013 CLK1.n278 GND 0.13fF $ **FLOATING
C3014 CLK1.n279 GND 0.14fF $ **FLOATING
C3015 CLK1.n280 GND 0.00fF $ **FLOATING
C3016 EESPFAL_s1_0/CLK1 GND 0.00fF $ **FLOATING
C3017 CLK1.n281 GND 0.01fF $ **FLOATING
C3018 CLK1.t24 GND 0.08fF
C3019 CLK1.n282 GND 0.34fF $ **FLOATING
C3020 CLK1.n283 GND 0.02fF $ **FLOATING
C3021 CLK1.n284 GND 0.03fF $ **FLOATING
C3022 CLK1.n285 GND 0.06fF $ **FLOATING
C3023 CLK1.n286 GND 0.03fF $ **FLOATING
C3024 CLK1.n287 GND 0.02fF $ **FLOATING
C3025 CLK1.t163 GND 0.03fF
C3026 CLK1.t187 GND 0.03fF
C3027 CLK1.n288 GND 0.15fF $ **FLOATING
C3028 CLK1.n289 GND 0.19fF $ **FLOATING
C3029 CLK1.n290 GND 0.02fF $ **FLOATING
C3030 CLK1.n291 GND 0.03fF $ **FLOATING
C3031 CLK1.n292 GND 0.14fF $ **FLOATING
C3032 CLK1.n293 GND 0.03fF $ **FLOATING
C3033 CLK1.n294 GND 0.02fF $ **FLOATING
C3034 CLK1.t138 GND 0.05fF
C3035 CLK1.n295 GND 0.29fF $ **FLOATING
C3036 CLK1.n296 GND 0.02fF $ **FLOATING
C3037 CLK1.n297 GND 0.03fF $ **FLOATING
C3038 CLK1.n298 GND 0.09fF $ **FLOATING
C3039 CLK1.n299 GND 0.03fF $ **FLOATING
C3040 CLK1.n300 GND 0.02fF $ **FLOATING
C3041 CLK1.t35 GND 0.03fF
C3042 CLK1.t136 GND 0.03fF
C3043 CLK1.n301 GND 0.10fF $ **FLOATING
C3044 CLK1.n302 GND 0.03fF $ **FLOATING
C3045 CLK1.n303 GND 0.02fF $ **FLOATING
C3046 CLK1.n304 GND 0.03fF $ **FLOATING
C3047 CLK1.t36 GND 0.09fF
C3048 CLK1.n305 GND 0.03fF $ **FLOATING
C3049 CLK1.n306 GND 0.02fF $ **FLOATING
C3050 CLK1.t37 GND 0.05fF
C3051 CLK1.n307 GND 0.03fF $ **FLOATING
C3052 CLK1.n308 GND 0.02fF $ **FLOATING
C3053 CLK1.n309 GND 0.03fF $ **FLOATING
C3054 CLK1.n310 GND 0.06fF $ **FLOATING
C3055 CLK1.n311 GND 0.03fF $ **FLOATING
C3056 CLK1.n312 GND 0.02fF $ **FLOATING
C3057 CLK1.n313 GND 0.03fF $ **FLOATING
C3058 CLK1.n314 GND 0.02fF $ **FLOATING
C3059 CLK1.n315 GND 0.03fF $ **FLOATING
C3060 CLK1.n316 GND 0.07fF $ **FLOATING
C3061 CLK1.n317 GND 0.03fF $ **FLOATING
C3062 CLK1.n318 GND 0.02fF $ **FLOATING
C3063 CLK1.n319 GND 0.02fF $ **FLOATING
C3064 CLK1.n320 GND 0.02fF $ **FLOATING
C3065 CLK1.n321 GND 0.02fF $ **FLOATING
C3066 CLK1.t170 GND 0.03fF
C3067 CLK1.t22 GND 0.07fF
C3068 CLK1.n322 GND 0.45fF $ **FLOATING
C3069 CLK1.n323 GND 0.02fF $ **FLOATING
C3070 CLK1.n324 GND 0.03fF $ **FLOATING
C3071 CLK1.n325 GND 0.14fF $ **FLOATING
C3072 CLK1.n326 GND 0.03fF $ **FLOATING
C3073 CLK1.n327 GND 0.02fF $ **FLOATING
C3074 CLK1.t105 GND 0.05fF
C3075 CLK1.n328 GND 0.29fF $ **FLOATING
C3076 CLK1.n329 GND 0.02fF $ **FLOATING
C3077 CLK1.n330 GND 0.03fF $ **FLOATING
C3078 CLK1.n331 GND 0.09fF $ **FLOATING
C3079 CLK1.n332 GND 0.03fF $ **FLOATING
C3080 CLK1.n333 GND 0.02fF $ **FLOATING
C3081 CLK1.t146 GND 0.03fF
C3082 CLK1.t103 GND 0.03fF
C3083 CLK1.n334 GND 0.10fF $ **FLOATING
C3084 CLK1.n335 GND 0.03fF $ **FLOATING
C3085 CLK1.n336 GND 0.02fF $ **FLOATING
C3086 CLK1.n337 GND 0.03fF $ **FLOATING
C3087 CLK1.t143 GND 0.09fF
C3088 CLK1.n338 GND 0.03fF $ **FLOATING
C3089 CLK1.n339 GND 0.02fF $ **FLOATING
C3090 CLK1.t144 GND 0.05fF
C3091 CLK1.n340 GND 0.03fF $ **FLOATING
C3092 CLK1.n341 GND 0.02fF $ **FLOATING
C3093 CLK1.n342 GND 0.03fF $ **FLOATING
C3094 CLK1.n343 GND 0.07fF $ **FLOATING
C3095 CLK1.n344 GND 0.03fF $ **FLOATING
C3096 CLK1.n345 GND 0.02fF $ **FLOATING
C3097 CLK1.t27 GND 0.07fF
C3098 CLK1.n346 GND 0.15fF $ **FLOATING
C3099 CLK1.n347 GND 0.47fF $ **FLOATING
C3100 CLK1.n348 GND 0.03fF $ **FLOATING
C3101 CLK1.n349 GND 0.03fF $ **FLOATING
C3102 CLK1.n350 GND 0.02fF $ **FLOATING
C3103 CLK1.n351 GND 0.03fF $ **FLOATING
C3104 CLK1.n352 GND 0.06fF $ **FLOATING
C3105 CLK1.n353 GND 0.14fF $ **FLOATING
C3106 CLK1.n354 GND 0.11fF $ **FLOATING
C3107 CLK1.n355 GND 0.18fF $ **FLOATING
C3108 CLK1.n356 GND 0.03fF $ **FLOATING
C3109 CLK1.n357 GND 0.02fF $ **FLOATING
C3110 CLK1.n358 GND 0.02fF $ **FLOATING
C3111 CLK1.n359 GND 0.29fF $ **FLOATING
C3112 CLK1.n360 GND 0.03fF $ **FLOATING
C3113 CLK1.n361 GND 0.03fF $ **FLOATING
C3114 CLK1.n362 GND 0.02fF $ **FLOATING
C3115 CLK1.n363 GND 0.03fF $ **FLOATING
C3116 CLK1.n364 GND 0.16fF $ **FLOATING
C3117 CLK1.n365 GND 0.09fF $ **FLOATING
C3118 CLK1.t145 GND 0.09fF
C3119 CLK1.t102 GND 0.09fF
C3120 CLK1.n366 GND 0.17fF $ **FLOATING
C3121 CLK1.n367 GND 0.03fF $ **FLOATING
C3122 CLK1.n368 GND 0.02fF $ **FLOATING
C3123 CLK1.n369 GND 0.17fF $ **FLOATING
C3124 EESPFAL_s2_0/EESPFAL_INV4_0/CLK GND 0.02fF $ **FLOATING
C3125 CLK1.n370 GND 0.03fF $ **FLOATING
C3126 CLK1.n371 GND 0.03fF $ **FLOATING
C3127 CLK1.n372 GND 0.03fF $ **FLOATING
C3128 CLK1.n373 GND 0.02fF $ **FLOATING
C3129 CLK1.n374 GND 0.03fF $ **FLOATING
C3130 CLK1.n375 GND 0.16fF $ **FLOATING
C3131 CLK1.t104 GND 0.09fF
C3132 CLK1.n376 GND 0.11fF $ **FLOATING
C3133 CLK1.n377 GND 0.18fF $ **FLOATING
C3134 CLK1.n378 GND 0.03fF $ **FLOATING
C3135 CLK1.n379 GND 0.02fF $ **FLOATING
C3136 CLK1.n380 GND 0.02fF $ **FLOATING
C3137 CLK1.n381 GND 0.03fF $ **FLOATING
C3138 CLK1.n382 GND 0.03fF $ **FLOATING
C3139 CLK1.n383 GND 0.03fF $ **FLOATING
C3140 CLK1.n384 GND 0.02fF $ **FLOATING
C3141 CLK1.n385 GND 0.03fF $ **FLOATING
C3142 CLK1.n386 GND 0.06fF $ **FLOATING
C3143 CLK1.n387 GND 0.07fF $ **FLOATING
C3144 CLK1.n388 GND 0.15fF $ **FLOATING
C3145 CLK1.n389 GND 0.08fF $ **FLOATING
C3146 CLK1.n390 GND 0.13fF $ **FLOATING
C3147 CLK1.n391 GND 0.07fF $ **FLOATING
C3148 CLK1.n392 GND 0.26fF $ **FLOATING
C3149 CLK1.n393 GND 0.07fF $ **FLOATING
C3150 CLK1.n394 GND 0.07fF $ **FLOATING
C3151 CLK1.n395 GND 0.10fF $ **FLOATING
C3152 CLK1.n396 GND 0.07fF $ **FLOATING
C3153 CLK1.n397 GND 0.07fF $ **FLOATING
C3154 CLK1.n398 GND 0.03fF $ **FLOATING
C3155 CLK1.n399 GND 0.02fF $ **FLOATING
C3156 CLK1.n400 GND 0.02fF $ **FLOATING
C3157 CLK1.t94 GND 0.03fF
C3158 CLK1.n401 GND 0.02fF $ **FLOATING
C3159 CLK1.n402 GND 0.03fF $ **FLOATING
C3160 CLK1.n403 GND 0.02fF $ **FLOATING
C3161 CLK1.n404 GND 0.02fF $ **FLOATING
C3162 CLK1.n405 GND 0.03fF $ **FLOATING
C3163 CLK1.n406 GND 0.03fF $ **FLOATING
C3164 CLK1.n407 GND 0.08fF $ **FLOATING
C3165 CLK1.n408 GND 0.03fF $ **FLOATING
C3166 CLK1.n409 GND 0.02fF $ **FLOATING
C3167 CLK1.t58 GND 0.07fF
C3168 CLK1.n410 GND 0.45fF $ **FLOATING
C3169 CLK1.n411 GND 0.02fF $ **FLOATING
C3170 CLK1.n412 GND 0.03fF $ **FLOATING
C3171 CLK1.n413 GND 0.14fF $ **FLOATING
C3172 CLK1.n414 GND 0.03fF $ **FLOATING
C3173 CLK1.n415 GND 0.02fF $ **FLOATING
C3174 CLK1.t11 GND 0.05fF
C3175 CLK1.n416 GND 0.29fF $ **FLOATING
C3176 CLK1.n417 GND 0.02fF $ **FLOATING
C3177 CLK1.n418 GND 0.03fF $ **FLOATING
C3178 CLK1.n419 GND 0.09fF $ **FLOATING
C3179 CLK1.n420 GND 0.03fF $ **FLOATING
C3180 CLK1.n421 GND 0.02fF $ **FLOATING
C3181 CLK1.t122 GND 0.03fF
C3182 CLK1.t9 GND 0.03fF
C3183 CLK1.n422 GND 0.10fF $ **FLOATING
C3184 CLK1.n423 GND 0.03fF $ **FLOATING
C3185 CLK1.n424 GND 0.02fF $ **FLOATING
C3186 CLK1.n425 GND 0.03fF $ **FLOATING
C3187 CLK1.t119 GND 0.09fF
C3188 CLK1.n426 GND 0.03fF $ **FLOATING
C3189 CLK1.n427 GND 0.02fF $ **FLOATING
C3190 CLK1.t120 GND 0.05fF
C3191 CLK1.n428 GND 0.03fF $ **FLOATING
C3192 CLK1.n429 GND 0.02fF $ **FLOATING
C3193 CLK1.n430 GND 0.03fF $ **FLOATING
C3194 CLK1.n431 GND 0.07fF $ **FLOATING
C3195 CLK1.n432 GND 0.03fF $ **FLOATING
C3196 CLK1.n433 GND 0.02fF $ **FLOATING
C3197 CLK1.t118 GND 0.07fF
C3198 CLK1.n434 GND 0.15fF $ **FLOATING
C3199 CLK1.n435 GND 0.47fF $ **FLOATING
C3200 CLK1.n436 GND 0.03fF $ **FLOATING
C3201 CLK1.n437 GND 0.03fF $ **FLOATING
C3202 CLK1.n438 GND 0.02fF $ **FLOATING
C3203 CLK1.n439 GND 0.03fF $ **FLOATING
C3204 CLK1.n440 GND 0.06fF $ **FLOATING
C3205 CLK1.n441 GND 0.14fF $ **FLOATING
C3206 CLK1.n442 GND 0.11fF $ **FLOATING
C3207 CLK1.n443 GND 0.18fF $ **FLOATING
C3208 CLK1.n444 GND 0.03fF $ **FLOATING
C3209 CLK1.n445 GND 0.02fF $ **FLOATING
C3210 CLK1.n446 GND 0.02fF $ **FLOATING
C3211 CLK1.n447 GND 0.29fF $ **FLOATING
C3212 CLK1.n448 GND 0.03fF $ **FLOATING
C3213 CLK1.n449 GND 0.03fF $ **FLOATING
C3214 CLK1.n450 GND 0.02fF $ **FLOATING
C3215 CLK1.n451 GND 0.03fF $ **FLOATING
C3216 CLK1.n452 GND 0.16fF $ **FLOATING
C3217 CLK1.n453 GND 0.09fF $ **FLOATING
C3218 CLK1.t121 GND 0.09fF
C3219 CLK1.t8 GND 0.09fF
C3220 CLK1.n454 GND 0.17fF $ **FLOATING
C3221 CLK1.n455 GND 0.03fF $ **FLOATING
C3222 CLK1.n456 GND 0.02fF $ **FLOATING
C3223 CLK1.n457 GND 0.17fF $ **FLOATING
C3224 EESPFAL_s2_0/EESPFAL_INV4_1/CLK GND 0.02fF $ **FLOATING
C3225 CLK1.n458 GND 0.03fF $ **FLOATING
C3226 CLK1.n459 GND 0.03fF $ **FLOATING
C3227 CLK1.n460 GND 0.03fF $ **FLOATING
C3228 CLK1.n461 GND 0.02fF $ **FLOATING
C3229 CLK1.n462 GND 0.03fF $ **FLOATING
C3230 CLK1.n463 GND 0.16fF $ **FLOATING
C3231 CLK1.t10 GND 0.09fF
C3232 CLK1.n464 GND 0.11fF $ **FLOATING
C3233 CLK1.n465 GND 0.18fF $ **FLOATING
C3234 CLK1.n466 GND 0.03fF $ **FLOATING
C3235 CLK1.n467 GND 0.02fF $ **FLOATING
C3236 CLK1.n468 GND 0.02fF $ **FLOATING
C3237 CLK1.n469 GND 0.03fF $ **FLOATING
C3238 CLK1.n470 GND 0.03fF $ **FLOATING
C3239 CLK1.n471 GND 0.03fF $ **FLOATING
C3240 CLK1.n472 GND 0.02fF $ **FLOATING
C3241 CLK1.n473 GND 0.03fF $ **FLOATING
C3242 CLK1.n474 GND 0.06fF $ **FLOATING
C3243 CLK1.n475 GND 0.07fF $ **FLOATING
C3244 CLK1.n476 GND 0.15fF $ **FLOATING
C3245 CLK1.n477 GND 0.10fF $ **FLOATING
C3246 CLK1.n478 GND 0.21fF $ **FLOATING
C3247 CLK1.n479 GND 0.12fF $ **FLOATING
C3248 CLK1.n480 GND 0.03fF $ **FLOATING
C3249 CLK1.n481 GND 0.03fF $ **FLOATING
C3250 CLK1.n482 GND 0.02fF $ **FLOATING
C3251 CLK1.n483 GND 0.03fF $ **FLOATING
C3252 CLK1.n484 GND 0.06fF $ **FLOATING
C3253 CLK1.n485 GND 0.06fF $ **FLOATING
C3254 CLK1.n486 GND 0.06fF $ **FLOATING
C3255 CLK1.n487 GND 0.03fF $ **FLOATING
C3256 CLK1.n488 GND 0.02fF $ **FLOATING
C3257 CLK1.n489 GND 0.02fF $ **FLOATING
C3258 CLK1.n490 GND 0.02fF $ **FLOATING
C3259 CLK1.n491 GND 0.03fF $ **FLOATING
C3260 CLK1.t193 GND 0.09fF
C3261 CLK1.n492 GND 0.03fF $ **FLOATING
C3262 CLK1.n493 GND 0.02fF $ **FLOATING
C3263 CLK1.t194 GND 0.05fF
C3264 CLK1.n494 GND 0.29fF $ **FLOATING
C3265 CLK1.t124 GND 0.03fF
C3266 CLK1.t142 GND 0.03fF
C3267 CLK1.n495 GND 0.10fF $ **FLOATING
C3268 CLK1.n496 GND 0.17fF $ **FLOATING
C3269 CLK1.n497 GND 0.02fF $ **FLOATING
C3270 CLK1.n498 GND 0.03fF $ **FLOATING
C3271 CLK1.n499 GND 0.16fF $ **FLOATING
C3272 CLK1.n500 GND 0.16fF $ **FLOATING
C3273 CLK1.n501 GND 0.03fF $ **FLOATING
C3274 CLK1.n502 GND 0.02fF $ **FLOATING
C3275 EESPFAL_s2_0/EESPFAL_XOR_v3_0/CLK GND 0.02fF $ **FLOATING
C3276 CLK1.t48 GND 0.05fF
C3277 CLK1.n503 GND 0.29fF $ **FLOATING
C3278 CLK1.n504 GND 0.02fF $ **FLOATING
C3279 CLK1.n505 GND 0.03fF $ **FLOATING
C3280 CLK1.t47 GND 0.09fF
C3281 CLK1.n506 GND 0.06fF $ **FLOATING
C3282 CLK1.n507 GND 0.03fF $ **FLOATING
C3283 CLK1.n508 GND 0.02fF $ **FLOATING
C3284 CLK1.n509 GND 0.02fF $ **FLOATING
C3285 CLK1.n510 GND 0.03fF $ **FLOATING
C3286 CLK1.n511 GND 0.02fF $ **FLOATING
C3287 CLK1.n512 GND 0.03fF $ **FLOATING
C3288 CLK1.n513 GND 0.06fF $ **FLOATING
C3289 CLK1.n514 GND 0.03fF $ **FLOATING
C3290 CLK1.n515 GND 0.02fF $ **FLOATING
C3291 CLK1.t129 GND 0.03fF
C3292 CLK1.t169 GND 0.03fF
C3293 CLK1.n516 GND 0.15fF $ **FLOATING
C3294 CLK1.n517 GND 0.03fF $ **FLOATING
C3295 CLK1.n518 GND 0.02fF $ **FLOATING
C3296 CLK1.n519 GND 0.03fF $ **FLOATING
C3297 CLK1.n520 GND 0.00fF $ **FLOATING
C3298 EESPFAL_s3_0/CLK1 GND 0.00fF $ **FLOATING
C3299 CLK1.n521 GND 0.01fF $ **FLOATING
C3300 CLK1.t116 GND 0.08fF
C3301 CLK1.n522 GND 0.34fF $ **FLOATING
C3302 CLK1.n523 GND 0.02fF $ **FLOATING
C3303 CLK1.n524 GND 0.03fF $ **FLOATING
C3304 CLK1.n525 GND 0.06fF $ **FLOATING
C3305 CLK1.n526 GND 0.03fF $ **FLOATING
C3306 CLK1.n527 GND 0.02fF $ **FLOATING
C3307 CLK1.t66 GND 0.03fF
C3308 CLK1.t196 GND 0.03fF
C3309 CLK1.n528 GND 0.15fF $ **FLOATING
C3310 CLK1.n529 GND 0.19fF $ **FLOATING
C3311 CLK1.n530 GND 0.02fF $ **FLOATING
C3312 CLK1.n531 GND 0.03fF $ **FLOATING
C3313 CLK1.n532 GND 0.14fF $ **FLOATING
C3314 CLK1.n533 GND 0.03fF $ **FLOATING
C3315 CLK1.n534 GND 0.02fF $ **FLOATING
C3316 CLK1.t155 GND 0.05fF
C3317 CLK1.n535 GND 0.29fF $ **FLOATING
C3318 CLK1.n536 GND 0.02fF $ **FLOATING
C3319 CLK1.n537 GND 0.03fF $ **FLOATING
C3320 CLK1.n538 GND 0.09fF $ **FLOATING
C3321 CLK1.n539 GND 0.03fF $ **FLOATING
C3322 CLK1.n540 GND 0.02fF $ **FLOATING
C3323 CLK1.t159 GND 0.03fF
C3324 CLK1.t157 GND 0.03fF
C3325 CLK1.n541 GND 0.10fF $ **FLOATING
C3326 CLK1.n542 GND 0.03fF $ **FLOATING
C3327 CLK1.n543 GND 0.02fF $ **FLOATING
C3328 CLK1.n544 GND 0.03fF $ **FLOATING
C3329 CLK1.t160 GND 0.09fF
C3330 CLK1.n545 GND 0.03fF $ **FLOATING
C3331 CLK1.n546 GND 0.02fF $ **FLOATING
C3332 CLK1.t161 GND 0.05fF
C3333 CLK1.n547 GND 0.03fF $ **FLOATING
C3334 CLK1.n548 GND 0.02fF $ **FLOATING
C3335 CLK1.n549 GND 0.03fF $ **FLOATING
C3336 CLK1.n550 GND 0.06fF $ **FLOATING
C3337 CLK1.n551 GND 0.03fF $ **FLOATING
C3338 CLK1.n552 GND 0.02fF $ **FLOATING
C3339 CLK1.n553 GND 0.03fF $ **FLOATING
C3340 CLK1.n554 GND 0.02fF $ **FLOATING
C3341 CLK1.n555 GND 0.03fF $ **FLOATING
C3342 CLK1.n556 GND 0.07fF $ **FLOATING
C3343 CLK1.n557 GND 0.03fF $ **FLOATING
C3344 CLK1.n558 GND 0.02fF $ **FLOATING
C3345 CLK1.t50 GND 0.08fF
C3346 CLK1.n559 GND 0.13fF $ **FLOATING
C3347 CLK1.n560 GND 0.36fF $ **FLOATING
C3348 CLK1.n561 GND 0.02fF $ **FLOATING
C3349 CLK1.n562 GND 0.03fF $ **FLOATING
C3350 CLK1.n563 GND 0.02fF $ **FLOATING
C3351 CLK1.n564 GND 0.03fF $ **FLOATING
C3352 CLK1.n565 GND 0.06fF $ **FLOATING
C3353 CLK1.n566 GND 0.06fF $ **FLOATING
C3354 CLK1.n567 GND 0.06fF $ **FLOATING
C3355 CLK1.n568 GND 0.03fF $ **FLOATING
C3356 CLK1.n569 GND 0.02fF $ **FLOATING
C3357 CLK1.n570 GND 0.03fF $ **FLOATING
C3358 CLK1.n571 GND 0.03fF $ **FLOATING
C3359 CLK1.n572 GND 0.03fF $ **FLOATING
C3360 CLK1.n573 GND 0.02fF $ **FLOATING
C3361 CLK1.n574 GND 0.03fF $ **FLOATING
C3362 CLK1.n575 GND 0.06fF $ **FLOATING
C3363 CLK1.n576 GND 0.14fF $ **FLOATING
C3364 CLK1.n577 GND 0.11fF $ **FLOATING
C3365 CLK1.n578 GND 0.18fF $ **FLOATING
C3366 CLK1.n579 GND 0.03fF $ **FLOATING
C3367 CLK1.n580 GND 0.02fF $ **FLOATING
C3368 CLK1.n581 GND 0.02fF $ **FLOATING
C3369 CLK1.n582 GND 0.29fF $ **FLOATING
C3370 CLK1.n583 GND 0.03fF $ **FLOATING
C3371 CLK1.n584 GND 0.03fF $ **FLOATING
C3372 CLK1.n585 GND 0.02fF $ **FLOATING
C3373 CLK1.n586 GND 0.03fF $ **FLOATING
C3374 CLK1.n587 GND 0.16fF $ **FLOATING
C3375 CLK1.n588 GND 0.09fF $ **FLOATING
C3376 CLK1.t158 GND 0.09fF
C3377 CLK1.t156 GND 0.09fF
C3378 CLK1.n589 GND 0.17fF $ **FLOATING
C3379 CLK1.n590 GND 0.03fF $ **FLOATING
C3380 CLK1.n591 GND 0.02fF $ **FLOATING
C3381 CLK1.n592 GND 0.17fF $ **FLOATING
C3382 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/CLK GND 0.02fF $ **FLOATING
C3383 CLK1.n593 GND 0.03fF $ **FLOATING
C3384 CLK1.n594 GND 0.03fF $ **FLOATING
C3385 CLK1.n595 GND 0.03fF $ **FLOATING
C3386 CLK1.n596 GND 0.02fF $ **FLOATING
C3387 CLK1.n597 GND 0.03fF $ **FLOATING
C3388 CLK1.n598 GND 0.16fF $ **FLOATING
C3389 CLK1.t154 GND 0.09fF
C3390 CLK1.n599 GND 0.11fF $ **FLOATING
C3391 CLK1.n600 GND 0.18fF $ **FLOATING
C3392 CLK1.n601 GND 0.03fF $ **FLOATING
C3393 CLK1.n602 GND 0.02fF $ **FLOATING
C3394 CLK1.n603 GND 0.02fF $ **FLOATING
C3395 CLK1.n604 GND 0.03fF $ **FLOATING
C3396 CLK1.n605 GND 0.03fF $ **FLOATING
C3397 CLK1.n606 GND 0.03fF $ **FLOATING
C3398 CLK1.n607 GND 0.02fF $ **FLOATING
C3399 CLK1.n608 GND 0.03fF $ **FLOATING
C3400 CLK1.n609 GND 0.06fF $ **FLOATING
C3401 CLK1.n610 GND 0.06fF $ **FLOATING
C3402 CLK1.n611 GND 0.06fF $ **FLOATING
C3403 CLK1.n612 GND 0.03fF $ **FLOATING
C3404 CLK1.n613 GND 0.02fF $ **FLOATING
C3405 CLK1.n614 GND 0.02fF $ **FLOATING
C3406 CLK1.n615 GND 0.03fF $ **FLOATING
C3407 CLK1.n616 GND 0.02fF $ **FLOATING
C3408 CLK1.n617 GND 0.03fF $ **FLOATING
C3409 CLK1.n618 GND 0.02fF $ **FLOATING
C3410 CLK1.n619 GND 0.03fF $ **FLOATING
C3411 CLK1.n620 GND 0.06fF $ **FLOATING
C3412 CLK1.n621 GND 0.07fF $ **FLOATING
C3413 CLK1.n622 GND 0.13fF $ **FLOATING
C3414 CLK1.n623 GND 0.08fF $ **FLOATING
C3415 CLK1.n624 GND 0.13fF $ **FLOATING
C3416 CLK1.n625 GND 0.02fF $ **FLOATING
C3417 CLK1.n626 GND 0.01fF $ **FLOATING
C3418 CLK1.n627 GND 0.03fF $ **FLOATING
C3419 CLK1.n628 GND 0.06fF $ **FLOATING
C3420 CLK1.n629 GND 0.03fF $ **FLOATING
C3421 CLK1.n630 GND 0.02fF $ **FLOATING
C3422 CLK1.n631 GND 0.02fF $ **FLOATING
C3423 CLK1.t65 GND 0.03fF
C3424 CLK1.t68 GND 0.03fF
C3425 CLK1.n632 GND 0.15fF $ **FLOATING
C3426 CLK1.n633 GND 0.03fF $ **FLOATING
C3427 CLK1.n634 GND 0.02fF $ **FLOATING
C3428 CLK1.n635 GND 0.03fF $ **FLOATING
C3429 CLK1.n636 GND 0.06fF $ **FLOATING
C3430 CLK1.n637 GND 0.03fF $ **FLOATING
C3431 CLK1.n638 GND 0.02fF $ **FLOATING
C3432 CLK1.n639 GND 0.02fF $ **FLOATING
C3433 CLK1.n640 GND 0.02fF $ **FLOATING
C3434 CLK1.n641 GND 0.03fF $ **FLOATING
C3435 CLK1.t139 GND 0.09fF
C3436 CLK1.n642 GND 0.03fF $ **FLOATING
C3437 CLK1.n643 GND 0.02fF $ **FLOATING
C3438 EESPFAL_s3_0/EESPFAL_XOR_v3_1/CLK GND 0.02fF $ **FLOATING
C3439 CLK1.n644 GND 0.02fF $ **FLOATING
C3440 CLK1.n645 GND 0.03fF $ **FLOATING
C3441 CLK1.n646 GND 0.16fF $ **FLOATING
C3442 CLK1.n647 GND 0.03fF $ **FLOATING
C3443 CLK1.n648 GND 0.02fF $ **FLOATING
C3444 CLK1.t93 GND 0.05fF
C3445 CLK1.n649 GND 0.29fF $ **FLOATING
C3446 CLK1.n650 GND 0.02fF $ **FLOATING
C3447 CLK1.n651 GND 0.03fF $ **FLOATING
C3448 CLK1.n652 GND 0.06fF $ **FLOATING
C3449 CLK1.n653 GND 0.03fF $ **FLOATING
C3450 CLK1.n654 GND 0.02fF $ **FLOATING
C3451 CLK1.n655 GND 0.03fF $ **FLOATING
C3452 CLK1.n656 GND 0.02fF $ **FLOATING
C3453 CLK1.n657 GND 0.03fF $ **FLOATING
C3454 CLK1.n658 GND 0.06fF $ **FLOATING
C3455 CLK1.n659 GND 0.03fF $ **FLOATING
C3456 CLK1.n660 GND 0.02fF $ **FLOATING
C3457 CLK1.t90 GND 0.03fF
C3458 CLK1.t195 GND 0.03fF
C3459 CLK1.n661 GND 0.15fF $ **FLOATING
C3460 CLK1.n662 GND 0.03fF $ **FLOATING
C3461 CLK1.n663 GND 0.02fF $ **FLOATING
C3462 CLK1.n664 GND 0.03fF $ **FLOATING
C3463 CLK1.t149 GND 0.07fF
C3464 CLK1.n665 GND 0.45fF $ **FLOATING
C3465 CLK1.n666 GND 0.02fF $ **FLOATING
C3466 CLK1.n667 GND 0.03fF $ **FLOATING
C3467 CLK1.n668 GND 0.14fF $ **FLOATING
C3468 CLK1.n669 GND 0.03fF $ **FLOATING
C3469 CLK1.n670 GND 0.02fF $ **FLOATING
C3470 CLK1.t46 GND 0.05fF
C3471 CLK1.n671 GND 0.29fF $ **FLOATING
C3472 CLK1.n672 GND 0.02fF $ **FLOATING
C3473 CLK1.n673 GND 0.03fF $ **FLOATING
C3474 CLK1.n674 GND 0.09fF $ **FLOATING
C3475 CLK1.n675 GND 0.03fF $ **FLOATING
C3476 CLK1.n676 GND 0.02fF $ **FLOATING
C3477 CLK1.t79 GND 0.03fF
C3478 CLK1.t44 GND 0.03fF
C3479 CLK1.n677 GND 0.10fF $ **FLOATING
C3480 CLK1.n678 GND 0.03fF $ **FLOATING
C3481 CLK1.n679 GND 0.02fF $ **FLOATING
C3482 CLK1.n680 GND 0.03fF $ **FLOATING
C3483 CLK1.t76 GND 0.09fF
C3484 CLK1.n681 GND 0.03fF $ **FLOATING
C3485 CLK1.n682 GND 0.02fF $ **FLOATING
C3486 CLK1.t77 GND 0.05fF
C3487 CLK1.n683 GND 0.03fF $ **FLOATING
C3488 CLK1.n684 GND 0.02fF $ **FLOATING
C3489 CLK1.n685 GND 0.03fF $ **FLOATING
C3490 CLK1.n686 GND 0.07fF $ **FLOATING
C3491 CLK1.n687 GND 0.03fF $ **FLOATING
C3492 CLK1.n688 GND 0.02fF $ **FLOATING
C3493 CLK1.t56 GND 0.07fF
C3494 CLK1.n689 GND 0.15fF $ **FLOATING
C3495 CLK1.n690 GND 0.47fF $ **FLOATING
C3496 CLK1.n691 GND 0.03fF $ **FLOATING
C3497 CLK1.n692 GND 0.03fF $ **FLOATING
C3498 CLK1.n693 GND 0.02fF $ **FLOATING
C3499 CLK1.n694 GND 0.03fF $ **FLOATING
C3500 CLK1.n695 GND 0.06fF $ **FLOATING
C3501 CLK1.n696 GND 0.14fF $ **FLOATING
C3502 CLK1.n697 GND 0.11fF $ **FLOATING
C3503 CLK1.n698 GND 0.18fF $ **FLOATING
C3504 CLK1.n699 GND 0.03fF $ **FLOATING
C3505 CLK1.n700 GND 0.02fF $ **FLOATING
C3506 CLK1.n701 GND 0.02fF $ **FLOATING
C3507 CLK1.n702 GND 0.29fF $ **FLOATING
C3508 CLK1.n703 GND 0.03fF $ **FLOATING
C3509 CLK1.n704 GND 0.03fF $ **FLOATING
C3510 CLK1.n705 GND 0.02fF $ **FLOATING
C3511 CLK1.n706 GND 0.03fF $ **FLOATING
C3512 CLK1.n707 GND 0.16fF $ **FLOATING
C3513 CLK1.n708 GND 0.09fF $ **FLOATING
C3514 CLK1.t78 GND 0.09fF
C3515 CLK1.t43 GND 0.09fF
C3516 CLK1.n709 GND 0.17fF $ **FLOATING
C3517 CLK1.n710 GND 0.03fF $ **FLOATING
C3518 CLK1.n711 GND 0.02fF $ **FLOATING
C3519 CLK1.n712 GND 0.17fF $ **FLOATING
C3520 EESPFAL_s3_0/EESPFAL_INV4_1/CLK GND 0.02fF $ **FLOATING
C3521 CLK1.n713 GND 0.03fF $ **FLOATING
C3522 CLK1.n714 GND 0.03fF $ **FLOATING
C3523 CLK1.n715 GND 0.03fF $ **FLOATING
C3524 CLK1.n716 GND 0.02fF $ **FLOATING
C3525 CLK1.n717 GND 0.03fF $ **FLOATING
C3526 CLK1.n718 GND 0.16fF $ **FLOATING
C3527 CLK1.t45 GND 0.09fF
C3528 CLK1.n719 GND 0.11fF $ **FLOATING
C3529 CLK1.n720 GND 0.18fF $ **FLOATING
C3530 CLK1.n721 GND 0.03fF $ **FLOATING
C3531 CLK1.n722 GND 0.02fF $ **FLOATING
C3532 CLK1.n723 GND 0.02fF $ **FLOATING
C3533 CLK1.n724 GND 0.03fF $ **FLOATING
C3534 CLK1.n725 GND 0.03fF $ **FLOATING
C3535 CLK1.n726 GND 0.03fF $ **FLOATING
C3536 CLK1.n727 GND 0.02fF $ **FLOATING
C3537 CLK1.n728 GND 0.03fF $ **FLOATING
C3538 CLK1.n729 GND 0.06fF $ **FLOATING
C3539 CLK1.n730 GND 0.07fF $ **FLOATING
C3540 CLK1.n731 GND 0.15fF $ **FLOATING
C3541 CLK1.n732 GND 0.10fF $ **FLOATING
C3542 CLK1.n733 GND 0.11fF $ **FLOATING
C3543 CLK1.n734 GND 0.21fF $ **FLOATING
C3544 CLK1.n735 GND 0.08fF $ **FLOATING
C3545 CLK1.n736 GND 0.06fF $ **FLOATING
C3546 CLK1.n737 GND 0.03fF $ **FLOATING
C3547 CLK1.n738 GND 0.02fF $ **FLOATING
C3548 CLK1.n739 GND 0.03fF $ **FLOATING
C3549 CLK1.n740 GND 0.02fF $ **FLOATING
C3550 CLK1.n741 GND 0.19fF $ **FLOATING
C3551 CLK1.n742 GND 0.03fF $ **FLOATING
C3552 CLK1.n743 GND 0.02fF $ **FLOATING
C3553 CLK1.n744 GND 0.03fF $ **FLOATING
C3554 CLK1.n745 GND 0.06fF $ **FLOATING
C3555 CLK1.n746 GND 0.06fF $ **FLOATING
C3556 CLK1.n747 GND 0.06fF $ **FLOATING
C3557 CLK1.n748 GND 0.03fF $ **FLOATING
C3558 CLK1.n749 GND 0.02fF $ **FLOATING
C3559 CLK1.n750 GND 0.03fF $ **FLOATING
C3560 CLK1.n751 GND 0.03fF $ **FLOATING
C3561 CLK1.n752 GND 0.02fF $ **FLOATING
C3562 CLK1.n753 GND 0.03fF $ **FLOATING
C3563 CLK1.n754 GND 0.02fF $ **FLOATING
C3564 CLK1.n755 GND 0.03fF $ **FLOATING
C3565 CLK1.n756 GND 0.14fF $ **FLOATING
C3566 CLK1.n757 GND 0.18fF $ **FLOATING
C3567 CLK1.t92 GND 0.09fF
C3568 CLK1.n758 GND 0.11fF $ **FLOATING
C3569 CLK1.n759 GND 0.03fF $ **FLOATING
C3570 CLK1.n760 GND 0.02fF $ **FLOATING
C3571 CLK1.n761 GND 0.03fF $ **FLOATING
C3572 CLK1.n762 GND 0.03fF $ **FLOATING
C3573 CLK1.t153 GND 0.03fF
C3574 CLK1.t180 GND 0.03fF
C3575 CLK1.n763 GND 0.10fF $ **FLOATING
C3576 CLK1.n764 GND 0.17fF $ **FLOATING
C3577 CLK1.n765 GND 0.03fF $ **FLOATING
C3578 CLK1.n766 GND 0.02fF $ **FLOATING
C3579 CLK1.n767 GND 0.03fF $ **FLOATING
C3580 CLK1.n768 GND 0.09fF $ **FLOATING
C3581 CLK1.t152 GND 0.09fF
C3582 CLK1.n769 GND 0.17fF $ **FLOATING
C3583 CLK1.t179 GND 0.09fF
C3584 CLK1.n770 GND 0.16fF $ **FLOATING
C3585 CLK1.n771 GND 0.09fF $ **FLOATING
C3586 CLK1.n772 GND 0.03fF $ **FLOATING
C3587 CLK1.n773 GND 0.02fF $ **FLOATING
C3588 CLK1.n774 GND 0.03fF $ **FLOATING
C3589 CLK1.n775 GND 0.03fF $ **FLOATING
C3590 CLK1.t140 GND 0.05fF
C3591 CLK1.n776 GND 0.29fF $ **FLOATING
C3592 CLK1.n777 GND 0.03fF $ **FLOATING
C3593 CLK1.n778 GND 0.02fF $ **FLOATING
C3594 CLK1.n779 GND 0.03fF $ **FLOATING
C3595 CLK1.n780 GND 0.11fF $ **FLOATING
C3596 CLK1.n781 GND 0.18fF $ **FLOATING
C3597 CLK1.n782 GND 0.14fF $ **FLOATING
C3598 CLK1.n783 GND 0.03fF $ **FLOATING
C3599 CLK1.n784 GND 0.02fF $ **FLOATING
C3600 CLK1.n785 GND 0.03fF $ **FLOATING
C3601 CLK1.n786 GND 0.03fF $ **FLOATING
C3602 CLK1.n787 GND 0.03fF $ **FLOATING
C3603 CLK1.n788 GND 0.02fF $ **FLOATING
C3604 CLK1.n789 GND 0.03fF $ **FLOATING
C3605 CLK1.n790 GND 0.06fF $ **FLOATING
C3606 CLK1.n791 GND 0.06fF $ **FLOATING
C3607 CLK1.n792 GND 0.06fF $ **FLOATING
C3608 CLK1.n793 GND 0.03fF $ **FLOATING
C3609 CLK1.n794 GND 0.02fF $ **FLOATING
C3610 CLK1.n795 GND 0.03fF $ **FLOATING
C3611 CLK1.n796 GND 0.19fF $ **FLOATING
C3612 CLK1.n797 GND 0.02fF $ **FLOATING
C3613 CLK1.n798 GND 0.03fF $ **FLOATING
C3614 CLK1.n799 GND 0.03fF $ **FLOATING
C3615 CLK1.n800 GND 0.02fF $ **FLOATING
C3616 CLK1.n801 GND 0.03fF $ **FLOATING
C3617 CLK1.n802 GND 0.06fF $ **FLOATING
C3618 CLK1.n803 GND 0.08fF $ **FLOATING
C3619 CLK1.n804 GND 0.19fF $ **FLOATING
C3620 CLK1.n805 GND 0.01fF $ **FLOATING
C3621 CLK1.n806 GND 0.00fF $ **FLOATING
C3622 CLK1.n807 GND 0.03fF $ **FLOATING
C3623 CLK1.n808 GND 0.36fF $ **FLOATING
C3624 CLK1.n809 GND 0.36fF $ **FLOATING
C3625 CLK1.n810 GND 0.02fF $ **FLOATING
C3626 CLK1.n811 GND 0.01fF $ **FLOATING
C3627 CLK1.n812 GND 0.03fF $ **FLOATING
C3628 CLK1.n813 GND 0.06fF $ **FLOATING
C3629 CLK1.n814 GND 0.03fF $ **FLOATING
C3630 CLK1.n815 GND 0.02fF $ **FLOATING
C3631 CLK1.n816 GND 0.02fF $ **FLOATING
C3632 CLK1.t54 GND 0.03fF
C3633 CLK1.t148 GND 0.03fF
C3634 CLK1.n817 GND 0.15fF $ **FLOATING
C3635 CLK1.n818 GND 0.03fF $ **FLOATING
C3636 CLK1.n819 GND 0.02fF $ **FLOATING
C3637 CLK1.n820 GND 0.03fF $ **FLOATING
C3638 CLK1.n821 GND 0.06fF $ **FLOATING
C3639 CLK1.n822 GND 0.03fF $ **FLOATING
C3640 CLK1.n823 GND 0.02fF $ **FLOATING
C3641 CLK1.n824 GND 0.02fF $ **FLOATING
C3642 CLK1.n825 GND 0.02fF $ **FLOATING
C3643 CLK1.n826 GND 0.03fF $ **FLOATING
C3644 CLK1.t184 GND 0.09fF
C3645 CLK1.n827 GND 0.03fF $ **FLOATING
C3646 CLK1.n828 GND 0.02fF $ **FLOATING
C3647 EESPFAL_s3_0/EESPFAL_XOR_v3_0/CLK GND 0.02fF $ **FLOATING
C3648 CLK1.n829 GND 0.02fF $ **FLOATING
C3649 CLK1.n830 GND 0.03fF $ **FLOATING
C3650 CLK1.n831 GND 0.16fF $ **FLOATING
C3651 CLK1.n832 GND 0.03fF $ **FLOATING
C3652 CLK1.n833 GND 0.02fF $ **FLOATING
C3653 CLK1.t21 GND 0.05fF
C3654 CLK1.n834 GND 0.29fF $ **FLOATING
C3655 CLK1.n835 GND 0.02fF $ **FLOATING
C3656 CLK1.n836 GND 0.03fF $ **FLOATING
C3657 CLK1.n837 GND 0.06fF $ **FLOATING
C3658 CLK1.n838 GND 0.03fF $ **FLOATING
C3659 CLK1.n839 GND 0.02fF $ **FLOATING
C3660 CLK1.n840 GND 0.03fF $ **FLOATING
C3661 CLK1.n841 GND 0.02fF $ **FLOATING
C3662 CLK1.n842 GND 0.03fF $ **FLOATING
C3663 CLK1.n843 GND 0.06fF $ **FLOATING
C3664 CLK1.n844 GND 0.03fF $ **FLOATING
C3665 CLK1.n845 GND 0.02fF $ **FLOATING
C3666 CLK1.t186 GND 0.03fF
C3667 CLK1.t61 GND 0.03fF
C3668 CLK1.n846 GND 0.15fF $ **FLOATING
C3669 CLK1.n847 GND 0.03fF $ **FLOATING
C3670 CLK1.n848 GND 0.02fF $ **FLOATING
C3671 CLK1.n849 GND 0.03fF $ **FLOATING
C3672 CLK1.t198 GND 0.07fF
C3673 CLK1.n850 GND 0.45fF $ **FLOATING
C3674 CLK1.n851 GND 0.02fF $ **FLOATING
C3675 CLK1.n852 GND 0.03fF $ **FLOATING
C3676 CLK1.n853 GND 0.14fF $ **FLOATING
C3677 CLK1.n854 GND 0.03fF $ **FLOATING
C3678 CLK1.n855 GND 0.02fF $ **FLOATING
C3679 CLK1.t126 GND 0.05fF
C3680 CLK1.n856 GND 0.29fF $ **FLOATING
C3681 CLK1.n857 GND 0.02fF $ **FLOATING
C3682 CLK1.n858 GND 0.03fF $ **FLOATING
C3683 CLK1.n859 GND 0.09fF $ **FLOATING
C3684 CLK1.n860 GND 0.03fF $ **FLOATING
C3685 CLK1.n861 GND 0.02fF $ **FLOATING
C3686 CLK1.t73 GND 0.03fF
C3687 CLK1.t128 GND 0.03fF
C3688 CLK1.n862 GND 0.10fF $ **FLOATING
C3689 CLK1.n863 GND 0.03fF $ **FLOATING
C3690 CLK1.n864 GND 0.02fF $ **FLOATING
C3691 CLK1.n865 GND 0.03fF $ **FLOATING
C3692 CLK1.t74 GND 0.09fF
C3693 CLK1.n866 GND 0.03fF $ **FLOATING
C3694 CLK1.n867 GND 0.02fF $ **FLOATING
C3695 CLK1.t75 GND 0.05fF
C3696 CLK1.n868 GND 0.03fF $ **FLOATING
C3697 CLK1.n869 GND 0.02fF $ **FLOATING
C3698 CLK1.n870 GND 0.03fF $ **FLOATING
C3699 CLK1.n871 GND 0.07fF $ **FLOATING
C3700 CLK1.n872 GND 0.03fF $ **FLOATING
C3701 CLK1.n873 GND 0.02fF $ **FLOATING
C3702 CLK1.t134 GND 0.07fF
C3703 CLK1.n874 GND 0.15fF $ **FLOATING
C3704 CLK1.n875 GND 0.47fF $ **FLOATING
C3705 CLK1.n876 GND 0.03fF $ **FLOATING
C3706 CLK1.n877 GND 0.03fF $ **FLOATING
C3707 CLK1.n878 GND 0.02fF $ **FLOATING
C3708 CLK1.n879 GND 0.03fF $ **FLOATING
C3709 CLK1.n880 GND 0.06fF $ **FLOATING
C3710 CLK1.n881 GND 0.14fF $ **FLOATING
C3711 CLK1.n882 GND 0.11fF $ **FLOATING
C3712 CLK1.n883 GND 0.18fF $ **FLOATING
C3713 CLK1.n884 GND 0.03fF $ **FLOATING
C3714 CLK1.n885 GND 0.02fF $ **FLOATING
C3715 CLK1.n886 GND 0.02fF $ **FLOATING
C3716 CLK1.n887 GND 0.29fF $ **FLOATING
C3717 CLK1.n888 GND 0.03fF $ **FLOATING
C3718 CLK1.n889 GND 0.03fF $ **FLOATING
C3719 CLK1.n890 GND 0.02fF $ **FLOATING
C3720 CLK1.n891 GND 0.03fF $ **FLOATING
C3721 CLK1.n892 GND 0.16fF $ **FLOATING
C3722 CLK1.n893 GND 0.09fF $ **FLOATING
C3723 CLK1.t72 GND 0.09fF
C3724 CLK1.t127 GND 0.09fF
C3725 CLK1.n894 GND 0.17fF $ **FLOATING
C3726 CLK1.n895 GND 0.03fF $ **FLOATING
C3727 CLK1.n896 GND 0.02fF $ **FLOATING
C3728 CLK1.n897 GND 0.17fF $ **FLOATING
C3729 EESPFAL_s3_0/EESPFAL_INV4_2/CLK GND 0.02fF $ **FLOATING
C3730 CLK1.n898 GND 0.03fF $ **FLOATING
C3731 CLK1.n899 GND 0.03fF $ **FLOATING
C3732 CLK1.n900 GND 0.03fF $ **FLOATING
C3733 CLK1.n901 GND 0.02fF $ **FLOATING
C3734 CLK1.n902 GND 0.03fF $ **FLOATING
C3735 CLK1.n903 GND 0.16fF $ **FLOATING
C3736 CLK1.t125 GND 0.09fF
C3737 CLK1.n904 GND 0.11fF $ **FLOATING
C3738 CLK1.n905 GND 0.18fF $ **FLOATING
C3739 CLK1.n906 GND 0.03fF $ **FLOATING
C3740 CLK1.n907 GND 0.02fF $ **FLOATING
C3741 CLK1.n908 GND 0.02fF $ **FLOATING
C3742 CLK1.n909 GND 0.03fF $ **FLOATING
C3743 CLK1.n910 GND 0.03fF $ **FLOATING
C3744 CLK1.n911 GND 0.03fF $ **FLOATING
C3745 CLK1.n912 GND 0.02fF $ **FLOATING
C3746 CLK1.n913 GND 0.03fF $ **FLOATING
C3747 CLK1.n914 GND 0.06fF $ **FLOATING
C3748 CLK1.n915 GND 0.07fF $ **FLOATING
C3749 CLK1.n916 GND 0.15fF $ **FLOATING
C3750 CLK1.n917 GND 0.10fF $ **FLOATING
C3751 CLK1.n918 GND 0.11fF $ **FLOATING
C3752 CLK1.n919 GND 0.21fF $ **FLOATING
C3753 CLK1.n920 GND 0.08fF $ **FLOATING
C3754 CLK1.n921 GND 0.06fF $ **FLOATING
C3755 CLK1.n922 GND 0.03fF $ **FLOATING
C3756 CLK1.n923 GND 0.02fF $ **FLOATING
C3757 CLK1.n924 GND 0.03fF $ **FLOATING
C3758 CLK1.n925 GND 0.02fF $ **FLOATING
C3759 CLK1.n926 GND 0.19fF $ **FLOATING
C3760 CLK1.n927 GND 0.03fF $ **FLOATING
C3761 CLK1.n928 GND 0.02fF $ **FLOATING
C3762 CLK1.n929 GND 0.03fF $ **FLOATING
C3763 CLK1.n930 GND 0.06fF $ **FLOATING
C3764 CLK1.n931 GND 0.06fF $ **FLOATING
C3765 CLK1.n932 GND 0.06fF $ **FLOATING
C3766 CLK1.n933 GND 0.03fF $ **FLOATING
C3767 CLK1.n934 GND 0.02fF $ **FLOATING
C3768 CLK1.n935 GND 0.03fF $ **FLOATING
C3769 CLK1.n936 GND 0.03fF $ **FLOATING
C3770 CLK1.n937 GND 0.02fF $ **FLOATING
C3771 CLK1.n938 GND 0.03fF $ **FLOATING
C3772 CLK1.n939 GND 0.02fF $ **FLOATING
C3773 CLK1.n940 GND 0.03fF $ **FLOATING
C3774 CLK1.n941 GND 0.14fF $ **FLOATING
C3775 CLK1.n942 GND 0.18fF $ **FLOATING
C3776 CLK1.t20 GND 0.09fF
C3777 CLK1.n943 GND 0.11fF $ **FLOATING
C3778 CLK1.n944 GND 0.03fF $ **FLOATING
C3779 CLK1.n945 GND 0.02fF $ **FLOATING
C3780 CLK1.n946 GND 0.03fF $ **FLOATING
C3781 CLK1.n947 GND 0.03fF $ **FLOATING
C3782 CLK1.t113 GND 0.03fF
C3783 CLK1.t39 GND 0.03fF
C3784 CLK1.n948 GND 0.10fF $ **FLOATING
C3785 CLK1.n949 GND 0.17fF $ **FLOATING
C3786 CLK1.n950 GND 0.03fF $ **FLOATING
C3787 CLK1.n951 GND 0.02fF $ **FLOATING
C3788 CLK1.n952 GND 0.03fF $ **FLOATING
C3789 CLK1.n953 GND 0.09fF $ **FLOATING
C3790 CLK1.t112 GND 0.09fF
C3791 CLK1.n954 GND 0.17fF $ **FLOATING
C3792 CLK1.t38 GND 0.09fF
C3793 CLK1.n955 GND 0.16fF $ **FLOATING
C3794 CLK1.n956 GND 0.09fF $ **FLOATING
C3795 CLK1.n957 GND 0.03fF $ **FLOATING
C3796 CLK1.n958 GND 0.02fF $ **FLOATING
C3797 CLK1.n959 GND 0.03fF $ **FLOATING
C3798 CLK1.n960 GND 0.03fF $ **FLOATING
C3799 CLK1.t185 GND 0.05fF
C3800 CLK1.n961 GND 0.29fF $ **FLOATING
C3801 CLK1.n962 GND 0.03fF $ **FLOATING
C3802 CLK1.n963 GND 0.02fF $ **FLOATING
C3803 CLK1.n964 GND 0.03fF $ **FLOATING
C3804 CLK1.n965 GND 0.11fF $ **FLOATING
C3805 CLK1.n966 GND 0.18fF $ **FLOATING
C3806 CLK1.n967 GND 0.14fF $ **FLOATING
C3807 CLK1.n968 GND 0.03fF $ **FLOATING
C3808 CLK1.n969 GND 0.02fF $ **FLOATING
C3809 CLK1.n970 GND 0.03fF $ **FLOATING
C3810 CLK1.n971 GND 0.03fF $ **FLOATING
C3811 CLK1.n972 GND 0.03fF $ **FLOATING
C3812 CLK1.n973 GND 0.02fF $ **FLOATING
C3813 CLK1.n974 GND 0.03fF $ **FLOATING
C3814 CLK1.n975 GND 0.06fF $ **FLOATING
C3815 CLK1.n976 GND 0.06fF $ **FLOATING
C3816 CLK1.n977 GND 0.06fF $ **FLOATING
C3817 CLK1.n978 GND 0.03fF $ **FLOATING
C3818 CLK1.n979 GND 0.02fF $ **FLOATING
C3819 CLK1.n980 GND 0.03fF $ **FLOATING
C3820 CLK1.n981 GND 0.19fF $ **FLOATING
C3821 CLK1.n982 GND 0.02fF $ **FLOATING
C3822 CLK1.n983 GND 0.03fF $ **FLOATING
C3823 CLK1.n984 GND 0.03fF $ **FLOATING
C3824 CLK1.n985 GND 0.02fF $ **FLOATING
C3825 CLK1.n986 GND 0.03fF $ **FLOATING
C3826 CLK1.n987 GND 0.06fF $ **FLOATING
C3827 CLK1.n988 GND 0.08fF $ **FLOATING
C3828 CLK1.n989 GND 0.19fF $ **FLOATING
C3829 CLK1.n990 GND 0.01fF $ **FLOATING
C3830 CLK1.n991 GND 0.00fF $ **FLOATING
C3831 CLK1.n992 GND 0.03fF $ **FLOATING
C3832 CLK1.n993 GND 0.07fF $ **FLOATING
C3833 CLK1.n994 GND 0.08fF $ **FLOATING
C3834 EESPFAL_s2_0/CLK1 GND 0.02fF $ **FLOATING
C3835 CLK1.n995 GND 0.01fF $ **FLOATING
C3836 CLK1.n996 GND 0.04fF $ **FLOATING
C3837 CLK1.n997 GND 0.21fF $ **FLOATING
C3838 CLK1.n998 GND 0.08fF $ **FLOATING
C3839 CLK1.n999 GND 0.06fF $ **FLOATING
C3840 CLK1.n1000 GND 0.03fF $ **FLOATING
C3841 CLK1.n1001 GND 0.02fF $ **FLOATING
C3842 CLK1.n1002 GND 0.03fF $ **FLOATING
C3843 CLK1.n1003 GND 0.02fF $ **FLOATING
C3844 CLK1.n1004 GND 0.19fF $ **FLOATING
C3845 CLK1.n1005 GND 0.03fF $ **FLOATING
C3846 CLK1.n1006 GND 0.02fF $ **FLOATING
C3847 CLK1.n1007 GND 0.03fF $ **FLOATING
C3848 CLK1.n1008 GND 0.06fF $ **FLOATING
C3849 CLK1.n1009 GND 0.06fF $ **FLOATING
C3850 CLK1.n1010 GND 0.06fF $ **FLOATING
C3851 CLK1.n1011 GND 0.03fF $ **FLOATING
C3852 CLK1.n1012 GND 0.02fF $ **FLOATING
C3853 CLK1.n1013 GND 0.03fF $ **FLOATING
C3854 CLK1.n1014 GND 0.03fF $ **FLOATING
C3855 CLK1.n1015 GND 0.03fF $ **FLOATING
C3856 CLK1.n1016 GND 0.02fF $ **FLOATING
C3857 CLK1.n1017 GND 0.03fF $ **FLOATING
C3858 CLK1.n1018 GND 0.14fF $ **FLOATING
C3859 CLK1.n1019 GND 0.18fF $ **FLOATING
C3860 CLK1.n1020 GND 0.11fF $ **FLOATING
C3861 CLK1.n1021 GND 0.03fF $ **FLOATING
C3862 CLK1.n1022 GND 0.02fF $ **FLOATING
C3863 CLK1.n1023 GND 0.03fF $ **FLOATING
C3864 CLK1.n1024 GND 0.03fF $ **FLOATING
C3865 CLK1.n1025 GND 0.03fF $ **FLOATING
C3866 CLK1.n1026 GND 0.02fF $ **FLOATING
C3867 CLK1.n1027 GND 0.03fF $ **FLOATING
C3868 CLK1.n1028 GND 0.09fF $ **FLOATING
C3869 CLK1.t141 GND 0.09fF
C3870 CLK1.n1029 GND 0.17fF $ **FLOATING
C3871 CLK1.t123 GND 0.09fF
C3872 CLK1.n1030 GND 0.09fF $ **FLOATING
C3873 CLK1.n1031 GND 0.03fF $ **FLOATING
C3874 CLK1.n1032 GND 0.02fF $ **FLOATING
C3875 CLK1.n1033 GND 0.03fF $ **FLOATING
C3876 CLK1.n1034 GND 0.03fF $ **FLOATING
C3877 CLK1.n1035 GND 0.03fF $ **FLOATING
C3878 CLK1.n1036 GND 0.02fF $ **FLOATING
C3879 CLK1.n1037 GND 0.03fF $ **FLOATING
C3880 CLK1.n1038 GND 0.11fF $ **FLOATING
C3881 CLK1.n1039 GND 0.18fF $ **FLOATING
C3882 CLK1.n1040 GND 0.14fF $ **FLOATING
C3883 CLK1.n1041 GND 0.03fF $ **FLOATING
C3884 CLK1.n1042 GND 0.02fF $ **FLOATING
C3885 CLK1.n1043 GND 0.03fF $ **FLOATING
C3886 CLK1.n1044 GND 0.03fF $ **FLOATING
C3887 CLK1.n1045 GND 0.03fF $ **FLOATING
C3888 CLK1.n1046 GND 0.02fF $ **FLOATING
C3889 CLK1.n1047 GND 0.03fF $ **FLOATING
C3890 CLK1.n1048 GND 0.06fF $ **FLOATING
C3891 CLK1.n1049 GND 0.06fF $ **FLOATING
C3892 CLK1.n1050 GND 0.06fF $ **FLOATING
C3893 CLK1.n1051 GND 0.03fF $ **FLOATING
C3894 CLK1.n1052 GND 0.02fF $ **FLOATING
C3895 CLK1.n1053 GND 0.03fF $ **FLOATING
C3896 CLK1.n1054 GND 0.07fF $ **FLOATING
C3897 CLK1.n1055 GND 0.09fF $ **FLOATING
C3898 CLK1.n1056 GND 0.02fF $ **FLOATING
C3899 CLK1.t162 GND 0.03fF
C3900 CLK1.n1057 GND 0.07fF $ **FLOATING
C3901 CLK1.n1058 GND 0.02fF $ **FLOATING
C3902 CLK1.n1059 GND 0.08fF $ **FLOATING
C3903 CLK1.n1060 GND 0.09fF $ **FLOATING
C3904 CLK1.t7 GND 0.03fF
C3905 CLK1.t59 GND 0.03fF
C3906 CLK1.n1061 GND 0.07fF $ **FLOATING
C3907 CLK1.n1062 GND 0.01fF $ **FLOATING
C3908 CLK1.n1063 GND 0.02fF $ **FLOATING
C3909 CLK1.n1064 GND 0.02fF $ **FLOATING
C3910 CLK1.n1065 GND 0.08fF $ **FLOATING
C3911 CLK1.n1066 GND 0.07fF $ **FLOATING
C3912 CLK1.n1067 GND 0.07fF $ **FLOATING
C3913 CLK1.n1068 GND 0.07fF $ **FLOATING
C3914 CLK1.n1069 GND 0.10fF $ **FLOATING
C3915 CLK1.n1070 GND 0.07fF $ **FLOATING
C3916 CLK1.n1071 GND 0.07fF $ **FLOATING
C3917 CLK1.n1072 GND 0.05fF $ **FLOATING
C3918 CLK1.n1073 GND 0.07fF $ **FLOATING
C3919 CLK1.n1074 GND 0.25fF $ **FLOATING
C3920 CLK1.n1075 GND 0.34fF $ **FLOATING
C3921 CLK1.n1076 GND 0.20fF $ **FLOATING
C3922 CLK1.n1077 GND 0.07fF $ **FLOATING
C3923 CLK1.n1078 GND 0.07fF $ **FLOATING
C3924 CLK1.t181 GND 0.05fF
C3925 CLK1.t85 GND 0.05fF
C3926 CLK1.n1079 GND 0.59fF $ **FLOATING
C3927 CLK1.t182 GND 0.03fF
C3928 CLK1.t107 GND 0.03fF
C3929 CLK1.n1080 GND 0.10fF $ **FLOATING
C3930 CLK1.t87 GND 0.03fF
C3931 CLK1.t99 GND 0.03fF
C3932 CLK1.n1081 GND 0.10fF $ **FLOATING
C3933 CLK1.n1082 GND 0.36fF $ **FLOATING
C3934 CLK1.n1083 GND 0.07fF $ **FLOATING
C3935 CLK1.t84 GND 0.17fF
C3936 CLK1.n1084 GND 0.31fF $ **FLOATING
C3937 CLK1.n1085 GND 0.18fF $ **FLOATING
C3938 CLK1.t86 GND 0.17fF
C3939 CLK1.n1086 GND 0.32fF $ **FLOATING
C3940 CLK1.t98 GND 0.17fF
C3941 CLK1.n1087 GND 0.18fF $ **FLOATING
C3942 CLK1.n1088 GND 0.07fF $ **FLOATING
C3943 CLK1.n1089 GND 0.07fF $ **FLOATING
C3944 EESPFAL_s2_0/EESPFAL_XOR_v3_1/CLK GND 0.04fF $ **FLOATING
C3945 CLK1.t106 GND 0.05fF
C3946 CLK1.t97 GND 0.05fF
C3947 CLK1.n1090 GND 0.59fF $ **FLOATING
C3948 CLK1.n1091 GND 0.07fF $ **FLOATING
C3949 CLK1.n1092 GND 0.31fF $ **FLOATING
C3950 CLK1.t96 GND 0.17fF
C3951 CLK1.n1093 GND 0.20fF $ **FLOATING
C3952 CLK1.n1094 GND 0.34fF $ **FLOATING
C3953 CLK1.n1095 GND 0.25fF $ **FLOATING
C3954 CLK1.n1096 GND 0.07fF $ **FLOATING
C3955 CLK1.n1097 GND 0.07fF $ **FLOATING
C3956 CLK1.n1098 GND 0.05fF $ **FLOATING
C3957 CLK1.t183 GND 0.03fF
C3958 CLK1.t6 GND 0.03fF
C3959 CLK1.n1099 GND 0.18fF $ **FLOATING
C3960 CLK1.n1100 GND 0.23fF $ **FLOATING
C3961 CLK1.n1101 GND 0.07fF $ **FLOATING
C3962 CLK1.n1102 GND 0.07fF $ **FLOATING
C3963 CLK1.n1103 GND 0.10fF $ **FLOATING
C3964 CLK1.n1104 GND 0.10fF $ **FLOATING
C3965 CLK1.n1105 GND 0.07fF $ **FLOATING
C3966 CLK1.n1106 GND 0.07fF $ **FLOATING
C3967 CLK1.n1107 GND 0.04fF $ **FLOATING
C3968 CLK1.t55 GND 0.03fF
C3969 CLK1.t31 GND 0.03fF
C3970 CLK1.n1108 GND 0.15fF $ **FLOATING
C3971 CLK1.t114 GND 0.03fF
C3972 CLK1.t28 GND 0.03fF
C3973 CLK1.n1109 GND 0.18fF $ **FLOATING
C3974 CLK1.n1110 GND 0.23fF $ **FLOATING
C3975 CLK1.n1111 GND 0.07fF $ **FLOATING
C3976 CLK1.n1112 GND 0.07fF $ **FLOATING
C3977 CLK1.n1113 GND 0.19fF $ **FLOATING
C3978 CLK1.n1114 GND 0.29fF $ **FLOATING
C3979 CLK1.n1115 GND 0.07fF $ **FLOATING
C3980 CLK1.n1116 GND 0.07fF $ **FLOATING
C3981 CLK1.n1117 GND 0.14fF $ **FLOATING
C3982 CLK1.n1118 GND 0.10fF $ **FLOATING
C3983 CLK1.n1119 GND 0.10fF $ **FLOATING
C3984 CLK1.n1120 GND 0.07fF $ **FLOATING
C3985 CLK1.n1121 GND 0.07fF $ **FLOATING
C3986 CLK1.n1122 GND 0.06fF $ **FLOATING
C3987 CLK1.n1123 GND 0.05fF $ **FLOATING
C3988 CLK1.n1124 GND 0.21fF $ **FLOATING
C3989 CLK1.n1125 GND 0.06fF $ **FLOATING
C3990 CLK1.n1126 GND 0.07fF $ **FLOATING
C3991 CLK1.n1127 GND 0.07fF $ **FLOATING
C3992 CLK1.n1128 GND 0.10fF $ **FLOATING
C3993 CLK1.n1129 GND 0.10fF $ **FLOATING
C3994 CLK1.n1130 GND 0.10fF $ **FLOATING
C3995 CLK1.n1131 GND 0.07fF $ **FLOATING
C3996 CLK1.n1132 GND 0.07fF $ **FLOATING
C3997 CLK1.n1133 GND 0.07fF $ **FLOATING
C3998 CLK1.n1134 GND 0.07fF $ **FLOATING
C3999 CLK1.n1135 GND 0.07fF $ **FLOATING
C4000 CLK1.n1136 GND 0.07fF $ **FLOATING
C4001 CLK1.n1137 GND 0.07fF $ **FLOATING
C4002 CLK1.n1138 GND 0.07fF $ **FLOATING
C4003 CLK1.n1139 GND 0.07fF $ **FLOATING
C4004 CLK1.n1140 GND 0.07fF $ **FLOATING
C4005 CLK1.n1141 GND 0.06fF $ **FLOATING
C4006 CLK1.n1142 GND 0.07fF $ **FLOATING
C4007 CLK1.n1143 GND 0.06fF $ **FLOATING
C4008 CLK1.n1144 GND 0.07fF $ **FLOATING
C4009 CLK1.n1145 GND 0.07fF $ **FLOATING
C4010 CLK1.n1146 GND 0.07fF $ **FLOATING
C4011 CLK1.n1147 GND 0.07fF $ **FLOATING
C4012 CLK1.n1148 GND 0.07fF $ **FLOATING
C4013 CLK1.n1149 GND 0.07fF $ **FLOATING
C4014 CLK1.n1150 GND 0.07fF $ **FLOATING
C4015 CLK1.n1151 GND 0.06fF $ **FLOATING
C4016 CLK1.n1152 GND 0.07fF $ **FLOATING
C4017 CLK1.n1153 GND 0.07fF $ **FLOATING
C4018 CLK1.n1154 GND 0.07fF $ **FLOATING
C4019 CLK1.n1155 GND 0.07fF $ **FLOATING
C4020 CLK1.n1156 GND 0.07fF $ **FLOATING
C4021 CLK1.n1157 GND 0.07fF $ **FLOATING
C4022 CLK1.n1158 GND 0.07fF $ **FLOATING
C4023 CLK1.n1159 GND 0.07fF $ **FLOATING
C4024 CLK1.n1160 GND 0.07fF $ **FLOATING
C4025 CLK1.n1161 GND 0.07fF $ **FLOATING
C4026 CLK1.n1162 GND 0.10fF $ **FLOATING
C4027 CLK1.n1163 GND 0.10fF $ **FLOATING
C4028 CLK1.n1164 GND 0.10fF $ **FLOATING
C4029 CLK1.n1165 GND 0.07fF $ **FLOATING
C4030 CLK1.n1166 GND 0.07fF $ **FLOATING
C4031 CLK1.n1167 GND 0.06fF $ **FLOATING
C4032 CLK1.n1168 GND 0.09fF $ **FLOATING
C4033 CLK1.n1169 GND 0.05fF $ **FLOATING
C4034 CLK1.n1170 GND 0.07fF $ **FLOATING
C4035 CLK1.n1171 GND 0.07fF $ **FLOATING
C4036 CLK1.n1172 GND 0.07fF $ **FLOATING
C4037 CLK1.n1173 GND 0.10fF $ **FLOATING
C4038 CLK1.n1174 GND 0.10fF $ **FLOATING
C4039 CLK1.n1175 GND 0.13fF $ **FLOATING
C4040 CLK1.n1176 GND 0.07fF $ **FLOATING
C4041 CLK1.n1177 GND 0.07fF $ **FLOATING
C4042 CLK1.n1178 GND 0.06fF $ **FLOATING
C4043 CLK1.n1179 GND 0.12fF $ **FLOATING
C4044 CLK1.n1180 GND 0.10fF $ **FLOATING
C4045 CLK1.n1181 GND 0.03fF $ **FLOATING
C4046 CLK1.n1182 GND 0.10fF $ **FLOATING
C4047 CLK1.n1183 GND 0.01fF $ **FLOATING
C4048 CLK1.n1184 GND 0.11fF $ **FLOATING
C4049 CLK1.n1185 GND 0.10fF $ **FLOATING
C4050 CLK1.t172 GND 0.03fF
C4051 CLK1.n1186 GND 0.10fF $ **FLOATING
C4052 CLK1.n1187 GND 0.02fF $ **FLOATING
C4053 CLK1.n1188 GND 0.02fF $ **FLOATING
C4054 CLK1.n1189 GND 0.02fF $ **FLOATING
C4055 CLK1.n1190 GND 0.09fF $ **FLOATING
C4056 CLK1.n1191 GND 0.13fF $ **FLOATING
C4057 CLK1.n1192 GND 0.09fF $ **FLOATING
C4058 CLK1.n1193 GND 0.02fF $ **FLOATING
C4059 CLK1.n1194 GND 0.03fF $ **FLOATING
C4060 CLK1.n1195 GND 0.02fF $ **FLOATING
C4061 CLK1.n1196 GND 0.03fF $ **FLOATING
C4062 CLK1.n1197 GND 0.06fF $ **FLOATING
C4063 CLK1.n1198 GND 0.06fF $ **FLOATING
C4064 CLK1.n1199 GND 0.06fF $ **FLOATING
C4065 CLK1.n1200 GND 0.03fF $ **FLOATING
C4066 CLK1.n1201 GND 0.02fF $ **FLOATING
C4067 CLK1.n1202 GND 0.03fF $ **FLOATING
C4068 CLK1.n1203 GND 0.03fF $ **FLOATING
C4069 CLK1.n1204 GND 0.03fF $ **FLOATING
C4070 CLK1.n1205 GND 0.02fF $ **FLOATING
C4071 CLK1.n1206 GND 0.03fF $ **FLOATING
C4072 CLK1.n1207 GND 0.06fF $ **FLOATING
C4073 CLK1.n1208 GND 0.14fF $ **FLOATING
C4074 CLK1.n1209 GND 0.11fF $ **FLOATING
C4075 CLK1.n1210 GND 0.18fF $ **FLOATING
C4076 CLK1.n1211 GND 0.03fF $ **FLOATING
C4077 CLK1.n1212 GND 0.02fF $ **FLOATING
C4078 CLK1.n1213 GND 0.02fF $ **FLOATING
C4079 CLK1.n1214 GND 0.29fF $ **FLOATING
C4080 CLK1.n1215 GND 0.03fF $ **FLOATING
C4081 CLK1.n1216 GND 0.03fF $ **FLOATING
C4082 CLK1.n1217 GND 0.02fF $ **FLOATING
C4083 CLK1.n1218 GND 0.03fF $ **FLOATING
C4084 CLK1.n1219 GND 0.16fF $ **FLOATING
C4085 CLK1.n1220 GND 0.09fF $ **FLOATING
C4086 CLK1.t34 GND 0.09fF
C4087 CLK1.t135 GND 0.09fF
C4088 CLK1.n1221 GND 0.17fF $ **FLOATING
C4089 CLK1.n1222 GND 0.03fF $ **FLOATING
C4090 CLK1.n1223 GND 0.02fF $ **FLOATING
C4091 CLK1.n1224 GND 0.17fF $ **FLOATING
C4092 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/CLK GND 0.02fF $ **FLOATING
C4093 CLK1.n1225 GND 0.03fF $ **FLOATING
C4094 CLK1.n1226 GND 0.03fF $ **FLOATING
C4095 CLK1.n1227 GND 0.03fF $ **FLOATING
C4096 CLK1.n1228 GND 0.02fF $ **FLOATING
C4097 CLK1.n1229 GND 0.03fF $ **FLOATING
C4098 CLK1.n1230 GND 0.16fF $ **FLOATING
C4099 CLK1.t137 GND 0.09fF
C4100 CLK1.n1231 GND 0.11fF $ **FLOATING
C4101 CLK1.n1232 GND 0.18fF $ **FLOATING
C4102 CLK1.n1233 GND 0.03fF $ **FLOATING
C4103 CLK1.n1234 GND 0.02fF $ **FLOATING
C4104 CLK1.n1235 GND 0.02fF $ **FLOATING
C4105 CLK1.n1236 GND 0.03fF $ **FLOATING
C4106 CLK1.n1237 GND 0.03fF $ **FLOATING
C4107 CLK1.n1238 GND 0.03fF $ **FLOATING
C4108 CLK1.n1239 GND 0.02fF $ **FLOATING
C4109 CLK1.n1240 GND 0.03fF $ **FLOATING
C4110 CLK1.n1241 GND 0.06fF $ **FLOATING
C4111 CLK1.n1242 GND 0.06fF $ **FLOATING
C4112 CLK1.n1243 GND 0.06fF $ **FLOATING
C4113 CLK1.n1244 GND 0.03fF $ **FLOATING
C4114 CLK1.n1245 GND 0.02fF $ **FLOATING
C4115 CLK1.n1246 GND 0.02fF $ **FLOATING
C4116 CLK1.n1247 GND 0.03fF $ **FLOATING
C4117 CLK1.n1248 GND 0.02fF $ **FLOATING
C4118 CLK1.n1249 GND 0.03fF $ **FLOATING
C4119 CLK1.n1250 GND 0.02fF $ **FLOATING
C4120 CLK1.n1251 GND 0.03fF $ **FLOATING
C4121 CLK1.n1252 GND 0.06fF $ **FLOATING
C4122 CLK1.n1253 GND 0.07fF $ **FLOATING
C4123 CLK1.n1254 GND 0.13fF $ **FLOATING
C4124 CLK1.n1255 GND 0.08fF $ **FLOATING
C4125 CLK1.n1256 GND 0.13fF $ **FLOATING
C4126 CLK1.n1257 GND 0.02fF $ **FLOATING
C4127 CLK1.n1258 GND 0.01fF $ **FLOATING
C4128 CLK1.n1259 GND 0.03fF $ **FLOATING
C4129 CLK1.n1260 GND 0.06fF $ **FLOATING
C4130 CLK1.n1261 GND 0.03fF $ **FLOATING
C4131 CLK1.n1262 GND 0.02fF $ **FLOATING
C4132 CLK1.n1263 GND 0.02fF $ **FLOATING
C4133 CLK1.t62 GND 0.03fF
C4134 CLK1.t101 GND 0.03fF
C4135 CLK1.n1264 GND 0.15fF $ **FLOATING
C4136 CLK1.n1265 GND 0.03fF $ **FLOATING
C4137 CLK1.n1266 GND 0.02fF $ **FLOATING
C4138 CLK1.n1267 GND 0.03fF $ **FLOATING
C4139 CLK1.n1268 GND 0.06fF $ **FLOATING
C4140 CLK1.n1269 GND 0.03fF $ **FLOATING
C4141 CLK1.n1270 GND 0.02fF $ **FLOATING
C4142 CLK1.n1271 GND 0.02fF $ **FLOATING
C4143 CLK1.n1272 GND 0.02fF $ **FLOATING
C4144 CLK1.n1273 GND 0.03fF $ **FLOATING
C4145 CLK1.t132 GND 0.09fF
C4146 CLK1.n1274 GND 0.03fF $ **FLOATING
C4147 CLK1.n1275 GND 0.02fF $ **FLOATING
C4148 EESPFAL_s1_0/EESPFAL_XOR_v3_1/CLK GND 0.02fF $ **FLOATING
C4149 CLK1.n1276 GND 0.02fF $ **FLOATING
C4150 CLK1.n1277 GND 0.03fF $ **FLOATING
C4151 CLK1.n1278 GND 0.16fF $ **FLOATING
C4152 CLK1.n1279 GND 0.03fF $ **FLOATING
C4153 CLK1.n1280 GND 0.02fF $ **FLOATING
C4154 CLK1.t70 GND 0.05fF
C4155 CLK1.n1281 GND 0.29fF $ **FLOATING
C4156 CLK1.n1282 GND 0.02fF $ **FLOATING
C4157 CLK1.n1283 GND 0.03fF $ **FLOATING
C4158 CLK1.n1284 GND 0.06fF $ **FLOATING
C4159 CLK1.n1285 GND 0.03fF $ **FLOATING
C4160 CLK1.n1286 GND 0.02fF $ **FLOATING
C4161 CLK1.n1287 GND 0.03fF $ **FLOATING
C4162 CLK1.n1288 GND 0.02fF $ **FLOATING
C4163 CLK1.n1289 GND 0.03fF $ **FLOATING
C4164 CLK1.n1290 GND 0.06fF $ **FLOATING
C4165 CLK1.n1291 GND 0.03fF $ **FLOATING
C4166 CLK1.n1292 GND 0.02fF $ **FLOATING
C4167 CLK1.t32 GND 0.03fF
C4168 CLK1.t53 GND 0.03fF
C4169 CLK1.n1293 GND 0.15fF $ **FLOATING
C4170 CLK1.n1294 GND 0.03fF $ **FLOATING
C4171 CLK1.n1295 GND 0.02fF $ **FLOATING
C4172 CLK1.n1296 GND 0.03fF $ **FLOATING
C4173 CLK1.t115 GND 0.07fF
C4174 CLK1.n1297 GND 0.45fF $ **FLOATING
C4175 CLK1.n1298 GND 0.02fF $ **FLOATING
C4176 CLK1.n1299 GND 0.03fF $ **FLOATING
C4177 CLK1.n1300 GND 0.14fF $ **FLOATING
C4178 CLK1.n1301 GND 0.03fF $ **FLOATING
C4179 CLK1.n1302 GND 0.02fF $ **FLOATING
C4180 CLK1.t13 GND 0.05fF
C4181 CLK1.n1303 GND 0.29fF $ **FLOATING
C4182 CLK1.n1304 GND 0.02fF $ **FLOATING
C4183 CLK1.n1305 GND 0.03fF $ **FLOATING
C4184 CLK1.n1306 GND 0.09fF $ **FLOATING
C4185 CLK1.n1307 GND 0.03fF $ **FLOATING
C4186 CLK1.n1308 GND 0.02fF $ **FLOATING
C4187 CLK1.t176 GND 0.03fF
C4188 CLK1.t15 GND 0.03fF
C4189 CLK1.n1309 GND 0.10fF $ **FLOATING
C4190 CLK1.n1310 GND 0.03fF $ **FLOATING
C4191 CLK1.n1311 GND 0.02fF $ **FLOATING
C4192 CLK1.n1312 GND 0.03fF $ **FLOATING
C4193 CLK1.t173 GND 0.09fF
C4194 CLK1.n1313 GND 0.03fF $ **FLOATING
C4195 CLK1.n1314 GND 0.02fF $ **FLOATING
C4196 CLK1.t174 GND 0.05fF
C4197 CLK1.n1315 GND 0.03fF $ **FLOATING
C4198 CLK1.n1316 GND 0.02fF $ **FLOATING
C4199 CLK1.n1317 GND 0.03fF $ **FLOATING
C4200 CLK1.n1318 GND 0.07fF $ **FLOATING
C4201 CLK1.n1319 GND 0.03fF $ **FLOATING
C4202 CLK1.n1320 GND 0.02fF $ **FLOATING
C4203 CLK1.t147 GND 0.07fF
C4204 CLK1.n1321 GND 0.15fF $ **FLOATING
C4205 CLK1.n1322 GND 0.47fF $ **FLOATING
C4206 CLK1.n1323 GND 0.03fF $ **FLOATING
C4207 CLK1.n1324 GND 0.03fF $ **FLOATING
C4208 CLK1.n1325 GND 0.02fF $ **FLOATING
C4209 CLK1.n1326 GND 0.03fF $ **FLOATING
C4210 CLK1.n1327 GND 0.06fF $ **FLOATING
C4211 CLK1.n1328 GND 0.14fF $ **FLOATING
C4212 CLK1.n1329 GND 0.11fF $ **FLOATING
C4213 CLK1.n1330 GND 0.18fF $ **FLOATING
C4214 CLK1.n1331 GND 0.03fF $ **FLOATING
C4215 CLK1.n1332 GND 0.02fF $ **FLOATING
C4216 CLK1.n1333 GND 0.02fF $ **FLOATING
C4217 CLK1.n1334 GND 0.29fF $ **FLOATING
C4218 CLK1.n1335 GND 0.03fF $ **FLOATING
C4219 CLK1.n1336 GND 0.03fF $ **FLOATING
C4220 CLK1.n1337 GND 0.02fF $ **FLOATING
C4221 CLK1.n1338 GND 0.03fF $ **FLOATING
C4222 CLK1.n1339 GND 0.16fF $ **FLOATING
C4223 CLK1.n1340 GND 0.09fF $ **FLOATING
C4224 CLK1.t175 GND 0.09fF
C4225 CLK1.t14 GND 0.09fF
C4226 CLK1.n1341 GND 0.17fF $ **FLOATING
C4227 CLK1.n1342 GND 0.03fF $ **FLOATING
C4228 CLK1.n1343 GND 0.02fF $ **FLOATING
C4229 CLK1.n1344 GND 0.17fF $ **FLOATING
C4230 EESPFAL_s1_0/EESPFAL_INV4_1/CLK GND 0.02fF $ **FLOATING
C4231 CLK1.n1345 GND 0.03fF $ **FLOATING
C4232 CLK1.n1346 GND 0.03fF $ **FLOATING
C4233 CLK1.n1347 GND 0.03fF $ **FLOATING
C4234 CLK1.n1348 GND 0.02fF $ **FLOATING
C4235 CLK1.n1349 GND 0.03fF $ **FLOATING
C4236 CLK1.n1350 GND 0.16fF $ **FLOATING
C4237 CLK1.t12 GND 0.09fF
C4238 CLK1.n1351 GND 0.11fF $ **FLOATING
C4239 CLK1.n1352 GND 0.18fF $ **FLOATING
C4240 CLK1.n1353 GND 0.03fF $ **FLOATING
C4241 CLK1.n1354 GND 0.02fF $ **FLOATING
C4242 CLK1.n1355 GND 0.02fF $ **FLOATING
C4243 CLK1.n1356 GND 0.03fF $ **FLOATING
C4244 CLK1.n1357 GND 0.03fF $ **FLOATING
C4245 CLK1.n1358 GND 0.03fF $ **FLOATING
C4246 CLK1.n1359 GND 0.02fF $ **FLOATING
C4247 CLK1.n1360 GND 0.03fF $ **FLOATING
C4248 CLK1.n1361 GND 0.06fF $ **FLOATING
C4249 CLK1.n1362 GND 0.07fF $ **FLOATING
C4250 CLK1.n1363 GND 0.15fF $ **FLOATING
C4251 CLK1.n1364 GND 0.10fF $ **FLOATING
C4252 CLK1.n1365 GND 0.11fF $ **FLOATING
C4253 CLK1.n1366 GND 0.21fF $ **FLOATING
C4254 CLK1.n1367 GND 0.08fF $ **FLOATING
C4255 CLK1.n1368 GND 0.06fF $ **FLOATING
C4256 CLK1.n1369 GND 0.03fF $ **FLOATING
C4257 CLK1.n1370 GND 0.02fF $ **FLOATING
C4258 CLK1.n1371 GND 0.03fF $ **FLOATING
C4259 CLK1.n1372 GND 0.02fF $ **FLOATING
C4260 CLK1.n1373 GND 0.19fF $ **FLOATING
C4261 CLK1.n1374 GND 0.03fF $ **FLOATING
C4262 CLK1.n1375 GND 0.02fF $ **FLOATING
C4263 CLK1.n1376 GND 0.03fF $ **FLOATING
C4264 CLK1.n1377 GND 0.06fF $ **FLOATING
C4265 CLK1.n1378 GND 0.06fF $ **FLOATING
C4266 CLK1.n1379 GND 0.06fF $ **FLOATING
C4267 CLK1.n1380 GND 0.03fF $ **FLOATING
C4268 CLK1.n1381 GND 0.02fF $ **FLOATING
C4269 CLK1.n1382 GND 0.03fF $ **FLOATING
C4270 CLK1.n1383 GND 0.03fF $ **FLOATING
C4271 CLK1.n1384 GND 0.02fF $ **FLOATING
C4272 CLK1.n1385 GND 0.03fF $ **FLOATING
C4273 CLK1.n1386 GND 0.02fF $ **FLOATING
C4274 CLK1.n1387 GND 0.03fF $ **FLOATING
C4275 CLK1.n1388 GND 0.14fF $ **FLOATING
C4276 CLK1.n1389 GND 0.18fF $ **FLOATING
C4277 CLK1.t69 GND 0.09fF
C4278 CLK1.n1390 GND 0.11fF $ **FLOATING
C4279 CLK1.n1391 GND 0.03fF $ **FLOATING
C4280 CLK1.n1392 GND 0.02fF $ **FLOATING
C4281 CLK1.n1393 GND 0.03fF $ **FLOATING
C4282 CLK1.n1394 GND 0.03fF $ **FLOATING
C4283 CLK1.t30 GND 0.03fF
C4284 CLK1.t131 GND 0.03fF
C4285 CLK1.n1395 GND 0.10fF $ **FLOATING
C4286 CLK1.n1396 GND 0.17fF $ **FLOATING
C4287 CLK1.n1397 GND 0.03fF $ **FLOATING
C4288 CLK1.n1398 GND 0.02fF $ **FLOATING
C4289 CLK1.n1399 GND 0.03fF $ **FLOATING
C4290 CLK1.n1400 GND 0.09fF $ **FLOATING
C4291 CLK1.t29 GND 0.09fF
C4292 CLK1.n1401 GND 0.17fF $ **FLOATING
C4293 CLK1.t130 GND 0.09fF
C4294 CLK1.n1402 GND 0.16fF $ **FLOATING
C4295 CLK1.n1403 GND 0.09fF $ **FLOATING
C4296 CLK1.n1404 GND 0.03fF $ **FLOATING
C4297 CLK1.n1405 GND 0.02fF $ **FLOATING
C4298 CLK1.n1406 GND 0.03fF $ **FLOATING
C4299 CLK1.n1407 GND 0.03fF $ **FLOATING
C4300 CLK1.t133 GND 0.05fF
C4301 CLK1.n1408 GND 0.29fF $ **FLOATING
C4302 CLK1.n1409 GND 0.03fF $ **FLOATING
C4303 CLK1.n1410 GND 0.02fF $ **FLOATING
C4304 CLK1.n1411 GND 0.03fF $ **FLOATING
C4305 CLK1.n1412 GND 0.11fF $ **FLOATING
C4306 CLK1.n1413 GND 0.18fF $ **FLOATING
C4307 CLK1.n1414 GND 0.14fF $ **FLOATING
C4308 CLK1.n1415 GND 0.03fF $ **FLOATING
C4309 CLK1.n1416 GND 0.02fF $ **FLOATING
C4310 CLK1.n1417 GND 0.03fF $ **FLOATING
C4311 CLK1.n1418 GND 0.03fF $ **FLOATING
C4312 CLK1.n1419 GND 0.03fF $ **FLOATING
C4313 CLK1.n1420 GND 0.02fF $ **FLOATING
C4314 CLK1.n1421 GND 0.03fF $ **FLOATING
C4315 CLK1.n1422 GND 0.06fF $ **FLOATING
C4316 CLK1.n1423 GND 0.06fF $ **FLOATING
C4317 CLK1.n1424 GND 0.06fF $ **FLOATING
C4318 CLK1.n1425 GND 0.03fF $ **FLOATING
C4319 CLK1.n1426 GND 0.02fF $ **FLOATING
C4320 CLK1.n1427 GND 0.03fF $ **FLOATING
C4321 CLK1.n1428 GND 0.19fF $ **FLOATING
C4322 CLK1.n1429 GND 0.02fF $ **FLOATING
C4323 CLK1.n1430 GND 0.03fF $ **FLOATING
C4324 CLK1.n1431 GND 0.03fF $ **FLOATING
C4325 CLK1.n1432 GND 0.02fF $ **FLOATING
C4326 CLK1.n1433 GND 0.03fF $ **FLOATING
C4327 CLK1.n1434 GND 0.06fF $ **FLOATING
C4328 CLK1.n1435 GND 0.08fF $ **FLOATING
C4329 CLK1.n1436 GND 0.19fF $ **FLOATING
C4330 CLK1.n1437 GND 0.01fF $ **FLOATING
C4331 CLK1.n1438 GND 0.00fF $ **FLOATING
C4332 CLK1.n1439 GND 0.03fF $ **FLOATING
C4333 CLK1.n1440 GND 0.36fF $ **FLOATING
C4334 CLK1.n1441 GND 0.36fF $ **FLOATING
C4335 CLK1.n1442 GND 0.02fF $ **FLOATING
C4336 CLK1.n1443 GND 0.01fF $ **FLOATING
C4337 CLK1.n1444 GND 0.03fF $ **FLOATING
C4338 CLK1.n1445 GND 0.06fF $ **FLOATING
C4339 CLK1.n1446 GND 0.03fF $ **FLOATING
C4340 CLK1.n1447 GND 0.02fF $ **FLOATING
C4341 CLK1.n1448 GND 0.02fF $ **FLOATING
C4342 CLK1.t168 GND 0.03fF
C4343 CLK1.t67 GND 0.03fF
C4344 CLK1.n1449 GND 0.15fF $ **FLOATING
C4345 CLK1.n1450 GND 0.03fF $ **FLOATING
C4346 CLK1.n1451 GND 0.02fF $ **FLOATING
C4347 CLK1.n1452 GND 0.03fF $ **FLOATING
C4348 CLK1.n1453 GND 0.06fF $ **FLOATING
C4349 CLK1.n1454 GND 0.03fF $ **FLOATING
C4350 CLK1.n1455 GND 0.02fF $ **FLOATING
C4351 CLK1.n1456 GND 0.02fF $ **FLOATING
C4352 CLK1.n1457 GND 0.02fF $ **FLOATING
C4353 CLK1.n1458 GND 0.03fF $ **FLOATING
C4354 CLK1.t51 GND 0.09fF
C4355 CLK1.n1459 GND 0.03fF $ **FLOATING
C4356 CLK1.n1460 GND 0.02fF $ **FLOATING
C4357 EESPFAL_s1_0/EESPFAL_XOR_v3_0/CLK GND 0.02fF $ **FLOATING
C4358 CLK1.n1461 GND 0.02fF $ **FLOATING
C4359 CLK1.n1462 GND 0.03fF $ **FLOATING
C4360 CLK1.n1463 GND 0.16fF $ **FLOATING
C4361 CLK1.n1464 GND 0.03fF $ **FLOATING
C4362 CLK1.n1465 GND 0.02fF $ **FLOATING
C4363 CLK1.t178 GND 0.05fF
C4364 CLK1.n1466 GND 0.29fF $ **FLOATING
C4365 CLK1.n1467 GND 0.02fF $ **FLOATING
C4366 CLK1.n1468 GND 0.03fF $ **FLOATING
C4367 CLK1.n1469 GND 0.06fF $ **FLOATING
C4368 CLK1.n1470 GND 0.03fF $ **FLOATING
C4369 CLK1.n1471 GND 0.02fF $ **FLOATING
C4370 CLK1.n1472 GND 0.03fF $ **FLOATING
C4371 CLK1.n1473 GND 0.02fF $ **FLOATING
C4372 CLK1.n1474 GND 0.03fF $ **FLOATING
C4373 CLK1.n1475 GND 0.06fF $ **FLOATING
C4374 CLK1.n1476 GND 0.03fF $ **FLOATING
C4375 CLK1.n1477 GND 0.02fF $ **FLOATING
C4376 CLK1.t91 GND 0.03fF
C4377 CLK1.t23 GND 0.03fF
C4378 CLK1.n1478 GND 0.15fF $ **FLOATING
C4379 CLK1.n1479 GND 0.03fF $ **FLOATING
C4380 CLK1.n1480 GND 0.02fF $ **FLOATING
C4381 CLK1.n1481 GND 0.03fF $ **FLOATING
C4382 CLK1.t171 GND 0.07fF
C4383 CLK1.n1482 GND 0.45fF $ **FLOATING
C4384 CLK1.n1483 GND 0.02fF $ **FLOATING
C4385 CLK1.n1484 GND 0.03fF $ **FLOATING
C4386 CLK1.n1485 GND 0.14fF $ **FLOATING
C4387 CLK1.n1486 GND 0.03fF $ **FLOATING
C4388 CLK1.n1487 GND 0.02fF $ **FLOATING
C4389 CLK1.t3 GND 0.05fF
C4390 CLK1.n1488 GND 0.29fF $ **FLOATING
C4391 CLK1.n1489 GND 0.02fF $ **FLOATING
C4392 CLK1.n1490 GND 0.03fF $ **FLOATING
C4393 CLK1.n1491 GND 0.09fF $ **FLOATING
C4394 CLK1.n1492 GND 0.03fF $ **FLOATING
C4395 CLK1.n1493 GND 0.02fF $ **FLOATING
C4396 CLK1.t83 GND 0.03fF
C4397 CLK1.t1 GND 0.03fF
C4398 CLK1.n1494 GND 0.10fF $ **FLOATING
C4399 CLK1.n1495 GND 0.03fF $ **FLOATING
C4400 CLK1.n1496 GND 0.02fF $ **FLOATING
C4401 CLK1.n1497 GND 0.03fF $ **FLOATING
C4402 CLK1.t80 GND 0.09fF
C4403 CLK1.n1498 GND 0.03fF $ **FLOATING
C4404 CLK1.n1499 GND 0.02fF $ **FLOATING
C4405 CLK1.t81 GND 0.05fF
C4406 CLK1.n1500 GND 0.03fF $ **FLOATING
C4407 CLK1.n1501 GND 0.02fF $ **FLOATING
C4408 CLK1.n1502 GND 0.03fF $ **FLOATING
C4409 CLK1.n1503 GND 0.07fF $ **FLOATING
C4410 CLK1.n1504 GND 0.03fF $ **FLOATING
C4411 CLK1.n1505 GND 0.02fF $ **FLOATING
C4412 CLK1.t192 GND 0.07fF
C4413 CLK1.n1506 GND 0.15fF $ **FLOATING
C4414 CLK1.n1507 GND 0.47fF $ **FLOATING
C4415 CLK1.n1508 GND 0.03fF $ **FLOATING
C4416 CLK1.n1509 GND 0.03fF $ **FLOATING
C4417 CLK1.n1510 GND 0.02fF $ **FLOATING
C4418 CLK1.n1511 GND 0.03fF $ **FLOATING
C4419 CLK1.n1512 GND 0.06fF $ **FLOATING
C4420 CLK1.n1513 GND 0.14fF $ **FLOATING
C4421 CLK1.n1514 GND 0.11fF $ **FLOATING
C4422 CLK1.n1515 GND 0.18fF $ **FLOATING
C4423 CLK1.n1516 GND 0.03fF $ **FLOATING
C4424 CLK1.n1517 GND 0.02fF $ **FLOATING
C4425 CLK1.n1518 GND 0.02fF $ **FLOATING
C4426 CLK1.n1519 GND 0.29fF $ **FLOATING
C4427 CLK1.n1520 GND 0.03fF $ **FLOATING
C4428 CLK1.n1521 GND 0.03fF $ **FLOATING
C4429 CLK1.n1522 GND 0.02fF $ **FLOATING
C4430 CLK1.n1523 GND 0.03fF $ **FLOATING
C4431 CLK1.n1524 GND 0.16fF $ **FLOATING
C4432 CLK1.n1525 GND 0.09fF $ **FLOATING
C4433 CLK1.t82 GND 0.09fF
C4434 CLK1.t0 GND 0.09fF
C4435 CLK1.n1526 GND 0.17fF $ **FLOATING
C4436 CLK1.n1527 GND 0.03fF $ **FLOATING
C4437 CLK1.n1528 GND 0.02fF $ **FLOATING
C4438 CLK1.n1529 GND 0.17fF $ **FLOATING
C4439 EESPFAL_s1_0/EESPFAL_INV4_2/CLK GND 0.02fF $ **FLOATING
C4440 CLK1.n1530 GND 0.03fF $ **FLOATING
C4441 CLK1.n1531 GND 0.03fF $ **FLOATING
C4442 CLK1.n1532 GND 0.03fF $ **FLOATING
C4443 CLK1.n1533 GND 0.02fF $ **FLOATING
C4444 CLK1.n1534 GND 0.03fF $ **FLOATING
C4445 CLK1.n1535 GND 0.16fF $ **FLOATING
C4446 CLK1.t2 GND 0.09fF
C4447 CLK1.n1536 GND 0.11fF $ **FLOATING
C4448 CLK1.n1537 GND 0.18fF $ **FLOATING
C4449 CLK1.n1538 GND 0.03fF $ **FLOATING
C4450 CLK1.n1539 GND 0.02fF $ **FLOATING
C4451 CLK1.n1540 GND 0.02fF $ **FLOATING
C4452 CLK1.n1541 GND 0.03fF $ **FLOATING
C4453 CLK1.n1542 GND 0.03fF $ **FLOATING
C4454 CLK1.n1543 GND 0.03fF $ **FLOATING
C4455 CLK1.n1544 GND 0.02fF $ **FLOATING
C4456 CLK1.n1545 GND 0.03fF $ **FLOATING
C4457 CLK1.n1546 GND 0.06fF $ **FLOATING
C4458 CLK1.n1547 GND 0.07fF $ **FLOATING
C4459 CLK1.n1548 GND 0.15fF $ **FLOATING
C4460 CLK1.n1549 GND 0.10fF $ **FLOATING
C4461 CLK1.n1550 GND 0.11fF $ **FLOATING
C4462 CLK1.n1551 GND 0.21fF $ **FLOATING
C4463 CLK1.n1552 GND 0.08fF $ **FLOATING
C4464 CLK1.n1553 GND 0.06fF $ **FLOATING
C4465 CLK1.n1554 GND 0.03fF $ **FLOATING
C4466 CLK1.n1555 GND 0.02fF $ **FLOATING
C4467 CLK1.n1556 GND 0.03fF $ **FLOATING
C4468 CLK1.n1557 GND 0.02fF $ **FLOATING
C4469 CLK1.n1558 GND 0.19fF $ **FLOATING
C4470 CLK1.n1559 GND 0.03fF $ **FLOATING
C4471 CLK1.n1560 GND 0.02fF $ **FLOATING
C4472 CLK1.n1561 GND 0.03fF $ **FLOATING
C4473 CLK1.n1562 GND 0.06fF $ **FLOATING
C4474 CLK1.n1563 GND 0.06fF $ **FLOATING
C4475 CLK1.n1564 GND 0.06fF $ **FLOATING
C4476 CLK1.n1565 GND 0.03fF $ **FLOATING
C4477 CLK1.n1566 GND 0.02fF $ **FLOATING
C4478 CLK1.n1567 GND 0.03fF $ **FLOATING
C4479 CLK1.n1568 GND 0.03fF $ **FLOATING
C4480 CLK1.n1569 GND 0.02fF $ **FLOATING
C4481 CLK1.n1570 GND 0.03fF $ **FLOATING
C4482 CLK1.n1571 GND 0.02fF $ **FLOATING
C4483 CLK1.n1572 GND 0.03fF $ **FLOATING
C4484 CLK1.n1573 GND 0.14fF $ **FLOATING
C4485 CLK1.n1574 GND 0.18fF $ **FLOATING
C4486 CLK1.t177 GND 0.09fF
C4487 CLK1.n1575 GND 0.11fF $ **FLOATING
C4488 CLK1.n1576 GND 0.03fF $ **FLOATING
C4489 CLK1.n1577 GND 0.02fF $ **FLOATING
C4490 CLK1.n1578 GND 0.03fF $ **FLOATING
C4491 CLK1.n1579 GND 0.03fF $ **FLOATING
C4492 CLK1.t42 GND 0.03fF
C4493 CLK1.t151 GND 0.03fF
C4494 CLK1.n1580 GND 0.10fF $ **FLOATING
C4495 CLK1.n1581 GND 0.17fF $ **FLOATING
C4496 CLK1.n1582 GND 0.03fF $ **FLOATING
C4497 CLK1.n1583 GND 0.02fF $ **FLOATING
C4498 CLK1.n1584 GND 0.03fF $ **FLOATING
C4499 CLK1.n1585 GND 0.09fF $ **FLOATING
C4500 CLK1.t41 GND 0.09fF
C4501 CLK1.n1586 GND 0.17fF $ **FLOATING
C4502 CLK1.t150 GND 0.09fF
C4503 CLK1.n1587 GND 0.16fF $ **FLOATING
C4504 CLK1.n1588 GND 0.09fF $ **FLOATING
C4505 CLK1.n1589 GND 0.03fF $ **FLOATING
C4506 CLK1.n1590 GND 0.02fF $ **FLOATING
C4507 CLK1.n1591 GND 0.03fF $ **FLOATING
C4508 CLK1.n1592 GND 0.03fF $ **FLOATING
C4509 CLK1.t52 GND 0.05fF
C4510 CLK1.n1593 GND 0.29fF $ **FLOATING
C4511 CLK1.n1594 GND 0.03fF $ **FLOATING
C4512 CLK1.n1595 GND 0.02fF $ **FLOATING
C4513 CLK1.n1596 GND 0.03fF $ **FLOATING
C4514 CLK1.n1597 GND 0.11fF $ **FLOATING
C4515 CLK1.n1598 GND 0.18fF $ **FLOATING
C4516 CLK1.n1599 GND 0.14fF $ **FLOATING
C4517 CLK1.n1600 GND 0.03fF $ **FLOATING
C4518 CLK1.n1601 GND 0.02fF $ **FLOATING
C4519 CLK1.n1602 GND 0.03fF $ **FLOATING
C4520 CLK1.n1603 GND 0.03fF $ **FLOATING
C4521 CLK1.n1604 GND 0.03fF $ **FLOATING
C4522 CLK1.n1605 GND 0.02fF $ **FLOATING
C4523 CLK1.n1606 GND 0.03fF $ **FLOATING
C4524 CLK1.n1607 GND 0.06fF $ **FLOATING
C4525 CLK1.n1608 GND 0.06fF $ **FLOATING
C4526 CLK1.n1609 GND 0.06fF $ **FLOATING
C4527 CLK1.n1610 GND 0.03fF $ **FLOATING
C4528 CLK1.n1611 GND 0.02fF $ **FLOATING
C4529 CLK1.n1612 GND 0.03fF $ **FLOATING
C4530 CLK1.n1613 GND 0.19fF $ **FLOATING
C4531 CLK1.n1614 GND 0.02fF $ **FLOATING
C4532 CLK1.n1615 GND 0.03fF $ **FLOATING
C4533 CLK1.n1616 GND 0.03fF $ **FLOATING
C4534 CLK1.n1617 GND 0.02fF $ **FLOATING
C4535 CLK1.n1618 GND 0.03fF $ **FLOATING
C4536 CLK1.n1619 GND 0.06fF $ **FLOATING
C4537 CLK1.n1620 GND 0.08fF $ **FLOATING
C4538 CLK1.n1621 GND 0.19fF $ **FLOATING
C4539 CLK1.n1622 GND 0.01fF $ **FLOATING
C4540 CLK1.n1623 GND 0.00fF $ **FLOATING
C4541 CLK1.n1624 GND 0.03fF $ **FLOATING
C4542 CLK1.n1625 GND 0.07fF $ **FLOATING
C4543 CLK1.n1626 GND 0.43fF $ **FLOATING
C4544 EESPFAL_s0_0/CLK1 GND 0.03fF $ **FLOATING
C4545 x1.t6 GND 0.45fF
C4546 EESPFAL_s0_0/x1 GND 4.91fF $ **FLOATING
C4547 x1.t4 GND 0.19fF
C4548 EESPFAL_s0_0/EESPFAL_NAND_v3_2/B_bar GND 0.71fF $ **FLOATING
C4549 x1.n0 GND 2.61fF $ **FLOATING
C4550 x1.t8 GND 0.32fF
C4551 x1.t3 GND 0.28fF
C4552 x1.n1 GND 2.43fF $ **FLOATING
C4553 EESPFAL_s1_0/EESPFAL_XOR_v3_1/A GND 0.44fF $ **FLOATING
C4554 x1.t9 GND 0.53fF
C4555 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/B GND 2.19fF $ **FLOATING
C4556 x1.t10 GND 0.36fF
C4557 EESPFAL_s2_0/EESPFAL_4in_NAND_0/B GND 2.91fF $ **FLOATING
C4558 x1.t7 GND 0.32fF
C4559 x1.t1 GND 0.28fF
C4560 x1.n2 GND 2.43fF $ **FLOATING
C4561 EESPFAL_s2_0/EESPFAL_XOR_v3_1/A GND 0.45fF $ **FLOATING
C4562 x1.t2 GND 0.16fF
C4563 EESPFAL_s2_0/EESPFAL_INV4_1/A_bar GND 0.58fF $ **FLOATING
C4564 x1.t5 GND 0.32fF
C4565 x1.t11 GND 0.28fF
C4566 x1.n3 GND 2.43fF $ **FLOATING
C4567 EESPFAL_s3_0/EESPFAL_XOR_v3_0/A GND 0.44fF $ **FLOATING
C4568 x1.t0 GND 0.22fF
C4569 EESPFAL_s3_0/EESPFAL_INV4_1/A GND 1.85fF $ **FLOATING
C4570 EESPFAL_s3_0/x1 GND 10.41fF $ **FLOATING
C4571 x1.n4 GND 0.95fF $ **FLOATING
C4572 EESPFAL_s2_0/x1 GND 1.09fF $ **FLOATING
C4573 x1.n5 GND 5.98fF $ **FLOATING
C4574 x1.n6 GND 1.82fF $ **FLOATING
C4575 x1.n7 GND 2.49fF $ **FLOATING
C4576 x1.n8 GND 2.73fF $ **FLOATING
C4577 x1.n9 GND 2.52fF $ **FLOATING
C4578 EESPFAL_s1_0/x1 GND 2.46fF $ **FLOATING
C4579 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t6 GND 0.04fF
C4580 EESPFAL_s3_0/EESPFAL_3in_NOR_v2_0/A_bar GND 0.53fF $ **FLOATING
C4581 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t3 GND 0.04fF
C4582 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t0 GND 0.04fF
C4583 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n0 GND 0.11fF $ **FLOATING
C4584 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t2 GND 0.13fF
C4585 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t1 GND 0.20fF
C4586 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n1 GND 0.19fF $ **FLOATING
C4587 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n2 GND 0.09fF $ **FLOATING
C4588 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t5 GND 0.04fF
C4589 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t4 GND 0.04fF
C4590 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n3 GND 0.09fF $ **FLOATING
C4591 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n4 GND 0.10fF $ **FLOATING
C4592 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t9 GND 0.05fF
C4593 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t8 GND 0.04fF
C4594 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.t7 GND 0.03fF
C4595 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n5 GND 0.05fF $ **FLOATING
C4596 EESPFAL_s3_0/EESPFAL_NAND_v3_0/OUT_bar.n6 GND 0.04fF $ **FLOATING
C4597 Dis1.t23 GND 0.21fF
C4598 Dis1.t4 GND 0.14fF
C4599 Dis1.n0 GND 0.53fF $ **FLOATING
C4600 Dis1.t6 GND 0.14fF
C4601 Dis1.n1 GND 0.92fF $ **FLOATING
C4602 Dis1.t13 GND 0.14fF
C4603 Dis1.n2 GND 0.28fF $ **FLOATING
C4604 EESPFAL_s0_0/EESPFAL_XOR_v3_0/Dis GND 0.28fF $ **FLOATING
C4605 Dis1.t20 GND 0.21fF
C4606 Dis1.t8 GND 0.14fF
C4607 Dis1.n3 GND 0.53fF $ **FLOATING
C4608 EESPFAL_s1_0/EESPFAL_3in_NAND_v2_0/Dis GND 0.27fF $ **FLOATING
C4609 Dis1.t27 GND 0.21fF
C4610 Dis1.t33 GND 0.14fF
C4611 Dis1.n4 GND 0.53fF $ **FLOATING
C4612 EESPFAL_s3_0/EESPFAL_3in_NAND_v2_0/Dis GND 0.31fF $ **FLOATING
C4613 Dis1.t14 GND 0.21fF
C4614 Dis1.t29 GND 0.14fF
C4615 Dis1.n5 GND 0.53fF $ **FLOATING
C4616 EESPFAL_s3_0/EESPFAL_INV4_1/Dis GND 0.60fF $ **FLOATING
C4617 Dis1.t30 GND 0.14fF
C4618 Dis1.n6 GND 0.87fF $ **FLOATING
C4619 Dis1.t1 GND 0.14fF
C4620 Dis1.n7 GND 0.28fF $ **FLOATING
C4621 EESPFAL_s3_0/EESPFAL_XOR_v3_1/Dis GND 0.26fF $ **FLOATING
C4622 Dis1.n8 GND 2.57fF $ **FLOATING
C4623 Dis1.t10 GND 0.21fF
C4624 Dis1.t26 GND 0.14fF
C4625 Dis1.n9 GND 0.53fF $ **FLOATING
C4626 EESPFAL_s3_0/EESPFAL_INV4_2/Dis GND 0.60fF $ **FLOATING
C4627 Dis1.t7 GND 0.14fF
C4628 Dis1.n10 GND 0.87fF $ **FLOATING
C4629 Dis1.t28 GND 0.14fF
C4630 Dis1.n11 GND 0.28fF $ **FLOATING
C4631 EESPFAL_s3_0/EESPFAL_XOR_v3_0/Dis GND 0.26fF $ **FLOATING
C4632 Dis1.n12 GND 0.80fF $ **FLOATING
C4633 EESPFAL_s3_0/Dis1 GND 0.58fF $ **FLOATING
C4634 EESPFAL_s2_0/Dis1 GND 0.59fF $ **FLOATING
C4635 Dis1.t24 GND 0.21fF
C4636 Dis1.t35 GND 0.14fF
C4637 Dis1.n13 GND 0.53fF $ **FLOATING
C4638 EESPFAL_s2_0/EESPFAL_INV4_1/Dis GND 0.60fF $ **FLOATING
C4639 Dis1.t5 GND 0.14fF
C4640 Dis1.n14 GND 0.88fF $ **FLOATING
C4641 Dis1.t21 GND 0.14fF
C4642 Dis1.n15 GND 0.28fF $ **FLOATING
C4643 EESPFAL_s2_0/EESPFAL_XOR_v3_0/Dis GND 0.17fF $ **FLOATING
C4644 Dis1.n16 GND 0.54fF $ **FLOATING
C4645 Dis1.t11 GND 0.21fF
C4646 Dis1.t18 GND 0.14fF
C4647 Dis1.n17 GND 0.53fF $ **FLOATING
C4648 EESPFAL_s2_0/EESPFAL_INV4_0/Dis GND 0.60fF $ **FLOATING
C4649 Dis1.t25 GND 0.14fF
C4650 Dis1.n18 GND 0.88fF $ **FLOATING
C4651 Dis1.t2 GND 0.14fF
C4652 Dis1.n19 GND 0.28fF $ **FLOATING
C4653 EESPFAL_s2_0/EESPFAL_XOR_v3_1/Dis GND 0.17fF $ **FLOATING
C4654 Dis1.n20 GND 1.16fF $ **FLOATING
C4655 Dis1.t34 GND 0.21fF
C4656 Dis1.t12 GND 0.14fF
C4657 Dis1.n21 GND 0.53fF $ **FLOATING
C4658 EESPFAL_s2_0/EESPFAL_4in_NAND_0/Dis GND 0.32fF $ **FLOATING
C4659 Dis1.n22 GND 1.64fF $ **FLOATING
C4660 Dis1.n23 GND 1.46fF $ **FLOATING
C4661 Dis1.t16 GND 0.21fF
C4662 Dis1.t0 GND 0.14fF
C4663 Dis1.n24 GND 0.53fF $ **FLOATING
C4664 EESPFAL_s1_0/EESPFAL_INV4_1/Dis GND 0.60fF $ **FLOATING
C4665 Dis1.t15 GND 0.14fF
C4666 Dis1.n25 GND 0.87fF $ **FLOATING
C4667 Dis1.t3 GND 0.14fF
C4668 Dis1.n26 GND 0.28fF $ **FLOATING
C4669 EESPFAL_s1_0/EESPFAL_XOR_v3_1/Dis GND 0.26fF $ **FLOATING
C4670 Dis1.n27 GND 1.28fF $ **FLOATING
C4671 Dis1.t32 GND 0.21fF
C4672 Dis1.t19 GND 0.14fF
C4673 Dis1.n28 GND 0.53fF $ **FLOATING
C4674 EESPFAL_s1_0/EESPFAL_INV4_2/Dis GND 0.60fF $ **FLOATING
C4675 Dis1.t31 GND 0.14fF
C4676 Dis1.n29 GND 0.87fF $ **FLOATING
C4677 Dis1.t22 GND 0.14fF
C4678 Dis1.n30 GND 0.28fF $ **FLOATING
C4679 EESPFAL_s1_0/EESPFAL_XOR_v3_0/Dis GND 0.26fF $ **FLOATING
C4680 Dis1.n31 GND 0.80fF $ **FLOATING
C4681 EESPFAL_s1_0/Dis1 GND 0.84fF $ **FLOATING
C4682 Dis1.t17 GND 0.21fF
C4683 Dis1.t9 GND 0.14fF
C4684 Dis1.n32 GND 0.53fF $ **FLOATING
C4685 EESPFAL_s0_0/EESPFAL_NAND_v3_2/Dis GND 0.28fF $ **FLOATING
C4686 Dis1.n33 GND 1.07fF $ **FLOATING
C4687 Dis1.n34 GND 0.82fF $ **FLOATING
C4688 EESPFAL_s0_0/Dis1 GND 0.05fF $ **FLOATING
C4689 CLK2.t29 GND 0.04fF
C4690 CLK2.t73 GND 0.03fF
C4691 CLK2.t27 GND 0.03fF
C4692 CLK2.n0 GND 0.08fF $ **FLOATING
C4693 CLK2.t71 GND 0.04fF
C4694 CLK2.t9 GND 0.06fF
C4695 CLK2.n1 GND 0.09fF $ **FLOATING
C4696 CLK2.n2 GND 0.26fF $ **FLOATING
C4697 CLK2.n3 GND 0.05fF $ **FLOATING
C4698 CLK2.n4 GND 0.02fF $ **FLOATING
C4699 CLK2.n5 GND 0.02fF $ **FLOATING
C4700 CLK2.n6 GND 0.02fF $ **FLOATING
C4701 CLK2.n7 GND 0.04fF $ **FLOATING
C4702 CLK2.n8 GND 0.02fF $ **FLOATING
C4703 CLK2.n9 GND 0.02fF $ **FLOATING
C4704 CLK2.n10 GND 0.02fF $ **FLOATING
C4705 CLK2.n11 GND 0.04fF $ **FLOATING
C4706 CLK2.n12 GND 0.02fF $ **FLOATING
C4707 CLK2.n13 GND 0.02fF $ **FLOATING
C4708 CLK2.n14 GND 0.02fF $ **FLOATING
C4709 CLK2.n15 GND 0.04fF $ **FLOATING
C4710 CLK2.n16 GND 0.02fF $ **FLOATING
C4711 CLK2.n17 GND 0.02fF $ **FLOATING
C4712 CLK2.n18 GND 0.02fF $ **FLOATING
C4713 CLK2.n19 GND 0.10fF $ **FLOATING
C4714 CLK2.n20 GND 0.02fF $ **FLOATING
C4715 CLK2.n21 GND 0.02fF $ **FLOATING
C4716 CLK2.n22 GND 0.02fF $ **FLOATING
C4717 CLK2.n23 GND 0.13fF $ **FLOATING
C4718 CLK2.n24 GND 0.02fF $ **FLOATING
C4719 CLK2.n25 GND 0.02fF $ **FLOATING
C4720 CLK2.n26 GND 0.01fF $ **FLOATING
C4721 CLK2.n27 GND 0.21fF $ **FLOATING
C4722 CLK2.t70 GND 0.06fF
C4723 CLK2.n28 GND 0.08fF $ **FLOATING
C4724 CLK2.n29 GND 0.02fF $ **FLOATING
C4725 CLK2.n30 GND 0.02fF $ **FLOATING
C4726 CLK2.n31 GND 0.02fF $ **FLOATING
C4727 CLK2.n32 GND 0.12fF $ **FLOATING
C4728 CLK2.n33 GND 0.02fF $ **FLOATING
C4729 CLK2.n34 GND 0.02fF $ **FLOATING
C4730 CLK2.n35 GND 0.02fF $ **FLOATING
C4731 CLK2.t72 GND 0.06fF
C4732 CLK2.n36 GND 0.07fF $ **FLOATING
C4733 CLK2.n37 GND 0.02fF $ **FLOATING
C4734 CLK2.n38 GND 0.02fF $ **FLOATING
C4735 CLK2.n39 GND 0.02fF $ **FLOATING
C4736 CLK2.n40 GND 0.13fF $ **FLOATING
C4737 CLK2.n41 GND 0.12fF $ **FLOATING
C4738 CLK2.n42 GND 0.02fF $ **FLOATING
C4739 CLK2.n43 GND 0.02fF $ **FLOATING
C4740 CLK2.t26 GND 0.06fF
C4741 CLK2.n44 GND 0.07fF $ **FLOATING
C4742 CLK2.n45 GND 0.02fF $ **FLOATING
C4743 CLK2.n46 GND 0.02fF $ **FLOATING
C4744 CLK2.n47 GND 0.02fF $ **FLOATING
C4745 CLK2.n48 GND 0.12fF $ **FLOATING
C4746 CLK2.n49 GND 0.02fF $ **FLOATING
C4747 CLK2.n50 GND 0.02fF $ **FLOATING
C4748 CLK2.n51 GND 0.02fF $ **FLOATING
C4749 CLK2.t28 GND 0.06fF
C4750 CLK2.n52 GND 0.08fF $ **FLOATING
C4751 CLK2.n53 GND 0.02fF $ **FLOATING
C4752 CLK2.n54 GND 0.02fF $ **FLOATING
C4753 CLK2.n55 GND 0.02fF $ **FLOATING
C4754 CLK2.n56 GND 0.21fF $ **FLOATING
C4755 CLK2.n57 GND 0.13fF $ **FLOATING
C4756 CLK2.n58 GND 0.02fF $ **FLOATING
C4757 CLK2.n59 GND 0.02fF $ **FLOATING
C4758 CLK2.n60 GND 0.01fF $ **FLOATING
C4759 CLK2.n61 GND 0.10fF $ **FLOATING
C4760 CLK2.n62 GND 0.02fF $ **FLOATING
C4761 CLK2.n63 GND 0.02fF $ **FLOATING
C4762 CLK2.n64 GND 0.02fF $ **FLOATING
C4763 CLK2.n65 GND 0.04fF $ **FLOATING
C4764 CLK2.n66 GND 0.02fF $ **FLOATING
C4765 CLK2.n67 GND 0.02fF $ **FLOATING
C4766 CLK2.n68 GND 0.02fF $ **FLOATING
C4767 CLK2.n69 GND 0.04fF $ **FLOATING
C4768 CLK2.n70 GND 0.02fF $ **FLOATING
C4769 CLK2.n71 GND 0.02fF $ **FLOATING
C4770 CLK2.n72 GND 0.02fF $ **FLOATING
C4771 CLK2.n73 GND 0.01fF $ **FLOATING
C4772 CLK2.n74 GND 0.02fF $ **FLOATING
C4773 CLK2.n75 GND 0.04fF $ **FLOATING
C4774 CLK2.n76 GND 0.02fF $ **FLOATING
C4775 CLK2.n77 GND 0.01fF $ **FLOATING
C4776 CLK2.n78 GND 0.05fF $ **FLOATING
C4777 CLK2.n79 GND 0.02fF $ **FLOATING
C4778 CLK2.t45 GND 0.03fF
C4779 CLK2.t22 GND 0.03fF
C4780 CLK2.n80 GND 0.11fF $ **FLOATING
C4781 CLK2.t5 GND 0.04fF
C4782 EESPFAL_s1_0/EESPFAL_NAND_v3_0/CLK GND 0.01fF $ **FLOATING
C4783 CLK2.n81 GND 0.12fF $ **FLOATING
C4784 CLK2.n82 GND 0.02fF $ **FLOATING
C4785 CLK2.t112 GND 0.03fF
C4786 CLK2.t7 GND 0.03fF
C4787 CLK2.n83 GND 0.08fF $ **FLOATING
C4788 CLK2.t42 GND 0.04fF
C4789 CLK2.t89 GND 0.03fF
C4790 CLK2.n84 GND 0.08fF $ **FLOATING
C4791 CLK2.n85 GND 0.01fF $ **FLOATING
C4792 CLK2.n86 GND 0.02fF $ **FLOATING
C4793 CLK2.n87 GND 0.02fF $ **FLOATING
C4794 CLK2.n88 GND 0.09fF $ **FLOATING
C4795 CLK2.t93 GND 0.04fF
C4796 CLK2.t95 GND 0.03fF
C4797 CLK2.t34 GND 0.03fF
C4798 CLK2.n89 GND 0.08fF $ **FLOATING
C4799 EESPFAL_s1_0/EESPFAL_NAND_v3_1/CLK GND 0.01fF $ **FLOATING
C4800 CLK2.t32 GND 0.04fF
C4801 CLK2.t115 GND 0.03fF
C4802 CLK2.t8 GND 0.03fF
C4803 CLK2.n90 GND 0.11fF $ **FLOATING
C4804 CLK2.n91 GND 0.09fF $ **FLOATING
C4805 CLK2.n92 GND 0.11fF $ **FLOATING
C4806 CLK2.t58 GND 0.03fF
C4807 CLK2.n93 GND 0.08fF $ **FLOATING
C4808 CLK2.n94 GND 0.01fF $ **FLOATING
C4809 CLK2.n95 GND 0.02fF $ **FLOATING
C4810 CLK2.t43 GND 0.03fF
C4811 CLK2.n96 GND 0.08fF $ **FLOATING
C4812 CLK2.n97 GND 0.01fF $ **FLOATING
C4813 CLK2.n98 GND 0.02fF $ **FLOATING
C4814 CLK2.n99 GND 0.11fF $ **FLOATING
C4815 CLK2.t23 GND 0.03fF
C4816 CLK2.t69 GND 0.03fF
C4817 CLK2.n100 GND 0.11fF $ **FLOATING
C4818 CLK2.t102 GND 0.04fF
C4819 EESPFAL_s2_0/EESPFAL_NAND_v3_0/CLK GND 0.01fF $ **FLOATING
C4820 CLK2.t36 GND 0.03fF
C4821 CLK2.t104 GND 0.03fF
C4822 CLK2.n101 GND 0.08fF $ **FLOATING
C4823 CLK2.t38 GND 0.04fF
C4824 CLK2.n102 GND 0.02fF $ **FLOATING
C4825 CLK2.n103 GND 0.02fF $ **FLOATING
C4826 CLK2.n104 GND 0.09fF $ **FLOATING
C4827 CLK2.t83 GND 0.04fF
C4828 CLK2.t57 GND 0.03fF
C4829 CLK2.t1 GND 0.03fF
C4830 CLK2.n105 GND 0.08fF $ **FLOATING
C4831 EESPFAL_s2_0/EESPFAL_NAND_v3_1/CLK GND 0.01fF $ **FLOATING
C4832 CLK2.t3 GND 0.04fF
C4833 CLK2.n106 GND 0.04fF $ **FLOATING
C4834 CLK2.n107 GND 0.02fF $ **FLOATING
C4835 CLK2.n108 GND 0.02fF $ **FLOATING
C4836 CLK2.n109 GND 0.01fF $ **FLOATING
C4837 CLK2.n110 GND 0.00fF $ **FLOATING
C4838 CLK2.n111 GND 0.01fF $ **FLOATING
C4839 CLK2.n112 GND 0.00fF $ **FLOATING
C4840 CLK2.n113 GND 0.00fF $ **FLOATING
C4841 CLK2.n114 GND 0.02fF $ **FLOATING
C4842 CLK2.n115 GND 0.02fF $ **FLOATING
C4843 CLK2.t90 GND 0.03fF
C4844 CLK2.t20 GND 0.03fF
C4845 CLK2.n116 GND 0.11fF $ **FLOATING
C4846 CLK2.n117 GND 0.05fF $ **FLOATING
C4847 CLK2.n118 GND 0.10fF $ **FLOATING
C4848 CLK2.n119 GND 0.02fF $ **FLOATING
C4849 CLK2.n120 GND 0.02fF $ **FLOATING
C4850 CLK2.n121 GND 0.01fF $ **FLOATING
C4851 CLK2.t108 GND 0.04fF
C4852 CLK2.n122 GND 0.02fF $ **FLOATING
C4853 CLK2.n123 GND 0.02fF $ **FLOATING
C4854 CLK2.n124 GND 0.02fF $ **FLOATING
C4855 CLK2.t109 GND 0.06fF
C4856 CLK2.n125 GND 0.02fF $ **FLOATING
C4857 CLK2.n126 GND 0.02fF $ **FLOATING
C4858 CLK2.t47 GND 0.03fF
C4859 CLK2.t110 GND 0.03fF
C4860 CLK2.n127 GND 0.08fF $ **FLOATING
C4861 CLK2.n128 GND 0.02fF $ **FLOATING
C4862 CLK2.n129 GND 0.02fF $ **FLOATING
C4863 CLK2.n130 GND 0.02fF $ **FLOATING
C4864 CLK2.n131 GND 0.13fF $ **FLOATING
C4865 CLK2.n132 GND 0.02fF $ **FLOATING
C4866 CLK2.n133 GND 0.02fF $ **FLOATING
C4867 CLK2.t55 GND 0.04fF
C4868 CLK2.n134 GND 0.02fF $ **FLOATING
C4869 CLK2.n135 GND 0.02fF $ **FLOATING
C4870 CLK2.n136 GND 0.02fF $ **FLOATING
C4871 CLK2.n137 GND 0.04fF $ **FLOATING
C4872 CLK2.n138 GND 0.02fF $ **FLOATING
C4873 CLK2.n139 GND 0.02fF $ **FLOATING
C4874 CLK2.n140 GND 0.01fF $ **FLOATING
C4875 CLK2.n141 GND 0.01fF $ **FLOATING
C4876 CLK2.n142 GND 0.02fF $ **FLOATING
C4877 CLK2.n143 GND 0.02fF $ **FLOATING
C4878 CLK2.t91 GND 0.03fF
C4879 CLK2.n144 GND 0.09fF $ **FLOATING
C4880 CLK2.n145 GND 0.02fF $ **FLOATING
C4881 CLK2.n146 GND 0.02fF $ **FLOATING
C4882 CLK2.n147 GND 0.02fF $ **FLOATING
C4883 CLK2.n148 GND 0.04fF $ **FLOATING
C4884 CLK2.n149 GND 0.02fF $ **FLOATING
C4885 CLK2.n150 GND 0.02fF $ **FLOATING
C4886 CLK2.n151 GND 0.01fF $ **FLOATING
C4887 CLK2.n152 GND 0.02fF $ **FLOATING
C4888 CLK2.n153 GND 0.02fF $ **FLOATING
C4889 CLK2.t86 GND 0.06fF
C4890 CLK2.n154 GND 0.02fF $ **FLOATING
C4891 CLK2.n155 GND 0.02fF $ **FLOATING
C4892 CLK2.t87 GND 0.04fF
C4893 CLK2.n156 GND 0.21fF $ **FLOATING
C4894 CLK2.t85 GND 0.03fF
C4895 CLK2.t18 GND 0.03fF
C4896 CLK2.n157 GND 0.08fF $ **FLOATING
C4897 CLK2.n158 GND 0.13fF $ **FLOATING
C4898 CLK2.n159 GND 0.02fF $ **FLOATING
C4899 CLK2.n160 GND 0.02fF $ **FLOATING
C4900 CLK2.n161 GND 0.12fF $ **FLOATING
C4901 CLK2.n162 GND 0.12fF $ **FLOATING
C4902 CLK2.n163 GND 0.02fF $ **FLOATING
C4903 CLK2.n164 GND 0.02fF $ **FLOATING
C4904 EESPFAL_s3_0/EESPFAL_NAND_v3_1/CLK GND 0.01fF $ **FLOATING
C4905 CLK2.t16 GND 0.04fF
C4906 CLK2.n165 GND 0.21fF $ **FLOATING
C4907 CLK2.n166 GND 0.02fF $ **FLOATING
C4908 CLK2.n167 GND 0.02fF $ **FLOATING
C4909 CLK2.t15 GND 0.06fF
C4910 CLK2.n168 GND 0.04fF $ **FLOATING
C4911 CLK2.n169 GND 0.02fF $ **FLOATING
C4912 CLK2.n170 GND 0.02fF $ **FLOATING
C4913 CLK2.n171 GND 0.01fF $ **FLOATING
C4914 CLK2.t10 GND 0.03fF
C4915 CLK2.t21 GND 0.03fF
C4916 CLK2.n172 GND 0.11fF $ **FLOATING
C4917 CLK2.n173 GND 0.14fF $ **FLOATING
C4918 CLK2.n174 GND 0.02fF $ **FLOATING
C4919 CLK2.n175 GND 0.02fF $ **FLOATING
C4920 CLK2.n176 GND 0.09fF $ **FLOATING
C4921 CLK2.n177 GND 0.01fF $ **FLOATING
C4922 CLK2.n178 GND 0.11fF $ **FLOATING
C4923 CLK2.t78 GND 0.05fF
C4924 CLK2.n179 GND 0.02fF $ **FLOATING
C4925 CLK2.n180 GND 0.02fF $ **FLOATING
C4926 CLK2.n181 GND 0.02fF $ **FLOATING
C4927 CLK2.n182 GND 0.13fF $ **FLOATING
C4928 CLK2.n183 GND 0.02fF $ **FLOATING
C4929 CLK2.n184 GND 0.02fF $ **FLOATING
C4930 CLK2.t62 GND 0.04fF
C4931 CLK2.n185 GND 0.02fF $ **FLOATING
C4932 CLK2.n186 GND 0.02fF $ **FLOATING
C4933 CLK2.n187 GND 0.02fF $ **FLOATING
C4934 CLK2.t116 GND 0.06fF
C4935 CLK2.n188 GND 0.02fF $ **FLOATING
C4936 CLK2.n189 GND 0.02fF $ **FLOATING
C4937 CLK2.t117 GND 0.03fF
C4938 CLK2.t68 GND 0.03fF
C4939 CLK2.n190 GND 0.08fF $ **FLOATING
C4940 CLK2.n191 GND 0.02fF $ **FLOATING
C4941 CLK2.n192 GND 0.02fF $ **FLOATING
C4942 CLK2.n193 GND 0.02fF $ **FLOATING
C4943 CLK2.n194 GND 0.12fF $ **FLOATING
C4944 CLK2.t67 GND 0.06fF
C4945 CLK2.n195 GND 0.13fF $ **FLOATING
C4946 CLK2.n196 GND 0.02fF $ **FLOATING
C4947 CLK2.n197 GND 0.02fF $ **FLOATING
C4948 CLK2.t14 GND 0.04fF
C4949 CLK2.n198 GND 0.02fF $ **FLOATING
C4950 CLK2.n199 GND 0.02fF $ **FLOATING
C4951 CLK2.n200 GND 0.02fF $ **FLOATING
C4952 CLK2.n201 GND 0.11fF $ **FLOATING
C4953 CLK2.t79 GND 0.05fF
C4954 CLK2.n202 GND 0.34fF $ **FLOATING
C4955 CLK2.n203 GND 0.02fF $ **FLOATING
C4956 CLK2.n204 GND 0.02fF $ **FLOATING
C4957 CLK2.n205 GND 0.02fF $ **FLOATING
C4958 CLK2.n206 GND 0.05fF $ **FLOATING
C4959 CLK2.n207 GND 0.04fF $ **FLOATING
C4960 CLK2.n208 GND 0.10fF $ **FLOATING
C4961 CLK2.n209 GND 0.02fF $ **FLOATING
C4962 CLK2.n210 GND 0.02fF $ **FLOATING
C4963 CLK2.n211 GND 0.02fF $ **FLOATING
C4964 CLK2.n212 GND 0.01fF $ **FLOATING
C4965 CLK2.n213 GND 0.21fF $ **FLOATING
C4966 CLK2.n214 GND 0.02fF $ **FLOATING
C4967 CLK2.n215 GND 0.02fF $ **FLOATING
C4968 CLK2.n216 GND 0.02fF $ **FLOATING
C4969 CLK2.n217 GND 0.08fF $ **FLOATING
C4970 CLK2.t13 GND 0.06fF
C4971 CLK2.n218 GND 0.12fF $ **FLOATING
C4972 CLK2.n219 GND 0.07fF $ **FLOATING
C4973 CLK2.n220 GND 0.02fF $ **FLOATING
C4974 CLK2.n221 GND 0.02fF $ **FLOATING
C4975 CLK2.n222 GND 0.02fF $ **FLOATING
C4976 EESPFAL_s3_0/EESPFAL_INV4_0/CLK GND 0.01fF $ **FLOATING
C4977 CLK2.n223 GND 0.13fF $ **FLOATING
C4978 CLK2.n224 GND 0.02fF $ **FLOATING
C4979 CLK2.n225 GND 0.02fF $ **FLOATING
C4980 CLK2.n226 GND 0.02fF $ **FLOATING
C4981 CLK2.n227 GND 0.07fF $ **FLOATING
C4982 CLK2.n228 GND 0.12fF $ **FLOATING
C4983 CLK2.t61 GND 0.06fF
C4984 CLK2.n229 GND 0.08fF $ **FLOATING
C4985 CLK2.n230 GND 0.02fF $ **FLOATING
C4986 CLK2.n231 GND 0.02fF $ **FLOATING
C4987 CLK2.n232 GND 0.02fF $ **FLOATING
C4988 CLK2.n233 GND 0.21fF $ **FLOATING
C4989 CLK2.n234 GND 0.01fF $ **FLOATING
C4990 CLK2.n235 GND 0.02fF $ **FLOATING
C4991 CLK2.n236 GND 0.02fF $ **FLOATING
C4992 CLK2.n237 GND 0.02fF $ **FLOATING
C4993 CLK2.n238 GND 0.10fF $ **FLOATING
C4994 CLK2.n239 GND 0.04fF $ **FLOATING
C4995 CLK2.n240 GND 0.05fF $ **FLOATING
C4996 CLK2.n241 GND 0.02fF $ **FLOATING
C4997 CLK2.n242 GND 0.02fF $ **FLOATING
C4998 CLK2.n243 GND 0.02fF $ **FLOATING
C4999 CLK2.n244 GND 0.32fF $ **FLOATING
C5000 CLK2.n245 GND 0.15fF $ **FLOATING
C5001 CLK2.n246 GND 0.15fF $ **FLOATING
C5002 CLK2.n247 GND 0.02fF $ **FLOATING
C5003 CLK2.n248 GND 0.02fF $ **FLOATING
C5004 CLK2.n249 GND 0.02fF $ **FLOATING
C5005 CLK2.n250 GND 0.05fF $ **FLOATING
C5006 CLK2.n251 GND 0.04fF $ **FLOATING
C5007 CLK2.n252 GND 0.04fF $ **FLOATING
C5008 CLK2.n253 GND 0.02fF $ **FLOATING
C5009 CLK2.n254 GND 0.02fF $ **FLOATING
C5010 CLK2.n255 GND 0.02fF $ **FLOATING
C5011 CLK2.n256 GND 0.02fF $ **FLOATING
C5012 CLK2.n257 GND 0.02fF $ **FLOATING
C5013 CLK2.n258 GND 0.02fF $ **FLOATING
C5014 CLK2.n259 GND 0.02fF $ **FLOATING
C5015 CLK2.n260 GND 0.10fF $ **FLOATING
C5016 CLK2.n261 GND 0.13fF $ **FLOATING
C5017 CLK2.n262 GND 0.08fF $ **FLOATING
C5018 CLK2.n263 GND 0.02fF $ **FLOATING
C5019 CLK2.n264 GND 0.02fF $ **FLOATING
C5020 CLK2.n265 GND 0.02fF $ **FLOATING
C5021 CLK2.n266 GND 0.02fF $ **FLOATING
C5022 CLK2.n267 GND 0.02fF $ **FLOATING
C5023 CLK2.n268 GND 0.02fF $ **FLOATING
C5024 CLK2.n269 GND 0.02fF $ **FLOATING
C5025 CLK2.n270 GND 0.07fF $ **FLOATING
C5026 CLK2.t17 GND 0.06fF
C5027 CLK2.n271 GND 0.12fF $ **FLOATING
C5028 CLK2.t84 GND 0.06fF
C5029 CLK2.n272 GND 0.07fF $ **FLOATING
C5030 CLK2.n273 GND 0.02fF $ **FLOATING
C5031 CLK2.n274 GND 0.02fF $ **FLOATING
C5032 CLK2.n275 GND 0.02fF $ **FLOATING
C5033 CLK2.n276 GND 0.02fF $ **FLOATING
C5034 CLK2.n277 GND 0.02fF $ **FLOATING
C5035 CLK2.n278 GND 0.02fF $ **FLOATING
C5036 CLK2.n279 GND 0.02fF $ **FLOATING
C5037 CLK2.n280 GND 0.08fF $ **FLOATING
C5038 CLK2.n281 GND 0.13fF $ **FLOATING
C5039 CLK2.n282 GND 0.10fF $ **FLOATING
C5040 CLK2.n283 GND 0.02fF $ **FLOATING
C5041 CLK2.n284 GND 0.02fF $ **FLOATING
C5042 CLK2.n285 GND 0.02fF $ **FLOATING
C5043 CLK2.n286 GND 0.02fF $ **FLOATING
C5044 CLK2.n287 GND 0.02fF $ **FLOATING
C5045 CLK2.n288 GND 0.02fF $ **FLOATING
C5046 CLK2.n289 GND 0.02fF $ **FLOATING
C5047 CLK2.n290 GND 0.04fF $ **FLOATING
C5048 CLK2.n291 GND 0.04fF $ **FLOATING
C5049 CLK2.n292 GND 0.05fF $ **FLOATING
C5050 CLK2.n293 GND 0.02fF $ **FLOATING
C5051 CLK2.n294 GND 0.02fF $ **FLOATING
C5052 CLK2.n295 GND 0.02fF $ **FLOATING
C5053 CLK2.n296 GND 0.06fF $ **FLOATING
C5054 CLK2.n297 GND 0.06fF $ **FLOATING
C5055 CLK2.n298 GND 0.02fF $ **FLOATING
C5056 CLK2.n299 GND 0.08fF $ **FLOATING
C5057 CLK2.n300 GND 0.01fF $ **FLOATING
C5058 CLK2.n301 GND 0.09fF $ **FLOATING
C5059 CLK2.n302 GND 0.08fF $ **FLOATING
C5060 CLK2.t44 GND 0.03fF
C5061 CLK2.n303 GND 0.08fF $ **FLOATING
C5062 CLK2.n304 GND 0.02fF $ **FLOATING
C5063 CLK2.n305 GND 0.02fF $ **FLOATING
C5064 CLK2.n306 GND 0.02fF $ **FLOATING
C5065 CLK2.n307 GND 0.07fF $ **FLOATING
C5066 CLK2.n308 GND 0.04fF $ **FLOATING
C5067 EESPFAL_s3_0/CLK2 GND 0.02fF $ **FLOATING
C5068 CLK2.n309 GND 0.01fF $ **FLOATING
C5069 CLK2.n310 GND 0.09fF $ **FLOATING
C5070 CLK2.n311 GND 0.05fF $ **FLOATING
C5071 CLK2.n312 GND 0.02fF $ **FLOATING
C5072 CLK2.n313 GND 0.02fF $ **FLOATING
C5073 CLK2.n314 GND 0.02fF $ **FLOATING
C5074 CLK2.n315 GND 0.02fF $ **FLOATING
C5075 CLK2.n316 GND 0.02fF $ **FLOATING
C5076 CLK2.n317 GND 0.02fF $ **FLOATING
C5077 CLK2.n318 GND 0.02fF $ **FLOATING
C5078 CLK2.n319 GND 0.04fF $ **FLOATING
C5079 CLK2.n320 GND 0.04fF $ **FLOATING
C5080 CLK2.n321 GND 0.10fF $ **FLOATING
C5081 CLK2.n322 GND 0.02fF $ **FLOATING
C5082 CLK2.n323 GND 0.02fF $ **FLOATING
C5083 CLK2.n324 GND 0.02fF $ **FLOATING
C5084 CLK2.n325 GND 0.01fF $ **FLOATING
C5085 CLK2.n326 GND 0.21fF $ **FLOATING
C5086 CLK2.n327 GND 0.02fF $ **FLOATING
C5087 CLK2.n328 GND 0.02fF $ **FLOATING
C5088 CLK2.n329 GND 0.02fF $ **FLOATING
C5089 CLK2.n330 GND 0.08fF $ **FLOATING
C5090 CLK2.t54 GND 0.06fF
C5091 CLK2.n331 GND 0.12fF $ **FLOATING
C5092 CLK2.n332 GND 0.12fF $ **FLOATING
C5093 CLK2.t46 GND 0.06fF
C5094 CLK2.n333 GND 0.07fF $ **FLOATING
C5095 CLK2.n334 GND 0.02fF $ **FLOATING
C5096 CLK2.n335 GND 0.02fF $ **FLOATING
C5097 CLK2.n336 GND 0.02fF $ **FLOATING
C5098 CLK2.n337 GND 0.13fF $ **FLOATING
C5099 EESPFAL_s3_0/EESPFAL_NAND_v3_0/CLK GND 0.01fF $ **FLOATING
C5100 CLK2.n338 GND 0.02fF $ **FLOATING
C5101 CLK2.n339 GND 0.02fF $ **FLOATING
C5102 CLK2.n340 GND 0.02fF $ **FLOATING
C5103 CLK2.n341 GND 0.07fF $ **FLOATING
C5104 CLK2.n342 GND 0.12fF $ **FLOATING
C5105 CLK2.t107 GND 0.06fF
C5106 CLK2.n343 GND 0.13fF $ **FLOATING
C5107 CLK2.n344 GND 0.08fF $ **FLOATING
C5108 CLK2.n345 GND 0.02fF $ **FLOATING
C5109 CLK2.n346 GND 0.02fF $ **FLOATING
C5110 CLK2.n347 GND 0.02fF $ **FLOATING
C5111 CLK2.n348 GND 0.21fF $ **FLOATING
C5112 CLK2.n349 GND 0.01fF $ **FLOATING
C5113 CLK2.n350 GND 0.01fF $ **FLOATING
C5114 CLK2.n351 GND 0.02fF $ **FLOATING
C5115 CLK2.n352 GND 0.02fF $ **FLOATING
C5116 CLK2.n353 GND 0.02fF $ **FLOATING
C5117 CLK2.n354 GND 0.02fF $ **FLOATING
C5118 CLK2.n355 GND 0.04fF $ **FLOATING
C5119 CLK2.n356 GND 0.04fF $ **FLOATING
C5120 CLK2.n357 GND 0.04fF $ **FLOATING
C5121 CLK2.n358 GND 0.02fF $ **FLOATING
C5122 CLK2.n359 GND 0.02fF $ **FLOATING
C5123 CLK2.n360 GND 0.02fF $ **FLOATING
C5124 CLK2.n361 GND 0.09fF $ **FLOATING
C5125 CLK2.n362 GND 0.05fF $ **FLOATING
C5126 CLK2.n363 GND 0.14fF $ **FLOATING
C5127 CLK2.n364 GND 0.02fF $ **FLOATING
C5128 CLK2.n365 GND 0.02fF $ **FLOATING
C5129 CLK2.n366 GND 0.01fF $ **FLOATING
C5130 CLK2.n367 GND 0.00fF $ **FLOATING
C5131 CLK2.n369 GND 0.01fF $ **FLOATING
C5132 CLK2.n370 GND 0.05fF $ **FLOATING
C5133 EESPFAL_s2_0/CLK2 GND 0.05fF $ **FLOATING
C5134 CLK2.n371 GND 0.00fF $ **FLOATING
C5135 CLK2.t12 GND 0.03fF
C5136 CLK2.t48 GND 0.03fF
C5137 CLK2.n372 GND 0.11fF $ **FLOATING
C5138 CLK2.n373 GND 0.05fF $ **FLOATING
C5139 CLK2.n374 GND 0.02fF $ **FLOATING
C5140 CLK2.n375 GND 0.02fF $ **FLOATING
C5141 CLK2.n376 GND 0.09fF $ **FLOATING
C5142 CLK2.n377 GND 0.04fF $ **FLOATING
C5143 CLK2.n378 GND 0.02fF $ **FLOATING
C5144 CLK2.n379 GND 0.02fF $ **FLOATING
C5145 CLK2.n380 GND 0.05fF $ **FLOATING
C5146 CLK2.n381 GND 0.14fF $ **FLOATING
C5147 CLK2.n382 GND 0.01fF $ **FLOATING
C5148 CLK2.n383 GND 0.04fF $ **FLOATING
C5149 CLK2.n384 GND 0.02fF $ **FLOATING
C5150 CLK2.n385 GND 0.02fF $ **FLOATING
C5151 CLK2.n386 GND 0.00fF $ **FLOATING
C5152 CLK2.n387 GND 0.00fF $ **FLOATING
C5153 CLK2.n388 GND 0.01fF $ **FLOATING
C5154 CLK2.n389 GND 0.02fF $ **FLOATING
C5155 CLK2.n390 GND 0.10fF $ **FLOATING
C5156 CLK2.n391 GND 0.02fF $ **FLOATING
C5157 CLK2.n392 GND 0.02fF $ **FLOATING
C5158 CLK2.n393 GND 0.02fF $ **FLOATING
C5159 CLK2.n394 GND 0.13fF $ **FLOATING
C5160 CLK2.n395 GND 0.02fF $ **FLOATING
C5161 CLK2.n396 GND 0.02fF $ **FLOATING
C5162 CLK2.n397 GND 0.01fF $ **FLOATING
C5163 CLK2.n398 GND 0.21fF $ **FLOATING
C5164 CLK2.t2 GND 0.06fF
C5165 CLK2.n399 GND 0.08fF $ **FLOATING
C5166 CLK2.n400 GND 0.02fF $ **FLOATING
C5167 CLK2.n401 GND 0.02fF $ **FLOATING
C5168 CLK2.n402 GND 0.02fF $ **FLOATING
C5169 CLK2.n403 GND 0.12fF $ **FLOATING
C5170 CLK2.n404 GND 0.02fF $ **FLOATING
C5171 CLK2.n405 GND 0.02fF $ **FLOATING
C5172 CLK2.n406 GND 0.02fF $ **FLOATING
C5173 CLK2.n407 GND 0.02fF $ **FLOATING
C5174 CLK2.t0 GND 0.06fF
C5175 CLK2.n408 GND 0.07fF $ **FLOATING
C5176 CLK2.n409 GND 0.02fF $ **FLOATING
C5177 CLK2.n410 GND 0.02fF $ **FLOATING
C5178 CLK2.n411 GND 0.12fF $ **FLOATING
C5179 CLK2.n412 GND 0.02fF $ **FLOATING
C5180 CLK2.n413 GND 0.02fF $ **FLOATING
C5181 CLK2.n414 GND 0.13fF $ **FLOATING
C5182 CLK2.t56 GND 0.06fF
C5183 CLK2.n415 GND 0.07fF $ **FLOATING
C5184 CLK2.n416 GND 0.02fF $ **FLOATING
C5185 CLK2.n417 GND 0.02fF $ **FLOATING
C5186 CLK2.n418 GND 0.02fF $ **FLOATING
C5187 CLK2.n419 GND 0.12fF $ **FLOATING
C5188 CLK2.n420 GND 0.02fF $ **FLOATING
C5189 CLK2.n421 GND 0.02fF $ **FLOATING
C5190 CLK2.n422 GND 0.02fF $ **FLOATING
C5191 CLK2.t82 GND 0.06fF
C5192 CLK2.n423 GND 0.08fF $ **FLOATING
C5193 CLK2.n424 GND 0.02fF $ **FLOATING
C5194 CLK2.n425 GND 0.02fF $ **FLOATING
C5195 CLK2.n426 GND 0.02fF $ **FLOATING
C5196 CLK2.n427 GND 0.21fF $ **FLOATING
C5197 CLK2.n428 GND 0.13fF $ **FLOATING
C5198 CLK2.n429 GND 0.02fF $ **FLOATING
C5199 CLK2.n430 GND 0.02fF $ **FLOATING
C5200 CLK2.n431 GND 0.01fF $ **FLOATING
C5201 CLK2.n432 GND 0.10fF $ **FLOATING
C5202 CLK2.n433 GND 0.02fF $ **FLOATING
C5203 CLK2.n434 GND 0.02fF $ **FLOATING
C5204 CLK2.n435 GND 0.02fF $ **FLOATING
C5205 CLK2.n436 GND 0.04fF $ **FLOATING
C5206 CLK2.n437 GND 0.02fF $ **FLOATING
C5207 CLK2.n438 GND 0.02fF $ **FLOATING
C5208 CLK2.n439 GND 0.02fF $ **FLOATING
C5209 CLK2.n440 GND 0.04fF $ **FLOATING
C5210 CLK2.n441 GND 0.02fF $ **FLOATING
C5211 CLK2.n442 GND 0.02fF $ **FLOATING
C5212 CLK2.n443 GND 0.02fF $ **FLOATING
C5213 CLK2.n444 GND 0.04fF $ **FLOATING
C5214 CLK2.n445 GND 0.02fF $ **FLOATING
C5215 CLK2.n446 GND 0.02fF $ **FLOATING
C5216 CLK2.n447 GND 0.02fF $ **FLOATING
C5217 CLK2.n448 GND 0.05fF $ **FLOATING
C5218 CLK2.n449 GND 0.02fF $ **FLOATING
C5219 CLK2.n450 GND 0.02fF $ **FLOATING
C5220 CLK2.n451 GND 0.02fF $ **FLOATING
C5221 CLK2.n452 GND 0.06fF $ **FLOATING
C5222 CLK2.n453 GND 0.02fF $ **FLOATING
C5223 CLK2.n454 GND 0.06fF $ **FLOATING
C5224 CLK2.n455 GND 0.02fF $ **FLOATING
C5225 CLK2.t106 GND 0.03fF
C5226 CLK2.n456 GND 0.08fF $ **FLOATING
C5227 CLK2.n457 GND 0.01fF $ **FLOATING
C5228 CLK2.n458 GND 0.09fF $ **FLOATING
C5229 CLK2.n459 GND 0.08fF $ **FLOATING
C5230 CLK2.n460 GND 0.02fF $ **FLOATING
C5231 CLK2.n461 GND 0.02fF $ **FLOATING
C5232 CLK2.t30 GND 0.03fF
C5233 CLK2.n462 GND 0.08fF $ **FLOATING
C5234 CLK2.n463 GND 0.01fF $ **FLOATING
C5235 CLK2.n464 GND 0.07fF $ **FLOATING
C5236 CLK2.n465 GND 0.09fF $ **FLOATING
C5237 CLK2.n466 GND 0.06fF $ **FLOATING
C5238 CLK2.n467 GND 0.05fF $ **FLOATING
C5239 CLK2.n468 GND 0.02fF $ **FLOATING
C5240 CLK2.n469 GND 0.02fF $ **FLOATING
C5241 CLK2.n470 GND 0.02fF $ **FLOATING
C5242 CLK2.n471 GND 0.04fF $ **FLOATING
C5243 CLK2.n472 GND 0.02fF $ **FLOATING
C5244 CLK2.n473 GND 0.02fF $ **FLOATING
C5245 CLK2.n474 GND 0.02fF $ **FLOATING
C5246 CLK2.n475 GND 0.04fF $ **FLOATING
C5247 CLK2.n476 GND 0.02fF $ **FLOATING
C5248 CLK2.n477 GND 0.02fF $ **FLOATING
C5249 CLK2.n478 GND 0.02fF $ **FLOATING
C5250 CLK2.n479 GND 0.04fF $ **FLOATING
C5251 CLK2.n480 GND 0.02fF $ **FLOATING
C5252 CLK2.n481 GND 0.02fF $ **FLOATING
C5253 CLK2.n482 GND 0.02fF $ **FLOATING
C5254 CLK2.n483 GND 0.10fF $ **FLOATING
C5255 CLK2.n484 GND 0.02fF $ **FLOATING
C5256 CLK2.n485 GND 0.02fF $ **FLOATING
C5257 CLK2.n486 GND 0.02fF $ **FLOATING
C5258 CLK2.n487 GND 0.13fF $ **FLOATING
C5259 CLK2.n488 GND 0.02fF $ **FLOATING
C5260 CLK2.n489 GND 0.02fF $ **FLOATING
C5261 CLK2.n490 GND 0.01fF $ **FLOATING
C5262 CLK2.n491 GND 0.21fF $ **FLOATING
C5263 CLK2.t37 GND 0.06fF
C5264 CLK2.n492 GND 0.08fF $ **FLOATING
C5265 CLK2.n493 GND 0.02fF $ **FLOATING
C5266 CLK2.n494 GND 0.02fF $ **FLOATING
C5267 CLK2.n495 GND 0.02fF $ **FLOATING
C5268 CLK2.n496 GND 0.12fF $ **FLOATING
C5269 CLK2.n497 GND 0.02fF $ **FLOATING
C5270 CLK2.n498 GND 0.02fF $ **FLOATING
C5271 CLK2.n499 GND 0.02fF $ **FLOATING
C5272 CLK2.t35 GND 0.06fF
C5273 CLK2.n500 GND 0.07fF $ **FLOATING
C5274 CLK2.n501 GND 0.02fF $ **FLOATING
C5275 CLK2.n502 GND 0.02fF $ **FLOATING
C5276 CLK2.n503 GND 0.02fF $ **FLOATING
C5277 CLK2.n504 GND 0.13fF $ **FLOATING
C5278 CLK2.n505 GND 0.12fF $ **FLOATING
C5279 CLK2.n506 GND 0.02fF $ **FLOATING
C5280 CLK2.n507 GND 0.02fF $ **FLOATING
C5281 CLK2.t103 GND 0.06fF
C5282 CLK2.n508 GND 0.07fF $ **FLOATING
C5283 CLK2.n509 GND 0.02fF $ **FLOATING
C5284 CLK2.n510 GND 0.02fF $ **FLOATING
C5285 CLK2.n511 GND 0.02fF $ **FLOATING
C5286 CLK2.n512 GND 0.12fF $ **FLOATING
C5287 CLK2.n513 GND 0.02fF $ **FLOATING
C5288 CLK2.n514 GND 0.02fF $ **FLOATING
C5289 CLK2.n515 GND 0.02fF $ **FLOATING
C5290 CLK2.t101 GND 0.06fF
C5291 CLK2.n516 GND 0.08fF $ **FLOATING
C5292 CLK2.n517 GND 0.02fF $ **FLOATING
C5293 CLK2.n518 GND 0.02fF $ **FLOATING
C5294 CLK2.n519 GND 0.02fF $ **FLOATING
C5295 CLK2.n520 GND 0.21fF $ **FLOATING
C5296 CLK2.n521 GND 0.13fF $ **FLOATING
C5297 CLK2.n522 GND 0.02fF $ **FLOATING
C5298 CLK2.n523 GND 0.02fF $ **FLOATING
C5299 CLK2.n524 GND 0.01fF $ **FLOATING
C5300 CLK2.n525 GND 0.10fF $ **FLOATING
C5301 CLK2.n526 GND 0.02fF $ **FLOATING
C5302 CLK2.n527 GND 0.02fF $ **FLOATING
C5303 CLK2.n528 GND 0.02fF $ **FLOATING
C5304 CLK2.n529 GND 0.04fF $ **FLOATING
C5305 CLK2.n530 GND 0.02fF $ **FLOATING
C5306 CLK2.n531 GND 0.02fF $ **FLOATING
C5307 CLK2.n532 GND 0.02fF $ **FLOATING
C5308 CLK2.n533 GND 0.04fF $ **FLOATING
C5309 CLK2.n534 GND 0.02fF $ **FLOATING
C5310 CLK2.n535 GND 0.02fF $ **FLOATING
C5311 CLK2.n536 GND 0.02fF $ **FLOATING
C5312 CLK2.n537 GND 0.14fF $ **FLOATING
C5313 CLK2.n538 GND 0.04fF $ **FLOATING
C5314 CLK2.n539 GND 0.02fF $ **FLOATING
C5315 CLK2.n540 GND 0.02fF $ **FLOATING
C5316 CLK2.n541 GND 0.01fF $ **FLOATING
C5317 CLK2.n542 GND 0.05fF $ **FLOATING
C5318 CLK2.n543 GND 0.02fF $ **FLOATING
C5319 CLK2.n544 GND 0.02fF $ **FLOATING
C5320 CLK2.n545 GND 0.02fF $ **FLOATING
C5321 CLK2.n546 GND 0.09fF $ **FLOATING
C5322 CLK2.n547 GND 0.15fF $ **FLOATING
C5323 CLK2.t60 GND 0.04fF
C5324 CLK2.t40 GND 0.03fF
C5325 CLK2.t25 GND 0.03fF
C5326 CLK2.n548 GND 0.08fF $ **FLOATING
C5327 EESPFAL_s2_0/EESPFAL_INV4_2/CLK GND 0.01fF $ **FLOATING
C5328 CLK2.t114 GND 0.04fF
C5329 CLK2.t96 GND 0.05fF
C5330 CLK2.n549 GND 0.11fF $ **FLOATING
C5331 CLK2.n550 GND 0.34fF $ **FLOATING
C5332 CLK2.n551 GND 0.05fF $ **FLOATING
C5333 CLK2.n552 GND 0.02fF $ **FLOATING
C5334 CLK2.n553 GND 0.02fF $ **FLOATING
C5335 CLK2.n554 GND 0.02fF $ **FLOATING
C5336 CLK2.n555 GND 0.04fF $ **FLOATING
C5337 CLK2.n556 GND 0.02fF $ **FLOATING
C5338 CLK2.n557 GND 0.02fF $ **FLOATING
C5339 CLK2.n558 GND 0.02fF $ **FLOATING
C5340 CLK2.n559 GND 0.10fF $ **FLOATING
C5341 CLK2.n560 GND 0.02fF $ **FLOATING
C5342 CLK2.n561 GND 0.02fF $ **FLOATING
C5343 CLK2.n562 GND 0.02fF $ **FLOATING
C5344 CLK2.n563 GND 0.13fF $ **FLOATING
C5345 CLK2.n564 GND 0.02fF $ **FLOATING
C5346 CLK2.n565 GND 0.02fF $ **FLOATING
C5347 CLK2.n566 GND 0.01fF $ **FLOATING
C5348 CLK2.n567 GND 0.21fF $ **FLOATING
C5349 CLK2.t113 GND 0.06fF
C5350 CLK2.n568 GND 0.08fF $ **FLOATING
C5351 CLK2.n569 GND 0.02fF $ **FLOATING
C5352 CLK2.n570 GND 0.02fF $ **FLOATING
C5353 CLK2.n571 GND 0.02fF $ **FLOATING
C5354 CLK2.n572 GND 0.12fF $ **FLOATING
C5355 CLK2.n573 GND 0.02fF $ **FLOATING
C5356 CLK2.n574 GND 0.02fF $ **FLOATING
C5357 CLK2.n575 GND 0.02fF $ **FLOATING
C5358 CLK2.n576 GND 0.02fF $ **FLOATING
C5359 CLK2.t24 GND 0.06fF
C5360 CLK2.n577 GND 0.07fF $ **FLOATING
C5361 CLK2.n578 GND 0.02fF $ **FLOATING
C5362 CLK2.n579 GND 0.02fF $ **FLOATING
C5363 CLK2.n580 GND 0.12fF $ **FLOATING
C5364 CLK2.n581 GND 0.02fF $ **FLOATING
C5365 CLK2.n582 GND 0.02fF $ **FLOATING
C5366 CLK2.n583 GND 0.13fF $ **FLOATING
C5367 CLK2.t39 GND 0.06fF
C5368 CLK2.n584 GND 0.07fF $ **FLOATING
C5369 CLK2.n585 GND 0.02fF $ **FLOATING
C5370 CLK2.n586 GND 0.02fF $ **FLOATING
C5371 CLK2.n587 GND 0.02fF $ **FLOATING
C5372 CLK2.n588 GND 0.12fF $ **FLOATING
C5373 CLK2.n589 GND 0.02fF $ **FLOATING
C5374 CLK2.n590 GND 0.02fF $ **FLOATING
C5375 CLK2.n591 GND 0.02fF $ **FLOATING
C5376 CLK2.t59 GND 0.06fF
C5377 CLK2.n592 GND 0.08fF $ **FLOATING
C5378 CLK2.n593 GND 0.02fF $ **FLOATING
C5379 CLK2.n594 GND 0.02fF $ **FLOATING
C5380 CLK2.n595 GND 0.02fF $ **FLOATING
C5381 CLK2.n596 GND 0.21fF $ **FLOATING
C5382 CLK2.n597 GND 0.13fF $ **FLOATING
C5383 CLK2.n598 GND 0.02fF $ **FLOATING
C5384 CLK2.n599 GND 0.02fF $ **FLOATING
C5385 CLK2.n600 GND 0.01fF $ **FLOATING
C5386 CLK2.n601 GND 0.10fF $ **FLOATING
C5387 CLK2.n602 GND 0.02fF $ **FLOATING
C5388 CLK2.n603 GND 0.02fF $ **FLOATING
C5389 CLK2.n604 GND 0.02fF $ **FLOATING
C5390 CLK2.n605 GND 0.04fF $ **FLOATING
C5391 CLK2.n606 GND 0.02fF $ **FLOATING
C5392 CLK2.n607 GND 0.02fF $ **FLOATING
C5393 CLK2.n608 GND 0.01fF $ **FLOATING
C5394 CLK2.n609 GND 0.15fF $ **FLOATING
C5395 CLK2.n610 GND 0.05fF $ **FLOATING
C5396 CLK2.n611 GND 0.02fF $ **FLOATING
C5397 CLK2.n612 GND 0.02fF $ **FLOATING
C5398 CLK2.n613 GND 0.02fF $ **FLOATING
C5399 CLK2.n614 GND 0.11fF $ **FLOATING
C5400 CLK2.n615 GND 0.02fF $ **FLOATING
C5401 CLK2.n616 GND 0.09fF $ **FLOATING
C5402 CLK2.n617 GND 0.02fF $ **FLOATING
C5403 CLK2.n618 GND 0.12fF $ **FLOATING
C5404 CLK2.n619 GND 0.11fF $ **FLOATING
C5405 CLK2.n620 GND 0.02fF $ **FLOATING
C5406 CLK2.n621 GND 0.02fF $ **FLOATING
C5407 CLK2.n622 GND 0.10fF $ **FLOATING
C5408 CLK2.t75 GND 0.04fF
C5409 CLK2.t77 GND 0.03fF
C5410 CLK2.t52 GND 0.03fF
C5411 CLK2.n623 GND 0.08fF $ **FLOATING
C5412 EESPFAL_s1_0/EESPFAL_INV4_0/CLK GND 0.01fF $ **FLOATING
C5413 CLK2.t50 GND 0.04fF
C5414 CLK2.t11 GND 0.05fF
C5415 CLK2.n624 GND 0.11fF $ **FLOATING
C5416 CLK2.n625 GND 0.34fF $ **FLOATING
C5417 CLK2.n626 GND 0.05fF $ **FLOATING
C5418 CLK2.n627 GND 0.02fF $ **FLOATING
C5419 CLK2.n628 GND 0.02fF $ **FLOATING
C5420 CLK2.n629 GND 0.02fF $ **FLOATING
C5421 CLK2.n630 GND 0.04fF $ **FLOATING
C5422 CLK2.n631 GND 0.02fF $ **FLOATING
C5423 CLK2.n632 GND 0.02fF $ **FLOATING
C5424 CLK2.n633 GND 0.02fF $ **FLOATING
C5425 CLK2.n634 GND 0.10fF $ **FLOATING
C5426 CLK2.n635 GND 0.02fF $ **FLOATING
C5427 CLK2.n636 GND 0.02fF $ **FLOATING
C5428 CLK2.n637 GND 0.02fF $ **FLOATING
C5429 CLK2.n638 GND 0.13fF $ **FLOATING
C5430 CLK2.n639 GND 0.02fF $ **FLOATING
C5431 CLK2.n640 GND 0.02fF $ **FLOATING
C5432 CLK2.n641 GND 0.01fF $ **FLOATING
C5433 CLK2.n642 GND 0.21fF $ **FLOATING
C5434 CLK2.t49 GND 0.06fF
C5435 CLK2.n643 GND 0.08fF $ **FLOATING
C5436 CLK2.n644 GND 0.02fF $ **FLOATING
C5437 CLK2.n645 GND 0.02fF $ **FLOATING
C5438 CLK2.n646 GND 0.02fF $ **FLOATING
C5439 CLK2.n647 GND 0.12fF $ **FLOATING
C5440 CLK2.n648 GND 0.02fF $ **FLOATING
C5441 CLK2.n649 GND 0.02fF $ **FLOATING
C5442 CLK2.n650 GND 0.02fF $ **FLOATING
C5443 CLK2.n651 GND 0.02fF $ **FLOATING
C5444 CLK2.t51 GND 0.06fF
C5445 CLK2.n652 GND 0.07fF $ **FLOATING
C5446 CLK2.n653 GND 0.02fF $ **FLOATING
C5447 CLK2.n654 GND 0.02fF $ **FLOATING
C5448 CLK2.n655 GND 0.12fF $ **FLOATING
C5449 CLK2.n656 GND 0.02fF $ **FLOATING
C5450 CLK2.n657 GND 0.02fF $ **FLOATING
C5451 CLK2.n658 GND 0.13fF $ **FLOATING
C5452 CLK2.t76 GND 0.06fF
C5453 CLK2.n659 GND 0.07fF $ **FLOATING
C5454 CLK2.n660 GND 0.02fF $ **FLOATING
C5455 CLK2.n661 GND 0.02fF $ **FLOATING
C5456 CLK2.n662 GND 0.02fF $ **FLOATING
C5457 CLK2.n663 GND 0.12fF $ **FLOATING
C5458 CLK2.n664 GND 0.02fF $ **FLOATING
C5459 CLK2.n665 GND 0.02fF $ **FLOATING
C5460 CLK2.n666 GND 0.02fF $ **FLOATING
C5461 CLK2.t74 GND 0.06fF
C5462 CLK2.n667 GND 0.08fF $ **FLOATING
C5463 CLK2.n668 GND 0.02fF $ **FLOATING
C5464 CLK2.n669 GND 0.02fF $ **FLOATING
C5465 CLK2.n670 GND 0.02fF $ **FLOATING
C5466 CLK2.n671 GND 0.21fF $ **FLOATING
C5467 CLK2.n672 GND 0.13fF $ **FLOATING
C5468 CLK2.n673 GND 0.02fF $ **FLOATING
C5469 CLK2.n674 GND 0.02fF $ **FLOATING
C5470 CLK2.n675 GND 0.01fF $ **FLOATING
C5471 CLK2.n676 GND 0.10fF $ **FLOATING
C5472 CLK2.n677 GND 0.02fF $ **FLOATING
C5473 CLK2.n678 GND 0.02fF $ **FLOATING
C5474 CLK2.n679 GND 0.02fF $ **FLOATING
C5475 CLK2.n680 GND 0.04fF $ **FLOATING
C5476 CLK2.n681 GND 0.02fF $ **FLOATING
C5477 CLK2.n682 GND 0.02fF $ **FLOATING
C5478 CLK2.n683 GND 0.02fF $ **FLOATING
C5479 CLK2.n684 GND 0.05fF $ **FLOATING
C5480 CLK2.n685 GND 0.02fF $ **FLOATING
C5481 CLK2.n686 GND 0.02fF $ **FLOATING
C5482 CLK2.n687 GND 0.02fF $ **FLOATING
C5483 CLK2.n688 GND 0.09fF $ **FLOATING
C5484 CLK2.n689 GND 0.15fF $ **FLOATING
C5485 CLK2.n690 GND 0.15fF $ **FLOATING
C5486 CLK2.n691 GND 0.05fF $ **FLOATING
C5487 CLK2.n692 GND 0.02fF $ **FLOATING
C5488 CLK2.n693 GND 0.02fF $ **FLOATING
C5489 CLK2.n694 GND 0.02fF $ **FLOATING
C5490 CLK2.n695 GND 0.04fF $ **FLOATING
C5491 CLK2.n696 GND 0.02fF $ **FLOATING
C5492 CLK2.n697 GND 0.02fF $ **FLOATING
C5493 CLK2.n698 GND 0.01fF $ **FLOATING
C5494 CLK2.n699 GND 0.14fF $ **FLOATING
C5495 CLK2.n700 GND 0.04fF $ **FLOATING
C5496 CLK2.n701 GND 0.02fF $ **FLOATING
C5497 CLK2.n702 GND 0.02fF $ **FLOATING
C5498 CLK2.n703 GND 0.02fF $ **FLOATING
C5499 CLK2.n704 GND 0.04fF $ **FLOATING
C5500 CLK2.n705 GND 0.02fF $ **FLOATING
C5501 CLK2.n706 GND 0.02fF $ **FLOATING
C5502 CLK2.n707 GND 0.02fF $ **FLOATING
C5503 CLK2.n708 GND 0.10fF $ **FLOATING
C5504 CLK2.n709 GND 0.02fF $ **FLOATING
C5505 CLK2.n710 GND 0.02fF $ **FLOATING
C5506 CLK2.n711 GND 0.02fF $ **FLOATING
C5507 CLK2.n712 GND 0.13fF $ **FLOATING
C5508 CLK2.n713 GND 0.02fF $ **FLOATING
C5509 CLK2.n714 GND 0.02fF $ **FLOATING
C5510 CLK2.n715 GND 0.01fF $ **FLOATING
C5511 CLK2.n716 GND 0.21fF $ **FLOATING
C5512 CLK2.t31 GND 0.06fF
C5513 CLK2.n717 GND 0.08fF $ **FLOATING
C5514 CLK2.n718 GND 0.02fF $ **FLOATING
C5515 CLK2.n719 GND 0.02fF $ **FLOATING
C5516 CLK2.n720 GND 0.02fF $ **FLOATING
C5517 CLK2.n721 GND 0.12fF $ **FLOATING
C5518 CLK2.n722 GND 0.02fF $ **FLOATING
C5519 CLK2.n723 GND 0.02fF $ **FLOATING
C5520 CLK2.n724 GND 0.02fF $ **FLOATING
C5521 CLK2.n725 GND 0.02fF $ **FLOATING
C5522 CLK2.t33 GND 0.06fF
C5523 CLK2.n726 GND 0.07fF $ **FLOATING
C5524 CLK2.n727 GND 0.02fF $ **FLOATING
C5525 CLK2.n728 GND 0.02fF $ **FLOATING
C5526 CLK2.n729 GND 0.12fF $ **FLOATING
C5527 CLK2.n730 GND 0.02fF $ **FLOATING
C5528 CLK2.n731 GND 0.02fF $ **FLOATING
C5529 CLK2.n732 GND 0.13fF $ **FLOATING
C5530 CLK2.t94 GND 0.06fF
C5531 CLK2.n733 GND 0.07fF $ **FLOATING
C5532 CLK2.n734 GND 0.02fF $ **FLOATING
C5533 CLK2.n735 GND 0.02fF $ **FLOATING
C5534 CLK2.n736 GND 0.02fF $ **FLOATING
C5535 CLK2.n737 GND 0.12fF $ **FLOATING
C5536 CLK2.n738 GND 0.02fF $ **FLOATING
C5537 CLK2.n739 GND 0.02fF $ **FLOATING
C5538 CLK2.n740 GND 0.02fF $ **FLOATING
C5539 CLK2.t92 GND 0.06fF
C5540 CLK2.n741 GND 0.08fF $ **FLOATING
C5541 CLK2.n742 GND 0.02fF $ **FLOATING
C5542 CLK2.n743 GND 0.02fF $ **FLOATING
C5543 CLK2.n744 GND 0.02fF $ **FLOATING
C5544 CLK2.n745 GND 0.21fF $ **FLOATING
C5545 CLK2.n746 GND 0.13fF $ **FLOATING
C5546 CLK2.n747 GND 0.02fF $ **FLOATING
C5547 CLK2.n748 GND 0.02fF $ **FLOATING
C5548 CLK2.n749 GND 0.01fF $ **FLOATING
C5549 CLK2.n750 GND 0.10fF $ **FLOATING
C5550 CLK2.n751 GND 0.02fF $ **FLOATING
C5551 CLK2.n752 GND 0.02fF $ **FLOATING
C5552 CLK2.n753 GND 0.02fF $ **FLOATING
C5553 CLK2.n754 GND 0.04fF $ **FLOATING
C5554 CLK2.n755 GND 0.02fF $ **FLOATING
C5555 CLK2.n756 GND 0.02fF $ **FLOATING
C5556 CLK2.n757 GND 0.02fF $ **FLOATING
C5557 CLK2.n758 GND 0.04fF $ **FLOATING
C5558 CLK2.n759 GND 0.02fF $ **FLOATING
C5559 CLK2.n760 GND 0.02fF $ **FLOATING
C5560 CLK2.n761 GND 0.02fF $ **FLOATING
C5561 CLK2.n762 GND 0.04fF $ **FLOATING
C5562 CLK2.n763 GND 0.02fF $ **FLOATING
C5563 CLK2.n764 GND 0.02fF $ **FLOATING
C5564 CLK2.n765 GND 0.02fF $ **FLOATING
C5565 CLK2.n766 GND 0.05fF $ **FLOATING
C5566 CLK2.n767 GND 0.02fF $ **FLOATING
C5567 CLK2.n768 GND 0.02fF $ **FLOATING
C5568 CLK2.n769 GND 0.02fF $ **FLOATING
C5569 CLK2.n770 GND 0.06fF $ **FLOATING
C5570 CLK2.n771 GND 0.02fF $ **FLOATING
C5571 CLK2.n772 GND 0.06fF $ **FLOATING
C5572 CLK2.n773 GND 0.02fF $ **FLOATING
C5573 CLK2.t81 GND 0.03fF
C5574 CLK2.n774 GND 0.08fF $ **FLOATING
C5575 CLK2.n775 GND 0.01fF $ **FLOATING
C5576 CLK2.n776 GND 0.09fF $ **FLOATING
C5577 CLK2.n777 GND 0.08fF $ **FLOATING
C5578 CLK2.n778 GND 0.02fF $ **FLOATING
C5579 CLK2.n779 GND 0.02fF $ **FLOATING
C5580 CLK2.n780 GND 0.07fF $ **FLOATING
C5581 CLK2.n781 GND 0.04fF $ **FLOATING
C5582 CLK2.n782 GND 0.09fF $ **FLOATING
C5583 CLK2.n783 GND 0.01fF $ **FLOATING
C5584 EESPFAL_s1_0/CLK2 GND 0.02fF $ **FLOATING
C5585 CLK2.n784 GND 0.01fF $ **FLOATING
C5586 CLK2.n785 GND 0.05fF $ **FLOATING
C5587 CLK2.n786 GND 0.02fF $ **FLOATING
C5588 CLK2.n787 GND 0.02fF $ **FLOATING
C5589 CLK2.n788 GND 0.02fF $ **FLOATING
C5590 CLK2.n789 GND 0.04fF $ **FLOATING
C5591 CLK2.n790 GND 0.02fF $ **FLOATING
C5592 CLK2.n791 GND 0.02fF $ **FLOATING
C5593 CLK2.n792 GND 0.02fF $ **FLOATING
C5594 CLK2.n793 GND 0.04fF $ **FLOATING
C5595 CLK2.n794 GND 0.02fF $ **FLOATING
C5596 CLK2.n795 GND 0.02fF $ **FLOATING
C5597 CLK2.n796 GND 0.02fF $ **FLOATING
C5598 CLK2.n797 GND 0.04fF $ **FLOATING
C5599 CLK2.n798 GND 0.02fF $ **FLOATING
C5600 CLK2.n799 GND 0.02fF $ **FLOATING
C5601 CLK2.n800 GND 0.02fF $ **FLOATING
C5602 CLK2.n801 GND 0.10fF $ **FLOATING
C5603 CLK2.n802 GND 0.02fF $ **FLOATING
C5604 CLK2.n803 GND 0.02fF $ **FLOATING
C5605 CLK2.n804 GND 0.02fF $ **FLOATING
C5606 CLK2.n805 GND 0.13fF $ **FLOATING
C5607 CLK2.n806 GND 0.02fF $ **FLOATING
C5608 CLK2.n807 GND 0.02fF $ **FLOATING
C5609 CLK2.n808 GND 0.01fF $ **FLOATING
C5610 CLK2.n809 GND 0.21fF $ **FLOATING
C5611 CLK2.t41 GND 0.06fF
C5612 CLK2.n810 GND 0.08fF $ **FLOATING
C5613 CLK2.n811 GND 0.02fF $ **FLOATING
C5614 CLK2.n812 GND 0.02fF $ **FLOATING
C5615 CLK2.n813 GND 0.02fF $ **FLOATING
C5616 CLK2.n814 GND 0.12fF $ **FLOATING
C5617 CLK2.n815 GND 0.02fF $ **FLOATING
C5618 CLK2.n816 GND 0.02fF $ **FLOATING
C5619 CLK2.n817 GND 0.02fF $ **FLOATING
C5620 CLK2.t111 GND 0.06fF
C5621 CLK2.n818 GND 0.07fF $ **FLOATING
C5622 CLK2.n819 GND 0.02fF $ **FLOATING
C5623 CLK2.n820 GND 0.02fF $ **FLOATING
C5624 CLK2.n821 GND 0.02fF $ **FLOATING
C5625 CLK2.n822 GND 0.13fF $ **FLOATING
C5626 CLK2.n823 GND 0.02fF $ **FLOATING
C5627 CLK2.t6 GND 0.06fF
C5628 CLK2.n824 GND 0.07fF $ **FLOATING
C5629 CLK2.n825 GND 0.02fF $ **FLOATING
C5630 CLK2.n826 GND 0.02fF $ **FLOATING
C5631 CLK2.n827 GND 0.02fF $ **FLOATING
C5632 CLK2.n828 GND 0.12fF $ **FLOATING
C5633 CLK2.n829 GND 0.02fF $ **FLOATING
C5634 CLK2.n830 GND 0.02fF $ **FLOATING
C5635 CLK2.n831 GND 0.02fF $ **FLOATING
C5636 CLK2.t4 GND 0.06fF
C5637 CLK2.n832 GND 0.08fF $ **FLOATING
C5638 CLK2.n833 GND 0.02fF $ **FLOATING
C5639 CLK2.n834 GND 0.02fF $ **FLOATING
C5640 CLK2.n835 GND 0.02fF $ **FLOATING
C5641 CLK2.n836 GND 0.21fF $ **FLOATING
C5642 CLK2.n837 GND 0.13fF $ **FLOATING
C5643 CLK2.n838 GND 0.02fF $ **FLOATING
C5644 CLK2.n839 GND 0.02fF $ **FLOATING
C5645 CLK2.n840 GND 0.01fF $ **FLOATING
C5646 CLK2.n841 GND 0.10fF $ **FLOATING
C5647 CLK2.n842 GND 0.02fF $ **FLOATING
C5648 CLK2.n843 GND 0.02fF $ **FLOATING
C5649 CLK2.n844 GND 0.02fF $ **FLOATING
C5650 CLK2.n845 GND 0.04fF $ **FLOATING
C5651 CLK2.n846 GND 0.02fF $ **FLOATING
C5652 CLK2.n847 GND 0.02fF $ **FLOATING
C5653 CLK2.n848 GND 0.02fF $ **FLOATING
C5654 CLK2.n849 GND 0.04fF $ **FLOATING
C5655 CLK2.n850 GND 0.02fF $ **FLOATING
C5656 CLK2.n851 GND 0.02fF $ **FLOATING
C5657 CLK2.n852 GND 0.02fF $ **FLOATING
C5658 CLK2.n853 GND 0.14fF $ **FLOATING
C5659 CLK2.n854 GND 0.05fF $ **FLOATING
C5660 CLK2.n855 GND 0.09fF $ **FLOATING
C5661 CLK2.n856 GND 0.01fF $ **FLOATING
C5662 CLK2.n857 GND 0.09fF $ **FLOATING
C5663 CLK2.n858 GND 0.16fF $ **FLOATING
C5664 CLK2.t64 GND 0.04fF
C5665 CLK2.t66 GND 0.03fF
C5666 CLK2.t98 GND 0.03fF
C5667 CLK2.n859 GND 0.08fF $ **FLOATING
C5668 EESPFAL_s0_0/EESPFAL_NAND_v3_1/CLK GND 0.01fF $ **FLOATING
C5669 CLK2.t100 GND 0.04fF
C5670 CLK2.t19 GND 0.03fF
C5671 CLK2.t80 GND 0.03fF
C5672 CLK2.n860 GND 0.11fF $ **FLOATING
C5673 CLK2.n861 GND 0.05fF $ **FLOATING
C5674 CLK2.n862 GND 0.02fF $ **FLOATING
C5675 CLK2.n863 GND 0.02fF $ **FLOATING
C5676 CLK2.n864 GND 0.09fF $ **FLOATING
C5677 CLK2.n865 GND 0.04fF $ **FLOATING
C5678 CLK2.n866 GND 0.02fF $ **FLOATING
C5679 CLK2.n867 GND 0.02fF $ **FLOATING
C5680 CLK2.n868 GND 0.05fF $ **FLOATING
C5681 CLK2.n869 GND 0.14fF $ **FLOATING
C5682 CLK2.n870 GND 0.04fF $ **FLOATING
C5683 CLK2.n871 GND 0.02fF $ **FLOATING
C5684 CLK2.n872 GND 0.02fF $ **FLOATING
C5685 CLK2.n873 GND 0.02fF $ **FLOATING
C5686 CLK2.n874 GND 0.04fF $ **FLOATING
C5687 CLK2.n875 GND 0.02fF $ **FLOATING
C5688 CLK2.n876 GND 0.02fF $ **FLOATING
C5689 CLK2.n877 GND 0.02fF $ **FLOATING
C5690 CLK2.n878 GND 0.10fF $ **FLOATING
C5691 CLK2.n879 GND 0.02fF $ **FLOATING
C5692 CLK2.n880 GND 0.02fF $ **FLOATING
C5693 CLK2.n881 GND 0.02fF $ **FLOATING
C5694 CLK2.n882 GND 0.13fF $ **FLOATING
C5695 CLK2.n883 GND 0.02fF $ **FLOATING
C5696 CLK2.n884 GND 0.02fF $ **FLOATING
C5697 CLK2.n885 GND 0.01fF $ **FLOATING
C5698 CLK2.n886 GND 0.21fF $ **FLOATING
C5699 CLK2.t99 GND 0.06fF
C5700 CLK2.n887 GND 0.08fF $ **FLOATING
C5701 CLK2.n888 GND 0.02fF $ **FLOATING
C5702 CLK2.n889 GND 0.02fF $ **FLOATING
C5703 CLK2.n890 GND 0.02fF $ **FLOATING
C5704 CLK2.n891 GND 0.12fF $ **FLOATING
C5705 CLK2.n892 GND 0.02fF $ **FLOATING
C5706 CLK2.n893 GND 0.02fF $ **FLOATING
C5707 CLK2.n894 GND 0.02fF $ **FLOATING
C5708 CLK2.n895 GND 0.02fF $ **FLOATING
C5709 CLK2.t97 GND 0.06fF
C5710 CLK2.n896 GND 0.07fF $ **FLOATING
C5711 CLK2.n897 GND 0.02fF $ **FLOATING
C5712 CLK2.n898 GND 0.02fF $ **FLOATING
C5713 CLK2.n899 GND 0.12fF $ **FLOATING
C5714 CLK2.n900 GND 0.02fF $ **FLOATING
C5715 CLK2.n901 GND 0.02fF $ **FLOATING
C5716 CLK2.n902 GND 0.13fF $ **FLOATING
C5717 CLK2.t65 GND 0.06fF
C5718 CLK2.n903 GND 0.07fF $ **FLOATING
C5719 CLK2.n904 GND 0.02fF $ **FLOATING
C5720 CLK2.n905 GND 0.02fF $ **FLOATING
C5721 CLK2.n906 GND 0.02fF $ **FLOATING
C5722 CLK2.n907 GND 0.12fF $ **FLOATING
C5723 CLK2.n908 GND 0.02fF $ **FLOATING
C5724 CLK2.n909 GND 0.02fF $ **FLOATING
C5725 CLK2.n910 GND 0.02fF $ **FLOATING
C5726 CLK2.t63 GND 0.06fF
C5727 CLK2.n911 GND 0.08fF $ **FLOATING
C5728 CLK2.n912 GND 0.02fF $ **FLOATING
C5729 CLK2.n913 GND 0.02fF $ **FLOATING
C5730 CLK2.n914 GND 0.02fF $ **FLOATING
C5731 CLK2.n915 GND 0.21fF $ **FLOATING
C5732 CLK2.n916 GND 0.13fF $ **FLOATING
C5733 CLK2.n917 GND 0.02fF $ **FLOATING
C5734 CLK2.n918 GND 0.02fF $ **FLOATING
C5735 CLK2.n919 GND 0.01fF $ **FLOATING
C5736 CLK2.n920 GND 0.10fF $ **FLOATING
C5737 CLK2.n921 GND 0.02fF $ **FLOATING
C5738 CLK2.n922 GND 0.02fF $ **FLOATING
C5739 CLK2.n923 GND 0.02fF $ **FLOATING
C5740 CLK2.n924 GND 0.04fF $ **FLOATING
C5741 CLK2.n925 GND 0.02fF $ **FLOATING
C5742 CLK2.n926 GND 0.02fF $ **FLOATING
C5743 CLK2.n927 GND 0.02fF $ **FLOATING
C5744 CLK2.n928 GND 0.04fF $ **FLOATING
C5745 CLK2.n929 GND 0.02fF $ **FLOATING
C5746 CLK2.n930 GND 0.02fF $ **FLOATING
C5747 CLK2.n931 GND 0.02fF $ **FLOATING
C5748 CLK2.n932 GND 0.04fF $ **FLOATING
C5749 CLK2.n933 GND 0.02fF $ **FLOATING
C5750 CLK2.n934 GND 0.02fF $ **FLOATING
C5751 CLK2.n935 GND 0.02fF $ **FLOATING
C5752 CLK2.n936 GND 0.05fF $ **FLOATING
C5753 CLK2.n937 GND 0.02fF $ **FLOATING
C5754 CLK2.n938 GND 0.02fF $ **FLOATING
C5755 CLK2.n939 GND 0.02fF $ **FLOATING
C5756 CLK2.n940 GND 0.06fF $ **FLOATING
C5757 CLK2.n941 GND 0.02fF $ **FLOATING
C5758 CLK2.n942 GND 0.06fF $ **FLOATING
C5759 CLK2.n943 GND 0.02fF $ **FLOATING
C5760 CLK2.n944 GND 0.01fF $ **FLOATING
C5761 CLK2.t53 GND 0.03fF
C5762 CLK2.n945 GND 0.08fF $ **FLOATING
C5763 CLK2.n946 GND 0.01fF $ **FLOATING
C5764 CLK2.n947 GND 0.11fF $ **FLOATING
C5765 CLK2.n948 GND 0.12fF $ **FLOATING
C5766 CLK2.t88 GND 0.03fF
C5767 CLK2.t105 GND 0.03fF
C5768 CLK2.n949 GND 0.05fF $ **FLOATING
C5769 CLK2.n950 GND 0.01fF $ **FLOATING
C5770 CLK2.n951 GND 0.02fF $ **FLOATING
C5771 CLK2.n952 GND 0.02fF $ **FLOATING
C5772 CLK2.n953 GND 0.06fF $ **FLOATING
C5773 CLK2.n954 GND 0.05fF $ **FLOATING
C5774 CLK2.n955 GND 0.02fF $ **FLOATING
C5775 CLK2.n956 GND 0.02fF $ **FLOATING
C5776 CLK2.n957 GND 0.09fF $ **FLOATING
C5777 CLK2.n958 GND 0.05fF $ **FLOATING
C5778 CLK2.n959 GND 0.04fF $ **FLOATING
C5779 CLK2.n960 GND 0.02fF $ **FLOATING
C5780 CLK2.n961 GND 0.01fF $ **FLOATING
C5781 CLK2.n962 GND 0.01fF $ **FLOATING
C5782 CLK2.n963 GND 0.00fF $ **FLOATING
C5783 CLK2.n964 GND 0.04fF $ **FLOATING
C5784 CLK2.n965 GND 0.00fF $ **FLOATING
C5785 EESPFAL_s0_0/CLK2 GND 0.01fF $ **FLOATING
C5786 EESPFAL_s1_0/EESPFAL_INV4_0/OUT GND 0.23fF $ **FLOATING
C5787 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t8 GND 0.03fF
C5788 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n0 GND 0.63fF $ **FLOATING
C5789 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t3 GND 0.04fF
C5790 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t2 GND 0.04fF
C5791 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n1 GND 0.11fF $ **FLOATING
C5792 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t1 GND 0.04fF
C5793 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t4 GND 0.04fF
C5794 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n2 GND 0.13fF $ **FLOATING
C5795 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t0 GND 0.25fF
C5796 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n3 GND 0.17fF $ **FLOATING
C5797 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n4 GND 0.12fF $ **FLOATING
C5798 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t7 GND 0.06fF
C5799 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t6 GND 0.05fF
C5800 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.t5 GND 0.04fF
C5801 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n5 GND 0.06fF $ **FLOATING
C5802 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C_bar.n6 GND 0.04fF $ **FLOATING
C5803 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t7 GND 0.05fF
C5804 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t4 GND 0.04fF
C5805 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t3 GND 0.04fF
C5806 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n0 GND 0.12fF $ **FLOATING
C5807 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t1 GND 0.04fF
C5808 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t0 GND 0.04fF
C5809 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n1 GND 0.13fF $ **FLOATING
C5810 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t6 GND 0.06fF
C5811 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t5 GND 0.06fF
C5812 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t8 GND 0.03fF
C5813 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n2 GND 0.06fF $ **FLOATING
C5814 EESPFAL_s1_0/EESPFAL_INV4_0/OUT_bar GND 0.01fF $ **FLOATING
C5815 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n3 GND 0.03fF $ **FLOATING
C5816 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n4 GND 0.11fF $ **FLOATING
C5817 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n5 GND 0.11fF $ **FLOATING
C5818 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.t2 GND 0.16fF
C5819 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n6 GND 0.18fF $ **FLOATING
C5820 EESPFAL_s1_0/EESPFAL_3in_NOR_v2_0/C.n7 GND 0.77fF $ **FLOATING
.ends

