magic
tech sky130A
timestamp 1671243859
<< nmoslvt >>
rect 980 -115 995 885
rect 1055 -115 1070 885
rect 1130 -115 1145 885
rect 1205 -115 1220 885
rect 1280 -115 1295 885
rect 1355 -115 1370 885
rect 1430 -115 1445 885
rect 1505 -115 1520 885
rect 1580 -115 1595 885
rect 1655 -115 1670 885
<< ndiff >>
rect 920 865 980 885
rect 920 -95 940 865
rect 960 -95 980 865
rect 920 -115 980 -95
rect 995 865 1055 885
rect 995 -95 1015 865
rect 1035 -95 1055 865
rect 995 -115 1055 -95
rect 1070 865 1130 885
rect 1070 -95 1090 865
rect 1110 -95 1130 865
rect 1070 -115 1130 -95
rect 1145 865 1205 885
rect 1145 -95 1165 865
rect 1185 -95 1205 865
rect 1145 -115 1205 -95
rect 1220 865 1280 885
rect 1220 -95 1240 865
rect 1260 -95 1280 865
rect 1220 -115 1280 -95
rect 1295 865 1355 885
rect 1295 -95 1315 865
rect 1335 -95 1355 865
rect 1295 -115 1355 -95
rect 1370 865 1430 885
rect 1370 -95 1390 865
rect 1410 -95 1430 865
rect 1370 -115 1430 -95
rect 1445 865 1505 885
rect 1445 -95 1465 865
rect 1485 -95 1505 865
rect 1445 -115 1505 -95
rect 1520 865 1580 885
rect 1520 -95 1540 865
rect 1560 -95 1580 865
rect 1520 -115 1580 -95
rect 1595 865 1655 885
rect 1595 -95 1615 865
rect 1635 -95 1655 865
rect 1595 -115 1655 -95
rect 1670 865 1730 885
rect 1670 -95 1690 865
rect 1710 -95 1730 865
rect 1670 -115 1730 -95
<< ndiffc >>
rect 940 -95 960 865
rect 1015 -95 1035 865
rect 1090 -95 1110 865
rect 1165 -95 1185 865
rect 1240 -95 1260 865
rect 1315 -95 1335 865
rect 1390 -95 1410 865
rect 1465 -95 1485 865
rect 1540 -95 1560 865
rect 1615 -95 1635 865
rect 1690 -95 1710 865
<< psubdiff >>
rect 860 865 920 885
rect 860 -95 880 865
rect 900 -95 920 865
rect 860 -115 920 -95
<< psubdiffcont >>
rect 880 -95 900 865
<< poly >>
rect 980 900 1670 915
rect 980 885 995 900
rect 1055 885 1070 900
rect 1130 885 1145 900
rect 1205 885 1220 900
rect 1280 885 1295 900
rect 1355 885 1370 900
rect 1430 885 1445 900
rect 1505 885 1520 900
rect 1580 885 1595 900
rect 1655 885 1670 900
rect 980 -130 995 -115
rect 1055 -130 1070 -115
rect 1130 -130 1145 -115
rect 1205 -130 1220 -115
rect 1280 -130 1295 -115
rect 1355 -130 1370 -115
rect 1430 -130 1445 -115
rect 1505 -130 1520 -115
rect 1580 -130 1595 -115
rect 1655 -130 1670 -115
<< locali >>
rect 1015 895 1635 915
rect 1015 875 1035 895
rect 1165 875 1185 895
rect 1315 875 1335 895
rect 1465 875 1485 895
rect 1615 875 1635 895
rect 870 865 970 875
rect 870 -95 880 865
rect 900 -95 940 865
rect 960 -95 970 865
rect 870 -105 970 -95
rect 1005 865 1045 875
rect 1005 -95 1015 865
rect 1035 -95 1045 865
rect 1005 -105 1045 -95
rect 1080 865 1120 875
rect 1080 -95 1090 865
rect 1110 -95 1120 865
rect 1080 -105 1120 -95
rect 1155 865 1195 875
rect 1155 -95 1165 865
rect 1185 -95 1195 865
rect 1155 -105 1195 -95
rect 1230 865 1270 875
rect 1230 -95 1240 865
rect 1260 -95 1270 865
rect 1230 -105 1270 -95
rect 1305 865 1345 875
rect 1305 -95 1315 865
rect 1335 -95 1345 865
rect 1305 -105 1345 -95
rect 1380 865 1420 875
rect 1380 -95 1390 865
rect 1410 -95 1420 865
rect 1380 -105 1420 -95
rect 1455 865 1495 875
rect 1455 -95 1465 865
rect 1485 -95 1495 865
rect 1455 -105 1495 -95
rect 1530 865 1570 875
rect 1530 -95 1540 865
rect 1560 -95 1570 865
rect 1530 -105 1570 -95
rect 1605 865 1645 875
rect 1605 -95 1615 865
rect 1635 -95 1645 865
rect 1605 -105 1645 -95
rect 1680 865 1720 875
rect 1680 -95 1690 865
rect 1710 -95 1720 865
rect 1680 -105 1720 -95
rect 940 -125 960 -105
rect 1090 -125 1110 -105
rect 1240 -125 1260 -105
rect 1390 -125 1410 -105
rect 1540 -125 1560 -105
rect 1690 -125 1710 -105
rect 940 -145 1710 -125
<< end >>
