* NGSPICE file created from CMOS_sbox_flat.ext - technology: sky130A

.subckt CMOS_sbox_flat x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar GND s0 s1 s2 s3 VDD
X0 a_275_n6086# CMOS_s2_0/CMOS_4in_AND_0/OUT.t2 a_575_n6996# VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X1 a_n787_n2858# x3.t0 GND.t64 GND.t63 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n432_n5418# x0_bar.t0 CMOS_s2_0/CMOS_XOR_0/XOR GND.t73 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 CMOS_s2_0/CMOS_3in_OR_0/B a_425_n4808# VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X4 s1.t1 a_275_n2858# VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X5 a_275_n9314# CMOS_s3_0/CMOS_3in_OR_0/B GND.t117 GND.t116 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X6 CMOS_s0_0/CMOS_AND_0/AND a_425_1648# GND.t90 GND.t87 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n2290_370# x3.t1 GND.t62 GND.t61 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 CMOS_s2_0/CMOS_XOR_0/XOR x0.t0 a_n732_n5418# GND.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X9 a_n2345_n6996# x3_bar.t0 a_n2045_n6086# GND.t69 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X10 a_n2495_n10224# x2_bar.t0 a_n2195_n9314# GND.t127 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X11 CMOS_s1_0/CMOS_3in_OR_0/A a_n787_n3768# GND.t93 GND.t92 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_n2345_n6996# x2.t0 VDD.t115 VDD.t114 sky130_fd_pr__pfet_01v8 ad=3.6e+12p pd=1.44e+07u as=0p ps=0u w=3e+06u l=150000u
X13 CMOS_s2_0/CMOS_3in_OR_0/B a_425_n4808# GND.t105 GND.t104 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_425_n4808# x2_bar.t1 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X15 a_n2195_n9314# x0.t1 a_n2345_n9314# GND.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X16 VDD.t65 CMOS_s2_0/CMOS_XOR_0/XOR a_425_n4808# VDD.t64 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X17 a_n787_n10224# CMOS_s3_0/CMOS_AND_1/A a_n787_n9314# GND.t81 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X18 a_n1990_n4808# x3_bar.t1 a_n2140_n5418# VDD.t45 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X19 CMOS_s0_0/CMOS_XOR_0/XOR x0.t2 a_n2290_1648# VDD.t39 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X20 CMOS_s1_0/CMOS_3in_OR_0/C.t0 a_n2495_n3768# GND.t51 GND.t50 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X21 a_n2290_1648# x3_bar.t2 VDD.t143 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X22 a_n787_1038# x2_bar.t2 a_n787_1648# VDD.t18 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X23 a_n787_n9314# x3_bar.t3 GND.t136 GND.t135 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X24 a_n787_1648# x1.t0 VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X25 a_425_n5418# x2_bar.t3 GND.t9 GND.t2 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X26 a_275_n9314# CMOS_s3_0/CMOS_3in_OR_0/C.t2 a_575_n10224# VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X27 CMOS_s2_0/CMOS_4in_AND_0/OUT.t0 a_n2345_n6996# GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X28 CMOS_s0_0/CMOS_AND_0/B a_n787_1038# GND.t49 GND.t35 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X29 a_425_n540# CMOS_s0_0/CMOS_AND_1/A a_425_370# GND.t11 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X30 a_n732_n1580# x3_bar.t4 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X31 a_425_n4808# CMOS_s2_0/CMOS_XOR_0/XOR a_425_n5418# GND.t12 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X32 VDD.t44 x3.t2 a_n2495_n10224# VDD.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X33 VDD.t38 x0.t3 a_n432_n4808# VDD.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X34 a_n1990_n5418# x2_bar.t4 a_n2140_n5418# GND.t99 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X35 VDD.t96 x2.t1 a_n1990_n4808# VDD.t95 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X36 s1.t0 a_275_n2858# GND.t75 GND.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X37 a_n1990_1038# x3_bar.t5 CMOS_s0_0/CMOS_XOR_0/XOR GND.t40 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X38 a_n2140_n540# x3.t3 a_n2290_n540# VDD.t30 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X39 CMOS_s0_0/CMOS_AND_1/AND a_425_n540# GND.t88 GND.t87 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X40 a_425_n10224# CMOS_s3_0/CMOS_3in_OR_0/A VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X41 CMOS_s3_0/CMOS_3in_OR_0/A a_n787_n10224# GND.t80 GND.t79 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X42 a_n2290_n540# x0_bar.t1 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X43 s0.t1 a_1637_1038# VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X44 VDD.t94 x2.t2 a_n787_n540# VDD.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X45 a_425_n6996# CMOS_s2_0/CMOS_3in_OR_0/A VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X46 a_n787_n540# x1_bar.t0 VDD.t103 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X47 GND.t122 CMOS_s2_0/CMOS_4in_AND_0/OUT.t3 a_275_n6086# GND.t121 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X48 a_n732_n2190# x1.t1 GND.t24 GND.t23 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X49 VDD.t57 x2_bar.t5 a_n2495_n10224# VDD.t56 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X50 a_575_n6996# CMOS_s2_0/CMOS_3in_OR_0/B a_425_n6996# VDD.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X51 a_n787_370# x1_bar.t1 GND.t67 GND.t65 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X52 GND.t119 x1_bar.t2 a_n432_n5418# GND.t118 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X53 CMOS_s3_0/CMOS_3in_OR_0/C.t0 a_n2495_n10224# GND.t83 GND.t82 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X54 GND.t126 x3_bar.t6 a_n1990_n5418# GND.t125 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X55 a_275_n2858# CMOS_s1_0/CMOS_3in_OR_0/C.t2 a_575_n3768# VDD.t129 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X56 a_425_1648# CMOS_s0_0/CMOS_AND_0/B VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X57 a_1637_1648# CMOS_s0_0/CMOS_AND_0/AND VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X58 VDD.t107 CMOS_s0_0/CMOS_XOR_0/XOR a_425_1648# VDD.t106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X59 a_n2140_n540# x0.t4 a_n2290_370# GND.t60 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X60 a_n2345_n6996# x1.t2 VDD.t92 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X61 CMOS_s3_0/CMOS_3in_OR_0/A a_n787_n10224# VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X62 VDD.t71 CMOS_s3_0/CMOS_AND_1/A a_n787_n10224# VDD.t70 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X63 a_n732_n8036# x3_bar.t7 VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X64 a_n2345_n6086# x2.t3 GND.t96 GND.t95 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X65 s3.t1 a_275_n9314# VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X66 a_n2140_n2190# x0.t5 a_n2290_n1580# VDD.t30 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X67 s3.t0 a_275_n9314# GND.t107 GND.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X68 VDD.t28 x0.t6 a_n2345_n6996# VDD.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X69 a_n732_n8646# x2.t4 GND.t98 GND.t97 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X70 VDD.t132 x0_bar.t2 a_n2495_n3768# VDD.t131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X71 VDD.t124 CMOS_s2_0/CMOS_AND_1/A a_n787_n6996# VDD.t123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X72 a_n2290_n1580# x2_bar.t6 VDD.t90 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X73 a_425_n540# CMOS_s0_0/CMOS_AND_1/B VDD.t118 VDD.t104 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X74 a_n787_n6996# x1_bar.t3 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X75 VDD.t8 CMOS_s0_0/CMOS_AND_1/A a_425_n540# VDD.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X76 CMOS_s1_0/CMOS_AND_1/A a_n2140_n2190# VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X77 a_n432_n1580# x1_bar.t4 CMOS_s1_0/CMOS_XOR_0/XOR VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X78 a_n2140_n2190# x2.t5 a_n2290_n2190# GND.t111 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X79 CMOS_s0_0/CMOS_XOR_0/XOR x3.t4 a_n2290_1038# GND.t60 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X80 GND.t19 x3_bar.t8 a_n1990_370# GND.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X81 a_n2290_1038# x0.t7 GND.t139 GND.t61 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X82 CMOS_s1_0/CMOS_XOR_0/XOR x1.t3 a_n732_n1580# VDD.t99 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X83 GND.t72 x2_bar.t7 a_n787_1038# GND.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X84 CMOS_s0_0/CMOS_AND_1/B a_n2140_n540# GND.t47 GND.t46 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X85 a_425_370# CMOS_s0_0/CMOS_AND_1/B GND.t108 GND.t44 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X86 a_n787_1038# x1.t4 GND.t66 GND.t65 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X87 a_n2290_n2190# x0.t8 GND.t30 GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X88 VDD.t17 x3.t5 a_n1990_1648# VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X89 CMOS_s1_0/CMOS_AND_1/A a_n2140_n2190# GND.t26 GND.t25 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X90 CMOS_s2_0/CMOS_3in_OR_0/A a_n787_n6996# VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X91 GND.t115 CMOS_s1_0/CMOS_3in_OR_0/C.t3 a_275_n2858# GND.t114 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X92 GND.t3 CMOS_s2_0/CMOS_3in_OR_0/A a_275_n6086# GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X93 CMOS_s1_0/CMOS_3in_OR_0/B a_425_n1580# VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X94 a_n432_n2190# x3_bar.t9 CMOS_s1_0/CMOS_XOR_0/XOR GND.t20 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X95 a_n2140_n8646# x1.t5 a_n2290_n8036# VDD.t35 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X96 CMOS_s0_0/CMOS_AND_1/A a_n787_n540# GND.t36 GND.t35 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X97 a_275_n6086# CMOS_s2_0/CMOS_3in_OR_0/B GND.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X98 CMOS_s1_0/CMOS_XOR_0/XOR x3.t6 a_n732_n2190# GND.t59 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X99 a_425_n3768# CMOS_s1_0/CMOS_3in_OR_0/A VDD.t80 VDD.t79 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X100 a_n2290_n8036# x0_bar.t3 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X101 a_1637_1038# CMOS_s0_0/CMOS_AND_1/AND a_1637_1648# VDD.t36 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X102 a_n2140_n8646# x0.t9 a_n2290_n8646# GND.t103 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X103 CMOS_s3_0/CMOS_AND_1/A a_n2140_n8646# VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X104 s0.t0 a_1637_1038# GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X105 a_n787_n540# x2.t6 a_n787_370# GND.t71 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X106 a_575_n3768# CMOS_s1_0/CMOS_3in_OR_0/B a_425_n3768# VDD.t134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X107 VDD.t148 x0.t10 a_n1990_n540# VDD.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X108 a_n2290_n8646# x1.t6 GND.t129 GND.t128 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X109 a_n2345_n2858# x0_bar.t4 GND.t131 GND.t130 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X110 a_n432_n8036# x2_bar.t8 CMOS_s3_0/CMOS_XOR_0/XOR VDD.t89 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X111 a_n2045_n6086# x1.t7 a_n2195_n6086# GND.t102 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X112 a_n732_n4808# x0_bar.t5 VDD.t150 VDD.t149 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X113 a_425_n1580# x2_bar.t9 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X114 CMOS_s1_0/CMOS_3in_OR_0/B a_425_n1580# GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X115 CMOS_s3_0/CMOS_AND_1/A a_n2140_n8646# GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X116 a_575_n10224# CMOS_s3_0/CMOS_3in_OR_0/B a_425_n10224# VDD.t133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X117 a_n432_n8646# x3_bar.t10 CMOS_s3_0/CMOS_XOR_0/XOR GND.t8 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X118 CMOS_s3_0/CMOS_XOR_0/XOR x2.t7 a_n732_n8036# VDD.t130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X119 a_n2195_n6086# x0.t11 a_n2345_n6086# GND.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X120 CMOS_s0_0/CMOS_AND_0/AND a_425_1648# VDD.t82 VDD.t81 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X121 VDD.t122 CMOS_s1_0/CMOS_XOR_0/XOR a_425_n1580# VDD.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X122 VDD.t63 x3_bar.t11 a_n2495_n3768# VDD.t62 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X123 s2.t1 a_275_n6086# VDD.t137 VDD.t136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X124 a_425_1038# CMOS_s0_0/CMOS_AND_0/B GND.t45 GND.t44 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X125 a_1637_1038# CMOS_s0_0/CMOS_AND_0/AND GND.t85 GND.t84 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X126 a_n2495_n10224# x0.t12 VDD.t141 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X127 a_n787_n6996# CMOS_s2_0/CMOS_AND_1/A a_n787_n6086# GND.t113 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X128 a_425_1648# CMOS_s0_0/CMOS_XOR_0/XOR a_425_1038# GND.t11 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X129 a_n1990_n1580# x0_bar.t6 a_n2140_n2190# VDD.t40 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X130 GND.t77 CMOS_s3_0/CMOS_3in_OR_0/C.t3 a_275_n9314# GND.t76 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X131 CMOS_s3_0/CMOS_XOR_0/XOR x3.t7 a_n732_n8646# GND.t58 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X132 a_n2495_n3768# x1.t8 VDD.t155 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X133 CMOS_s3_0/CMOS_3in_OR_0/B a_425_n8036# VDD.t120 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X134 a_n787_n6086# x1_bar.t5 GND.t34 GND.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X135 a_n732_n5418# x1.t9 GND.t101 GND.t100 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X136 a_425_n2190# x2_bar.t10 GND.t22 GND.t21 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X137 VDD.t77 CMOS_s1_0/CMOS_AND_1/A a_n787_n3768# VDD.t76 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X138 CMOS_s3_0/CMOS_3in_OR_0/B a_425_n8036# GND.t110 GND.t109 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X139 a_425_n1580# CMOS_s1_0/CMOS_XOR_0/XOR a_425_n2190# GND.t112 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X140 a_n787_n3768# x3.t8 VDD.t113 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X141 CMOS_s0_0/CMOS_AND_1/AND a_425_n540# VDD.t78 VDD.t10 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X142 VDD.t86 x3.t9 a_n432_n1580# VDD.t85 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X143 a_n787_n10224# x3_bar.t12 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X144 VDD.t88 x3_bar.t13 a_n2345_n6996# VDD.t87 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X145 VDD.t117 x2.t8 a_n1990_n1580# VDD.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X146 a_n1990_n2190# x2_bar.t11 a_n2140_n2190# GND.t70 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X147 a_n2345_n9314# x3.t10 GND.t57 GND.t56 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X148 a_425_n8036# x1.t10 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X149 CMOS_s2_0/CMOS_3in_OR_0/A a_n787_n6996# GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X150 GND.t89 CMOS_s1_0/CMOS_3in_OR_0/A a_275_n2858# GND.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X151 CMOS_s0_0/CMOS_AND_0/B a_n787_1038# VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X152 a_n2140_n5418# x3.t11 a_n2290_n4808# VDD.t53 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X153 VDD.t147 CMOS_s3_0/CMOS_XOR_0/XOR a_425_n8036# VDD.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X154 a_275_n2858# CMOS_s1_0/CMOS_3in_OR_0/B GND.t120 GND.t112 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X155 a_425_n8646# x1.t11 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X156 CMOS_s1_0/CMOS_3in_OR_0/A a_n787_n3768# VDD.t84 VDD.t83 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X157 CMOS_s3_0/CMOS_3in_OR_0/C.t1 a_n2495_n10224# VDD.t73 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X158 CMOS_s0_0/CMOS_AND_1/B a_n2140_n540# VDD.t46 VDD.t19 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X159 GND.t138 x1_bar.t6 a_n432_n2190# GND.t137 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X160 a_n1990_n8036# x1_bar.t7 a_n2140_n8646# VDD.t26 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X161 a_n2290_n4808# x2_bar.t12 VDD.t98 VDD.t97 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X162 GND.t134 x0_bar.t7 a_n1990_n2190# GND.t133 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X163 a_425_n8036# CMOS_s3_0/CMOS_XOR_0/XOR a_425_n8646# GND.t116 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X164 CMOS_s2_0/CMOS_AND_1/A a_n2140_n5418# VDD.t52 VDD.t51 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X165 a_n1990_1648# x0_bar.t8 CMOS_s0_0/CMOS_XOR_0/XOR VDD.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X166 GND.t91 x0_bar.t9 a_n1990_1038# GND.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X167 CMOS_s2_0/CMOS_4in_AND_0/OUT.t1 a_n2345_n6996# VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X168 a_n1990_n8646# x0_bar.t10 a_n2140_n8646# GND.t41 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X169 a_n2495_n3768# x3_bar.t14 a_n2195_n2858# GND.t68 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X170 a_n432_n4808# x1_bar.t8 CMOS_s2_0/CMOS_XOR_0/XOR VDD.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X171 CMOS_s1_0/CMOS_3in_OR_0/C.t1 a_n2495_n3768# VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X172 a_n2140_n5418# x2.t9 a_n2290_n5418# GND.t94 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X173 a_n1990_370# x0_bar.t11 a_n2140_n540# GND.t40 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X174 CMOS_s0_0/CMOS_AND_1/A a_n787_n540# VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X175 a_n2195_n2858# x1.t12 a_n2345_n2858# GND.t132 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X176 VDD.t61 x3.t12 a_n432_n8036# VDD.t60 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X177 CMOS_s2_0/CMOS_XOR_0/XOR x1.t13 a_n732_n4808# VDD.t151 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X178 GND.t38 CMOS_s0_0/CMOS_AND_1/AND a_1637_1038# GND.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X179 VDD.t126 x0.t13 a_n1990_n8036# VDD.t125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X180 a_n2290_n5418# x3.t13 GND.t55 GND.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X181 s2.t0 a_275_n6086# GND.t124 GND.t123 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X182 a_n787_n3768# CMOS_s1_0/CMOS_AND_1/A a_n787_n2858# GND.t86 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X183 CMOS_s2_0/CMOS_AND_1/A a_n2140_n5418# GND.t53 GND.t52 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X184 a_n1990_n540# x3_bar.t15 a_n2140_n540# VDD.t40 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X185 GND.t78 CMOS_s3_0/CMOS_3in_OR_0/A a_275_n9314# GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X186 GND.t32 x2_bar.t13 a_n432_n8646# GND.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X187 GND.t43 x1_bar.t9 a_n1990_n8646# GND.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
R0 CMOS_s2_0/CMOS_4in_AND_0/OUT.t2 CMOS_s2_0/CMOS_4in_AND_0/OUT.t3 1221.07
R1 CMOS_s2_0/CMOS_3in_OR_0/C CMOS_s2_0/CMOS_4in_AND_0/OUT.n0 739.238
R2 CMOS_s2_0/CMOS_3in_OR_0/C CMOS_s2_0/CMOS_4in_AND_0/OUT.t2 633.02
R3 CMOS_s2_0/CMOS_4in_AND_0/OUT CMOS_s2_0/CMOS_4in_AND_0/OUT.t0 114.438
R4 CMOS_s2_0/CMOS_4in_AND_0/OUT.n0 CMOS_s2_0/CMOS_4in_AND_0/OUT 95.237
R5 CMOS_s2_0/CMOS_4in_AND_0/OUT.n0 CMOS_s2_0/CMOS_4in_AND_0/OUT.t1 45.156
R6 VDD.t125 VDD.t12 552.101
R7 VDD.n453 VDD.t51 535.897
R8 VDD.n480 VDD.t49 451.594
R9 VDD.n187 VDD.t119 371.739
R10 VDD.n369 VDD.t108 371.739
R11 VDD.t89 VDD.t60 206.521
R12 VDD.t130 VDD.t138 206.521
R13 VDD.t26 VDD.t35 206.521
R14 VDD.t35 VDD.t144 206.521
R15 VDD.t146 VDD.t152 206.521
R16 VDD.t29 VDD.t37 206.521
R17 VDD.t151 VDD.t149 206.521
R18 VDD.t62 VDD.t154 206.521
R19 VDD.t154 VDD.t131 206.521
R20 VDD.t64 VDD.t14 206.521
R21 VDD.t121 VDD.t85 206.521
R22 VDD.t99 VDD.t31 206.521
R23 VDD.n187 VDD.t146 165.217
R24 VDD.n369 VDD.t64 165.217
R25 VDD.n296 VDD.t26 112.898
R26 VDD.n230 VDD.t130 110.144
R27 VDD.n412 VDD.t151 110.144
R28 VDD.n582 VDD.t99 110.144
R29 VDD.n230 VDD.t89 96.376
R30 VDD.n412 VDD.t29 96.376
R31 VDD.n582 VDD.t121 96.376
R32 VDD.n296 VDD.t125 93.623
R33 VDD.n480 VDD.t62 85.362
R34 VDD.n454 VDD.n453 63.333
R35 VDD.n844 VDD.t39 38.206
R36 VDD.n494 VDD.t53 33.476
R37 VDD.n852 VDD.t142 32.01
R38 VDD.n834 VDD.t21 29.945
R39 VDD.n503 VDD.t97 28.047
R40 VDD.n188 VDD.n187 27.142
R41 VDD.n370 VDD.n369 27.142
R42 VDD.n808 VDD.t100 24.782
R43 VDD.n762 VDD.t41 24.782
R44 VDD.n715 VDD.t74 24.782
R45 VDD.n42 VDD.t66 24.782
R46 VDD.n89 VDD.t54 24.782
R47 VDD.n145 VDD.t43 24.782
R48 VDD.n231 VDD.n230 24.428
R49 VDD.n413 VDD.n412 24.428
R50 VDD.n583 VDD.n582 24.428
R51 VDD.n826 VDD.t16 23.75
R52 VDD.n207 VDD.t153 22.029
R53 VDD.n327 VDD.t145 22.029
R54 VDD.n290 VDD.t126 22.029
R55 VDD.n272 VDD.t13 22.029
R56 VDD.n252 VDD.t139 22.029
R57 VDD.n216 VDD.t61 22.029
R58 VDD.n185 VDD.t147 22.029
R59 VDD.n172 VDD.t120 22.029
R60 VDD.n389 VDD.t15 22.029
R61 VDD.n507 VDD.t98 22.029
R62 VDD.n471 VDD.t96 22.029
R63 VDD.n452 VDD.t52 22.029
R64 VDD.n434 VDD.t150 22.029
R65 VDD.n398 VDD.t38 22.029
R66 VDD.n367 VDD.t65 22.029
R67 VDD.n354 VDD.t109 22.029
R68 VDD.n525 VDD.t11 22.029
R69 VDD.n538 VDD.t122 22.029
R70 VDD.n559 VDD.t105 22.029
R71 VDD.n622 VDD.t20 22.029
R72 VDD.n639 VDD.t117 22.029
R73 VDD.n672 VDD.t90 22.029
R74 VDD.n604 VDD.t32 22.029
R75 VDD.n568 VDD.t86 22.029
R76 VDD.n856 VDD.t143 22.029
R77 VDD.n825 VDD.t17 22.029
R78 VDD.n816 VDD.t101 22.029
R79 VDD.n783 VDD.t48 22.029
R80 VDD.n770 VDD.t42 22.029
R81 VDD.n749 VDD.t107 22.029
R82 VDD.n736 VDD.t82 22.029
R83 VDD.n723 VDD.t75 22.029
R84 VDD.n690 VDD.t4 22.029
R85 VDD.n9 VDD.t111 22.029
R86 VDD.n50 VDD.t67 22.029
R87 VDD.n63 VDD.t69 22.029
R88 VDD.n76 VDD.t71 22.029
R89 VDD.n97 VDD.t55 22.029
R90 VDD.n110 VDD.t73 22.029
R91 VDD.n127 VDD.t57 22.029
R92 VDD.n163 VDD.t137 22.029
R93 VDD.n207 VDD.t2 22.029
R94 VDD.n221 VDD.t25 22.029
R95 VDD.n235 VDD.t124 22.029
R96 VDD.n257 VDD.t128 22.029
R97 VDD.n277 VDD.t6 22.029
R98 VDD.n295 VDD.t88 22.029
R99 VDD.n332 VDD.t115 22.029
R100 VDD.n345 VDD.t59 22.029
R101 VDD.n389 VDD.t80 22.029
R102 VDD.n403 VDD.t84 22.029
R103 VDD.n417 VDD.t77 22.029
R104 VDD.n439 VDD.t113 22.029
R105 VDD.n466 VDD.t50 22.029
R106 VDD.n485 VDD.t63 22.029
R107 VDD.n525 VDD.t78 22.029
R108 VDD.n538 VDD.t8 22.029
R109 VDD.n559 VDD.t118 22.029
R110 VDD.n573 VDD.t34 22.029
R111 VDD.n587 VDD.t94 22.029
R112 VDD.n609 VDD.t103 22.029
R113 VDD.n622 VDD.t46 22.029
R114 VDD.n639 VDD.t148 22.029
R115 VDD.n672 VDD.t23 22.029
R116 VDD.n248 VDD.t127 21.714
R117 VDD.n273 VDD.t5 21.714
R118 VDD.n323 VDD.t114 21.714
R119 VDD.n199 VDD.t1 21.714
R120 VDD.n430 VDD.t112 21.714
R121 VDD.n381 VDD.t79 21.714
R122 VDD.n600 VDD.t102 21.714
R123 VDD.n472 VDD.t95 20.809
R124 VDD.n660 VDD.t30 20.201
R125 VDD.n481 VDD.n480 19.904
R126 VDD.n0 VDD.t141 19.7
R127 VDD.n0 VDD.t44 19.7
R128 VDD.n309 VDD.t92 19.7
R129 VDD.n309 VDD.t28 19.7
R130 VDD.n336 VDD.t155 19.7
R131 VDD.n336 VDD.t132 19.7
R132 VDD.n800 VDD.t18 18.586
R133 VDD.n754 VDD.t106 18.586
R134 VDD.n707 VDD.t36 18.586
R135 VDD.n5 VDD.t110 18.586
R136 VDD.n34 VDD.t133 18.586
R137 VDD.n81 VDD.t70 18.586
R138 VDD.n106 VDD.t72 18.586
R139 VDD.n136 VDD.t140 18.586
R140 VDD.n668 VDD.t22 16.925
R141 VDD.n240 VDD.t123 16.285
R142 VDD.n315 VDD.t27 16.285
R143 VDD.n159 VDD.t136 16.285
R144 VDD.n191 VDD.t9 16.285
R145 VDD.n422 VDD.t76 16.285
R146 VDD.n341 VDD.t58 16.285
R147 VDD.n373 VDD.t134 16.285
R148 VDD.n592 VDD.t93 16.285
R149 VDD.n648 VDD.t40 15.833
R150 VDD.n551 VDD.t104 13.103
R151 VDD.n640 VDD.t116 12.557
R152 VDD.n779 VDD.t47 12.391
R153 VDD.n732 VDD.t81 12.391
R154 VDD.n686 VDD.t3 12.391
R155 VDD.n26 VDD.t0 12.391
R156 VDD.n59 VDD.t68 12.391
R157 VDD.n128 VDD.t56 12.391
R158 VDD.t87 VDD.n296 11.761
R159 VDD.n846 VDD.n843 11.52
R160 VDD.n802 VDD.n799 11.52
R161 VDD.n756 VDD.n753 11.52
R162 VDD.n709 VDD.n706 11.52
R163 VDD.n36 VDD.n33 11.52
R164 VDD.n83 VDD.n80 11.52
R165 VDD.n138 VDD.n135 11.52
R166 VDD.n217 VDD.t24 10.857
R167 VDD.n305 VDD.t91 10.857
R168 VDD.n181 VDD.t135 10.857
R169 VDD.n399 VDD.t83 10.857
R170 VDD.n363 VDD.t129 10.857
R171 VDD.n569 VDD.t33 10.857
R172 VDD.n543 VDD.t7 9.827
R173 VDD.n618 VDD.t19 9.827
R174 VDD.n3 VDD.n2 8.855
R175 VDD.n57 VDD.n56 8.855
R176 VDD.n104 VDD.n103 8.855
R177 VDD.n108 VDD.n107 8.855
R178 VDD.n107 VDD.n106 8.855
R179 VDD.n113 VDD.n112 8.855
R180 VDD.n112 VDD.n111 8.855
R181 VDD.n117 VDD.n116 8.855
R182 VDD.n116 VDD.n115 8.855
R183 VDD.n121 VDD.n120 8.855
R184 VDD.n120 VDD.n119 8.855
R185 VDD.n125 VDD.n124 8.855
R186 VDD.n124 VDD.n123 8.855
R187 VDD.n130 VDD.n129 8.855
R188 VDD.n129 VDD.n128 8.855
R189 VDD.n135 VDD.n134 8.855
R190 VDD.n134 VDD.n133 8.855
R191 VDD.n138 VDD.n137 8.855
R192 VDD.n137 VDD.n136 8.855
R193 VDD.n142 VDD.n141 8.855
R194 VDD.n141 VDD.n140 8.855
R195 VDD.n147 VDD.n146 8.855
R196 VDD.n146 VDD.n145 8.855
R197 VDD.n151 VDD.n150 8.855
R198 VDD.n61 VDD.n60 8.855
R199 VDD.n60 VDD.n59 8.855
R200 VDD.n66 VDD.n65 8.855
R201 VDD.n65 VDD.n64 8.855
R202 VDD.n70 VDD.n69 8.855
R203 VDD.n69 VDD.n68 8.855
R204 VDD.n74 VDD.n73 8.855
R205 VDD.n73 VDD.n72 8.855
R206 VDD.n80 VDD.n79 8.855
R207 VDD.n79 VDD.n78 8.855
R208 VDD.n83 VDD.n82 8.855
R209 VDD.n82 VDD.n81 8.855
R210 VDD.n87 VDD.n86 8.855
R211 VDD.n86 VDD.n85 8.855
R212 VDD.n91 VDD.n90 8.855
R213 VDD.n90 VDD.n89 8.855
R214 VDD.n95 VDD.n94 8.855
R215 VDD.n7 VDD.n6 8.855
R216 VDD.n6 VDD.n5 8.855
R217 VDD.n12 VDD.n11 8.855
R218 VDD.n11 VDD.n10 8.855
R219 VDD.n16 VDD.n15 8.855
R220 VDD.n15 VDD.n14 8.855
R221 VDD.n20 VDD.n19 8.855
R222 VDD.n19 VDD.n18 8.855
R223 VDD.n24 VDD.n23 8.855
R224 VDD.n23 VDD.n22 8.855
R225 VDD.n28 VDD.n27 8.855
R226 VDD.n27 VDD.n26 8.855
R227 VDD.n33 VDD.n32 8.855
R228 VDD.n32 VDD.n31 8.855
R229 VDD.n36 VDD.n35 8.855
R230 VDD.n35 VDD.n34 8.855
R231 VDD.n40 VDD.n39 8.855
R232 VDD.n39 VDD.n38 8.855
R233 VDD.n44 VDD.n43 8.855
R234 VDD.n43 VDD.n42 8.855
R235 VDD.n48 VDD.n47 8.855
R236 VDD.n262 VDD.n261 8.855
R237 VDD.n261 VDD.n260 8.855
R238 VDD.n157 VDD.n156 8.855
R239 VDD.n447 VDD.n446 8.855
R240 VDD.n339 VDD.n338 8.855
R241 VDD.n450 VDD.n449 8.855
R242 VDD.n684 VDD.n683 8.855
R243 VDD.n688 VDD.n687 8.855
R244 VDD.n687 VDD.n686 8.855
R245 VDD.n693 VDD.n692 8.855
R246 VDD.n692 VDD.n691 8.855
R247 VDD.n697 VDD.n696 8.855
R248 VDD.n696 VDD.n695 8.855
R249 VDD.n701 VDD.n700 8.855
R250 VDD.n700 VDD.n699 8.855
R251 VDD.n706 VDD.n705 8.855
R252 VDD.n705 VDD.n704 8.855
R253 VDD.n709 VDD.n708 8.855
R254 VDD.n708 VDD.n707 8.855
R255 VDD.n713 VDD.n712 8.855
R256 VDD.n712 VDD.n711 8.855
R257 VDD.n717 VDD.n716 8.855
R258 VDD.n716 VDD.n715 8.855
R259 VDD.n721 VDD.n720 8.855
R260 VDD.n730 VDD.n729 8.855
R261 VDD.n734 VDD.n733 8.855
R262 VDD.n733 VDD.n732 8.855
R263 VDD.n739 VDD.n738 8.855
R264 VDD.n738 VDD.n737 8.855
R265 VDD.n743 VDD.n742 8.855
R266 VDD.n742 VDD.n741 8.855
R267 VDD.n747 VDD.n746 8.855
R268 VDD.n746 VDD.n745 8.855
R269 VDD.n753 VDD.n752 8.855
R270 VDD.n752 VDD.n751 8.855
R271 VDD.n756 VDD.n755 8.855
R272 VDD.n755 VDD.n754 8.855
R273 VDD.n760 VDD.n759 8.855
R274 VDD.n759 VDD.n758 8.855
R275 VDD.n764 VDD.n763 8.855
R276 VDD.n763 VDD.n762 8.855
R277 VDD.n768 VDD.n767 8.855
R278 VDD.n777 VDD.n776 8.855
R279 VDD.n781 VDD.n780 8.855
R280 VDD.n780 VDD.n779 8.855
R281 VDD.n786 VDD.n785 8.855
R282 VDD.n785 VDD.n784 8.855
R283 VDD.n790 VDD.n789 8.855
R284 VDD.n789 VDD.n788 8.855
R285 VDD.n794 VDD.n793 8.855
R286 VDD.n793 VDD.n792 8.855
R287 VDD.n799 VDD.n798 8.855
R288 VDD.n798 VDD.n797 8.855
R289 VDD.n802 VDD.n801 8.855
R290 VDD.n801 VDD.n800 8.855
R291 VDD.n806 VDD.n805 8.855
R292 VDD.n805 VDD.n804 8.855
R293 VDD.n810 VDD.n809 8.855
R294 VDD.n809 VDD.n808 8.855
R295 VDD.n814 VDD.n813 8.855
R296 VDD.n823 VDD.n822 8.855
R297 VDD.n828 VDD.n827 8.855
R298 VDD.n827 VDD.n826 8.855
R299 VDD.n832 VDD.n831 8.855
R300 VDD.n831 VDD.n830 8.855
R301 VDD.n836 VDD.n835 8.855
R302 VDD.n835 VDD.n834 8.855
R303 VDD.n840 VDD.n839 8.855
R304 VDD.n839 VDD.n838 8.855
R305 VDD.n843 VDD.n681 8.855
R306 VDD.n681 VDD.n680 8.855
R307 VDD.n846 VDD.n845 8.855
R308 VDD.n845 VDD.n844 8.855
R309 VDD.n850 VDD.n849 8.855
R310 VDD.n849 VDD.n848 8.855
R311 VDD.n854 VDD.n853 8.855
R312 VDD.n853 VDD.n852 8.855
R313 VDD.n859 VDD.n858 8.855
R314 VDD.n446 VDD.n445 7.349
R315 VDD.n521 VDD.t10 6.551
R316 VDD.n480 VDD.t45 6.333
R317 VDD.n242 VDD.n239 6.063
R318 VDD.n317 VDD.n314 6.063
R319 VDD.n193 VDD.n190 6.063
R320 VDD.n424 VDD.n421 6.063
R321 VDD.n496 VDD.n493 6.063
R322 VDD.n375 VDD.n372 6.063
R323 VDD.n545 VDD.n542 6.063
R324 VDD.n594 VDD.n591 6.063
R325 VDD.n662 VDD.n659 6.063
R326 VDD.n297 VDD.t87 5.428
R327 VDD.n335 VDD.n154 4.91
R328 VDD.n516 VDD.n335 4.775
R329 VDD.n679 VDD.n516 4.775
R330 VDD.n863 VDD.n679 4.775
R331 VDD.n154 VDD.n153 4.65
R332 VDD.n105 VDD.n104 4.65
R333 VDD.n109 VDD.n108 4.65
R334 VDD.n114 VDD.n113 4.65
R335 VDD.n118 VDD.n117 4.65
R336 VDD.n122 VDD.n121 4.65
R337 VDD.n126 VDD.n125 4.65
R338 VDD.n131 VDD.n130 4.65
R339 VDD.n135 VDD.n132 4.65
R340 VDD.n139 VDD.n138 4.65
R341 VDD.n143 VDD.n142 4.65
R342 VDD.n148 VDD.n147 4.65
R343 VDD.n152 VDD.n151 4.65
R344 VDD.n101 VDD.n100 4.65
R345 VDD.n99 VDD.n98 4.65
R346 VDD.n58 VDD.n57 4.65
R347 VDD.n62 VDD.n61 4.65
R348 VDD.n67 VDD.n66 4.65
R349 VDD.n71 VDD.n70 4.65
R350 VDD.n75 VDD.n74 4.65
R351 VDD.n80 VDD.n77 4.65
R352 VDD.n84 VDD.n83 4.65
R353 VDD.n88 VDD.n87 4.65
R354 VDD.n92 VDD.n91 4.65
R355 VDD.n96 VDD.n95 4.65
R356 VDD.n54 VDD.n53 4.65
R357 VDD.n52 VDD.n51 4.65
R358 VDD.n8 VDD.n7 4.65
R359 VDD.n13 VDD.n12 4.65
R360 VDD.n17 VDD.n16 4.65
R361 VDD.n21 VDD.n20 4.65
R362 VDD.n25 VDD.n24 4.65
R363 VDD.n29 VDD.n28 4.65
R364 VDD.n33 VDD.n30 4.65
R365 VDD.n37 VDD.n36 4.65
R366 VDD.n41 VDD.n40 4.65
R367 VDD.n45 VDD.n44 4.65
R368 VDD.n49 VDD.n48 4.65
R369 VDD.n263 VDD.n262 4.65
R370 VDD.n448 VDD.n447 4.65
R371 VDD.n451 VDD.n450 4.65
R372 VDD.n443 VDD.n442 4.65
R373 VDD.n689 VDD.n688 4.65
R374 VDD.n694 VDD.n693 4.65
R375 VDD.n698 VDD.n697 4.65
R376 VDD.n702 VDD.n701 4.65
R377 VDD.n706 VDD.n703 4.65
R378 VDD.n710 VDD.n709 4.65
R379 VDD.n714 VDD.n713 4.65
R380 VDD.n718 VDD.n717 4.65
R381 VDD.n722 VDD.n721 4.65
R382 VDD.n725 VDD.n724 4.65
R383 VDD.n727 VDD.n726 4.65
R384 VDD.n731 VDD.n730 4.65
R385 VDD.n735 VDD.n734 4.65
R386 VDD.n740 VDD.n739 4.65
R387 VDD.n744 VDD.n743 4.65
R388 VDD.n748 VDD.n747 4.65
R389 VDD.n753 VDD.n750 4.65
R390 VDD.n757 VDD.n756 4.65
R391 VDD.n761 VDD.n760 4.65
R392 VDD.n765 VDD.n764 4.65
R393 VDD.n769 VDD.n768 4.65
R394 VDD.n772 VDD.n771 4.65
R395 VDD.n774 VDD.n773 4.65
R396 VDD.n778 VDD.n777 4.65
R397 VDD.n782 VDD.n781 4.65
R398 VDD.n787 VDD.n786 4.65
R399 VDD.n791 VDD.n790 4.65
R400 VDD.n795 VDD.n794 4.65
R401 VDD.n799 VDD.n796 4.65
R402 VDD.n803 VDD.n802 4.65
R403 VDD.n807 VDD.n806 4.65
R404 VDD.n811 VDD.n810 4.65
R405 VDD.n815 VDD.n814 4.65
R406 VDD.n818 VDD.n817 4.65
R407 VDD.n820 VDD.n819 4.65
R408 VDD.n824 VDD.n823 4.65
R409 VDD.n829 VDD.n828 4.65
R410 VDD.n833 VDD.n832 4.65
R411 VDD.n837 VDD.n836 4.65
R412 VDD.n841 VDD.n840 4.65
R413 VDD.n843 VDD.n842 4.65
R414 VDD.n847 VDD.n846 4.65
R415 VDD.n851 VDD.n850 4.65
R416 VDD.n855 VDD.n854 4.65
R417 VDD.n860 VDD.n859 4.65
R418 VDD.n862 VDD.n861 4.65
R419 VDD.n266 VDD.n265 4.427
R420 VDD.n270 VDD.n269 4.427
R421 VDD.n275 VDD.n274 4.427
R422 VDD.n280 VDD.n279 4.427
R423 VDD.n284 VDD.n283 4.427
R424 VDD.n288 VDD.n287 4.427
R425 VDD.n293 VDD.n292 4.427
R426 VDD.n299 VDD.n298 4.427
R427 VDD.n303 VDD.n302 4.427
R428 VDD.n307 VDD.n306 4.427
R429 VDD.n314 VDD.n313 4.427
R430 VDD.n317 VDD.n316 4.427
R431 VDD.n321 VDD.n320 4.427
R432 VDD.n325 VDD.n324 4.427
R433 VDD.n330 VDD.n329 4.427
R434 VDD.n214 VDD.n213 4.427
R435 VDD.n219 VDD.n218 4.427
R436 VDD.n224 VDD.n223 4.427
R437 VDD.n228 VDD.n227 4.427
R438 VDD.n233 VDD.n232 4.427
R439 VDD.n239 VDD.n238 4.427
R440 VDD.n242 VDD.n241 4.427
R441 VDD.n246 VDD.n245 4.427
R442 VDD.n250 VDD.n249 4.427
R443 VDD.n255 VDD.n254 4.427
R444 VDD.n166 VDD.n165 4.427
R445 VDD.n170 VDD.n169 4.427
R446 VDD.n175 VDD.n174 4.427
R447 VDD.n179 VDD.n178 4.427
R448 VDD.n183 VDD.n182 4.427
R449 VDD.n190 VDD.n189 4.427
R450 VDD.n193 VDD.n192 4.427
R451 VDD.n197 VDD.n196 4.427
R452 VDD.n201 VDD.n200 4.427
R453 VDD.n205 VDD.n204 4.427
R454 VDD.n456 VDD.n455 4.427
R455 VDD.n460 VDD.n459 4.427
R456 VDD.n464 VDD.n463 4.427
R457 VDD.n469 VDD.n468 4.427
R458 VDD.n474 VDD.n473 4.427
R459 VDD.n478 VDD.n477 4.427
R460 VDD.n483 VDD.n482 4.427
R461 VDD.n488 VDD.n487 4.427
R462 VDD.n493 VDD.n492 4.427
R463 VDD.n496 VDD.n495 4.427
R464 VDD.n500 VDD.n499 4.427
R465 VDD.n505 VDD.n504 4.427
R466 VDD.n510 VDD.n509 4.427
R467 VDD.n396 VDD.n395 4.427
R468 VDD.n401 VDD.n400 4.427
R469 VDD.n406 VDD.n405 4.427
R470 VDD.n410 VDD.n409 4.427
R471 VDD.n415 VDD.n414 4.427
R472 VDD.n421 VDD.n420 4.427
R473 VDD.n424 VDD.n423 4.427
R474 VDD.n428 VDD.n427 4.427
R475 VDD.n432 VDD.n431 4.427
R476 VDD.n437 VDD.n436 4.427
R477 VDD.n348 VDD.n347 4.427
R478 VDD.n352 VDD.n351 4.427
R479 VDD.n357 VDD.n356 4.427
R480 VDD.n361 VDD.n360 4.427
R481 VDD.n365 VDD.n364 4.427
R482 VDD.n372 VDD.n371 4.427
R483 VDD.n375 VDD.n374 4.427
R484 VDD.n379 VDD.n378 4.427
R485 VDD.n383 VDD.n382 4.427
R486 VDD.n387 VDD.n386 4.427
R487 VDD.n616 VDD.n615 4.427
R488 VDD.n620 VDD.n619 4.427
R489 VDD.n625 VDD.n624 4.427
R490 VDD.n629 VDD.n628 4.427
R491 VDD.n633 VDD.n632 4.427
R492 VDD.n637 VDD.n636 4.427
R493 VDD.n642 VDD.n641 4.427
R494 VDD.n646 VDD.n645 4.427
R495 VDD.n650 VDD.n649 4.427
R496 VDD.n654 VDD.n653 4.427
R497 VDD.n659 VDD.n658 4.427
R498 VDD.n662 VDD.n661 4.427
R499 VDD.n666 VDD.n665 4.427
R500 VDD.n670 VDD.n669 4.427
R501 VDD.n675 VDD.n674 4.427
R502 VDD.n566 VDD.n565 4.427
R503 VDD.n571 VDD.n570 4.427
R504 VDD.n576 VDD.n575 4.427
R505 VDD.n580 VDD.n579 4.427
R506 VDD.n585 VDD.n584 4.427
R507 VDD.n591 VDD.n590 4.427
R508 VDD.n594 VDD.n593 4.427
R509 VDD.n598 VDD.n597 4.427
R510 VDD.n602 VDD.n601 4.427
R511 VDD.n607 VDD.n606 4.427
R512 VDD.n519 VDD.n518 4.427
R513 VDD.n523 VDD.n522 4.427
R514 VDD.n528 VDD.n527 4.427
R515 VDD.n532 VDD.n531 4.427
R516 VDD.n536 VDD.n535 4.427
R517 VDD.n542 VDD.n541 4.427
R518 VDD.n545 VDD.n544 4.427
R519 VDD.n549 VDD.n548 4.427
R520 VDD.n553 VDD.n552 4.427
R521 VDD.n557 VDD.n556 4.427
R522 VDD.n161 VDD.n160 4.427
R523 VDD.n160 VDD.n159 4.427
R524 VDD.n265 VDD.n264 4.427
R525 VDD.n269 VDD.n268 4.427
R526 VDD.n274 VDD.n273 4.427
R527 VDD.n279 VDD.n278 4.427
R528 VDD.n283 VDD.n282 4.427
R529 VDD.n287 VDD.n286 4.427
R530 VDD.n292 VDD.n291 4.427
R531 VDD.n298 VDD.n297 4.427
R532 VDD.n302 VDD.n301 4.427
R533 VDD.n306 VDD.n305 4.427
R534 VDD.n313 VDD.n312 4.427
R535 VDD.n316 VDD.n315 4.427
R536 VDD.n320 VDD.n319 4.427
R537 VDD.n324 VDD.n323 4.427
R538 VDD.n218 VDD.n217 4.427
R539 VDD.n223 VDD.n222 4.427
R540 VDD.n227 VDD.n226 4.427
R541 VDD.n232 VDD.n231 4.427
R542 VDD.n238 VDD.n237 4.427
R543 VDD.n241 VDD.n240 4.427
R544 VDD.n245 VDD.n244 4.427
R545 VDD.n249 VDD.n248 4.427
R546 VDD.n165 VDD.n164 4.427
R547 VDD.n169 VDD.n168 4.427
R548 VDD.n174 VDD.n173 4.427
R549 VDD.n178 VDD.n177 4.427
R550 VDD.n182 VDD.n181 4.427
R551 VDD.n189 VDD.n188 4.427
R552 VDD.n192 VDD.n191 4.427
R553 VDD.n196 VDD.n195 4.427
R554 VDD.n200 VDD.n199 4.427
R555 VDD.n514 VDD.n513 4.427
R556 VDD.n343 VDD.n342 4.427
R557 VDD.n342 VDD.n341 4.427
R558 VDD.n455 VDD.n454 4.427
R559 VDD.n459 VDD.n458 4.427
R560 VDD.n463 VDD.n462 4.427
R561 VDD.n468 VDD.n467 4.427
R562 VDD.n473 VDD.n472 4.427
R563 VDD.n477 VDD.n476 4.427
R564 VDD.n482 VDD.n481 4.427
R565 VDD.n487 VDD.n486 4.427
R566 VDD.n492 VDD.n491 4.427
R567 VDD.n495 VDD.n494 4.427
R568 VDD.n499 VDD.n498 4.427
R569 VDD.n504 VDD.n503 4.427
R570 VDD.n509 VDD.n508 4.427
R571 VDD.n513 VDD.n512 4.427
R572 VDD.n400 VDD.n399 4.427
R573 VDD.n405 VDD.n404 4.427
R574 VDD.n409 VDD.n408 4.427
R575 VDD.n414 VDD.n413 4.427
R576 VDD.n420 VDD.n419 4.427
R577 VDD.n423 VDD.n422 4.427
R578 VDD.n427 VDD.n426 4.427
R579 VDD.n431 VDD.n430 4.427
R580 VDD.n347 VDD.n346 4.427
R581 VDD.n351 VDD.n350 4.427
R582 VDD.n356 VDD.n355 4.427
R583 VDD.n360 VDD.n359 4.427
R584 VDD.n364 VDD.n363 4.427
R585 VDD.n371 VDD.n370 4.427
R586 VDD.n374 VDD.n373 4.427
R587 VDD.n378 VDD.n377 4.427
R588 VDD.n382 VDD.n381 4.427
R589 VDD.n619 VDD.n618 4.427
R590 VDD.n624 VDD.n623 4.427
R591 VDD.n628 VDD.n627 4.427
R592 VDD.n632 VDD.n631 4.427
R593 VDD.n636 VDD.n635 4.427
R594 VDD.n641 VDD.n640 4.427
R595 VDD.n645 VDD.n644 4.427
R596 VDD.n649 VDD.n648 4.427
R597 VDD.n653 VDD.n652 4.427
R598 VDD.n658 VDD.n657 4.427
R599 VDD.n661 VDD.n660 4.427
R600 VDD.n665 VDD.n664 4.427
R601 VDD.n669 VDD.n668 4.427
R602 VDD.n570 VDD.n569 4.427
R603 VDD.n575 VDD.n574 4.427
R604 VDD.n579 VDD.n578 4.427
R605 VDD.n584 VDD.n583 4.427
R606 VDD.n590 VDD.n589 4.427
R607 VDD.n593 VDD.n592 4.427
R608 VDD.n597 VDD.n596 4.427
R609 VDD.n601 VDD.n600 4.427
R610 VDD.n522 VDD.n521 4.427
R611 VDD.n527 VDD.n526 4.427
R612 VDD.n531 VDD.n530 4.427
R613 VDD.n535 VDD.n534 4.427
R614 VDD.n541 VDD.n540 4.427
R615 VDD.n544 VDD.n543 4.427
R616 VDD.n548 VDD.n547 4.427
R617 VDD.n552 VDD.n551 4.427
R618 VDD.n683 VDD.n682 4.288
R619 VDD.n729 VDD.n728 4.288
R620 VDD.n776 VDD.n775 4.288
R621 VDD.n822 VDD.n821 4.288
R622 VDD.n2 VDD.n1 4.288
R623 VDD.n56 VDD.n55 4.288
R624 VDD.n103 VDD.n102 4.288
R625 VDD.n150 VDD.n149 4.288
R626 VDD.n94 VDD.n93 4.288
R627 VDD.n47 VDD.n46 4.288
R628 VDD.n720 VDD.n719 4.288
R629 VDD.n767 VDD.n766 4.288
R630 VDD.n813 VDD.n812 4.288
R631 VDD.n858 VDD.n857 4.288
R632 VDD.n685 VDD.n684 2.562
R633 VDD.n4 VDD.n3 2.562
R634 VDD.n158 VDD.n157 2.562
R635 VDD.n340 VDD.n339 2.562
R636 VDD.n144 VDD.n0 2.329
R637 VDD.n310 VDD.n309 2.329
R638 VDD.n502 VDD.n336 2.329
R639 VDD.n334 VDD.n333 2.325
R640 VDD.n259 VDD.n258 2.325
R641 VDD.n267 VDD.n266 2.325
R642 VDD.n271 VDD.n270 2.325
R643 VDD.n276 VDD.n275 2.325
R644 VDD.n281 VDD.n280 2.325
R645 VDD.n285 VDD.n284 2.325
R646 VDD.n289 VDD.n288 2.325
R647 VDD.n294 VDD.n293 2.325
R648 VDD.n300 VDD.n299 2.325
R649 VDD.n304 VDD.n303 2.325
R650 VDD.n308 VDD.n307 2.325
R651 VDD.n314 VDD.n311 2.325
R652 VDD.n318 VDD.n317 2.325
R653 VDD.n322 VDD.n321 2.325
R654 VDD.n326 VDD.n325 2.325
R655 VDD.n331 VDD.n330 2.325
R656 VDD.n215 VDD.n214 2.325
R657 VDD.n220 VDD.n219 2.325
R658 VDD.n225 VDD.n224 2.325
R659 VDD.n229 VDD.n228 2.325
R660 VDD.n234 VDD.n233 2.325
R661 VDD.n239 VDD.n236 2.325
R662 VDD.n243 VDD.n242 2.325
R663 VDD.n247 VDD.n246 2.325
R664 VDD.n251 VDD.n250 2.325
R665 VDD.n256 VDD.n255 2.325
R666 VDD.n211 VDD.n210 2.325
R667 VDD.n167 VDD.n166 2.325
R668 VDD.n171 VDD.n170 2.325
R669 VDD.n176 VDD.n175 2.325
R670 VDD.n180 VDD.n179 2.325
R671 VDD.n184 VDD.n183 2.325
R672 VDD.n190 VDD.n186 2.325
R673 VDD.n194 VDD.n193 2.325
R674 VDD.n198 VDD.n197 2.325
R675 VDD.n202 VDD.n201 2.325
R676 VDD.n206 VDD.n205 2.325
R677 VDD.n209 VDD.n208 2.325
R678 VDD.n162 VDD.n161 2.325
R679 VDD.n515 VDD.n514 2.325
R680 VDD.n441 VDD.n440 2.325
R681 VDD.n457 VDD.n456 2.325
R682 VDD.n461 VDD.n460 2.325
R683 VDD.n465 VDD.n464 2.325
R684 VDD.n470 VDD.n469 2.325
R685 VDD.n475 VDD.n474 2.325
R686 VDD.n479 VDD.n478 2.325
R687 VDD.n484 VDD.n483 2.325
R688 VDD.n489 VDD.n488 2.325
R689 VDD.n493 VDD.n490 2.325
R690 VDD.n497 VDD.n496 2.325
R691 VDD.n501 VDD.n500 2.325
R692 VDD.n506 VDD.n505 2.325
R693 VDD.n511 VDD.n510 2.325
R694 VDD.n397 VDD.n396 2.325
R695 VDD.n402 VDD.n401 2.325
R696 VDD.n407 VDD.n406 2.325
R697 VDD.n411 VDD.n410 2.325
R698 VDD.n416 VDD.n415 2.325
R699 VDD.n421 VDD.n418 2.325
R700 VDD.n425 VDD.n424 2.325
R701 VDD.n429 VDD.n428 2.325
R702 VDD.n433 VDD.n432 2.325
R703 VDD.n438 VDD.n437 2.325
R704 VDD.n393 VDD.n392 2.325
R705 VDD.n349 VDD.n348 2.325
R706 VDD.n353 VDD.n352 2.325
R707 VDD.n358 VDD.n357 2.325
R708 VDD.n362 VDD.n361 2.325
R709 VDD.n366 VDD.n365 2.325
R710 VDD.n372 VDD.n368 2.325
R711 VDD.n376 VDD.n375 2.325
R712 VDD.n380 VDD.n379 2.325
R713 VDD.n384 VDD.n383 2.325
R714 VDD.n388 VDD.n387 2.325
R715 VDD.n391 VDD.n390 2.325
R716 VDD.n344 VDD.n343 2.325
R717 VDD.n678 VDD.n677 2.325
R718 VDD.n611 VDD.n610 2.325
R719 VDD.n561 VDD.n560 2.325
R720 VDD.n617 VDD.n616 2.325
R721 VDD.n621 VDD.n620 2.325
R722 VDD.n626 VDD.n625 2.325
R723 VDD.n630 VDD.n629 2.325
R724 VDD.n634 VDD.n633 2.325
R725 VDD.n638 VDD.n637 2.325
R726 VDD.n643 VDD.n642 2.325
R727 VDD.n647 VDD.n646 2.325
R728 VDD.n651 VDD.n650 2.325
R729 VDD.n655 VDD.n654 2.325
R730 VDD.n659 VDD.n656 2.325
R731 VDD.n663 VDD.n662 2.325
R732 VDD.n667 VDD.n666 2.325
R733 VDD.n671 VDD.n670 2.325
R734 VDD.n676 VDD.n675 2.325
R735 VDD.n613 VDD.n612 2.325
R736 VDD.n567 VDD.n566 2.325
R737 VDD.n572 VDD.n571 2.325
R738 VDD.n577 VDD.n576 2.325
R739 VDD.n581 VDD.n580 2.325
R740 VDD.n586 VDD.n585 2.325
R741 VDD.n591 VDD.n588 2.325
R742 VDD.n595 VDD.n594 2.325
R743 VDD.n599 VDD.n598 2.325
R744 VDD.n603 VDD.n602 2.325
R745 VDD.n608 VDD.n607 2.325
R746 VDD.n563 VDD.n562 2.325
R747 VDD.n524 VDD.n523 2.325
R748 VDD.n529 VDD.n528 2.325
R749 VDD.n533 VDD.n532 2.325
R750 VDD.n537 VDD.n536 2.325
R751 VDD.n542 VDD.n539 2.325
R752 VDD.n546 VDD.n545 2.325
R753 VDD.n550 VDD.n549 2.325
R754 VDD.n554 VDD.n553 2.325
R755 VDD.n558 VDD.n557 2.325
R756 VDD.n615 VDD.n614 2.261
R757 VDD.n518 VDD.n517 2.261
R758 VDD.n674 VDD.n673 2.261
R759 VDD.n556 VDD.n555 2.261
R760 VDD.n213 VDD.n212 1.791
R761 VDD.n395 VDD.n394 1.791
R762 VDD.n565 VDD.n564 1.791
R763 VDD.n329 VDD.n328 1.791
R764 VDD.n254 VDD.n253 1.791
R765 VDD.n204 VDD.n203 1.791
R766 VDD.n436 VDD.n435 1.791
R767 VDD.n386 VDD.n385 1.791
R768 VDD.n606 VDD.n605 1.791
R769 VDD.n520 VDD.n519 1.31
R770 VDD.n689 VDD.n685 1.145
R771 VDD.n8 VDD.n4 1.145
R772 VDD.n162 VDD.n158 1.119
R773 VDD.n344 VDD.n340 1.119
R774 VDD.n820 VDD.n818 0.957
R775 VDD.n101 VDD.n99 0.777
R776 VDD.n445 VDD.n444 0.754
R777 VDD.n524 VDD.n520 0.566
R778 VDD.n54 VDD.n52 0.525
R779 VDD.n727 VDD.n725 0.525
R780 VDD.n774 VDD.n772 0.525
R781 VDD.n211 VDD.n209 0.305
R782 VDD.n393 VDD.n391 0.305
R783 VDD.n563 VDD.n561 0.305
R784 VDD.n263 VDD.n259 0.295
R785 VDD.n443 VDD.n441 0.295
R786 VDD.n613 VDD.n611 0.295
R787 VDD.n156 VDD.n155 0.227
R788 VDD.n338 VDD.n337 0.227
R789 VDD.n863 VDD.n862 0.135
R790 VDD.n17 VDD.n13 0.09
R791 VDD.n21 VDD.n17 0.09
R792 VDD.n25 VDD.n21 0.09
R793 VDD.n29 VDD.n25 0.09
R794 VDD.n30 VDD.n29 0.09
R795 VDD.n41 VDD.n37 0.09
R796 VDD.n45 VDD.n41 0.09
R797 VDD.n49 VDD.n45 0.09
R798 VDD.n58 VDD.n54 0.09
R799 VDD.n62 VDD.n58 0.09
R800 VDD.n71 VDD.n67 0.09
R801 VDD.n75 VDD.n71 0.09
R802 VDD.n77 VDD.n75 0.09
R803 VDD.n88 VDD.n84 0.09
R804 VDD.n92 VDD.n88 0.09
R805 VDD.n96 VDD.n92 0.09
R806 VDD.n105 VDD.n101 0.09
R807 VDD.n109 VDD.n105 0.09
R808 VDD.n118 VDD.n114 0.09
R809 VDD.n122 VDD.n118 0.09
R810 VDD.n126 VDD.n122 0.09
R811 VDD.n132 VDD.n131 0.09
R812 VDD.n143 VDD.n139 0.09
R813 VDD.n152 VDD.n148 0.09
R814 VDD.n154 VDD.n152 0.09
R815 VDD.n698 VDD.n694 0.09
R816 VDD.n702 VDD.n698 0.09
R817 VDD.n703 VDD.n702 0.09
R818 VDD.n714 VDD.n710 0.09
R819 VDD.n718 VDD.n714 0.09
R820 VDD.n722 VDD.n718 0.09
R821 VDD.n731 VDD.n727 0.09
R822 VDD.n735 VDD.n731 0.09
R823 VDD.n744 VDD.n740 0.09
R824 VDD.n748 VDD.n744 0.09
R825 VDD.n750 VDD.n748 0.09
R826 VDD.n761 VDD.n757 0.09
R827 VDD.n765 VDD.n761 0.09
R828 VDD.n769 VDD.n765 0.09
R829 VDD.n778 VDD.n774 0.09
R830 VDD.n782 VDD.n778 0.09
R831 VDD.n791 VDD.n787 0.09
R832 VDD.n795 VDD.n791 0.09
R833 VDD.n796 VDD.n795 0.09
R834 VDD.n807 VDD.n803 0.09
R835 VDD.n811 VDD.n807 0.09
R836 VDD.n815 VDD.n811 0.09
R837 VDD.n824 VDD.n820 0.09
R838 VDD.n833 VDD.n829 0.09
R839 VDD.n837 VDD.n833 0.09
R840 VDD.n841 VDD.n837 0.09
R841 VDD.n842 VDD.n841 0.09
R842 VDD.n851 VDD.n847 0.09
R843 VDD.n855 VDD.n851 0.09
R844 VDD.n862 VDD.n860 0.09
R845 VDD.n63 VDD.n62 0.078
R846 VDD.n131 VDD.n127 0.078
R847 VDD.n335 VDD.n334 0.078
R848 VDD.n516 VDD.n515 0.078
R849 VDD.n679 VDD.n678 0.078
R850 VDD.n690 VDD.n689 0.078
R851 VDD.n736 VDD.n735 0.078
R852 VDD.n783 VDD.n782 0.078
R853 VDD.n110 VDD.n109 0.071
R854 VDD.n9 VDD.n8 0.07
R855 VDD.n37 VDD 0.065
R856 VDD.n84 CMOS_s3_0/CMOS_AND_1/VDD 0.065
R857 VDD.n139 CMOS_s3_0/CMOS_3in_AND_0/VDD 0.065
R858 VDD.n710 CMOS_s0_0/CMOS_OR_0/VDD 0.065
R859 VDD.n757 CMOS_s0_0/CMOS_AND_0/VDD 0.065
R860 VDD.n803 CMOS_s0_0/CMOS_OR_1/VDD 0.065
R861 VDD.n829 VDD.n825 0.065
R862 VDD.n847 CMOS_s0_0/CMOS_XOR_0/VDD 0.065
R863 VDD.n148 VDD.n144 0.063
R864 VDD.n52 VDD.n50 0.056
R865 VDD.n99 VDD.n97 0.056
R866 VDD.n725 VDD.n723 0.056
R867 VDD.n772 VDD.n770 0.056
R868 VDD.n818 VDD.n816 0.056
R869 VDD.n856 VDD.n855 0.055
R870 VDD.n171 VDD.n167 0.052
R871 VDD.n180 VDD.n176 0.052
R872 VDD.n184 VDD.n180 0.052
R873 VDD.n186 VDD.n184 0.052
R874 VDD.n198 VDD.n194 0.052
R875 VDD.n202 VDD.n198 0.052
R876 VDD.n206 VDD.n202 0.052
R877 VDD.n215 VDD.n211 0.052
R878 VDD.n229 VDD.n225 0.052
R879 VDD.n234 VDD.n229 0.052
R880 VDD.n236 VDD.n234 0.052
R881 VDD.n247 VDD.n243 0.052
R882 VDD.n251 VDD.n247 0.052
R883 VDD.n267 VDD.n263 0.052
R884 VDD.n271 VDD.n267 0.052
R885 VDD.n285 VDD.n281 0.052
R886 VDD.n289 VDD.n285 0.052
R887 VDD.n304 VDD.n300 0.052
R888 VDD.n308 VDD.n304 0.052
R889 VDD.n311 VDD.n308 0.052
R890 VDD.n322 VDD.n318 0.052
R891 VDD.n326 VDD.n322 0.052
R892 VDD.n353 VDD.n349 0.052
R893 VDD.n362 VDD.n358 0.052
R894 VDD.n366 VDD.n362 0.052
R895 VDD.n368 VDD.n366 0.052
R896 VDD.n380 VDD.n376 0.052
R897 VDD.n384 VDD.n380 0.052
R898 VDD.n388 VDD.n384 0.052
R899 VDD.n397 VDD.n393 0.052
R900 VDD.n411 VDD.n407 0.052
R901 VDD.n416 VDD.n411 0.052
R902 VDD.n418 VDD.n416 0.052
R903 VDD.n429 VDD.n425 0.052
R904 VDD.n433 VDD.n429 0.052
R905 VDD.n448 VDD.n443 0.052
R906 VDD.n451 VDD.n448 0.052
R907 VDD.n461 VDD.n457 0.052
R908 VDD.n465 VDD.n461 0.052
R909 VDD.n479 VDD.n475 0.052
R910 VDD.n484 VDD.n479 0.052
R911 VDD.n490 VDD.n489 0.052
R912 VDD.n501 VDD.n497 0.052
R913 VDD.n515 VDD.n511 0.052
R914 VDD.n533 VDD.n529 0.052
R915 VDD.n537 VDD.n533 0.052
R916 VDD.n539 VDD.n537 0.052
R917 VDD.n550 VDD.n546 0.052
R918 VDD.n554 VDD.n550 0.052
R919 VDD.n558 VDD.n554 0.052
R920 VDD.n567 VDD.n563 0.052
R921 VDD.n581 VDD.n577 0.052
R922 VDD.n586 VDD.n581 0.052
R923 VDD.n588 VDD.n586 0.052
R924 VDD.n599 VDD.n595 0.052
R925 VDD.n603 VDD.n599 0.052
R926 VDD.n617 VDD.n613 0.052
R927 VDD.n621 VDD.n617 0.052
R928 VDD.n630 VDD.n626 0.052
R929 VDD.n634 VDD.n630 0.052
R930 VDD.n638 VDD.n634 0.052
R931 VDD.n647 VDD.n643 0.052
R932 VDD.n651 VDD.n647 0.052
R933 VDD.n655 VDD.n651 0.052
R934 VDD.n656 VDD.n655 0.052
R935 VDD.n667 VDD.n663 0.052
R936 VDD.n671 VDD.n667 0.052
R937 VDD.n678 VDD.n676 0.052
R938 VDD.n300 VDD.n295 0.05
R939 VDD.n172 VDD.n171 0.045
R940 VDD.n221 VDD.n220 0.045
R941 VDD.n354 VDD.n353 0.045
R942 VDD.n403 VDD.n402 0.045
R943 VDD.n489 VDD.n485 0.045
R944 VDD.n525 VDD.n524 0.045
R945 VDD.n573 VDD.n572 0.045
R946 VDD.n272 VDD.n271 0.041
R947 VDD.n452 VDD.n451 0.041
R948 VDD.n466 VDD.n465 0.041
R949 VDD.n622 VDD.n621 0.041
R950 VDD.n163 VDD.n162 0.04
R951 VDD.n345 VDD.n344 0.04
R952 VDD.n194 CMOS_s3_0/CMOS_AND_0/VDD 0.037
R953 VDD.n220 VDD.n216 0.037
R954 VDD.n243 CMOS_s3_0/CMOS_XOR_0/VDD 0.037
R955 VDD.n277 VDD.n276 0.037
R956 VDD.n294 VDD.n290 0.037
R957 VDD.n318 CMOS_s3_0/CMOS_XNOR_0/VDD 0.037
R958 VDD.n376 CMOS_s2_0/CMOS_AND_0/VDD 0.037
R959 VDD.n402 VDD.n398 0.037
R960 VDD.n425 CMOS_s2_0/CMOS_XOR_0/VDD 0.037
R961 VDD.n475 VDD.n471 0.037
R962 VDD.n497 CMOS_s2_0/CMOS_XNOR_0/VDD 0.037
R963 VDD.n506 VDD.n502 0.037
R964 VDD.n546 CMOS_s1_0/CMOS_AND_0/VDD 0.037
R965 VDD.n572 VDD.n568 0.037
R966 VDD.n595 CMOS_s1_0/CMOS_XOR_0/VDD 0.037
R967 VDD.n643 VDD.n639 0.037
R968 VDD.n663 CMOS_s1_0/CMOS_XNOR_0/VDD 0.037
R969 VDD.n860 VDD.n856 0.035
R970 VDD.n50 VDD.n49 0.033
R971 VDD.n97 VDD.n96 0.033
R972 VDD.n723 VDD.n722 0.033
R973 VDD.n770 VDD.n769 0.033
R974 VDD.n816 VDD.n815 0.033
R975 VDD.n209 VDD.n207 0.032
R976 VDD.n259 VDD.n257 0.032
R977 VDD.n334 VDD.n332 0.032
R978 VDD.n391 VDD.n389 0.032
R979 VDD.n441 VDD.n439 0.032
R980 VDD.n561 VDD.n559 0.032
R981 VDD.n611 VDD.n609 0.032
R982 VDD.n252 VDD.n251 0.031
R983 VDD.n327 VDD.n326 0.031
R984 VDD.n434 VDD.n433 0.031
R985 VDD.n507 VDD.n506 0.031
R986 VDD.n604 VDD.n603 0.031
R987 VDD.n672 VDD.n671 0.031
R988 CMOS_s0_0/VDD VDD.n863 0.027
R989 VDD.n144 VDD.n143 0.026
R990 VDD.n30 VDD 0.025
R991 VDD.n132 CMOS_s3_0/CMOS_3in_AND_0/VDD 0.025
R992 VDD.n703 CMOS_s0_0/CMOS_OR_0/VDD 0.025
R993 VDD.n796 CMOS_s0_0/CMOS_OR_1/VDD 0.025
R994 VDD.n825 VDD.n824 0.025
R995 VDD.n842 CMOS_s0_0/CMOS_XOR_0/VDD 0.025
R996 VDD.n13 VDD.n9 0.02
R997 VDD.n256 VDD.n252 0.02
R998 VDD.n331 VDD.n327 0.02
R999 VDD.n438 VDD.n434 0.02
R1000 VDD.n511 VDD.n507 0.02
R1001 VDD.n608 VDD.n604 0.02
R1002 VDD.n676 VDD.n672 0.02
R1003 VDD.n207 VDD.n206 0.019
R1004 VDD.n257 VDD.n256 0.019
R1005 VDD.n332 VDD.n331 0.019
R1006 VDD.n389 VDD.n388 0.019
R1007 VDD.n439 VDD.n438 0.019
R1008 VDD.n559 VDD.n558 0.019
R1009 VDD.n609 VDD.n608 0.019
R1010 VDD.n114 VDD.n110 0.018
R1011 VDD.n77 VDD.n76 0.017
R1012 VDD.n750 VDD.n749 0.017
R1013 VDD.n281 VDD.n277 0.015
R1014 VDD.n335 CMOS_s3_0/VDD 0.015
R1015 VDD.n502 VDD.n501 0.015
R1016 VDD.n516 CMOS_s2_0/VDD 0.015
R1017 VDD.n679 CMOS_s1_0/VDD 0.015
R1018 VDD.n216 VDD.n215 0.014
R1019 VDD.n290 VDD.n289 0.014
R1020 VDD.n398 VDD.n397 0.014
R1021 VDD.n471 VDD.n470 0.014
R1022 VDD.n490 CMOS_s2_0/CMOS_XNOR_0/VDD 0.014
R1023 VDD.n568 VDD.n567 0.014
R1024 VDD.n639 VDD.n638 0.014
R1025 VDD.n656 CMOS_s1_0/CMOS_XNOR_0/VDD 0.014
R1026 VDD.n67 VDD.n63 0.011
R1027 VDD.n127 VDD.n126 0.011
R1028 VDD.n167 VDD.n163 0.011
R1029 VDD.n349 VDD.n345 0.011
R1030 VDD.n694 VDD.n690 0.011
R1031 VDD.n740 VDD.n736 0.011
R1032 VDD.n787 VDD.n783 0.011
R1033 VDD.n186 VDD.n185 0.01
R1034 VDD.n236 VDD.n235 0.01
R1035 VDD.n276 VDD.n272 0.01
R1036 VDD.n311 VDD.n310 0.01
R1037 VDD.n368 VDD.n367 0.01
R1038 VDD.n418 VDD.n417 0.01
R1039 VDD.n457 VDD.n452 0.01
R1040 VDD.n470 VDD.n466 0.01
R1041 VDD.n539 VDD.n538 0.01
R1042 VDD.n588 VDD.n587 0.01
R1043 VDD.n626 VDD.n622 0.01
R1044 CMOS_s0_0/VDD VDD 0.008
R1045 VDD.n76 CMOS_s3_0/CMOS_AND_1/VDD 0.007
R1046 VDD.n749 CMOS_s0_0/CMOS_AND_0/VDD 0.007
R1047 VDD.n176 VDD.n172 0.006
R1048 VDD.n225 VDD.n221 0.006
R1049 VDD.n358 VDD.n354 0.006
R1050 VDD.n407 VDD.n403 0.006
R1051 VDD.n485 VDD.n484 0.006
R1052 VDD.n529 VDD.n525 0.006
R1053 VDD.n577 VDD.n573 0.006
R1054 VDD.n185 CMOS_s3_0/CMOS_AND_0/VDD 0.004
R1055 VDD.n235 CMOS_s3_0/CMOS_XOR_0/VDD 0.004
R1056 VDD.n367 CMOS_s2_0/CMOS_AND_0/VDD 0.004
R1057 VDD.n417 CMOS_s2_0/CMOS_XOR_0/VDD 0.004
R1058 VDD.n538 CMOS_s1_0/CMOS_AND_0/VDD 0.004
R1059 VDD.n587 CMOS_s1_0/CMOS_XOR_0/VDD 0.004
R1060 VDD.n310 CMOS_s3_0/CMOS_XNOR_0/VDD 0.003
R1061 VDD.n295 VDD.n294 0.002
R1062 x3.n2 x3.t11 993.097
R1063 x3.n8 x3.t3 993.097
R1064 x3.t12 x3.t7 924.95
R1065 x3.t9 x3.t6 924.95
R1066 x3.t5 x3.t4 924.95
R1067 CMOS_s3_0/CMOS_XOR_0/B x3.t12 633.02
R1068 CMOS_s1_0/CMOS_XOR_0/B x3.t9 633.02
R1069 CMOS_s0_0/CMOS_XOR_0/B x3.t5 633.02
R1070 x3.n4 x3.t0 579.86
R1071 x3.n0 x3.t10 570.366
R1072 x3.n0 x3.t2 570.366
R1073 x3.n4 x3.t8 547.727
R1074 x3.n2 x3.t13 356.59
R1075 x3.n8 x3.t1 356.59
R1076 x3.n10 CMOS_s0_0/CMOS_XOR_0/B 317
R1077 x3.n3 CMOS_s2_0/CMOS_XNOR_0/A 173
R1078 x3.n9 CMOS_s0_0/CMOS_XNOR_0/A 173
R1079 x3.n1 x3 158.792
R1080 x3 x3.n0 78.72
R1081 CMOS_s2_0/CMOS_XNOR_0/A x3.n2 78.72
R1082 CMOS_s0_0/CMOS_XNOR_0/A x3.n8 78.72
R1083 x3.n1 CMOS_s3_0/CMOS_XOR_0/B 42.892
R1084 x3.n7 CMOS_s1_0/CMOS_XOR_0/B 42.892
R1085 x3.n6 x3.n5 10.794
R1086 x3.n5 x3.n4 8.764
R1087 x3.n3 CMOS_s3_0/x3 3.443
R1088 x3.n7 x3.n6 3.406
R1089 x3.n10 x3.n9 3.128
R1090 x3.n5 CMOS_s1_0/CMOS_AND_1/B 2.72
R1091 x3.n9 CMOS_s1_0/x3 1.758
R1092 CMOS_s2_0/x3 x3.n3 1.599
R1093 x3.n6 CMOS_s2_0/x3 1.464
R1094 CMOS_s1_0/x3 x3.n7 0.157
R1095 CMOS_s3_0/x3 x3.n1 0.157
R1096 x3 x3.n10 0.151
R1097 CMOS_s0_0/x3 x3 0.003
R1098 GND.n324 GND.t16 2383.33
R1099 GND.n675 GND.t25 2383.33
R1100 GND.n163 GND.t46 1283.79
R1101 GND.n164 GND.n163 284.705
R1102 GND.n37 GND.t84 180.204
R1103 GND.n361 GND.t103 159.607
R1104 GND.n292 GND.t58 159.607
R1105 GND.n535 GND.t94 159.607
R1106 GND.n468 GND.t10 159.607
R1107 GND.n712 GND.t111 159.607
R1108 GND.n643 GND.t59 159.607
R1109 GND.n189 GND.t60 159.607
R1110 GND.n325 GND.n324 150.98
R1111 GND.n676 GND.n675 150.98
R1112 GND.n29 GND.t37 135.153
R1113 GND.n369 GND.t128 133.725
R1114 GND.n300 GND.t97 133.725
R1115 GND.n543 GND.t54 133.725
R1116 GND.n476 GND.t100 133.725
R1117 GND.n720 GND.t29 133.725
R1118 GND.n651 GND.t23 133.725
R1119 GND.n197 GND.t61 133.725
R1120 GND.n351 GND.t41 125.098
R1121 GND.n280 GND.t8 125.098
R1122 GND.n525 GND.t99 125.098
R1123 GND.n456 GND.t73 125.098
R1124 GND.n702 GND.t70 125.098
R1125 GND.n631 GND.t20 125.098
R1126 GND.n177 GND.t40 125.098
R1127 GND.n369 GND.t56 103.529
R1128 GND.n300 GND.t135 103.529
R1129 GND.n253 GND.t0 103.529
R1130 GND.n499 GND.t6 103.529
R1131 GND.n543 GND.t95 103.529
R1132 GND.n476 GND.t33 103.529
R1133 GND.n429 GND.t2 103.529
R1134 GND.n720 GND.t130 103.529
R1135 GND.n651 GND.t63 103.529
R1136 GND.n604 GND.t21 103.529
R1137 GND.n83 GND.t44 103.529
R1138 GND.n130 GND.t65 103.529
R1139 GND.n343 GND.t42 99.215
R1140 GND.n271 GND.t31 99.215
R1141 GND.n517 GND.t125 99.215
R1142 GND.n447 GND.t118 99.215
R1143 GND.n694 GND.t133 99.215
R1144 GND.n622 GND.t137 99.215
R1145 GND.n169 GND.t18 99.215
R1146 GND.n7 GND.t4 90.102
R1147 GND.n333 GND.t82 77.647
R1148 GND.n361 GND.t48 77.647
R1149 GND.n292 GND.t81 77.647
R1150 GND.n213 GND.t106 77.647
R1151 GND.n244 GND.t116 77.647
R1152 GND.n494 GND.t52 77.647
R1153 GND.n535 GND.t39 77.647
R1154 GND.n468 GND.t113 77.647
R1155 GND.n389 GND.t123 77.647
R1156 GND.n420 GND.t12 77.647
R1157 GND.n684 GND.t50 77.647
R1158 GND.n712 GND.t132 77.647
R1159 GND.n643 GND.t86 77.647
R1160 GND.n564 GND.t74 77.647
R1161 GND.n595 GND.t112 77.647
R1162 GND.n75 GND.t11 77.647
R1163 GND.n122 GND.t71 77.647
R1164 GND.n355 GND.t127 51.764
R1165 GND.n271 GND.t79 51.764
R1166 GND.n222 GND.t109 51.764
R1167 GND.n236 GND.t76 51.764
R1168 GND.n529 GND.t102 51.764
R1169 GND.n447 GND.t27 51.764
R1170 GND.n398 GND.t104 51.764
R1171 GND.n412 GND.t121 51.764
R1172 GND.n706 GND.t68 51.764
R1173 GND.n622 GND.t92 51.764
R1174 GND.n573 GND.t14 51.764
R1175 GND.n587 GND.t114 51.764
R1176 GND.n54 GND.t87 51.764
R1177 GND.n100 GND.t35 51.764
R1178 GND.n380 GND.n379 37.883
R1179 GND.n554 GND.n553 35.52
R1180 GND.n731 GND.n730 35.52
R1181 GND.n204 GND.n203 35.52
R1182 GND.n201 GND.t139 30.21
R1183 GND.n378 GND.t57 30.21
R1184 GND.n337 GND.t83 30.21
R1185 GND.n309 GND.t136 30.21
R1186 GND.n275 GND.t80 30.21
R1187 GND.n235 GND.t77 30.21
R1188 GND.n217 GND.t107 30.21
R1189 GND.n552 GND.t96 30.21
R1190 GND.n503 GND.t7 30.21
R1191 GND.n485 GND.t34 30.21
R1192 GND.n451 GND.t28 30.21
R1193 GND.n411 GND.t122 30.21
R1194 GND.n393 GND.t124 30.21
R1195 GND.n729 GND.t131 30.21
R1196 GND.n688 GND.t51 30.21
R1197 GND.n660 GND.t64 30.21
R1198 GND.n626 GND.t93 30.21
R1199 GND.n586 GND.t115 30.21
R1200 GND.n568 GND.t75 30.21
R1201 GND.n58 GND.t88 30.21
R1202 GND.n91 GND.t108 30.21
R1203 GND.n104 GND.t36 30.21
R1204 GND.n138 GND.t67 30.21
R1205 GND.n168 GND.t19 30.21
R1206 GND.n201 GND.t62 30.21
R1207 GND.n150 GND.t47 30.21
R1208 GND.n226 GND.t110 30.21
R1209 GND.n261 GND.t1 30.21
R1210 GND.n270 GND.t32 30.21
R1211 GND.n304 GND.t98 30.21
R1212 GND.n323 GND.t17 30.21
R1213 GND.n342 GND.t43 30.21
R1214 GND.n373 GND.t129 30.21
R1215 GND.n402 GND.t105 30.21
R1216 GND.n437 GND.t9 30.21
R1217 GND.n446 GND.t119 30.21
R1218 GND.n480 GND.t101 30.21
R1219 GND.n498 GND.t53 30.21
R1220 GND.n516 GND.t126 30.21
R1221 GND.n547 GND.t55 30.21
R1222 GND.n577 GND.t15 30.21
R1223 GND.n612 GND.t22 30.21
R1224 GND.n621 GND.t138 30.21
R1225 GND.n655 GND.t24 30.21
R1226 GND.n674 GND.t26 30.21
R1227 GND.n693 GND.t134 30.21
R1228 GND.n724 GND.t30 30.21
R1229 GND.n11 GND.t5 30.21
R1230 GND.n24 GND.t38 30.21
R1231 GND.n45 GND.t85 30.21
R1232 GND.n58 GND.t90 30.21
R1233 GND.n91 GND.t45 30.21
R1234 GND.n104 GND.t49 30.21
R1235 GND.n117 GND.t72 30.21
R1236 GND.n138 GND.t66 30.21
R1237 GND.n168 GND.t91 30.21
R1238 GND.n521 GND.t69 25.882
R1239 GND.n208 GND.t117 24
R1240 GND.n208 GND.t78 24
R1241 GND.n384 GND.t13 24
R1242 GND.n384 GND.t3 24
R1243 GND.n559 GND.t120 24
R1244 GND.n559 GND.t89 24
R1245 GND.n294 GND.n291 11.52
R1246 GND.n246 GND.n243 11.52
R1247 GND.n363 GND.n360 11.52
R1248 GND.n470 GND.n467 11.52
R1249 GND.n422 GND.n419 11.52
R1250 GND.n537 GND.n534 11.52
R1251 GND.n645 GND.n642 11.52
R1252 GND.n597 GND.n594 11.52
R1253 GND.n714 GND.n711 11.52
R1254 GND.n31 GND.n28 11.52
R1255 GND.n77 GND.n74 11.52
R1256 GND.n124 GND.n121 11.52
R1257 GND.n191 GND.n188 11.52
R1258 GND.n554 GND.n381 9.77
R1259 GND.n731 GND.n556 9.77
R1260 GND.n211 GND.n210 9.154
R1261 GND.n215 GND.n214 9.154
R1262 GND.n214 GND.n213 9.154
R1263 GND.n220 GND.n219 9.154
R1264 GND.n219 GND.n218 9.154
R1265 GND.n224 GND.n223 9.154
R1266 GND.n223 GND.n222 9.154
R1267 GND.n229 GND.n228 9.154
R1268 GND.n228 GND.n227 9.154
R1269 GND.n233 GND.n232 9.154
R1270 GND.n232 GND.n231 9.154
R1271 GND.n238 GND.n237 9.154
R1272 GND.n237 GND.n236 9.154
R1273 GND.n243 GND.n242 9.154
R1274 GND.n242 GND.n241 9.154
R1275 GND.n246 GND.n245 9.154
R1276 GND.n245 GND.n244 9.154
R1277 GND.n250 GND.n249 9.154
R1278 GND.n249 GND.n248 9.154
R1279 GND.n255 GND.n254 9.154
R1280 GND.n254 GND.n253 9.154
R1281 GND.n259 GND.n258 9.154
R1282 GND.n268 GND.n267 9.154
R1283 GND.n273 GND.n272 9.154
R1284 GND.n272 GND.n271 9.154
R1285 GND.n278 GND.n277 9.154
R1286 GND.n277 GND.n276 9.154
R1287 GND.n282 GND.n281 9.154
R1288 GND.n281 GND.n280 9.154
R1289 GND.n286 GND.n285 9.154
R1290 GND.n285 GND.n284 9.154
R1291 GND.n291 GND.n290 9.154
R1292 GND.n290 GND.n289 9.154
R1293 GND.n294 GND.n293 9.154
R1294 GND.n293 GND.n292 9.154
R1295 GND.n298 GND.n297 9.154
R1296 GND.n297 GND.n296 9.154
R1297 GND.n302 GND.n301 9.154
R1298 GND.n301 GND.n300 9.154
R1299 GND.n307 GND.n306 9.154
R1300 GND.n313 GND.n312 9.154
R1301 GND.n316 GND.n315 9.154
R1302 GND.n321 GND.n320 9.154
R1303 GND.n327 GND.n326 9.154
R1304 GND.n326 GND.n325 9.154
R1305 GND.n331 GND.n330 9.154
R1306 GND.n330 GND.n329 9.154
R1307 GND.n335 GND.n334 9.154
R1308 GND.n334 GND.n333 9.154
R1309 GND.n340 GND.n339 9.154
R1310 GND.n339 GND.n338 9.154
R1311 GND.n345 GND.n344 9.154
R1312 GND.n344 GND.n343 9.154
R1313 GND.n349 GND.n348 9.154
R1314 GND.n348 GND.n347 9.154
R1315 GND.n353 GND.n352 9.154
R1316 GND.n352 GND.n351 9.154
R1317 GND.n357 GND.n356 9.154
R1318 GND.n356 GND.n355 9.154
R1319 GND.n360 GND.n207 9.154
R1320 GND.n207 GND.n206 9.154
R1321 GND.n363 GND.n362 9.154
R1322 GND.n362 GND.n361 9.154
R1323 GND.n367 GND.n366 9.154
R1324 GND.n366 GND.n365 9.154
R1325 GND.n371 GND.n370 9.154
R1326 GND.n370 GND.n369 9.154
R1327 GND.n376 GND.n375 9.154
R1328 GND.n387 GND.n386 9.154
R1329 GND.n391 GND.n390 9.154
R1330 GND.n390 GND.n389 9.154
R1331 GND.n396 GND.n395 9.154
R1332 GND.n395 GND.n394 9.154
R1333 GND.n400 GND.n399 9.154
R1334 GND.n399 GND.n398 9.154
R1335 GND.n405 GND.n404 9.154
R1336 GND.n404 GND.n403 9.154
R1337 GND.n409 GND.n408 9.154
R1338 GND.n408 GND.n407 9.154
R1339 GND.n414 GND.n413 9.154
R1340 GND.n413 GND.n412 9.154
R1341 GND.n419 GND.n418 9.154
R1342 GND.n418 GND.n417 9.154
R1343 GND.n422 GND.n421 9.154
R1344 GND.n421 GND.n420 9.154
R1345 GND.n426 GND.n425 9.154
R1346 GND.n425 GND.n424 9.154
R1347 GND.n431 GND.n430 9.154
R1348 GND.n430 GND.n429 9.154
R1349 GND.n435 GND.n434 9.154
R1350 GND.n444 GND.n443 9.154
R1351 GND.n449 GND.n448 9.154
R1352 GND.n448 GND.n447 9.154
R1353 GND.n454 GND.n453 9.154
R1354 GND.n453 GND.n452 9.154
R1355 GND.n458 GND.n457 9.154
R1356 GND.n457 GND.n456 9.154
R1357 GND.n462 GND.n461 9.154
R1358 GND.n461 GND.n460 9.154
R1359 GND.n467 GND.n466 9.154
R1360 GND.n466 GND.n465 9.154
R1361 GND.n470 GND.n469 9.154
R1362 GND.n469 GND.n468 9.154
R1363 GND.n474 GND.n473 9.154
R1364 GND.n473 GND.n472 9.154
R1365 GND.n478 GND.n477 9.154
R1366 GND.n477 GND.n476 9.154
R1367 GND.n483 GND.n482 9.154
R1368 GND.n492 GND.n491 9.154
R1369 GND.n496 GND.n495 9.154
R1370 GND.n495 GND.n494 9.154
R1371 GND.n501 GND.n500 9.154
R1372 GND.n500 GND.n499 9.154
R1373 GND.n506 GND.n505 9.154
R1374 GND.n505 GND.n504 9.154
R1375 GND.n510 GND.n509 9.154
R1376 GND.n509 GND.n508 9.154
R1377 GND.n514 GND.n513 9.154
R1378 GND.n513 GND.n512 9.154
R1379 GND.n519 GND.n518 9.154
R1380 GND.n518 GND.n517 9.154
R1381 GND.n523 GND.n522 9.154
R1382 GND.n522 GND.n521 9.154
R1383 GND.n527 GND.n526 9.154
R1384 GND.n526 GND.n525 9.154
R1385 GND.n531 GND.n530 9.154
R1386 GND.n530 GND.n529 9.154
R1387 GND.n534 GND.n383 9.154
R1388 GND.n383 GND.n382 9.154
R1389 GND.n537 GND.n536 9.154
R1390 GND.n536 GND.n535 9.154
R1391 GND.n541 GND.n540 9.154
R1392 GND.n540 GND.n539 9.154
R1393 GND.n545 GND.n544 9.154
R1394 GND.n544 GND.n543 9.154
R1395 GND.n550 GND.n549 9.154
R1396 GND.n562 GND.n561 9.154
R1397 GND.n566 GND.n565 9.154
R1398 GND.n565 GND.n564 9.154
R1399 GND.n571 GND.n570 9.154
R1400 GND.n570 GND.n569 9.154
R1401 GND.n575 GND.n574 9.154
R1402 GND.n574 GND.n573 9.154
R1403 GND.n580 GND.n579 9.154
R1404 GND.n579 GND.n578 9.154
R1405 GND.n584 GND.n583 9.154
R1406 GND.n583 GND.n582 9.154
R1407 GND.n589 GND.n588 9.154
R1408 GND.n588 GND.n587 9.154
R1409 GND.n594 GND.n593 9.154
R1410 GND.n593 GND.n592 9.154
R1411 GND.n597 GND.n596 9.154
R1412 GND.n596 GND.n595 9.154
R1413 GND.n601 GND.n600 9.154
R1414 GND.n600 GND.n599 9.154
R1415 GND.n606 GND.n605 9.154
R1416 GND.n605 GND.n604 9.154
R1417 GND.n610 GND.n609 9.154
R1418 GND.n619 GND.n618 9.154
R1419 GND.n624 GND.n623 9.154
R1420 GND.n623 GND.n622 9.154
R1421 GND.n629 GND.n628 9.154
R1422 GND.n628 GND.n627 9.154
R1423 GND.n633 GND.n632 9.154
R1424 GND.n632 GND.n631 9.154
R1425 GND.n637 GND.n636 9.154
R1426 GND.n636 GND.n635 9.154
R1427 GND.n642 GND.n641 9.154
R1428 GND.n641 GND.n640 9.154
R1429 GND.n645 GND.n644 9.154
R1430 GND.n644 GND.n643 9.154
R1431 GND.n649 GND.n648 9.154
R1432 GND.n648 GND.n647 9.154
R1433 GND.n653 GND.n652 9.154
R1434 GND.n652 GND.n651 9.154
R1435 GND.n658 GND.n657 9.154
R1436 GND.n664 GND.n663 9.154
R1437 GND.n667 GND.n666 9.154
R1438 GND.n672 GND.n671 9.154
R1439 GND.n678 GND.n677 9.154
R1440 GND.n677 GND.n676 9.154
R1441 GND.n682 GND.n681 9.154
R1442 GND.n681 GND.n680 9.154
R1443 GND.n686 GND.n685 9.154
R1444 GND.n685 GND.n684 9.154
R1445 GND.n691 GND.n690 9.154
R1446 GND.n690 GND.n689 9.154
R1447 GND.n696 GND.n695 9.154
R1448 GND.n695 GND.n694 9.154
R1449 GND.n700 GND.n699 9.154
R1450 GND.n699 GND.n698 9.154
R1451 GND.n704 GND.n703 9.154
R1452 GND.n703 GND.n702 9.154
R1453 GND.n708 GND.n707 9.154
R1454 GND.n707 GND.n706 9.154
R1455 GND.n711 GND.n558 9.154
R1456 GND.n558 GND.n557 9.154
R1457 GND.n714 GND.n713 9.154
R1458 GND.n713 GND.n712 9.154
R1459 GND.n718 GND.n717 9.154
R1460 GND.n717 GND.n716 9.154
R1461 GND.n722 GND.n721 9.154
R1462 GND.n721 GND.n720 9.154
R1463 GND.n727 GND.n726 9.154
R1464 GND.n5 GND.n4 9.154
R1465 GND.n52 GND.n51 9.154
R1466 GND.n98 GND.n97 9.154
R1467 GND.n102 GND.n101 9.154
R1468 GND.n101 GND.n100 9.154
R1469 GND.n107 GND.n106 9.154
R1470 GND.n106 GND.n105 9.154
R1471 GND.n111 GND.n110 9.154
R1472 GND.n110 GND.n109 9.154
R1473 GND.n115 GND.n114 9.154
R1474 GND.n114 GND.n113 9.154
R1475 GND.n121 GND.n120 9.154
R1476 GND.n120 GND.n119 9.154
R1477 GND.n124 GND.n123 9.154
R1478 GND.n123 GND.n122 9.154
R1479 GND.n128 GND.n127 9.154
R1480 GND.n127 GND.n126 9.154
R1481 GND.n132 GND.n131 9.154
R1482 GND.n131 GND.n130 9.154
R1483 GND.n136 GND.n135 9.154
R1484 GND.n56 GND.n55 9.154
R1485 GND.n55 GND.n54 9.154
R1486 GND.n61 GND.n60 9.154
R1487 GND.n60 GND.n59 9.154
R1488 GND.n65 GND.n64 9.154
R1489 GND.n64 GND.n63 9.154
R1490 GND.n69 GND.n68 9.154
R1491 GND.n68 GND.n67 9.154
R1492 GND.n74 GND.n73 9.154
R1493 GND.n73 GND.n72 9.154
R1494 GND.n77 GND.n76 9.154
R1495 GND.n76 GND.n75 9.154
R1496 GND.n81 GND.n80 9.154
R1497 GND.n80 GND.n79 9.154
R1498 GND.n85 GND.n84 9.154
R1499 GND.n84 GND.n83 9.154
R1500 GND.n89 GND.n88 9.154
R1501 GND.n9 GND.n8 9.154
R1502 GND.n8 GND.n7 9.154
R1503 GND.n14 GND.n13 9.154
R1504 GND.n13 GND.n12 9.154
R1505 GND.n18 GND.n17 9.154
R1506 GND.n17 GND.n16 9.154
R1507 GND.n22 GND.n21 9.154
R1508 GND.n21 GND.n20 9.154
R1509 GND.n28 GND.n27 9.154
R1510 GND.n27 GND.n26 9.154
R1511 GND.n31 GND.n30 9.154
R1512 GND.n30 GND.n29 9.154
R1513 GND.n35 GND.n34 9.154
R1514 GND.n34 GND.n33 9.154
R1515 GND.n39 GND.n38 9.154
R1516 GND.n38 GND.n37 9.154
R1517 GND.n43 GND.n42 9.154
R1518 GND.n145 GND.n144 9.154
R1519 GND.n148 GND.n147 9.154
R1520 GND.n153 GND.n152 9.154
R1521 GND.n156 GND.n155 9.154
R1522 GND.n161 GND.n160 9.154
R1523 GND.n166 GND.n165 9.154
R1524 GND.n165 GND.n164 9.154
R1525 GND.n171 GND.n170 9.154
R1526 GND.n170 GND.n169 9.154
R1527 GND.n175 GND.n174 9.154
R1528 GND.n174 GND.n173 9.154
R1529 GND.n179 GND.n178 9.154
R1530 GND.n178 GND.n177 9.154
R1531 GND.n183 GND.n182 9.154
R1532 GND.n182 GND.n181 9.154
R1533 GND.n188 GND.n187 9.154
R1534 GND.n187 GND.n186 9.154
R1535 GND.n191 GND.n190 9.154
R1536 GND.n190 GND.n189 9.154
R1537 GND.n195 GND.n194 9.154
R1538 GND.n194 GND.n193 9.154
R1539 GND.n199 GND.n198 9.154
R1540 GND.n198 GND.n197 9.154
R1541 GND.n2 GND.n1 9.154
R1542 GND.n320 GND.n319 8.108
R1543 GND.n210 GND.n209 8.108
R1544 GND.n386 GND.n385 8.108
R1545 GND.n671 GND.n670 8.108
R1546 GND.n561 GND.n560 8.108
R1547 GND.n152 GND.n151 8.108
R1548 GND.n160 GND.n159 8.108
R1549 GND.n144 GND.n143 8.108
R1550 GND.n252 GND.n208 6.21
R1551 GND.n428 GND.n384 6.21
R1552 GND.n603 GND.n559 6.21
R1553 GND.n381 GND.n380 4.909
R1554 GND.n733 GND.n732 4.894
R1555 GND.n556 GND.n555 4.894
R1556 GND.n379 GND.n378 4.706
R1557 GND.n553 GND.n552 4.706
R1558 GND.n730 GND.n729 4.706
R1559 GND.n216 GND.n215 4.65
R1560 GND.n221 GND.n220 4.65
R1561 GND.n225 GND.n224 4.65
R1562 GND.n230 GND.n229 4.65
R1563 GND.n234 GND.n233 4.65
R1564 GND.n239 GND.n238 4.65
R1565 GND.n243 GND.n240 4.65
R1566 GND.n247 GND.n246 4.65
R1567 GND.n251 GND.n250 4.65
R1568 GND.n256 GND.n255 4.65
R1569 GND.n260 GND.n259 4.65
R1570 GND.n263 GND.n262 4.65
R1571 GND.n265 GND.n264 4.65
R1572 GND.n269 GND.n268 4.65
R1573 GND.n274 GND.n273 4.65
R1574 GND.n279 GND.n278 4.65
R1575 GND.n283 GND.n282 4.65
R1576 GND.n287 GND.n286 4.65
R1577 GND.n291 GND.n288 4.65
R1578 GND.n295 GND.n294 4.65
R1579 GND.n299 GND.n298 4.65
R1580 GND.n303 GND.n302 4.65
R1581 GND.n308 GND.n307 4.65
R1582 GND.n311 GND.n310 4.65
R1583 GND.n314 GND.n313 4.65
R1584 GND.n317 GND.n316 4.65
R1585 GND.n322 GND.n321 4.65
R1586 GND.n328 GND.n327 4.65
R1587 GND.n332 GND.n331 4.65
R1588 GND.n336 GND.n335 4.65
R1589 GND.n341 GND.n340 4.65
R1590 GND.n346 GND.n345 4.65
R1591 GND.n350 GND.n349 4.65
R1592 GND.n354 GND.n353 4.65
R1593 GND.n358 GND.n357 4.65
R1594 GND.n360 GND.n359 4.65
R1595 GND.n364 GND.n363 4.65
R1596 GND.n368 GND.n367 4.65
R1597 GND.n372 GND.n371 4.65
R1598 GND.n377 GND.n376 4.65
R1599 GND.n392 GND.n391 4.65
R1600 GND.n397 GND.n396 4.65
R1601 GND.n401 GND.n400 4.65
R1602 GND.n406 GND.n405 4.65
R1603 GND.n410 GND.n409 4.65
R1604 GND.n415 GND.n414 4.65
R1605 GND.n419 GND.n416 4.65
R1606 GND.n423 GND.n422 4.65
R1607 GND.n427 GND.n426 4.65
R1608 GND.n432 GND.n431 4.65
R1609 GND.n436 GND.n435 4.65
R1610 GND.n439 GND.n438 4.65
R1611 GND.n441 GND.n440 4.65
R1612 GND.n445 GND.n444 4.65
R1613 GND.n450 GND.n449 4.65
R1614 GND.n455 GND.n454 4.65
R1615 GND.n459 GND.n458 4.65
R1616 GND.n463 GND.n462 4.65
R1617 GND.n467 GND.n464 4.65
R1618 GND.n471 GND.n470 4.65
R1619 GND.n475 GND.n474 4.65
R1620 GND.n479 GND.n478 4.65
R1621 GND.n484 GND.n483 4.65
R1622 GND.n487 GND.n486 4.65
R1623 GND.n489 GND.n488 4.65
R1624 GND.n493 GND.n492 4.65
R1625 GND.n497 GND.n496 4.65
R1626 GND.n502 GND.n501 4.65
R1627 GND.n507 GND.n506 4.65
R1628 GND.n511 GND.n510 4.65
R1629 GND.n515 GND.n514 4.65
R1630 GND.n520 GND.n519 4.65
R1631 GND.n524 GND.n523 4.65
R1632 GND.n528 GND.n527 4.65
R1633 GND.n532 GND.n531 4.65
R1634 GND.n534 GND.n533 4.65
R1635 GND.n538 GND.n537 4.65
R1636 GND.n542 GND.n541 4.65
R1637 GND.n546 GND.n545 4.65
R1638 GND.n551 GND.n550 4.65
R1639 GND.n567 GND.n566 4.65
R1640 GND.n572 GND.n571 4.65
R1641 GND.n576 GND.n575 4.65
R1642 GND.n581 GND.n580 4.65
R1643 GND.n585 GND.n584 4.65
R1644 GND.n590 GND.n589 4.65
R1645 GND.n594 GND.n591 4.65
R1646 GND.n598 GND.n597 4.65
R1647 GND.n602 GND.n601 4.65
R1648 GND.n607 GND.n606 4.65
R1649 GND.n611 GND.n610 4.65
R1650 GND.n614 GND.n613 4.65
R1651 GND.n616 GND.n615 4.65
R1652 GND.n620 GND.n619 4.65
R1653 GND.n625 GND.n624 4.65
R1654 GND.n630 GND.n629 4.65
R1655 GND.n634 GND.n633 4.65
R1656 GND.n638 GND.n637 4.65
R1657 GND.n642 GND.n639 4.65
R1658 GND.n646 GND.n645 4.65
R1659 GND.n650 GND.n649 4.65
R1660 GND.n654 GND.n653 4.65
R1661 GND.n659 GND.n658 4.65
R1662 GND.n662 GND.n661 4.65
R1663 GND.n665 GND.n664 4.65
R1664 GND.n668 GND.n667 4.65
R1665 GND.n673 GND.n672 4.65
R1666 GND.n679 GND.n678 4.65
R1667 GND.n683 GND.n682 4.65
R1668 GND.n687 GND.n686 4.65
R1669 GND.n692 GND.n691 4.65
R1670 GND.n697 GND.n696 4.65
R1671 GND.n701 GND.n700 4.65
R1672 GND.n705 GND.n704 4.65
R1673 GND.n709 GND.n708 4.65
R1674 GND.n711 GND.n710 4.65
R1675 GND.n715 GND.n714 4.65
R1676 GND.n719 GND.n718 4.65
R1677 GND.n723 GND.n722 4.65
R1678 GND.n728 GND.n727 4.65
R1679 GND.n140 GND.n139 4.65
R1680 GND.n99 GND.n98 4.65
R1681 GND.n103 GND.n102 4.65
R1682 GND.n108 GND.n107 4.65
R1683 GND.n112 GND.n111 4.65
R1684 GND.n116 GND.n115 4.65
R1685 GND.n121 GND.n118 4.65
R1686 GND.n125 GND.n124 4.65
R1687 GND.n129 GND.n128 4.65
R1688 GND.n133 GND.n132 4.65
R1689 GND.n137 GND.n136 4.65
R1690 GND.n95 GND.n94 4.65
R1691 GND.n93 GND.n92 4.65
R1692 GND.n53 GND.n52 4.65
R1693 GND.n57 GND.n56 4.65
R1694 GND.n62 GND.n61 4.65
R1695 GND.n66 GND.n65 4.65
R1696 GND.n70 GND.n69 4.65
R1697 GND.n74 GND.n71 4.65
R1698 GND.n78 GND.n77 4.65
R1699 GND.n82 GND.n81 4.65
R1700 GND.n86 GND.n85 4.65
R1701 GND.n90 GND.n89 4.65
R1702 GND.n49 GND.n48 4.65
R1703 GND.n47 GND.n46 4.65
R1704 GND.n10 GND.n9 4.65
R1705 GND.n15 GND.n14 4.65
R1706 GND.n19 GND.n18 4.65
R1707 GND.n23 GND.n22 4.65
R1708 GND.n28 GND.n25 4.65
R1709 GND.n32 GND.n31 4.65
R1710 GND.n36 GND.n35 4.65
R1711 GND.n40 GND.n39 4.65
R1712 GND.n44 GND.n43 4.65
R1713 GND.n146 GND.n145 4.65
R1714 GND.n149 GND.n148 4.65
R1715 GND.n154 GND.n153 4.65
R1716 GND.n157 GND.n156 4.65
R1717 GND.n162 GND.n161 4.65
R1718 GND.n167 GND.n166 4.65
R1719 GND.n172 GND.n171 4.65
R1720 GND.n176 GND.n175 4.65
R1721 GND.n180 GND.n179 4.65
R1722 GND.n184 GND.n183 4.65
R1723 GND.n188 GND.n185 4.65
R1724 GND.n192 GND.n191 4.65
R1725 GND.n196 GND.n195 4.65
R1726 GND.n200 GND.n199 4.65
R1727 GND.n142 GND.n141 4.65
R1728 GND.n732 GND.n731 3.127
R1729 GND.n555 GND.n554 3.127
R1730 GND.n205 GND.n204 3.127
R1731 GND.n258 GND.n257 2.759
R1732 GND.n434 GND.n433 2.759
R1733 GND.n609 GND.n608 2.759
R1734 GND.n51 GND.n50 2.759
R1735 GND.n97 GND.n96 2.759
R1736 GND.n135 GND.n134 2.759
R1737 GND.n88 GND.n87 2.759
R1738 GND.n203 GND.n202 2.612
R1739 GND.n212 GND.n211 2.562
R1740 GND.n388 GND.n387 2.562
R1741 GND.n563 GND.n562 2.562
R1742 GND.n6 GND.n5 2.562
R1743 GND.n202 GND.n2 2.562
R1744 GND.n205 GND 2.382
R1745 GND.n4 GND.n3 1.853
R1746 GND.n42 GND.n41 1.853
R1747 GND.n1 GND.n0 1.593
R1748 GND.n216 GND.n212 1.145
R1749 GND.n392 GND.n388 1.145
R1750 GND.n567 GND.n563 1.145
R1751 GND.n10 GND.n6 1.145
R1752 GND.n202 GND.n201 1.09
R1753 GND.n265 GND.n263 0.525
R1754 GND.n441 GND.n439 0.525
R1755 GND.n616 GND.n614 0.525
R1756 GND.n49 GND.n47 0.525
R1757 GND.n95 GND.n93 0.525
R1758 GND.n319 GND.n318 0.524
R1759 GND.n670 GND.n669 0.524
R1760 GND.n159 GND.n158 0.524
R1761 GND.n314 GND.n311 0.507
R1762 GND.n489 GND.n487 0.507
R1763 GND.n665 GND.n662 0.507
R1764 GND.n142 GND.n140 0.507
R1765 GND.n225 GND.n221 0.09
R1766 GND.n234 GND.n230 0.09
R1767 GND.n240 GND.n239 0.09
R1768 GND.n251 GND.n247 0.09
R1769 GND.n260 GND.n256 0.09
R1770 GND.n269 GND.n265 0.09
R1771 GND.n283 GND.n279 0.09
R1772 GND.n287 GND.n283 0.09
R1773 GND.n288 GND.n287 0.09
R1774 GND.n299 GND.n295 0.09
R1775 GND.n303 GND.n299 0.09
R1776 GND.n317 GND.n314 0.09
R1777 GND.n322 GND.n317 0.09
R1778 GND.n332 GND.n328 0.09
R1779 GND.n336 GND.n332 0.09
R1780 GND.n350 GND.n346 0.09
R1781 GND.n354 GND.n350 0.09
R1782 GND.n358 GND.n354 0.09
R1783 GND.n359 GND.n358 0.09
R1784 GND.n368 GND.n364 0.09
R1785 GND.n372 GND.n368 0.09
R1786 GND.n401 GND.n397 0.09
R1787 GND.n410 GND.n406 0.09
R1788 GND.n416 GND.n415 0.09
R1789 GND.n427 GND.n423 0.09
R1790 GND.n436 GND.n432 0.09
R1791 GND.n445 GND.n441 0.09
R1792 GND.n459 GND.n455 0.09
R1793 GND.n463 GND.n459 0.09
R1794 GND.n464 GND.n463 0.09
R1795 GND.n475 GND.n471 0.09
R1796 GND.n479 GND.n475 0.09
R1797 GND.n493 GND.n489 0.09
R1798 GND.n497 GND.n493 0.09
R1799 GND.n511 GND.n507 0.09
R1800 GND.n515 GND.n511 0.09
R1801 GND.n524 GND.n520 0.09
R1802 GND.n528 GND.n524 0.09
R1803 GND.n532 GND.n528 0.09
R1804 GND.n533 GND.n532 0.09
R1805 GND.n542 GND.n538 0.09
R1806 GND.n546 GND.n542 0.09
R1807 GND.n576 GND.n572 0.09
R1808 GND.n585 GND.n581 0.09
R1809 GND.n591 GND.n590 0.09
R1810 GND.n602 GND.n598 0.09
R1811 GND.n611 GND.n607 0.09
R1812 GND.n620 GND.n616 0.09
R1813 GND.n634 GND.n630 0.09
R1814 GND.n638 GND.n634 0.09
R1815 GND.n639 GND.n638 0.09
R1816 GND.n650 GND.n646 0.09
R1817 GND.n654 GND.n650 0.09
R1818 GND.n668 GND.n665 0.09
R1819 GND.n673 GND.n668 0.09
R1820 GND.n683 GND.n679 0.09
R1821 GND.n687 GND.n683 0.09
R1822 GND.n701 GND.n697 0.09
R1823 GND.n705 GND.n701 0.09
R1824 GND.n709 GND.n705 0.09
R1825 GND.n710 GND.n709 0.09
R1826 GND.n719 GND.n715 0.09
R1827 GND.n723 GND.n719 0.09
R1828 GND.n19 GND.n15 0.09
R1829 GND.n23 GND.n19 0.09
R1830 GND.n25 GND.n23 0.09
R1831 GND.n36 GND.n32 0.09
R1832 GND.n40 GND.n36 0.09
R1833 GND.n44 GND.n40 0.09
R1834 GND.n53 GND.n49 0.09
R1835 GND.n57 GND.n53 0.09
R1836 GND.n66 GND.n62 0.09
R1837 GND.n70 GND.n66 0.09
R1838 GND.n71 GND.n70 0.09
R1839 GND.n82 GND.n78 0.09
R1840 GND.n86 GND.n82 0.09
R1841 GND.n90 GND.n86 0.09
R1842 GND.n99 GND.n95 0.09
R1843 GND.n103 GND.n99 0.09
R1844 GND.n112 GND.n108 0.09
R1845 GND.n116 GND.n112 0.09
R1846 GND.n118 GND.n116 0.09
R1847 GND.n129 GND.n125 0.09
R1848 GND.n133 GND.n129 0.09
R1849 GND.n137 GND.n133 0.09
R1850 GND.n146 GND.n142 0.09
R1851 GND.n149 GND.n146 0.09
R1852 GND.n157 GND.n154 0.09
R1853 GND.n162 GND.n157 0.09
R1854 GND.n167 GND.n162 0.09
R1855 GND.n176 GND.n172 0.09
R1856 GND.n180 GND.n176 0.09
R1857 GND.n184 GND.n180 0.09
R1858 GND.n185 GND.n184 0.09
R1859 GND.n196 GND.n192 0.09
R1860 GND.n200 GND.n196 0.09
R1861 GND.n491 GND.n490 0.089
R1862 CMOS_s0_0/GND GND.n733 0.085
R1863 GND.n556 CMOS_s1_0/GND 0.085
R1864 GND.n381 CMOS_s2_0/GND 0.085
R1865 GND.n226 GND.n225 0.078
R1866 GND.n239 GND.n235 0.078
R1867 GND.n275 GND.n274 0.078
R1868 GND.n402 GND.n401 0.078
R1869 GND.n415 GND.n411 0.078
R1870 GND.n451 GND.n450 0.078
R1871 GND.n577 GND.n576 0.078
R1872 GND.n590 GND.n586 0.078
R1873 GND.n626 GND.n625 0.078
R1874 GND.n11 GND.n10 0.078
R1875 GND.n58 GND.n57 0.078
R1876 GND.n104 GND.n103 0.078
R1877 GND.n306 GND.n305 0.074
R1878 GND.n375 GND.n374 0.074
R1879 GND.n482 GND.n481 0.074
R1880 GND.n549 GND.n548 0.074
R1881 GND.n657 GND.n656 0.074
R1882 GND.n726 GND.n725 0.074
R1883 GND.n217 GND.n216 0.072
R1884 GND.n393 GND.n392 0.072
R1885 GND.n568 GND.n567 0.072
R1886 GND.n323 GND.n322 0.071
R1887 GND.n337 GND.n336 0.071
R1888 GND.n498 GND.n497 0.071
R1889 GND.n674 GND.n673 0.071
R1890 GND.n688 GND.n687 0.071
R1891 GND.n150 GND.n149 0.071
R1892 GND.n247 GND 0.065
R1893 GND.n274 GND.n270 0.065
R1894 GND.n295 CMOS_s3_0/CMOS_XOR_0/GND 0.065
R1895 GND.n346 GND.n342 0.065
R1896 GND.n364 CMOS_s3_0/CMOS_3in_AND_0/GND 0.065
R1897 GND.n423 CMOS_s2_0/CMOS_3in_OR_0/GND 0.065
R1898 GND.n450 GND.n446 0.065
R1899 GND.n471 CMOS_s2_0/CMOS_XOR_0/GND 0.065
R1900 GND.n520 GND.n516 0.065
R1901 GND.n538 CMOS_s2_0/CMOS_4in_AND_0/GND 0.065
R1902 GND.n598 CMOS_s1_0/CMOS_3in_OR_0/GND 0.065
R1903 GND.n625 GND.n621 0.065
R1904 GND.n646 CMOS_s1_0/CMOS_XOR_0/GND 0.065
R1905 GND.n697 GND.n693 0.065
R1906 GND.n715 CMOS_s1_0/CMOS_3in_AND_0/GND 0.065
R1907 GND.n32 CMOS_s0_0/CMOS_OR_0/GND 0.065
R1908 GND.n78 CMOS_s0_0/CMOS_AND_0/GND 0.065
R1909 GND.n125 CMOS_s0_0/CMOS_AND_2/GND 0.065
R1910 GND.n172 GND.n168 0.065
R1911 GND.n192 CMOS_s0_0/CMOS_XOR_0/GND 0.065
R1912 GND.n256 GND.n252 0.063
R1913 GND.n432 GND.n428 0.063
R1914 GND.n503 GND.n502 0.063
R1915 GND.n607 GND.n603 0.063
R1916 CMOS_s0_0/GND GND.n205 0.062
R1917 GND.n732 CMOS_s1_0/GND 0.062
R1918 GND.n555 CMOS_s2_0/GND 0.062
R1919 GND.n263 GND.n261 0.056
R1920 GND.n311 GND.n309 0.056
R1921 GND.n439 GND.n437 0.056
R1922 GND.n487 GND.n485 0.056
R1923 GND.n614 GND.n612 0.056
R1924 GND.n662 GND.n660 0.056
R1925 GND.n47 GND.n45 0.056
R1926 GND.n93 GND.n91 0.056
R1927 GND.n140 GND.n138 0.056
R1928 GND.n304 GND.n303 0.055
R1929 GND.n373 GND.n372 0.055
R1930 GND.n480 GND.n479 0.055
R1931 GND.n547 GND.n546 0.055
R1932 GND.n655 GND.n654 0.055
R1933 GND.n724 GND.n723 0.055
R1934 GND.n201 GND.n200 0.055
R1935 GND.n380 CMOS_s3_0/GND 0.048
R1936 GND.n267 GND.n266 0.047
R1937 GND.n443 GND.n442 0.047
R1938 GND.n618 GND.n617 0.047
R1939 GND.n308 GND.n304 0.035
R1940 GND.n377 GND.n373 0.035
R1941 GND.n484 GND.n480 0.035
R1942 GND.n551 GND.n547 0.035
R1943 GND.n659 GND.n655 0.035
R1944 GND.n728 GND.n724 0.035
R1945 GND.n261 GND.n260 0.033
R1946 GND.n309 GND.n308 0.033
R1947 GND.n378 GND.n377 0.033
R1948 GND.n437 GND.n436 0.033
R1949 GND.n485 GND.n484 0.033
R1950 GND.n552 GND.n551 0.033
R1951 GND.n612 GND.n611 0.033
R1952 GND.n660 GND.n659 0.033
R1953 GND.n729 GND.n728 0.033
R1954 GND.n45 GND.n44 0.033
R1955 GND.n91 GND.n90 0.033
R1956 GND.n138 GND.n137 0.033
R1957 GND.n252 GND.n251 0.026
R1958 GND.n428 GND.n427 0.026
R1959 GND.n507 GND.n503 0.026
R1960 GND.n603 GND.n602 0.026
R1961 GND.n240 GND 0.025
R1962 GND.n270 GND.n269 0.025
R1963 GND.n288 CMOS_s3_0/CMOS_XOR_0/GND 0.025
R1964 GND.n342 GND.n341 0.025
R1965 GND.n359 CMOS_s3_0/CMOS_3in_AND_0/GND 0.025
R1966 GND.n416 CMOS_s2_0/CMOS_3in_OR_0/GND 0.025
R1967 GND.n446 GND.n445 0.025
R1968 GND.n464 CMOS_s2_0/CMOS_XOR_0/GND 0.025
R1969 GND.n516 GND.n515 0.025
R1970 GND.n533 CMOS_s2_0/CMOS_4in_AND_0/GND 0.025
R1971 GND.n591 CMOS_s1_0/CMOS_3in_OR_0/GND 0.025
R1972 GND.n621 GND.n620 0.025
R1973 GND.n639 CMOS_s1_0/CMOS_XOR_0/GND 0.025
R1974 GND.n693 GND.n692 0.025
R1975 GND.n710 CMOS_s1_0/CMOS_3in_AND_0/GND 0.025
R1976 GND.n71 CMOS_s0_0/CMOS_AND_0/GND 0.025
R1977 GND.n168 GND.n167 0.025
R1978 GND.n185 CMOS_s0_0/CMOS_XOR_0/GND 0.025
R1979 GND.n328 GND.n323 0.018
R1980 GND.n341 GND.n337 0.018
R1981 GND.n502 GND.n498 0.018
R1982 GND.n679 GND.n674 0.018
R1983 GND.n692 GND.n688 0.018
R1984 GND.n25 GND.n24 0.018
R1985 GND.n118 GND.n117 0.018
R1986 GND.n154 GND.n150 0.018
R1987 GND.n221 GND.n217 0.017
R1988 GND.n397 GND.n393 0.017
R1989 GND.n572 GND.n568 0.017
R1990 GND.n230 GND.n226 0.011
R1991 GND.n235 GND.n234 0.011
R1992 GND.n279 GND.n275 0.011
R1993 GND.n406 GND.n402 0.011
R1994 GND.n411 GND.n410 0.011
R1995 GND.n455 GND.n451 0.011
R1996 GND.n581 GND.n577 0.011
R1997 GND.n586 GND.n585 0.011
R1998 GND.n630 GND.n626 0.011
R1999 GND.n15 GND.n11 0.011
R2000 GND.n62 GND.n58 0.011
R2001 GND.n108 GND.n104 0.011
R2002 GND.n24 CMOS_s0_0/CMOS_OR_0/GND 0.006
R2003 GND.n117 CMOS_s0_0/CMOS_AND_2/GND 0.006
R2004 x0_bar.t7 x0_bar.t6 1345.61
R2005 x0_bar.t9 x0_bar.t8 1345.61
R2006 x0_bar.n3 x0_bar.t3 683.32
R2007 x0_bar.n1 x0_bar.t1 681.713
R2008 x0_bar.n4 x0_bar.t5 616.084
R2009 x0_bar.n6 x0_bar.t4 570.366
R2010 x0_bar.n6 x0_bar.t2 570.366
R2011 x0_bar.n3 x0_bar.t10 528.72
R2012 x0_bar.n4 x0_bar.t0 528.72
R2013 x0_bar.n1 x0_bar.t11 528.72
R2014 x0_bar.n8 CMOS_s1_0/CMOS_XNOR_0/A_bar 507.08
R2015 x0_bar.n0 CMOS_s0_0/CMOS_XOR_0/A_bar 507.08
R2016 CMOS_s1_0/CMOS_XNOR_0/A_bar x0_bar.t7 392.02
R2017 CMOS_s0_0/CMOS_XOR_0/A_bar x0_bar.t9 392.02
R2018 CMOS_s3_0/x0_bar x0_bar 346.044
R2019 x0_bar.n2 CMOS_s0_0/CMOS_XNOR_0/B_bar 344.84
R2020 x0_bar.n7 CMOS_s1_0/CMOS_3in_AND_0/C 337.8
R2021 CMOS_s1_0/CMOS_3in_AND_0/C x0_bar.n6 78.72
R2022 x0_bar.n5 x0_bar.n4 14.546
R2023 x0_bar x0_bar.n3 3.68
R2024 x0_bar.n4 CMOS_s2_0/CMOS_XOR_0/B_bar 3.68
R2025 CMOS_s0_0/CMOS_XNOR_0/B_bar x0_bar.n1 3.68
R2026 x0_bar.n5 CMOS_s3_0/x0_bar 2.872
R2027 x0_bar.n0 CMOS_s0_0/x0_bar 2.169
R2028 CMOS_s1_0/x0_bar x0_bar.n8 2.166
R2029 CMOS_s2_0/x0_bar x0_bar.n5 2.163
R2030 x0_bar.n7 CMOS_s2_0/x0_bar 1.582
R2031 CMOS_s1_0/x0_bar x0_bar.n2 1.557
R2032 x0_bar.n2 x0_bar.n0 1.317
R2033 x0_bar.n8 x0_bar.n7 1.292
R2034 s1.n2 s1.t1 120.552
R2035 s1.n1 s1.t0 98.438
R2036 s1 s1.n2 7.84
R2037 s1 s1.n1 3.68
R2038 s1.n1 s1.n0 3.084
R2039 s1.n0 CMOS_s1_0/s1 0.374
R2040 x0.t1 x0.t12 1221.07
R2041 x0.n7 x0.t5 993.097
R2042 x0.n0 x0.t2 993.097
R2043 x0.t13 x0.t9 924.95
R2044 x0.t3 x0.t0 924.95
R2045 x0.t10 x0.t4 923.343
R2046 CMOS_s3_0/CMOS_XNOR_0/B x0.t13 633.02
R2047 CMOS_s2_0/CMOS_XOR_0/B x0.t3 633.02
R2048 CMOS_s0_0/CMOS_XNOR_0/B x0.t10 633.02
R2049 x0.n4 x0.t11 570.366
R2050 x0.n4 x0.t6 570.366
R2051 x0.n3 CMOS_s3_0/CMOS_XNOR_0/B 535.88
R2052 x0.n2 CMOS_s0_0/CMOS_XNOR_0/B 535.88
R2053 x0.n3 x0 428.025
R2054 x0.n5 CMOS_s2_0/CMOS_4in_AND_0/C 422.28
R2055 x0 x0.t1 392.02
R2056 x0.n8 CMOS_s1_0/CMOS_XNOR_0/A 391.88
R2057 x0.n1 CMOS_s0_0/CMOS_XOR_0/A 391.88
R2058 x0.n7 x0.t8 356.59
R2059 x0.n0 x0.t7 356.59
R2060 CMOS_s2_0/CMOS_4in_AND_0/C x0.n4 78.72
R2061 CMOS_s1_0/CMOS_XNOR_0/A x0.n7 78.72
R2062 CMOS_s0_0/CMOS_XOR_0/A x0.n0 78.72
R2063 x0.n6 CMOS_s2_0/CMOS_XOR_0/B 45.03
R2064 x0.n8 CMOS_s2_0/x0 3.444
R2065 x0.n6 x0.n5 3.393
R2066 x0.n2 x0.n1 3.128
R2067 x0.n1 CMOS_s0_0/x0 1.597
R2068 CMOS_s1_0/x0 x0.n8 1.597
R2069 x0.n5 CMOS_s3_0/x0 1.487
R2070 CMOS_s1_0/x0 x0.n2 0.315
R2071 CMOS_s2_0/x0 x0.n6 0.156
R2072 CMOS_s3_0/x0 x0.n3 0.152
R2073 x3_bar.t6 x3_bar.t1 1345.61
R2074 x3_bar.t8 x3_bar.t15 1345.61
R2075 x3_bar.t11 x3_bar.t14 1221.07
R2076 x3_bar.n7 x3_bar.t13 811.366
R2077 x3_bar.n0 x3_bar.t2 683.32
R2078 x3_bar.n10 x3_bar.t11 630.3
R2079 x3_bar.n5 x3_bar.t7 616.084
R2080 x3_bar.n12 x3_bar.t4 616.084
R2081 x3_bar.n3 x3_bar.t3 579.86
R2082 x3_bar.n3 x3_bar.t12 547.727
R2083 x3_bar.n5 x3_bar.t10 528.72
R2084 x3_bar.n12 x3_bar.t9 528.72
R2085 x3_bar.n0 x3_bar.t5 528.72
R2086 CMOS_s2_0/CMOS_XNOR_0/A_bar x3_bar.t6 392.02
R2087 CMOS_s0_0/CMOS_XNOR_0/A_bar x3_bar.t8 392.02
R2088 x3_bar.n7 x3_bar.t0 329.366
R2089 x3_bar.n9 CMOS_s2_0/CMOS_XNOR_0/A_bar 286.14
R2090 x3_bar.n2 CMOS_s0_0/CMOS_XNOR_0/A_bar 286.14
R2091 x3_bar.n8 CMOS_s2_0/CMOS_4in_AND_0/A 264.208
R2092 x3_bar.n1 CMOS_s0_0/CMOS_XOR_0/B_bar 125.96
R2093 CMOS_s2_0/CMOS_4in_AND_0/A x3_bar.n7 78.72
R2094 x3_bar.n11 x3_bar.n10 38.547
R2095 x3_bar.n6 x3_bar.n5 12.409
R2096 x3_bar.n13 x3_bar.n12 12.409
R2097 x3_bar.n6 x3_bar.n4 11.74
R2098 x3_bar.n4 x3_bar.n3 8.764
R2099 x3_bar.n5 x3_bar 3.68
R2100 x3_bar.n12 CMOS_s1_0/CMOS_XOR_0/B_bar 3.68
R2101 CMOS_s0_0/CMOS_XOR_0/B_bar x3_bar.n0 3.68
R2102 x3_bar.n4 CMOS_s3_0/CMOS_AND_1/B 2.72
R2103 x3_bar.n10 CMOS_s1_0/CMOS_3in_AND_0/A 2.72
R2104 CMOS_s1_0/x3_bar x3_bar.n2 2.459
R2105 x3_bar.n13 x3_bar.n11 2.458
R2106 CMOS_s1_0/x3_bar x3_bar.n13 2.167
R2107 CMOS_s3_0/x3_bar x3_bar.n6 2.167
R2108 CMOS_s2_0/x3_bar x3_bar.n9 2.112
R2109 x3_bar.n8 CMOS_s3_0/x3_bar 1.82
R2110 x3_bar.n2 x3_bar.n1 1.375
R2111 x3_bar.n1 CMOS_s0_0/x3_bar 1.205
R2112 x3_bar.n9 x3_bar.n8 1.109
R2113 x3_bar.n11 CMOS_s2_0/x3_bar 0.403
R2114 x2_bar.t13 x2_bar.t8 1345.61
R2115 x2_bar.t5 x2_bar.t0 1221.07
R2116 x2_bar.t7 x2_bar.t2 1221.07
R2117 x2_bar.n8 x2_bar.t12 683.32
R2118 x2_bar.n11 x2_bar.t6 683.32
R2119 x2_bar.n5 x2_bar.t5 630.3
R2120 x2_bar.n3 x2_bar.t3 579.86
R2121 x2_bar.n1 x2_bar.t10 579.86
R2122 x2_bar.n3 x2_bar.t1 547.727
R2123 x2_bar.n1 x2_bar.t9 547.727
R2124 x2_bar.n8 x2_bar.t4 528.72
R2125 x2_bar.n11 x2_bar.t11 528.72
R2126 CMOS_s3_0/CMOS_XOR_0/A_bar x2_bar.t13 392.02
R2127 CMOS_s0_0/CMOS_OR_1/B x2_bar.t7 392.02
R2128 x2_bar.n0 CMOS_s0_0/CMOS_OR_1/B 285.69
R2129 x2_bar.n9 CMOS_s2_0/CMOS_XNOR_0/B_bar 198.92
R2130 x2_bar.n12 CMOS_s1_0/CMOS_XNOR_0/B_bar 198.92
R2131 x2_bar.n6 CMOS_s3_0/CMOS_XOR_0/A_bar 44.234
R2132 x2_bar.n6 x2_bar.n5 41.121
R2133 x2_bar.n7 x2_bar.n4 17.994
R2134 x2_bar.n10 x2_bar.n2 17.994
R2135 x2_bar.n4 x2_bar.n3 8.764
R2136 x2_bar.n2 x2_bar.n1 8.764
R2137 CMOS_s2_0/CMOS_XNOR_0/B_bar x2_bar.n8 3.68
R2138 CMOS_s1_0/CMOS_XNOR_0/B_bar x2_bar.n11 3.68
R2139 CMOS_s1_0/x2_bar x2_bar.n0 2.877
R2140 CMOS_s3_0/x2_bar x2_bar.n6 2.762
R2141 x2_bar.n5 x2_bar 2.72
R2142 x2_bar.n4 CMOS_s2_0/CMOS_AND_0/B 2.72
R2143 x2_bar.n2 CMOS_s1_0/CMOS_AND_0/B 2.72
R2144 x2_bar.n0 CMOS_s0_0/x2_bar 2.16
R2145 x2_bar.n10 CMOS_s2_0/x2_bar 2.132
R2146 x2_bar.n7 CMOS_s3_0/x2_bar 2.132
R2147 x2_bar.n12 x2_bar.n10 1.697
R2148 x2_bar.n9 x2_bar.n7 1.697
R2149 CMOS_s1_0/x2_bar x2_bar.n12 1.205
R2150 CMOS_s2_0/x2_bar x2_bar.n9 1.205
R2151 x2.t0 x2.t3 1221.07
R2152 x2.t6 x2.t2 1221.07
R2153 x2.n0 x2.t7 993.097
R2154 x2.t1 x2.t9 924.95
R2155 x2.t8 x2.t5 924.95
R2156 CMOS_s2_0/CMOS_4in_AND_0/D x2.t0 633.02
R2157 CMOS_s2_0/CMOS_XNOR_0/B x2.t1 633.02
R2158 CMOS_s1_0/CMOS_XNOR_0/B x2.t8 633.02
R2159 CMOS_s0_0/CMOS_AND_2/A x2.t6 392.02
R2160 x2.n3 CMOS_s2_0/CMOS_XNOR_0/B 389.96
R2161 x2.n4 CMOS_s1_0/CMOS_XNOR_0/B 389.96
R2162 x2.n0 x2.t4 356.59
R2163 x2.n2 CMOS_s2_0/CMOS_4in_AND_0/D 228.36
R2164 x2.n5 CMOS_s0_0/CMOS_AND_2/A 214.75
R2165 CMOS_s3_0/x2 x2.n1 16.257
R2166 x2.n1 x2.n0 8.764
R2167 x2.n4 CMOS_s2_0/x2 4.888
R2168 x2.n3 x2.n2 4.574
R2169 x2.n1 x2 2.72
R2170 x2 x2.n5 2.621
R2171 x2.n5 CMOS_s1_0/x2 2.412
R2172 x2.n2 CMOS_s3_0/x2 0.313
R2173 CMOS_s1_0/x2 x2.n4 0.154
R2174 CMOS_s2_0/x2 x2.n3 0.154
R2175 CMOS_s0_0/x2 x2 0.001
R2176 CMOS_s1_0/CMOS_3in_OR_0/C.t2 CMOS_s1_0/CMOS_3in_OR_0/C.t3 1221.07
R2177 CMOS_s1_0/CMOS_3in_OR_0/C CMOS_s1_0/CMOS_3in_OR_0/C.n0 787.238
R2178 CMOS_s1_0/CMOS_3in_OR_0/C CMOS_s1_0/CMOS_3in_OR_0/C.t2 633.02
R2179 CMOS_s1_0/CMOS_3in_AND_0/OUT CMOS_s1_0/CMOS_3in_OR_0/C.t0 117.958
R2180 CMOS_s1_0/CMOS_3in_OR_0/C.n0 CMOS_s1_0/CMOS_3in_AND_0/OUT 91.717
R2181 CMOS_s1_0/CMOS_3in_OR_0/C.n0 CMOS_s1_0/CMOS_3in_OR_0/C.t1 45.156
R2182 x1.t7 x1.t2 1221.07
R2183 x1.t12 x1.t8 1221.07
R2184 x1.n2 x1.t5 993.097
R2185 x1.n4 x1.t13 993.097
R2186 x1.n8 x1.t3 993.097
R2187 x1.n0 x1.t11 579.86
R2188 x1.n12 x1.t4 579.86
R2189 x1.n0 x1.t10 547.727
R2190 x1.n12 x1.t0 547.727
R2191 x1.n13 CMOS_s0_0/CMOS_OR_1/A 451.88
R2192 x1.n7 CMOS_s2_0/CMOS_4in_AND_0/B 400.52
R2193 x1.n6 x1.t7 389.3
R2194 x1.n10 x1.t12 389.3
R2195 x1.n2 x1.t6 356.59
R2196 x1.n4 x1.t9 356.59
R2197 x1.n8 x1.t1 356.59
R2198 x1.n11 CMOS_s1_0/CMOS_3in_AND_0/B 352.52
R2199 x1.n3 CMOS_s3_0/CMOS_XNOR_0/A 318.92
R2200 x1.n10 x1.n9 211.594
R2201 x1.n6 x1.n5 183.874
R2202 CMOS_s3_0/CMOS_XNOR_0/A x1.n2 78.72
R2203 CMOS_s0_0/CMOS_OR_1/A x1.n12 78.72
R2204 x1.n3 x1.n1 20.982
R2205 x1.n1 x1.n0 8.764
R2206 x1.n5 x1.n4 8.764
R2207 x1.n9 x1.n8 8.764
R2208 x1.n13 CMOS_s1_0/x1 4.88
R2209 x1.n1 x1 2.72
R2210 x1.n5 CMOS_s2_0/CMOS_XOR_0/A 2.72
R2211 CMOS_s2_0/CMOS_4in_AND_0/B x1.n6 2.72
R2212 x1.n9 CMOS_s1_0/CMOS_XOR_0/A 2.72
R2213 CMOS_s1_0/CMOS_3in_AND_0/B x1.n10 2.72
R2214 CMOS_s1_0/x1 x1.n11 2.699
R2215 CMOS_s2_0/x1 x1.n7 2.699
R2216 x1.n11 CMOS_s2_0/x1 2.343
R2217 x1.n7 CMOS_s3_0/x1 2.343
R2218 CMOS_s3_0/x1 x1.n3 1.597
R2219 x1 x1.n13 0.154
R2220 CMOS_s0_0/x1 x1 0.001
R2221 CMOS_s3_0/CMOS_3in_OR_0/C.t2 CMOS_s3_0/CMOS_3in_OR_0/C.t3 1221.07
R2222 CMOS_s3_0/CMOS_3in_OR_0/C CMOS_s3_0/CMOS_3in_OR_0/C.n0 787.238
R2223 CMOS_s3_0/CMOS_3in_OR_0/C CMOS_s3_0/CMOS_3in_OR_0/C.t2 633.02
R2224 CMOS_s3_0/CMOS_3in_AND_0/OUT CMOS_s3_0/CMOS_3in_OR_0/C.t0 117.958
R2225 CMOS_s3_0/CMOS_3in_OR_0/C.n0 CMOS_s3_0/CMOS_3in_AND_0/OUT 91.717
R2226 CMOS_s3_0/CMOS_3in_OR_0/C.n0 CMOS_s3_0/CMOS_3in_OR_0/C.t1 45.156
R2227 s0 s0.t1 117.353
R2228 s0.n0 s0.t0 95.65
R2229 s0 s0.n0 10.009
R2230 s0.n0 CMOS_s0_0/s0 0.913
R2231 x1_bar.t9 x1_bar.t7 1345.61
R2232 x1_bar.t2 x1_bar.t8 1345.61
R2233 x1_bar.t6 x1_bar.t4 1345.61
R2234 x1_bar.n2 x1_bar.t5 579.86
R2235 x1_bar.n0 x1_bar.t1 579.86
R2236 x1_bar.n2 x1_bar.t3 547.727
R2237 x1_bar.n0 x1_bar.t0 547.727
R2238 CMOS_s3_0/x1_bar x1_bar 436.286
R2239 x1_bar x1_bar.t9 392.02
R2240 CMOS_s2_0/CMOS_XOR_0/A_bar x1_bar.t2 392.02
R2241 CMOS_s1_0/CMOS_XOR_0/A_bar x1_bar.t6 392.02
R2242 x1_bar.n1 CMOS_s0_0/CMOS_AND_2/B 380.225
R2243 CMOS_s0_0/CMOS_AND_2/B x1_bar.n0 78.72
R2244 x1_bar.n5 CMOS_s2_0/CMOS_XOR_0/A_bar 44.915
R2245 x1_bar.n6 CMOS_s1_0/CMOS_XOR_0/A_bar 44.915
R2246 x1_bar.n4 x1_bar.n3 11.862
R2247 x1_bar.n3 x1_bar.n2 8.764
R2248 x1_bar.n1 CMOS_s0_0/x1_bar 4.631
R2249 x1_bar.n3 CMOS_s2_0/CMOS_AND_1/B 2.72
R2250 CMOS_s1_0/x1_bar x1_bar.n6 2.663
R2251 CMOS_s2_0/x1_bar x1_bar.n5 2.663
R2252 x1_bar.n6 CMOS_s2_0/x1_bar 2.372
R2253 x1_bar.n4 CMOS_s3_0/x1_bar 1.561
R2254 x1_bar.n5 x1_bar.n4 0.803
R2255 CMOS_s1_0/x1_bar x1_bar.n1 0.406
R2256 s3.n2 s3.t1 120.552
R2257 s3.n1 s3.t0 98.438
R2258 s3 s3.n2 7.84
R2259 s3 s3.n1 3.68
R2260 s3.n1 s3.n0 3.084
R2261 s3.n0 CMOS_s3_0/s3 0.374
R2262 s2.n2 s2.t1 120.552
R2263 s2.n1 s2.t0 98.438
R2264 s2 s2.n2 7.84
R2265 s2 s2.n1 3.68
R2266 s2.n1 s2.n0 3.084
R2267 s2.n0 CMOS_s2_0/s2 0.374
C0 a_n1990_n1580# x1 0.00fF
C1 CMOS_s1_0/CMOS_3in_OR_0/B CMOS_s1_0/CMOS_3in_OR_0/C 0.06fF
C2 CMOS_s3_0/CMOS_XOR_0/XOR CMOS_s3_0/CMOS_3in_OR_0/A 0.02fF
C3 VDD a_n2195_n9314# 0.01fF
C4 a_n2345_n6996# x3 0.06fF
C5 VDD a_n1990_n540# 0.04fF
C6 a_n787_n6996# CMOS_s2_0/CMOS_3in_OR_0/A 0.07fF
C7 a_n2140_n5418# CMOS_s2_0/CMOS_AND_1/A 0.08fF
C8 CMOS_s3_0/CMOS_3in_OR_0/B a_575_n10224# 0.00fF
C9 a_n732_n1580# CMOS_s1_0/CMOS_AND_1/A 0.01fF
C10 CMOS_s3_0/CMOS_3in_OR_0/B a_n732_n8646# 0.00fF
C11 CMOS_s0_0/CMOS_AND_1/B a_425_n540# 0.04fF
C12 a_n787_n6996# a_n732_n5418# 0.00fF
C13 a_n432_n2190# x3 0.01fF
C14 a_n2290_n8036# a_n2140_n8646# 0.02fF
C15 VDD CMOS_s2_0/CMOS_3in_OR_0/A 0.56fF
C16 CMOS_s0_0/CMOS_AND_0/B x1 0.00fF
C17 VDD a_n732_n5418# 0.01fF
C18 a_n2290_1648# CMOS_s0_0/CMOS_XOR_0/XOR 0.02fF
C19 a_n2345_n9314# CMOS_s3_0/CMOS_3in_OR_0/C 0.00fF
C20 VDD CMOS_s0_0/CMOS_XOR_0/XOR 1.15fF
C21 a_n732_n1580# CMOS_s0_0/CMOS_AND_1/B 0.00fF
C22 a_n787_n540# CMOS_s0_0/CMOS_AND_1/AND 0.00fF
C23 a_n732_n8646# x2 0.00fF
C24 a_n1990_n2190# CMOS_s1_0/CMOS_XOR_0/XOR 0.00fF
C25 a_n732_n2190# a_n2140_n2190# 0.00fF
C26 a_n2495_n10224# x2 0.02fF
C27 CMOS_s2_0/CMOS_4in_AND_0/OUT a_n432_n8646# 0.00fF
C28 a_n2345_n6996# a_n787_n6086# 0.00fF
C29 CMOS_s0_0/CMOS_AND_0/AND a_1637_1038# 0.05fF
C30 VDD a_n1990_n2190# 0.01fF
C31 a_n2290_n5418# x2 0.01fF
C32 a_n732_n8646# x3 0.01fF
C33 a_425_n5418# x1 0.00fF
C34 a_n2495_n10224# x3 0.09fF
C35 VDD a_n787_370# 0.01fF
C36 a_425_n8036# a_n432_n8646# 0.00fF
C37 VDD a_425_n4808# 0.82fF
C38 a_n2290_n2190# VDD 0.01fF
C39 VDD CMOS_s3_0/CMOS_3in_OR_0/C 2.11fF
C40 a_n2290_n5418# x3 0.00fF
C41 a_n2495_n3768# CMOS_s1_0/CMOS_3in_OR_0/A 0.00fF
C42 a_n2140_n5418# x1 0.05fF
C43 a_275_n2858# CMOS_s2_0/CMOS_3in_OR_0/B 0.01fF
C44 a_n732_n8036# CMOS_s3_0/CMOS_3in_OR_0/B 0.00fF
C45 a_n2140_n8646# x2 0.05fF
C46 CMOS_s2_0/CMOS_4in_AND_0/OUT a_275_n6086# 0.05fF
C47 VDD a_425_1038# 0.01fF
C48 VDD a_n1990_1648# 0.05fF
C49 a_275_n9314# a_n787_n10224# 0.01fF
C50 a_n2140_n8646# x3 0.17fF
C51 a_425_n8036# a_275_n6086# 0.00fF
C52 a_n787_n540# a_n2290_n540# 0.00fF
C53 x1 a_425_n8646# 0.01fF
C54 CMOS_s0_0/CMOS_AND_1/AND a_425_370# 0.00fF
C55 a_n732_n8036# x3 0.01fF
C56 a_n732_n8646# a_n787_n10224# 0.00fF
C57 a_425_n10224# CMOS_s3_0/CMOS_3in_OR_0/A 0.01fF
C58 a_575_n10224# a_n787_n10224# 0.00fF
C59 a_425_n3768# a_275_n2858# 0.02fF
C60 a_n2495_n10224# a_n787_n10224# 0.00fF
C61 a_n787_n540# CMOS_s1_0/CMOS_XOR_0/XOR 0.00fF
C62 a_425_n5418# CMOS_s1_0/CMOS_3in_OR_0/C 0.00fF
C63 CMOS_s0_0/CMOS_AND_1/A a_425_1648# 0.00fF
C64 VDD a_n787_n540# 0.83fF
C65 VDD a_n2495_n3768# 1.44fF
C66 a_575_n3768# a_275_n2858# 0.02fF
C67 a_n2140_n5418# CMOS_s1_0/CMOS_3in_OR_0/C 0.01fF
C68 CMOS_s3_0/CMOS_AND_1/A CMOS_s3_0/CMOS_3in_OR_0/C 0.02fF
C69 a_n2345_n2858# a_n2495_n3768# 0.01fF
C70 a_n732_n4808# a_425_n4808# 0.00fF
C71 VDD a_n1990_n4808# 0.05fF
C72 CMOS_s0_0/CMOS_AND_0/AND CMOS_s0_0/CMOS_XOR_0/XOR 0.00fF
C73 a_n1990_n5418# CMOS_s2_0/CMOS_AND_1/A 0.00fF
C74 CMOS_s3_0/CMOS_XOR_0/XOR a_425_n10224# 0.00fF
C75 a_n432_n5418# a_425_n4808# 0.00fF
C76 CMOS_s3_0/CMOS_XOR_0/XOR a_425_n8646# 0.01fF
C77 CMOS_s1_0/CMOS_AND_1/A a_275_n2858# 0.00fF
C78 VDD a_n2290_n8036# 0.05fF
C79 a_425_n2190# x1 0.00fF
C80 a_n787_n9314# x1 0.01fF
C81 a_n732_n8036# a_n787_n10224# 0.00fF
C82 a_275_n6086# CMOS_s2_0/CMOS_AND_1/A 0.00fF
C83 a_n2345_n6996# a_n1990_n8646# 0.00fF
C84 CMOS_s1_0/CMOS_3in_OR_0/B a_425_n2190# 0.01fF
C85 a_n2140_n540# a_n2140_n2190# 0.02fF
C86 CMOS_s1_0/CMOS_3in_OR_0/A x3 0.02fF
C87 x1 a_425_1648# 0.00fF
C88 CMOS_s0_0/CMOS_AND_1/AND a_425_n540# 0.05fF
C89 a_n787_n9314# CMOS_s3_0/CMOS_3in_OR_0/A 0.00fF
C90 a_n1990_370# CMOS_s0_0/CMOS_AND_1/B 0.00fF
C91 a_n787_1648# CMOS_s0_0/CMOS_XOR_0/XOR 0.02fF
C92 a_n2345_n9314# x2 0.00fF
C93 VDD a_425_370# 0.01fF
C94 CMOS_s1_0/CMOS_AND_1/A CMOS_s0_0/CMOS_AND_1/B 0.00fF
C95 a_n2290_n540# x2 0.01fF
C96 a_n2195_n6086# a_n2345_n6996# 0.01fF
C97 CMOS_s0_0/CMOS_AND_0/AND a_425_1038# 0.00fF
C98 x1 a_n432_n8646# 0.01fF
C99 VDD CMOS_s3_0/CMOS_3in_OR_0/B 0.51fF
C100 a_n787_1038# a_n2290_1648# 0.00fF
C101 CMOS_s1_0/CMOS_3in_OR_0/A CMOS_s2_0/CMOS_XOR_0/XOR 0.00fF
C102 VDD a_n787_1038# 0.51fF
C103 a_n2290_1038# CMOS_s0_0/CMOS_XOR_0/XOR 0.01fF
C104 a_n2345_n9314# x3 0.00fF
C105 VDD a_n1990_1038# 0.01fF
C106 a_n2290_n540# x3 0.00fF
C107 a_n787_n6996# x2 0.00fF
C108 CMOS_s2_0/CMOS_4in_AND_0/OUT CMOS_s2_0/CMOS_3in_OR_0/A 0.10fF
C109 a_n1990_n5418# x1 0.00fF
C110 VDD a_n2290_n1580# 0.05fF
C111 CMOS_s1_0/CMOS_XOR_0/XOR x2 0.00fF
C112 a_n2290_1648# x2 0.00fF
C113 a_n732_n5418# a_n787_n3768# 0.00fF
C114 a_n1990_n8646# a_n2495_n10224# 0.00fF
C115 VDD x2 3.33fF
C116 a_n787_n6996# x3 0.03fF
C117 CMOS_s1_0/CMOS_XOR_0/XOR x3 0.35fF
C118 a_n2290_1648# x3 0.02fF
C119 a_n2290_n4808# a_n2495_n3768# 0.00fF
C120 a_n787_n540# a_n732_n2190# 0.00fF
C121 CMOS_s1_0/CMOS_AND_1/A a_n432_n2190# 0.00fF
C122 VDD x3 5.44fF
C123 a_275_n6086# x1 0.00fF
C124 VDD a_n2195_n2858# 0.01fF
C125 a_n2345_n2858# x2 0.00fF
C126 CMOS_s3_0/CMOS_AND_1/A a_n2290_n8036# 0.00fF
C127 a_n787_n6996# CMOS_s2_0/CMOS_XOR_0/XOR 0.01fF
C128 CMOS_s2_0/CMOS_4in_AND_0/OUT a_425_n4808# 0.00fF
C129 a_n2345_n2858# x3 0.00fF
C130 a_n787_n6996# a_n787_n6086# 0.01fF
C131 VDD CMOS_s2_0/CMOS_XOR_0/XOR 1.07fF
C132 CMOS_s3_0/CMOS_XOR_0/XOR a_n432_n8646# 0.01fF
C133 a_n1990_n8646# a_n2140_n8646# 0.01fF
C134 a_n2140_n540# a_n1990_n540# 0.03fF
C135 VDD a_n787_n6086# 0.00fF
C136 a_425_n540# CMOS_s1_0/CMOS_XOR_0/XOR 0.00fF
C137 a_425_n8036# CMOS_s3_0/CMOS_3in_OR_0/C 0.00fF
C138 a_n2140_n2190# x1 0.04fF
C139 CMOS_s3_0/CMOS_AND_1/A CMOS_s3_0/CMOS_3in_OR_0/B 0.01fF
C140 VDD a_425_n540# 0.83fF
C141 a_n2195_n6086# a_n2140_n8646# 0.00fF
C142 CMOS_s0_0/CMOS_AND_0/B a_425_1648# 0.04fF
C143 a_n787_n540# a_n787_1648# 0.00fF
C144 a_n732_n1580# CMOS_s1_0/CMOS_XOR_0/XOR 0.02fF
C145 a_n2140_n540# CMOS_s0_0/CMOS_XOR_0/XOR 0.03fF
C146 VDD a_n732_n1580# 0.06fF
C147 CMOS_s3_0/CMOS_XOR_0/XOR a_275_n6086# 0.00fF
C148 CMOS_s3_0/CMOS_AND_1/A x2 0.07fF
C149 VDD a_n787_n10224# 0.75fF
C150 CMOS_s3_0/CMOS_AND_1/A x3 0.03fF
C151 a_n2140_n540# a_n787_370# 0.00fF
C152 CMOS_s2_0/CMOS_3in_OR_0/A CMOS_s2_0/CMOS_AND_1/A 0.00fF
C153 a_425_n6996# a_n787_n6996# 0.00fF
C154 a_n732_n5418# CMOS_s2_0/CMOS_AND_1/A 0.00fF
C155 a_n2495_n3768# a_n787_n3768# 0.00fF
C156 CMOS_s0_0/CMOS_AND_0/AND a_n787_1038# 0.00fF
C157 CMOS_s0_0/CMOS_AND_1/A CMOS_s0_0/CMOS_XOR_0/XOR 0.07fF
C158 a_425_n6996# VDD 0.06fF
C159 a_n2290_n4808# x2 0.02fF
C160 a_n2140_n2190# CMOS_s1_0/CMOS_3in_OR_0/C 0.01fF
C161 a_n2345_n6996# a_n2290_n5418# 0.00fF
C162 a_275_n9314# a_575_n10224# 0.02fF
C163 a_n1990_n1580# a_n2140_n2190# 0.03fF
C164 CMOS_s0_0/CMOS_AND_1/A a_n787_370# 0.00fF
C165 a_n732_n4808# CMOS_s2_0/CMOS_XOR_0/XOR 0.02fF
C166 a_n2140_n540# a_n1990_1648# 0.00fF
C167 a_n2290_n4808# x3 0.00fF
C168 a_425_n3768# CMOS_s1_0/CMOS_3in_OR_0/A 0.01fF
C169 a_n787_n6996# CMOS_s2_0/CMOS_3in_OR_0/B 0.00fF
C170 a_n732_n2190# x3 0.01fF
C171 a_n2140_n5418# a_n1990_n5418# 0.01fF
C172 a_n432_n5418# CMOS_s2_0/CMOS_XOR_0/XOR 0.01fF
C173 a_n2195_n9314# x1 0.01fF
C174 a_425_n5418# a_275_n6086# 0.00fF
C175 a_n1990_n540# x1 0.00fF
C176 a_n2345_n6996# a_n2140_n8646# 0.01fF
C177 VDD CMOS_s2_0/CMOS_3in_OR_0/B 0.52fF
C178 a_n432_n8036# CMOS_s3_0/CMOS_3in_OR_0/B 0.00fF
C179 a_n787_1038# a_n787_1648# 0.01fF
C180 a_575_n3768# CMOS_s1_0/CMOS_3in_OR_0/A 0.00fF
C181 CMOS_s0_0/CMOS_AND_0/B a_1637_1038# 0.00fF
C182 a_425_n1580# a_425_370# 0.00fF
C183 CMOS_s3_0/CMOS_AND_1/A a_n787_n10224# 0.05fF
C184 CMOS_s0_0/CMOS_AND_1/A a_425_1038# 0.00fF
C185 CMOS_s2_0/CMOS_3in_OR_0/A x1 0.00fF
C186 a_n787_1038# a_n2290_1038# 0.00fF
C187 a_n787_n540# a_n2140_n540# 0.02fF
C188 a_n732_n5418# x1 0.00fF
C189 x2 a_n787_1648# 0.00fF
C190 x1 CMOS_s0_0/CMOS_XOR_0/XOR 0.21fF
C191 a_n432_n4808# a_425_n4808# 0.00fF
C192 a_275_n2858# CMOS_s1_0/CMOS_3in_OR_0/A 0.10fF
C193 CMOS_s0_0/CMOS_AND_1/AND CMOS_s0_0/CMOS_AND_1/B 0.00fF
C194 a_n1990_n2190# x1 0.00fF
C195 a_n2290_1038# x2 0.00fF
C196 a_425_n3768# CMOS_s1_0/CMOS_XOR_0/XOR 0.00fF
C197 CMOS_s1_0/CMOS_AND_1/A CMOS_s1_0/CMOS_3in_OR_0/A 0.00fF
C198 a_n432_n8036# x3 0.03fF
C199 a_n732_n8646# a_n2140_n8646# 0.00fF
C200 VDD a_425_n3768# 0.06fF
C201 x1 a_425_n4808# 0.00fF
C202 a_n2140_n8646# a_n2495_n10224# 0.01fF
C203 a_425_n8036# CMOS_s3_0/CMOS_3in_OR_0/B 0.08fF
C204 VDD a_n1990_n8646# 0.01fF
C205 a_n2290_1038# x3 0.01fF
C206 a_n2290_n2190# x1 0.00fF
C207 a_n2195_n6086# a_n787_n6996# 0.00fF
C208 a_n787_n540# CMOS_s0_0/CMOS_AND_1/A 0.05fF
C209 CMOS_s3_0/CMOS_3in_OR_0/C x1 0.03fF
C210 CMOS_s2_0/CMOS_4in_AND_0/OUT x2 0.01fF
C211 a_425_n1580# x3 0.01fF
C212 CMOS_s1_0/CMOS_3in_OR_0/B a_425_n4808# 0.00fF
C213 a_n2195_n6086# VDD 0.01fF
C214 VDD a_575_n3768# 0.06fF
C215 CMOS_s2_0/CMOS_4in_AND_0/OUT x3 0.05fF
C216 a_n787_n3768# x3 0.06fF
C217 a_425_n8036# x2 0.00fF
C218 CMOS_s3_0/CMOS_3in_OR_0/C CMOS_s3_0/CMOS_3in_OR_0/A 0.10fF
C219 a_n787_n3768# a_n2195_n2858# 0.00fF
C220 a_n2495_n3768# a_n787_n2858# 0.00fF
C221 CMOS_s3_0/CMOS_XOR_0/XOR CMOS_s2_0/CMOS_3in_OR_0/A 0.00fF
C222 a_n1990_n4808# CMOS_s2_0/CMOS_AND_1/A 0.00fF
C223 a_275_n2858# CMOS_s1_0/CMOS_XOR_0/XOR 0.01fF
C224 a_275_n6086# a_575_n6996# 0.02fF
C225 a_n732_n5418# CMOS_s1_0/CMOS_3in_OR_0/C 0.00fF
C226 x1 a_n1990_1648# 0.01fF
C227 a_425_n8036# x3 0.01fF
C228 VDD a_275_n2858# 0.59fF
C229 CMOS_s2_0/CMOS_4in_AND_0/OUT CMOS_s2_0/CMOS_XOR_0/XOR 0.00fF
C230 CMOS_s1_0/CMOS_AND_1/A CMOS_s1_0/CMOS_XOR_0/XOR 0.05fF
C231 CMOS_s0_0/CMOS_AND_1/B a_n2290_n540# 0.00fF
C232 a_n787_n3768# CMOS_s2_0/CMOS_XOR_0/XOR 0.00fF
C233 CMOS_s2_0/CMOS_3in_OR_0/B a_n732_n4808# 0.00fF
C234 VDD a_n1990_370# 0.00fF
C235 a_n2045_n6086# x2 0.00fF
C236 a_425_n540# a_425_n1580# 0.01fF
C237 VDD CMOS_s1_0/CMOS_AND_1/A 0.52fF
C238 CMOS_s2_0/CMOS_4in_AND_0/OUT a_n787_n6086# 0.01fF
C239 a_n1990_n8036# x2 0.00fF
C240 a_n432_n8036# a_n787_n10224# 0.00fF
C241 a_n432_n5418# CMOS_s2_0/CMOS_3in_OR_0/B 0.00fF
C242 a_n732_n8036# a_n2140_n8646# 0.00fF
C243 a_n2140_n540# a_n1990_1038# 0.00fF
C244 a_n2045_n6086# x3 0.00fF
C245 CMOS_s1_0/CMOS_3in_OR_0/C a_425_n4808# 0.01fF
C246 CMOS_s0_0/CMOS_AND_1/B CMOS_s1_0/CMOS_XOR_0/XOR 0.00fF
C247 CMOS_s3_0/CMOS_XOR_0/XOR CMOS_s3_0/CMOS_3in_OR_0/C 0.00fF
C248 a_n787_n540# x1 0.00fF
C249 a_n1990_n8036# x3 0.01fF
C250 a_n2495_n3768# x1 0.13fF
C251 a_n732_n1580# a_425_n1580# 0.00fF
C252 VDD CMOS_s0_0/CMOS_AND_1/B 0.85fF
C253 CMOS_s0_0/CMOS_AND_0/B CMOS_s0_0/CMOS_XOR_0/XOR 0.32fF
C254 a_n2140_n540# x2 0.21fF
C255 CMOS_s3_0/CMOS_AND_1/A a_n1990_n8646# 0.00fF
C256 CMOS_s0_0/CMOS_AND_1/A a_425_370# 0.01fF
C257 a_n432_n1580# a_n787_n540# 0.00fF
C258 a_n732_n1580# a_n787_n3768# 0.00fF
C259 a_n2140_n540# x3 0.07fF
C260 a_n2345_n6996# a_n787_n6996# 0.01fF
C261 a_n1990_n4808# x1 0.00fF
C262 VDD a_n2345_n6996# 1.65fF
C263 CMOS_s1_0/CMOS_XOR_0/XOR a_n432_n2190# 0.01fF
C264 CMOS_s2_0/CMOS_AND_1/A x2 0.01fF
C265 CMOS_s0_0/CMOS_AND_1/A x2 0.01fF
C266 a_n2290_n8036# x1 0.00fF
C267 a_425_n6996# CMOS_s2_0/CMOS_4in_AND_0/OUT 0.01fF
C268 VDD a_n432_n2190# 0.01fF
C269 a_n2140_n5418# a_n732_n5418# 0.00fF
C270 a_n2345_n9314# a_n2495_n10224# 0.01fF
C271 CMOS_s2_0/CMOS_AND_1/A x3 0.01fF
C272 CMOS_s0_0/CMOS_AND_1/A x3 0.00fF
C273 a_425_n5418# a_425_n4808# 0.01fF
C274 VDD a_275_n9314# 0.54fF
C275 a_1637_1038# a_425_1648# 0.01fF
C276 CMOS_s0_0/CMOS_AND_0/B a_425_1038# 0.00fF
C277 a_n2495_n3768# CMOS_s1_0/CMOS_3in_OR_0/C 0.05fF
C278 a_425_n6996# a_425_n8036# 0.00fF
C279 a_n787_n540# a_n2290_370# 0.00fF
C280 a_n787_n6996# a_n732_n8646# 0.00fF
C281 a_n1990_n1580# a_n2495_n3768# 0.00fF
C282 CMOS_s2_0/CMOS_AND_1/A CMOS_s2_0/CMOS_XOR_0/XOR 0.05fF
C283 VDD a_n732_n8646# 0.01fF
C284 VDD a_575_n10224# 0.06fF
C285 CMOS_s3_0/CMOS_3in_OR_0/B x1 0.06fF
C286 VDD a_n2495_n10224# 1.40fF
C287 CMOS_s2_0/CMOS_4in_AND_0/OUT CMOS_s2_0/CMOS_3in_OR_0/B 0.06fF
C288 a_n787_1038# x1 0.04fF
C289 a_n787_n6086# CMOS_s2_0/CMOS_AND_1/A 0.01fF
C290 a_n1990_1038# x1 0.00fF
C291 VDD a_n2290_n5418# 0.01fF
C292 CMOS_s0_0/CMOS_AND_1/A a_425_n540# 0.07fF
C293 x1 a_n2290_n1580# 0.00fF
C294 CMOS_s3_0/CMOS_3in_OR_0/B CMOS_s3_0/CMOS_3in_OR_0/A 0.04fF
C295 CMOS_s1_0/CMOS_AND_1/A a_n732_n2190# 0.00fF
C296 a_425_n8036# CMOS_s2_0/CMOS_3in_OR_0/B 0.00fF
C297 x1 x2 0.27fF
C298 CMOS_s3_0/CMOS_3in_OR_0/C a_425_n10224# 0.01fF
C299 CMOS_s2_0/CMOS_3in_OR_0/A a_575_n6996# 0.00fF
C300 a_425_n3768# a_425_n1580# 0.00fF
C301 a_n432_n4808# CMOS_s2_0/CMOS_XOR_0/XOR 0.03fF
C302 x1 x3 0.53fF
C303 VDD a_n2140_n8646# 1.10fF
C304 x1 a_n2195_n2858# 0.01fF
C305 a_n2290_n8646# x2 0.00fF
C306 a_425_n3768# a_n787_n3768# 0.00fF
C307 a_n732_n8036# a_n787_n6996# 0.00fF
C308 CMOS_s1_0/CMOS_3in_OR_0/B x3 0.00fF
C309 a_1637_1648# CMOS_s0_0/CMOS_AND_1/AND 0.01fF
C310 a_n432_n1580# x3 0.03fF
C311 a_575_n3768# a_425_n1580# 0.00fF
C312 CMOS_s3_0/CMOS_AND_1/A a_275_n9314# 0.00fF
C313 CMOS_s3_0/CMOS_3in_OR_0/A x3 0.00fF
C314 a_n2290_n8646# x3 0.00fF
C315 x1 CMOS_s2_0/CMOS_XOR_0/XOR 0.09fF
C316 a_575_n6996# a_425_n4808# 0.00fF
C317 a_n2345_n6086# x2 0.00fF
C318 VDD a_n732_n8036# 0.06fF
C319 CMOS_s3_0/CMOS_XOR_0/XOR CMOS_s3_0/CMOS_3in_OR_0/B 0.04fF
C320 a_n2195_n6086# CMOS_s2_0/CMOS_4in_AND_0/OUT 0.00fF
C321 a_n2140_n5418# a_n2495_n3768# 0.01fF
C322 a_575_n3768# a_n787_n3768# 0.00fF
C323 a_n787_n6086# x1 0.00fF
C324 CMOS_s1_0/CMOS_3in_OR_0/B CMOS_s2_0/CMOS_XOR_0/XOR 0.00fF
C325 a_275_n2858# a_425_n1580# 0.01fF
C326 a_n2345_n6086# x3 0.00fF
C327 CMOS_s3_0/CMOS_AND_1/A a_n732_n8646# 0.00fF
C328 CMOS_s3_0/CMOS_AND_1/A a_n2495_n10224# 0.00fF
C329 CMOS_s3_0/CMOS_XOR_0/XOR x2 0.09fF
C330 CMOS_s1_0/CMOS_3in_OR_0/C x2 0.00fF
C331 a_n2290_370# x2 0.01fF
C332 CMOS_s0_0/CMOS_AND_1/B a_n787_1648# 0.00fF
C333 CMOS_s0_0/CMOS_XOR_0/XOR a_425_1648# 0.06fF
C334 a_275_n2858# a_n787_n3768# 0.01fF
C335 a_n2140_n5418# a_n1990_n4808# 0.03fF
C336 a_n1990_n1580# x2 0.03fF
C337 CMOS_s3_0/CMOS_XOR_0/XOR x3 0.35fF
C338 CMOS_s1_0/CMOS_AND_1/A a_n787_n3768# 0.05fF
C339 VDD CMOS_s0_0/CMOS_AND_1/AND 0.44fF
C340 CMOS_s1_0/CMOS_3in_OR_0/C x3 0.06fF
C341 x1 a_n787_n10224# 0.03fF
C342 a_n2290_370# x3 0.00fF
C343 CMOS_s1_0/CMOS_3in_OR_0/C a_n2195_n2858# 0.00fF
C344 a_n787_1038# CMOS_s0_0/CMOS_AND_0/B 0.07fF
C345 CMOS_s2_0/CMOS_3in_OR_0/B CMOS_s2_0/CMOS_AND_1/A 0.01fF
C346 a_n787_n9314# CMOS_s3_0/CMOS_3in_OR_0/C 0.01fF
C347 CMOS_s1_0/CMOS_3in_OR_0/B a_n732_n1580# 0.00fF
C348 a_n1990_n1580# x3 0.01fF
C349 CMOS_s3_0/CMOS_AND_1/A a_n2140_n8646# 0.08fF
C350 a_n787_n10224# CMOS_s3_0/CMOS_3in_OR_0/A 0.07fF
C351 CMOS_s1_0/CMOS_3in_OR_0/C CMOS_s2_0/CMOS_XOR_0/XOR 0.03fF
C352 CMOS_s1_0/CMOS_XOR_0/XOR CMOS_s1_0/CMOS_3in_OR_0/A 0.02fF
C353 a_275_n6086# CMOS_s2_0/CMOS_3in_OR_0/A 0.10fF
C354 VDD CMOS_s1_0/CMOS_3in_OR_0/A 0.55fF
C355 CMOS_s0_0/CMOS_AND_0/B x3 0.00fF
C356 CMOS_s3_0/CMOS_AND_1/A a_n732_n8036# 0.01fF
C357 a_1637_1648# VDD 0.06fF
C358 a_425_1038# a_425_1648# 0.01fF
C359 a_n432_n4808# CMOS_s2_0/CMOS_3in_OR_0/B 0.00fF
C360 a_n432_n2190# a_425_n1580# 0.00fF
C361 a_n2345_n6996# CMOS_s2_0/CMOS_4in_AND_0/OUT 0.05fF
C362 a_n1990_n540# a_n2140_n2190# 0.00fF
C363 CMOS_s3_0/CMOS_XOR_0/XOR a_n787_n10224# 0.01fF
C364 a_n2140_n540# a_n1990_370# 0.01fF
C365 VDD a_n2345_n9314# 0.01fF
C366 VDD a_n2290_n540# 0.03fF
C367 a_n432_n2190# a_n787_n3768# 0.00fF
C368 a_275_n6086# a_425_n4808# 0.01fF
C369 CMOS_s3_0/CMOS_3in_OR_0/B a_425_n10224# 0.00fF
C370 x1 CMOS_s2_0/CMOS_3in_OR_0/B 0.00fF
C371 CMOS_s3_0/CMOS_3in_OR_0/B a_425_n8646# 0.01fF
C372 a_n2140_n5418# x2 0.34fF
C373 VDD a_n787_n6996# 0.78fF
C374 a_425_n5418# CMOS_s2_0/CMOS_XOR_0/XOR 0.01fF
C375 a_n2140_n5418# x3 0.06fF
C376 VDD CMOS_s1_0/CMOS_XOR_0/XOR 1.07fF
C377 a_1637_1038# CMOS_s0_0/CMOS_XOR_0/XOR 0.00fF
C378 VDD a_n2290_1648# 0.04fF
C379 a_n2140_n5418# a_n2195_n2858# 0.00fF
C380 a_n2140_n540# CMOS_s0_0/CMOS_AND_1/B 0.12fF
C381 a_425_n8036# a_275_n9314# 0.01fF
C382 a_n1990_n2190# a_n2140_n2190# 0.01fF
C383 a_425_n8646# x2 0.00fF
C384 CMOS_s2_0/CMOS_4in_AND_0/OUT a_n732_n8646# 0.00fF
C385 a_n2345_n6996# a_n2045_n6086# 0.01fF
C386 a_n2345_n6996# a_n1990_n8036# 0.00fF
C387 a_n2140_n5418# CMOS_s2_0/CMOS_XOR_0/XOR 0.04fF
C388 a_n2290_n2190# a_n2140_n2190# 0.01fF
C389 VDD a_n2345_n2858# 0.01fF
C390 a_275_n2858# a_n787_n2858# 0.00fF
C391 a_425_n8036# a_n732_n8646# 0.00fF
C392 a_n1990_n8646# x1 0.00fF
C393 a_425_n8036# a_575_n10224# 0.00fF
C394 CMOS_s0_0/CMOS_AND_0/AND CMOS_s0_0/CMOS_AND_1/AND 0.09fF
C395 CMOS_s1_0/CMOS_AND_1/A a_n787_n2858# 0.01fF
C396 CMOS_s1_0/CMOS_3in_OR_0/B a_425_n3768# 0.00fF
C397 CMOS_s0_0/CMOS_AND_1/A CMOS_s0_0/CMOS_AND_1/B 0.18fF
C398 a_n2195_n6086# x1 0.00fF
C399 CMOS_s3_0/CMOS_XOR_0/XOR CMOS_s2_0/CMOS_3in_OR_0/B 0.00fF
C400 CMOS_s2_0/CMOS_4in_AND_0/OUT a_n2140_n8646# 0.01fF
C401 a_1637_1038# a_425_1038# 0.00fF
C402 CMOS_s1_0/CMOS_3in_OR_0/B a_575_n3768# 0.00fF
C403 a_n1990_n8036# a_n2495_n10224# 0.00fF
C404 a_425_370# a_425_1648# 0.00fF
C405 a_n2345_n6996# CMOS_s2_0/CMOS_AND_1/A 0.00fF
C406 a_n1990_370# x1 0.00fF
C407 a_n732_n8036# CMOS_s2_0/CMOS_4in_AND_0/OUT 0.01fF
C408 a_1637_1648# CMOS_s0_0/CMOS_AND_0/AND 0.01fF
C409 CMOS_s1_0/CMOS_AND_1/A x1 0.08fF
C410 CMOS_s1_0/CMOS_3in_OR_0/B a_275_n2858# 0.12fF
C411 a_n787_1038# a_425_1648# 0.01fF
C412 a_n787_n6996# a_n732_n4808# 0.00fF
C413 VDD CMOS_s3_0/CMOS_AND_1/A 0.51fF
C414 a_425_n10224# a_n787_n10224# 0.00fF
C415 a_n787_n9314# x2 0.00fF
C416 a_n1990_n540# CMOS_s0_0/CMOS_XOR_0/XOR 0.00fF
C417 a_425_n3768# CMOS_s1_0/CMOS_3in_OR_0/C 0.01fF
C418 CMOS_s3_0/CMOS_XOR_0/XOR a_n1990_n8646# 0.00fF
C419 a_425_n8036# a_n732_n8036# 0.00fF
C420 a_n2140_n2190# a_n2495_n3768# 0.01fF
C421 CMOS_s1_0/CMOS_3in_OR_0/B CMOS_s1_0/CMOS_AND_1/A 0.01fF
C422 CMOS_s3_0/CMOS_3in_OR_0/B a_n432_n8646# 0.00fF
C423 a_n432_n1580# CMOS_s1_0/CMOS_AND_1/A 0.00fF
C424 a_n2045_n6086# a_n2140_n8646# 0.00fF
C425 VDD a_n732_n4808# 0.06fF
C426 a_n787_n6996# a_n432_n5418# 0.00fF
C427 a_n1990_n8036# a_n2140_n8646# 0.03fF
C428 CMOS_s0_0/CMOS_AND_1/B x1 0.01fF
C429 VDD a_n432_n5418# 0.01fF
C430 a_575_n3768# CMOS_s1_0/CMOS_3in_OR_0/C 0.01fF
C431 a_425_n5418# CMOS_s2_0/CMOS_3in_OR_0/B 0.01fF
C432 a_n2195_n9314# CMOS_s3_0/CMOS_3in_OR_0/C 0.00fF
C433 a_n432_n1580# CMOS_s0_0/CMOS_AND_1/B 0.00fF
C434 a_n432_n8646# x2 0.00fF
C435 a_n732_n2190# CMOS_s1_0/CMOS_XOR_0/XOR 0.01fF
C436 VDD a_n2290_n4808# 0.05fF
C437 VDD a_n732_n2190# 0.01fF
C438 VDD CMOS_s0_0/CMOS_AND_0/AND 0.58fF
C439 a_n2290_n5418# CMOS_s2_0/CMOS_AND_1/A 0.00fF
C440 a_n732_n5418# a_425_n4808# 0.00fF
C441 a_n432_n8646# x3 0.01fF
C442 a_275_n6086# CMOS_s3_0/CMOS_3in_OR_0/B 0.01fF
C443 a_n1990_n5418# x2 0.01fF
C444 a_275_n2858# CMOS_s1_0/CMOS_3in_OR_0/C 0.05fF
C445 a_n787_370# CMOS_s0_0/CMOS_XOR_0/XOR 0.00fF
C446 a_n2345_n6996# x1 0.10fF
C447 a_425_n540# a_425_n2190# 0.00fF
C448 CMOS_s1_0/CMOS_AND_1/A CMOS_s1_0/CMOS_3in_OR_0/C 0.02fF
C449 a_n432_n2190# x1 0.00fF
C450 a_n1990_n5418# x3 0.00fF
C451 a_n787_n3768# CMOS_s1_0/CMOS_3in_OR_0/A 0.07fF
C452 a_n1990_n1580# CMOS_s1_0/CMOS_AND_1/A 0.00fF
C453 a_275_n9314# x1 0.04fF
C454 a_425_n540# a_425_1648# 0.01fF
C455 CMOS_s1_0/CMOS_3in_OR_0/B a_n432_n2190# 0.00fF
C456 a_n2345_n6996# a_n2290_n8646# 0.00fF
C457 a_n787_n6996# a_n432_n8036# 0.00fF
C458 a_n787_n9314# a_n787_n10224# 0.01fF
C459 a_425_1038# CMOS_s0_0/CMOS_XOR_0/XOR 0.01fF
C460 a_n2290_370# CMOS_s0_0/CMOS_AND_1/B 0.00fF
C461 a_n1990_n5418# CMOS_s2_0/CMOS_XOR_0/XOR 0.00fF
C462 a_n1990_1648# CMOS_s0_0/CMOS_XOR_0/XOR 0.03fF
C463 a_n2345_n6086# a_n2345_n6996# 0.00fF
C464 VDD a_n787_1648# 0.05fF
C465 a_275_n9314# CMOS_s3_0/CMOS_3in_OR_0/A 0.10fF
C466 a_n787_n540# a_n1990_n540# 0.00fF
C467 x1 a_n732_n8646# 0.01fF
C468 VDD a_n432_n8036# 0.06fF
C469 x1 a_n2495_n10224# 0.04fF
C470 VDD a_n2290_1038# 0.01fF
C471 a_n2140_n2190# a_n2290_n1580# 0.02fF
C472 CMOS_s1_0/CMOS_XOR_0/XOR a_425_n1580# 0.09fF
C473 a_275_n6086# CMOS_s2_0/CMOS_XOR_0/XOR 0.01fF
C474 a_n2290_n5418# x1 0.00fF
C475 CMOS_s2_0/CMOS_4in_AND_0/OUT a_n787_n6996# 0.10fF
C476 VDD a_425_n1580# 0.82fF
C477 a_n2140_n2190# x2 0.34fF
C478 a_n432_n8646# a_n787_n10224# 0.00fF
C479 a_n2195_n6086# a_n2140_n5418# 0.00fF
C480 a_575_n6996# CMOS_s2_0/CMOS_3in_OR_0/B 0.00fF
C481 a_575_n10224# CMOS_s3_0/CMOS_3in_OR_0/A 0.00fF
C482 a_n2495_n10224# CMOS_s3_0/CMOS_3in_OR_0/A 0.00fF
C483 CMOS_s0_0/CMOS_AND_0/B CMOS_s0_0/CMOS_AND_1/B 0.01fF
C484 a_n2290_n8646# a_n2495_n10224# 0.00fF
C485 CMOS_s1_0/CMOS_XOR_0/XOR a_n787_n3768# 0.01fF
C486 a_275_n6086# a_n787_n6086# 0.00fF
C487 VDD CMOS_s2_0/CMOS_4in_AND_0/OUT 2.47fF
C488 a_n787_n540# CMOS_s0_0/CMOS_XOR_0/XOR 0.01fF
C489 VDD a_n787_n3768# 0.78fF
C490 a_n2140_n2190# x3 0.17fF
C491 a_n2140_n2190# a_n2195_n2858# 0.00fF
C492 a_n1990_n2190# a_n2495_n3768# 0.00fF
C493 CMOS_s3_0/CMOS_XOR_0/XOR a_275_n9314# 0.01fF
C494 CMOS_s0_0/CMOS_AND_1/AND CMOS_s0_0/CMOS_AND_1/A 0.01fF
C495 x1 a_n2140_n8646# 0.06fF
C496 a_425_n8036# VDD 0.82fF
C497 a_n787_n540# a_n787_370# 0.01fF
C498 a_n2290_n2190# a_n2495_n3768# 0.00fF
C499 a_n787_n6996# a_n2045_n6086# 0.00fF
C500 CMOS_s3_0/CMOS_XOR_0/XOR a_n732_n8646# 0.01fF
C501 a_n732_n8036# x1 0.00fF
C502 a_n2290_n8646# a_n2140_n8646# 0.01fF
C503 a_n2140_n540# a_n2290_n540# 0.02fF
C504 VDD a_n2045_n6086# 0.01fF
C505 VDD a_n1990_n8036# 0.05fF
C506 CMOS_s3_0/CMOS_AND_1/A a_n432_n8036# 0.00fF
C507 a_425_n6996# a_275_n6086# 0.02fF
C508 a_n732_n1580# a_n2140_n2190# 0.00fF
C509 CMOS_s1_0/CMOS_3in_OR_0/A a_n787_n2858# 0.00fF
C510 VDD a_n2140_n540# 1.07fF
C511 a_425_370# CMOS_s0_0/CMOS_XOR_0/XOR 0.00fF
C512 a_n2195_n9314# x2 0.00fF
C513 CMOS_s3_0/CMOS_XOR_0/XOR a_n2140_n8646# 0.04fF
C514 a_n2345_n6996# a_n2140_n5418# 0.01fF
C515 a_n1990_n540# x2 0.01fF
C516 CMOS_s3_0/CMOS_AND_1/A CMOS_s2_0/CMOS_4in_AND_0/OUT 0.01fF
C517 a_n787_1038# CMOS_s0_0/CMOS_XOR_0/XOR 0.07fF
C518 CMOS_s1_0/CMOS_3in_OR_0/B CMOS_s0_0/CMOS_AND_1/AND 0.00fF
C519 a_n787_n6996# CMOS_s2_0/CMOS_AND_1/A 0.05fF
C520 a_n1990_1038# CMOS_s0_0/CMOS_XOR_0/XOR 0.01fF
C521 a_n2195_n9314# x3 0.00fF
C522 a_n1990_n540# x3 0.00fF
C523 a_n787_n3768# a_n732_n4808# 0.00fF
C524 CMOS_s3_0/CMOS_XOR_0/XOR a_n732_n8036# 0.02fF
C525 CMOS_s0_0/CMOS_AND_1/A CMOS_s1_0/CMOS_XOR_0/XOR 0.00fF
C526 a_275_n6086# CMOS_s2_0/CMOS_3in_OR_0/B 0.12fF
C527 VDD CMOS_s0_0/CMOS_AND_1/A 0.54fF
C528 VDD CMOS_s2_0/CMOS_AND_1/A 0.52fF
C529 x2 CMOS_s0_0/CMOS_XOR_0/XOR 0.05fF
C530 a_n787_1038# a_n787_370# 0.00fF
C531 a_n732_n2190# a_425_n1580# 0.00fF
C532 CMOS_s3_0/CMOS_3in_OR_0/C CMOS_s3_0/CMOS_3in_OR_0/B 0.06fF
C533 CMOS_s2_0/CMOS_3in_OR_0/A x3 0.00fF
C534 a_275_n2858# a_425_n2190# 0.00fF
C535 a_n1990_n2190# x2 0.01fF
C536 a_n1990_n4808# a_n2495_n3768# 0.00fF
C537 a_275_n9314# a_425_n10224# 0.02fF
C538 x3 CMOS_s0_0/CMOS_XOR_0/XOR 0.32fF
C539 a_n732_n2190# a_n787_n3768# 0.00fF
C540 CMOS_s1_0/CMOS_3in_OR_0/B CMOS_s1_0/CMOS_3in_OR_0/A 0.04fF
C541 a_275_n9314# a_425_n8646# 0.00fF
C542 VDD a_n787_n2858# 0.00fF
C543 a_n787_370# x2 0.01fF
C544 CMOS_s3_0/CMOS_AND_1/A a_n1990_n8036# 0.00fF
C545 a_n2290_n2190# x2 0.01fF
C546 CMOS_s2_0/CMOS_3in_OR_0/A CMOS_s2_0/CMOS_XOR_0/XOR 0.02fF
C547 a_n787_n6996# a_n432_n4808# 0.00fF
C548 a_n1990_n2190# x3 0.00fF
C549 CMOS_s3_0/CMOS_3in_OR_0/C x2 0.03fF
C550 a_n732_n5418# CMOS_s2_0/CMOS_XOR_0/XOR 0.01fF
C551 a_n2140_n5418# a_n2290_n5418# 0.01fF
C552 a_n2345_n9314# x1 0.01fF
C553 a_n2290_n540# x1 0.00fF
C554 CMOS_s2_0/CMOS_3in_OR_0/A a_n787_n6086# 0.00fF
C555 a_n787_1038# a_425_1038# 0.00fF
C556 a_n787_370# x3 0.00fF
C557 VDD a_n432_n4808# 0.06fF
C558 a_n2290_n2190# x3 0.00fF
C559 a_n787_1038# a_n1990_1648# 0.00fF
C560 CMOS_s3_0/CMOS_3in_OR_0/C x3 0.00fF
C561 a_n787_n6996# x1 0.01fF
C562 a_n2195_n9314# a_n787_n10224# 0.00fF
C563 a_425_n540# CMOS_s0_0/CMOS_XOR_0/XOR 0.00fF
C564 CMOS_s1_0/CMOS_XOR_0/XOR x1 0.09fF
C565 x2 a_n1990_1648# 0.00fF
C566 CMOS_s2_0/CMOS_XOR_0/XOR a_425_n4808# 0.09fF
C567 a_n2290_1648# x1 0.01fF
C568 a_n787_n540# a_425_370# 0.00fF
C569 VDD x1 2.45fF
C570 CMOS_s2_0/CMOS_4in_AND_0/OUT a_n432_n8036# 0.01fF
C571 CMOS_s1_0/CMOS_3in_OR_0/B CMOS_s1_0/CMOS_XOR_0/XOR 0.04fF
C572 CMOS_s1_0/CMOS_3in_OR_0/A CMOS_s1_0/CMOS_3in_OR_0/C 0.10fF
C573 a_n432_n1580# CMOS_s1_0/CMOS_XOR_0/XOR 0.03fF
C574 CMOS_s0_0/CMOS_AND_1/AND CMOS_s0_0/CMOS_AND_0/B 0.00fF
C575 x3 a_n1990_1648# 0.03fF
C576 a_n787_n540# a_n787_1038# 0.01fF
C577 CMOS_s1_0/CMOS_3in_OR_0/B VDD 0.51fF
C578 a_425_n540# a_n787_370# 0.00fF
C579 VDD a_n432_n1580# 0.06fF
C580 a_n2345_n2858# x1 0.01fF
C581 VDD CMOS_s3_0/CMOS_3in_OR_0/A 0.52fF
C582 VDD a_n2290_n8646# 0.01fF
C583 a_425_n8036# a_n432_n8036# 0.00fF
C584 CMOS_s2_0/CMOS_AND_1/A a_n732_n4808# 0.01fF
C585 a_n787_n540# x2 0.05fF
C586 a_n2495_n3768# x2 0.05fF
C587 a_n787_n9314# a_275_n9314# 0.00fF
C588 a_425_n6996# CMOS_s2_0/CMOS_3in_OR_0/A 0.01fF
C589 a_n432_n5418# CMOS_s2_0/CMOS_AND_1/A 0.00fF
C590 a_n2345_n6086# VDD 0.01fF
C591 CMOS_s3_0/CMOS_3in_OR_0/C a_n787_n10224# 0.10fF
C592 a_n2495_n3768# x3 0.11fF
C593 a_425_n540# a_425_1038# 0.00fF
C594 a_n787_n540# x3 0.01fF
C595 CMOS_s3_0/CMOS_XOR_0/XOR a_n787_n6996# 0.00fF
C596 a_n2495_n3768# a_n2195_n2858# 0.01fF
C597 a_425_n8036# CMOS_s2_0/CMOS_4in_AND_0/OUT 0.01fF
C598 a_n2290_n4808# CMOS_s2_0/CMOS_AND_1/A 0.00fF
C599 a_n1990_n4808# x2 0.03fF
C600 CMOS_s1_0/CMOS_XOR_0/XOR CMOS_s1_0/CMOS_3in_OR_0/C 0.00fF
C601 a_n2345_n6996# a_n1990_n5418# 0.00fF
C602 a_n787_n9314# a_n2495_n10224# 0.00fF
C603 CMOS_s3_0/CMOS_XOR_0/XOR VDD 1.07fF
C604 CMOS_s1_0/CMOS_AND_1/A a_n2140_n2190# 0.08fF
C605 VDD CMOS_s1_0/CMOS_3in_OR_0/C 2.54fF
C606 a_n1990_n1580# CMOS_s1_0/CMOS_XOR_0/XOR 0.00fF
C607 VDD a_n2290_370# 0.00fF
C608 a_425_n6996# a_425_n4808# 0.00fF
C609 a_n1990_n4808# x3 0.00fF
C610 VDD a_n1990_n1580# 0.05fF
C611 CMOS_s2_0/CMOS_3in_OR_0/A CMOS_s2_0/CMOS_3in_OR_0/B 0.04fF
C612 CMOS_s2_0/CMOS_4in_AND_0/OUT a_n2045_n6086# 0.00fF
C613 a_n2290_n8036# x2 0.00fF
C614 a_n732_n5418# CMOS_s2_0/CMOS_3in_OR_0/B 0.00fF
C615 CMOS_s3_0/CMOS_AND_1/A x1 0.03fF
C616 a_n2345_n2858# CMOS_s1_0/CMOS_3in_OR_0/C 0.00fF
C617 a_n787_n540# a_425_n540# 0.01fF
C618 a_n2290_n8036# x3 0.01fF
C619 a_n1990_n4808# CMOS_s2_0/CMOS_XOR_0/XOR 0.00fF
C620 CMOS_s3_0/CMOS_AND_1/A CMOS_s3_0/CMOS_3in_OR_0/A 0.00fF
C621 VDD CMOS_s0_0/CMOS_AND_0/B 0.58fF
C622 CMOS_s3_0/CMOS_AND_1/A a_n2290_n8646# 0.00fF
C623 a_n787_1038# a_n1990_1038# 0.00fF
C624 a_n432_n5418# x1 0.00fF
C625 a_n732_n1580# a_n787_n540# 0.00fF
C626 CMOS_s2_0/CMOS_3in_OR_0/B a_425_n4808# 0.08fF
C627 CMOS_s3_0/CMOS_3in_OR_0/B x2 0.00fF
C628 a_n2290_n4808# x1 0.00fF
C629 a_n787_1038# x2 0.00fF
C630 a_n732_n2190# x1 0.00fF
C631 a_n1990_1038# x2 0.00fF
C632 CMOS_s0_0/CMOS_AND_1/A a_425_n1580# 0.00fF
C633 CMOS_s3_0/CMOS_3in_OR_0/B x3 0.00fF
C634 a_n2290_n1580# x2 0.02fF
C635 VDD a_425_n5418# 0.01fF
C636 CMOS_s1_0/CMOS_3in_OR_0/B a_n732_n2190# 0.00fF
C637 a_n787_1038# x3 0.01fF
C638 a_n1990_1038# x3 0.01fF
C639 CMOS_s2_0/CMOS_4in_AND_0/OUT CMOS_s2_0/CMOS_AND_1/A 0.02fF
C640 CMOS_s3_0/CMOS_XOR_0/XOR CMOS_s3_0/CMOS_AND_1/A 0.05fF
C641 a_n2290_n1580# x3 0.01fF
C642 a_425_n3768# a_425_n4808# 0.00fF
C643 x2 x3 0.62fF
C644 VDD a_n2140_n5418# 1.09fF
C645 a_n2195_n2858# x2 0.00fF
C646 CMOS_s1_0/CMOS_3in_OR_0/C a_n732_n4808# 0.01fF
C647 a_425_n540# a_425_370# 0.01fF
C648 a_n787_n3768# a_n787_n2858# 0.01fF
C649 a_n2195_n2858# x3 0.00fF
C650 a_n432_n5418# CMOS_s1_0/CMOS_3in_OR_0/C 0.00fF
C651 x1 a_n787_1648# 0.01fF
C652 a_575_n3768# a_425_n4808# 0.00fF
C653 a_n432_n8036# x1 0.00fF
C654 x2 CMOS_s2_0/CMOS_XOR_0/XOR 0.00fF
C655 VDD a_425_n10224# 0.06fF
C656 CMOS_s0_0/CMOS_AND_1/AND a_425_1648# 0.00fF
C657 VDD a_425_n8646# 0.01fF
C658 a_n1990_370# CMOS_s0_0/CMOS_XOR_0/XOR 0.00fF
C659 CMOS_s0_0/CMOS_AND_1/B a_n1990_n540# 0.00fF
C660 a_n787_n3768# a_n432_n4808# 0.00fF
C661 a_n2290_1038# x1 0.00fF
C662 CMOS_s2_0/CMOS_XOR_0/XOR x3 0.00fF
C663 x1 a_425_n1580# 0.00fF
C664 CMOS_s3_0/CMOS_3in_OR_0/B a_n787_n10224# 0.00fF
C665 a_425_n540# x2 0.00fF
C666 CMOS_s1_0/CMOS_AND_1/A a_n1990_n2190# 0.00fF
C667 a_275_n2858# a_425_n4808# 0.00fF
C668 a_n787_n6086# x3 0.00fF
C669 CMOS_s1_0/CMOS_3in_OR_0/B a_425_n1580# 0.08fF
C670 CMOS_s2_0/CMOS_4in_AND_0/OUT x1 0.04fF
C671 a_n787_n6996# a_575_n6996# 0.00fF
C672 a_n432_n1580# a_425_n1580# 0.00fF
C673 a_n787_n3768# x1 0.01fF
C674 CMOS_s0_0/CMOS_AND_1/B CMOS_s0_0/CMOS_XOR_0/XOR 0.01fF
C675 a_n2290_n2190# CMOS_s1_0/CMOS_AND_1/A 0.00fF
C676 CMOS_s0_0/CMOS_AND_1/A a_n2140_n540# 0.00fF
C677 x2 a_n787_n10224# 0.00fF
C678 VDD a_575_n6996# 0.06fF
C679 a_1637_1648# a_425_1648# 0.00fF
C680 CMOS_s1_0/CMOS_3in_OR_0/B a_n787_n3768# 0.00fF
C681 a_n432_n1580# a_n787_n3768# 0.00fF
C682 a_425_n8036# x1 0.05fF
C683 CMOS_s0_0/CMOS_AND_0/AND CMOS_s0_0/CMOS_AND_0/B 0.01fF
C684 CMOS_s0_0/CMOS_AND_1/B a_n787_370# 0.01fF
C685 a_n2345_n6996# CMOS_s2_0/CMOS_3in_OR_0/A 0.00fF
C686 a_n732_n1580# x3 0.01fF
C687 a_n787_n10224# x3 0.02fF
C688 CMOS_s3_0/CMOS_XOR_0/XOR a_n432_n8036# 0.03fF
C689 a_n2345_n6086# CMOS_s2_0/CMOS_4in_AND_0/OUT 0.00fF
C690 a_n2140_n5418# a_n732_n4808# 0.00fF
C691 CMOS_s1_0/CMOS_XOR_0/XOR a_425_n2190# 0.01fF
C692 a_n2045_n6086# x1 0.00fF
C693 a_n1990_n8036# x1 0.00fF
C694 VDD a_425_n2190# 0.01fF
C695 a_n787_n9314# VDD 0.00fF
C696 CMOS_s1_0/CMOS_3in_OR_0/C a_425_n1580# 0.00fF
C697 a_n2195_n9314# a_n2495_n10224# 0.01fF
C698 CMOS_s3_0/CMOS_XOR_0/XOR CMOS_s2_0/CMOS_4in_AND_0/OUT 0.03fF
C699 VDD a_425_1648# 0.81fF
C700 CMOS_s0_0/CMOS_AND_0/B a_n787_1648# 0.00fF
C701 a_n2140_n5418# a_n2290_n4808# 0.02fF
C702 a_n787_n3768# CMOS_s1_0/CMOS_3in_OR_0/C 0.10fF
C703 a_n787_n540# a_n1990_370# 0.00fF
C704 a_n2140_n540# x1 0.01fF
C705 CMOS_s0_0/CMOS_AND_1/AND a_1637_1038# 0.08fF
C706 CMOS_s1_0/CMOS_AND_1/A a_n2495_n3768# 0.00fF
C707 a_n432_n4808# CMOS_s2_0/CMOS_AND_1/A 0.00fF
C708 CMOS_s3_0/CMOS_XOR_0/XOR a_425_n8036# 0.09fF
C709 a_425_n6996# CMOS_s2_0/CMOS_XOR_0/XOR 0.00fF
C710 VDD a_n432_n8646# 0.01fF
C711 CMOS_s3_0/CMOS_3in_OR_0/C a_275_n9314# 0.05fF
C712 a_n2195_n9314# a_n2140_n8646# 0.00fF
C713 a_n787_n540# CMOS_s0_0/CMOS_AND_1/B 0.09fF
C714 VDD a_n1990_n5418# 0.01fF
C715 x1 CMOS_s2_0/CMOS_AND_1/A 0.08fF
C716 a_275_n6086# a_n787_n6996# 0.01fF
C717 CMOS_s3_0/CMOS_3in_OR_0/C a_575_n10224# 0.01fF
C718 CMOS_s3_0/CMOS_XOR_0/XOR a_n1990_n8036# 0.00fF
C719 a_1637_1648# a_1637_1038# 0.01fF
C720 CMOS_s3_0/CMOS_3in_OR_0/C a_n2495_n10224# 0.05fF
C721 CMOS_s2_0/CMOS_3in_OR_0/B CMOS_s2_0/CMOS_XOR_0/XOR 0.04fF
C722 VDD a_275_n6086# 0.59fF
C723 x1 a_n787_n2858# 0.00fF
C724 a_n1990_n8646# x2 0.00fF
C725 a_n787_n9314# CMOS_s3_0/CMOS_AND_1/A 0.01fF
C726 a_n2140_n540# a_n2290_370# 0.01fF
C727 a_n1990_n1580# a_n2140_n540# 0.00fF
C728 a_n1990_n8646# x3 0.00fF
C729 a_n2195_n6086# x2 0.00fF
C730 a_n2140_n5418# CMOS_s2_0/CMOS_4in_AND_0/OUT 0.01fF
C731 CMOS_s3_0/CMOS_3in_OR_0/C a_n2140_n8646# 0.01fF
C732 a_n2140_n2190# CMOS_s1_0/CMOS_XOR_0/XOR 0.04fF
C733 a_n2345_n6996# a_n1990_n4808# 0.00fF
C734 VDD a_n2140_n2190# 1.09fF
C735 a_n2195_n6086# x3 0.00fF
C736 CMOS_s3_0/CMOS_AND_1/A a_n432_n8646# 0.00fF
C737 VDD a_1637_1038# 0.50fF
C738 CMOS_s1_0/CMOS_3in_OR_0/C CMOS_s2_0/CMOS_AND_1/A 0.01fF
C739 CMOS_s1_0/CMOS_AND_1/A a_n2290_n1580# 0.00fF
C740 a_n1990_370# x2 0.01fF
C741 CMOS_s2_0/CMOS_4in_AND_0/OUT a_425_n8646# 0.00fF
C742 a_n2345_n6996# a_n2290_n8036# 0.00fF
C743 CMOS_s1_0/CMOS_AND_1/A x2 0.01fF
C744 CMOS_s1_0/CMOS_3in_OR_0/B x1 0.00fF
C745 a_n787_1038# CMOS_s0_0/CMOS_AND_1/B 0.01fF
C746 a_275_n2858# x3 0.00fF
C747 CMOS_s0_0/CMOS_AND_0/AND a_425_1648# 0.07fF
C748 CMOS_s0_0/CMOS_AND_1/AND CMOS_s0_0/CMOS_XOR_0/XOR 0.01fF
C749 x1 CMOS_s3_0/CMOS_3in_OR_0/A 0.03fF
C750 a_n2290_n8646# x1 0.01fF
C751 a_n1990_370# x3 0.00fF
C752 a_n2290_n5418# a_n2495_n3768# 0.00fF
C753 CMOS_s1_0/CMOS_3in_OR_0/C a_n787_n2858# 0.01fF
C754 a_425_n8036# a_425_n10224# 0.00fF
C755 a_425_n8036# a_425_n8646# 0.01fF
C756 a_425_n6996# CMOS_s2_0/CMOS_3in_OR_0/B 0.00fF
C757 a_n2140_n5418# a_n2045_n6086# 0.00fF
C758 CMOS_s1_0/CMOS_AND_1/A x3 0.09fF
C759 CMOS_s1_0/CMOS_3in_OR_0/B a_n432_n1580# 0.00fF
C760 CMOS_s0_0/CMOS_AND_1/B x2 0.17fF
C761 CMOS_s0_0/CMOS_AND_1/A CMOS_s0_0/CMOS_AND_0/B 0.01fF
C762 a_n2345_n6086# x1 0.00fF
C763 a_275_n2858# CMOS_s2_0/CMOS_XOR_0/XOR 0.00fF
C764 a_n432_n4808# CMOS_s1_0/CMOS_3in_OR_0/C 0.01fF
C765 CMOS_s2_0/CMOS_4in_AND_0/OUT a_575_n6996# 0.01fF
C766 CMOS_s0_0/CMOS_AND_1/B x3 0.02fF
C767 CMOS_s3_0/CMOS_XOR_0/XOR x1 0.23fF
C768 a_n787_1648# a_425_1648# 0.00fF
C769 x1 CMOS_s1_0/CMOS_3in_OR_0/C 0.09fF
C770 a_425_n8036# a_575_n6996# 0.00fF
C771 a_275_n9314# CMOS_s3_0/CMOS_3in_OR_0/B 0.12fF
C772 a_n2290_370# x1 0.00fF
C773 a_425_n2190# a_425_n1580# 0.01fF
C774 a_n2345_n6996# x2 0.03fF
C775 a_575_n10224# GND 0.02fF
C776 a_425_n10224# GND 0.02fF
C777 a_n787_n9314# GND 0.03fF
C778 a_n2195_n9314# GND 0.03fF
C779 a_n2345_n9314# GND 0.03fF
C780 a_275_n9314# GND 0.94fF
C781 CMOS_s3_0/CMOS_3in_OR_0/C GND 1.11fF $ **FLOATING
C782 CMOS_s3_0/CMOS_3in_OR_0/A GND 0.58fF
C783 a_n787_n10224# GND 0.50fF
C784 a_n2495_n10224# GND 0.71fF
C785 a_425_n8646# GND 0.03fF
C786 a_n432_n8646# GND 0.03fF
C787 a_n732_n8646# GND 0.02fF
C788 a_n1990_n8646# GND 0.02fF
C789 a_n2290_n8646# GND 0.02fF
C790 CMOS_s3_0/CMOS_3in_OR_0/B GND 1.98fF
C791 a_n432_n8036# GND 0.01fF
C792 a_n732_n8036# GND 0.01fF
C793 CMOS_s3_0/CMOS_AND_1/A GND 1.10fF
C794 a_n1990_n8036# GND 0.01fF
C795 a_n2290_n8036# GND 0.01fF
C796 a_425_n8036# GND 0.52fF
C797 CMOS_s3_0/CMOS_XOR_0/XOR GND 1.13fF
C798 a_n2140_n8646# GND 0.58fF
C799 a_575_n6996# GND 0.02fF
C800 a_425_n6996# GND 0.02fF
C801 a_n787_n6086# GND 0.03fF
C802 a_n2045_n6086# GND 0.03fF
C803 a_n2195_n6086# GND 0.03fF
C804 a_n2345_n6086# GND 0.03fF
C805 a_275_n6086# GND 0.90fF
C806 CMOS_s2_0/CMOS_4in_AND_0/OUT GND 0.85fF $ **FLOATING
C807 CMOS_s2_0/CMOS_3in_OR_0/A GND 0.56fF
C808 a_n787_n6996# GND 0.46fF
C809 a_n2345_n6996# GND 0.47fF
C810 a_425_n5418# GND 0.03fF
C811 a_n432_n5418# GND 0.03fF
C812 a_n732_n5418# GND 0.02fF
C813 a_n1990_n5418# GND 0.02fF
C814 a_n2290_n5418# GND 0.02fF
C815 CMOS_s2_0/CMOS_3in_OR_0/B GND 1.97fF
C816 a_n432_n4808# GND 0.01fF
C817 a_n732_n4808# GND 0.01fF
C818 CMOS_s2_0/CMOS_AND_1/A GND 1.08fF
C819 a_n1990_n4808# GND 0.01fF
C820 a_n2290_n4808# GND 0.01fF
C821 a_425_n4808# GND 0.52fF
C822 CMOS_s2_0/CMOS_XOR_0/XOR GND 1.12fF
C823 a_n2140_n5418# GND 0.59fF
C824 a_575_n3768# GND 0.02fF
C825 a_425_n3768# GND 0.02fF
C826 a_n787_n2858# GND 0.03fF
C827 a_n2195_n2858# GND 0.03fF
C828 a_n2345_n2858# GND 0.03fF
C829 a_275_n2858# GND 0.90fF
C830 CMOS_s1_0/CMOS_3in_OR_0/C GND 1.18fF $ **FLOATING
C831 CMOS_s1_0/CMOS_3in_OR_0/A GND 0.56fF
C832 a_n787_n3768# GND 0.47fF
C833 a_n2495_n3768# GND 0.63fF
C834 a_425_n2190# GND 0.02fF
C835 a_n432_n2190# GND 0.03fF
C836 a_n732_n2190# GND 0.02fF
C837 a_n1990_n2190# GND 0.02fF
C838 a_n2290_n2190# GND 0.02fF
C839 CMOS_s1_0/CMOS_3in_OR_0/B GND 1.95fF
C840 a_n432_n1580# GND 0.01fF
C841 a_n732_n1580# GND 0.01fF
C842 CMOS_s1_0/CMOS_AND_1/A GND 1.08fF
C843 a_n1990_n1580# GND 0.01fF
C844 a_n2290_n1580# GND 0.01fF
C845 a_425_n1580# GND 0.50fF
C846 CMOS_s1_0/CMOS_XOR_0/XOR GND 1.12fF
C847 a_n2140_n2190# GND 0.58fF
C848 a_n1990_n540# GND 0.00fF
C849 a_n2290_n540# GND 0.00fF
C850 a_425_370# GND 0.03fF
C851 a_n787_370# GND 0.03fF
C852 a_n1990_370# GND 0.02fF
C853 a_n2290_370# GND 0.01fF
C854 a_425_n540# GND 0.52fF
C855 CMOS_s0_0/CMOS_AND_1/B GND 0.86fF
C856 a_n787_n540# GND 0.46fF
C857 a_n2140_n540# GND 0.54fF
C858 CMOS_s0_0/CMOS_AND_1/A GND 0.95fF
C859 x2 GND 5.93fF
C860 a_425_1038# GND 0.03fF
C861 a_n1990_1038# GND 0.02fF
C862 a_n2290_1038# GND 0.01fF
C863 a_1637_1648# GND 0.02fF
C864 a_n787_1648# GND 0.01fF
C865 a_n1990_1648# GND 0.00fF
C866 a_n2290_1648# GND 0.00fF
C867 a_1637_1038# GND 0.67fF
C868 CMOS_s0_0/CMOS_AND_1/AND GND 1.28fF
C869 CMOS_s0_0/CMOS_AND_0/AND GND 0.64fF
C870 a_425_1648# GND 0.50fF
C871 CMOS_s0_0/CMOS_XOR_0/XOR GND 1.60fF
C872 CMOS_s0_0/CMOS_AND_0/B GND 0.57fF
C873 a_n787_1038# GND 0.61fF
C874 x1 GND 7.76fF
C875 x3 GND 3.72fF
C876 VDD GND 89.82fF
C877 CMOS_s0_0/x1_bar GND 2.51fF $ **FLOATING
C878 x1_bar.t1 GND 0.18fF
C879 x1_bar.t0 GND 0.26fF
C880 x1_bar.n0 GND 0.37fF $ **FLOATING
C881 CMOS_s0_0/CMOS_AND_2/B GND 0.62fF $ **FLOATING
C882 x1_bar.n1 GND 5.36fF $ **FLOATING
C883 x1_bar.t7 GND 0.42fF
C884 x1_bar.t9 GND 0.37fF
C885 CMOS_s3_0/x1_bar GND 6.56fF $ **FLOATING
C886 x1_bar.t5 GND 0.18fF
C887 x1_bar.t3 GND 0.26fF
C888 x1_bar.n2 GND 0.36fF $ **FLOATING
C889 CMOS_s2_0/CMOS_AND_1/B GND 0.05fF $ **FLOATING
C890 x1_bar.n3 GND 0.95fF $ **FLOATING
C891 x1_bar.n4 GND 2.73fF $ **FLOATING
C892 x1_bar.t8 GND 0.42fF
C893 x1_bar.t2 GND 0.37fF
C894 CMOS_s2_0/CMOS_XOR_0/A_bar GND 0.69fF $ **FLOATING
C895 x1_bar.n5 GND 4.45fF $ **FLOATING
C896 CMOS_s2_0/x1_bar GND 2.52fF $ **FLOATING
C897 x1_bar.t4 GND 0.42fF
C898 x1_bar.t6 GND 0.37fF
C899 CMOS_s1_0/CMOS_XOR_0/A_bar GND 0.69fF $ **FLOATING
C900 x1_bar.n6 GND 5.24fF $ **FLOATING
C901 CMOS_s1_0/x1_bar GND 1.55fF $ **FLOATING
C902 CMOS_s3_0/CMOS_3in_OR_0/C.t3 GND 0.10fF
C903 CMOS_s3_0/CMOS_3in_OR_0/C.t2 GND 0.12fF
C904 CMOS_s3_0/CMOS_3in_OR_0/C.t1 GND 0.31fF
C905 CMOS_s3_0/CMOS_3in_OR_0/C.t0 GND 0.29fF
C906 CMOS_s3_0/CMOS_3in_AND_0/OUT GND 0.19fF $ **FLOATING
C907 CMOS_s3_0/CMOS_3in_OR_0/C.n0 GND 0.70fF $ **FLOATING
C908 x1.t10 GND 0.19fF
C909 x1.t11 GND 0.13fF
C910 x1.n0 GND 0.27fF $ **FLOATING
C911 x1.n1 GND 1.68fF $ **FLOATING
C912 x1.t5 GND 0.26fF
C913 x1.t6 GND 0.10fF
C914 x1.n2 GND 0.29fF $ **FLOATING
C915 CMOS_s3_0/CMOS_XNOR_0/A GND 0.38fF $ **FLOATING
C916 x1.n3 GND 5.28fF $ **FLOATING
C917 CMOS_s3_0/x1 GND 1.48fF $ **FLOATING
C918 x1.t13 GND 0.26fF
C919 x1.t9 GND 0.10fF
C920 x1.n4 GND 0.28fF $ **FLOATING
C921 CMOS_s2_0/CMOS_XOR_0/A GND 0.04fF $ **FLOATING
C922 x1.n5 GND 1.38fF $ **FLOATING
C923 x1.t2 GND 0.28fF
C924 x1.t7 GND 0.24fF
C925 x1.n6 GND 0.36fF $ **FLOATING
C926 CMOS_s2_0/CMOS_4in_AND_0/B GND 0.41fF $ **FLOATING
C927 x1.n7 GND 2.50fF $ **FLOATING
C928 CMOS_s2_0/x1 GND 1.89fF $ **FLOATING
C929 x1.t3 GND 0.26fF
C930 x1.t1 GND 0.10fF
C931 x1.n8 GND 0.28fF $ **FLOATING
C932 CMOS_s1_0/CMOS_XOR_0/A GND 0.04fF $ **FLOATING
C933 x1.n9 GND 1.45fF $ **FLOATING
C934 x1.t8 GND 0.28fF
C935 x1.t12 GND 0.24fF
C936 x1.n10 GND 0.38fF $ **FLOATING
C937 CMOS_s1_0/CMOS_3in_AND_0/B GND 0.37fF $ **FLOATING
C938 x1.n11 GND 2.46fF $ **FLOATING
C939 CMOS_s1_0/x1 GND 2.83fF $ **FLOATING
C940 x1.t0 GND 0.19fF
C941 x1.t4 GND 0.13fF
C942 x1.n12 GND 0.27fF $ **FLOATING
C943 CMOS_s0_0/CMOS_OR_1/A GND 0.52fF $ **FLOATING
C944 x1.n13 GND 3.99fF $ **FLOATING
C945 CMOS_s0_0/x1 GND 0.08fF $ **FLOATING
C946 CMOS_s1_0/CMOS_3in_OR_0/C.t3 GND 0.12fF
C947 CMOS_s1_0/CMOS_3in_OR_0/C.t2 GND 0.14fF
C948 CMOS_s1_0/CMOS_3in_OR_0/C.t1 GND 0.37fF
C949 CMOS_s1_0/CMOS_3in_OR_0/C.t0 GND 0.34fF
C950 CMOS_s1_0/CMOS_3in_AND_0/OUT GND 0.23fF $ **FLOATING
C951 CMOS_s1_0/CMOS_3in_OR_0/C.n0 GND 0.84fF $ **FLOATING
C952 x2.t7 GND 0.31fF
C953 x2.t4 GND 0.12fF
C954 x2.n0 GND 0.34fF $ **FLOATING
C955 x2.n1 GND 1.93fF $ **FLOATING
C956 CMOS_s3_0/x2 GND 5.54fF $ **FLOATING
C957 x2.t3 GND 0.26fF
C958 x2.t0 GND 0.32fF
C959 CMOS_s2_0/CMOS_4in_AND_0/D GND 0.52fF $ **FLOATING
C960 x2.n2 GND 2.71fF $ **FLOATING
C961 x2.t9 GND 0.89fF
C962 x2.t1 GND 0.60fF
C963 CMOS_s2_0/CMOS_XNOR_0/B GND 0.70fF $ **FLOATING
C964 x2.n3 GND 2.78fF $ **FLOATING
C965 CMOS_s2_0/x2 GND 2.33fF $ **FLOATING
C966 x2.t5 GND 0.89fF
C967 x2.t8 GND 0.60fF
C968 CMOS_s1_0/CMOS_XNOR_0/B GND 0.70fF $ **FLOATING
C969 x2.n4 GND 2.92fF $ **FLOATING
C970 CMOS_s1_0/x2 GND 1.22fF $ **FLOATING
C971 x2.t2 GND 0.34fF
C972 x2.t6 GND 0.28fF
C973 CMOS_s0_0/CMOS_AND_2/A GND 0.50fF $ **FLOATING
C974 x2.n5 GND 4.51fF $ **FLOATING
C975 CMOS_s0_0/x2 GND 0.09fF $ **FLOATING
C976 CMOS_s0_0/x2_bar GND 1.22fF $ **FLOATING
C977 x2_bar.t2 GND 0.36fF
C978 x2_bar.t7 GND 0.30fF
C979 CMOS_s0_0/CMOS_OR_1/B GND 0.60fF $ **FLOATING
C980 x2_bar.n0 GND 4.65fF $ **FLOATING
C981 x2_bar.t9 GND 0.25fF
C982 x2_bar.t10 GND 0.17fF
C983 x2_bar.n1 GND 0.35fF $ **FLOATING
C984 CMOS_s1_0/CMOS_AND_0/B GND 0.05fF $ **FLOATING
C985 x2_bar.n2 GND 1.62fF $ **FLOATING
C986 x2_bar.t1 GND 0.25fF
C987 x2_bar.t3 GND 0.17fF
C988 x2_bar.n3 GND 0.35fF $ **FLOATING
C989 CMOS_s2_0/CMOS_AND_0/B GND 0.05fF $ **FLOATING
C990 x2_bar.n4 GND 1.62fF $ **FLOATING
C991 x2_bar.t8 GND 0.40fF
C992 x2_bar.t13 GND 0.35fF
C993 CMOS_s3_0/CMOS_XOR_0/A_bar GND 0.62fF $ **FLOATING
C994 x2_bar.t0 GND 0.28fF
C995 x2_bar.t5 GND 0.33fF
C996 x2_bar.n5 GND 0.50fF $ **FLOATING
C997 x2_bar.n6 GND 7.07fF $ **FLOATING
C998 CMOS_s3_0/x2_bar GND 2.34fF $ **FLOATING
C999 x2_bar.n7 GND 4.06fF $ **FLOATING
C1000 x2_bar.t4 GND 0.29fF
C1001 x2_bar.t12 GND 0.28fF
C1002 x2_bar.n8 GND 0.76fF $ **FLOATING
C1003 CMOS_s2_0/CMOS_XNOR_0/B_bar GND 0.27fF $ **FLOATING
C1004 x2_bar.n9 GND 1.93fF $ **FLOATING
C1005 CMOS_s2_0/x2_bar GND 1.60fF $ **FLOATING
C1006 x2_bar.n10 GND 4.06fF $ **FLOATING
C1007 x2_bar.t11 GND 0.29fF
C1008 x2_bar.t6 GND 0.28fF
C1009 x2_bar.n11 GND 0.76fF $ **FLOATING
C1010 CMOS_s1_0/CMOS_XNOR_0/B_bar GND 0.27fF $ **FLOATING
C1011 x2_bar.n12 GND 1.93fF $ **FLOATING
C1012 CMOS_s1_0/x2_bar GND 1.96fF $ **FLOATING
C1013 CMOS_s0_0/x3_bar GND 0.56fF $ **FLOATING
C1014 x3_bar.t5 GND 0.21fF
C1015 x3_bar.t2 GND 0.21fF
C1016 x3_bar.n0 GND 0.56fF $ **FLOATING
C1017 CMOS_s0_0/CMOS_XOR_0/B_bar GND 0.14fF $ **FLOATING
C1018 x3_bar.n1 GND 1.24fF $ **FLOATING
C1019 x3_bar.t15 GND 0.29fF
C1020 x3_bar.t8 GND 0.26fF
C1021 CMOS_s0_0/CMOS_XNOR_0/A_bar GND 0.42fF $ **FLOATING
C1022 x3_bar.n2 GND 1.82fF $ **FLOATING
C1023 x3_bar.t1 GND 0.29fF
C1024 x3_bar.t6 GND 0.26fF
C1025 CMOS_s2_0/CMOS_XNOR_0/A_bar GND 0.42fF $ **FLOATING
C1026 x3_bar.t3 GND 0.12fF
C1027 x3_bar.t12 GND 0.18fF
C1028 x3_bar.n3 GND 0.25fF $ **FLOATING
C1029 CMOS_s3_0/CMOS_AND_1/B GND 0.03fF $ **FLOATING
C1030 x3_bar.n4 GND 0.81fF $ **FLOATING
C1031 x3_bar.t10 GND 0.21fF
C1032 x3_bar.t7 GND 0.19fF
C1033 x3_bar.n5 GND 1.24fF $ **FLOATING
C1034 x3_bar.n6 GND 4.45fF $ **FLOATING
C1035 CMOS_s3_0/x3_bar GND 1.39fF $ **FLOATING
C1036 x3_bar.t0 GND 0.09fF
C1037 x3_bar.t13 GND 0.21fF
C1038 x3_bar.n7 GND 0.22fF $ **FLOATING
C1039 CMOS_s2_0/CMOS_4in_AND_0/A GND 0.30fF $ **FLOATING
C1040 x3_bar.n8 GND 1.48fF $ **FLOATING
C1041 x3_bar.n9 GND 1.61fF $ **FLOATING
C1042 CMOS_s2_0/x3_bar GND 0.88fF $ **FLOATING
C1043 x3_bar.t14 GND 0.20fF
C1044 x3_bar.t11 GND 0.24fF
C1045 CMOS_s1_0/CMOS_3in_AND_0/A GND 0.03fF $ **FLOATING
C1046 x3_bar.n10 GND 0.27fF $ **FLOATING
C1047 x3_bar.n11 GND 1.89fF $ **FLOATING
C1048 x3_bar.t9 GND 0.21fF
C1049 x3_bar.t4 GND 0.19fF
C1050 CMOS_s1_0/CMOS_XOR_0/B_bar GND 0.03fF $ **FLOATING
C1051 x3_bar.n12 GND 1.24fF $ **FLOATING
C1052 x3_bar.n13 GND 2.74fF $ **FLOATING
C1053 CMOS_s1_0/x3_bar GND 1.61fF $ **FLOATING
C1054 CMOS_s0_0/x0 GND 0.51fF $ **FLOATING
C1055 x0.t2 GND 0.19fF
C1056 x0.t7 GND 0.08fF
C1057 x0.n0 GND 0.22fF $ **FLOATING
C1058 CMOS_s0_0/CMOS_XOR_0/A GND 0.33fF $ **FLOATING
C1059 x0.n1 GND 1.79fF $ **FLOATING
C1060 x0.t4 GND 0.56fF
C1061 x0.t10 GND 0.38fF
C1062 CMOS_s0_0/CMOS_XNOR_0/B GND 0.54fF $ **FLOATING
C1063 x0.n2 GND 1.51fF $ **FLOATING
C1064 x0.t12 GND 0.21fF
C1065 x0.t1 GND 0.18fF
C1066 x0.t9 GND 0.56fF
C1067 x0.t13 GND 0.38fF
C1068 CMOS_s3_0/CMOS_XNOR_0/B GND 0.54fF $ **FLOATING
C1069 x0.n3 GND 3.76fF $ **FLOATING
C1070 CMOS_s3_0/x0 GND 0.51fF $ **FLOATING
C1071 x0.t11 GND 0.10fF
C1072 x0.t6 GND 0.15fF
C1073 x0.n4 GND 0.18fF $ **FLOATING
C1074 CMOS_s2_0/CMOS_4in_AND_0/C GND 0.35fF $ **FLOATING
C1075 x0.n5 GND 1.85fF $ **FLOATING
C1076 x0.t0 GND 0.56fF
C1077 x0.t3 GND 0.38fF
C1078 CMOS_s2_0/CMOS_XOR_0/B GND 0.42fF $ **FLOATING
C1079 x0.n6 GND 2.52fF $ **FLOATING
C1080 CMOS_s2_0/x0 GND 1.03fF $ **FLOATING
C1081 x0.t5 GND 0.19fF
C1082 x0.t8 GND 0.08fF
C1083 x0.n7 GND 0.22fF $ **FLOATING
C1084 CMOS_s1_0/CMOS_XNOR_0/A GND 0.33fF $ **FLOATING
C1085 x0.n8 GND 1.88fF $ **FLOATING
C1086 CMOS_s1_0/x0 GND 0.56fF $ **FLOATING
C1087 CMOS_s0_0/x0_bar GND 0.92fF $ **FLOATING
C1088 x0_bar.t8 GND 0.30fF
C1089 x0_bar.t9 GND 0.26fF
C1090 CMOS_s0_0/CMOS_XOR_0/A_bar GND 0.64fF $ **FLOATING
C1091 x0_bar.n0 GND 1.95fF $ **FLOATING
C1092 x0_bar.t11 GND 0.21fF
C1093 x0_bar.t1 GND 0.21fF
C1094 x0_bar.n1 GND 0.57fF $ **FLOATING
C1095 CMOS_s0_0/CMOS_XNOR_0/B_bar GND 0.33fF $ **FLOATING
C1096 x0_bar.n2 GND 1.56fF $ **FLOATING
C1097 x0_bar.t10 GND 0.21fF
C1098 x0_bar.t3 GND 0.21fF
C1099 x0_bar.n3 GND 0.57fF $ **FLOATING
C1100 CMOS_s3_0/x0_bar GND 5.05fF $ **FLOATING
C1101 x0_bar.t0 GND 0.21fF
C1102 x0_bar.t5 GND 0.20fF
C1103 CMOS_s2_0/CMOS_XOR_0/B_bar GND 0.03fF $ **FLOATING
C1104 x0_bar.n4 GND 1.45fF $ **FLOATING
C1105 x0_bar.n5 GND 3.16fF $ **FLOATING
C1106 CMOS_s2_0/x0_bar GND 1.34fF $ **FLOATING
C1107 x0_bar.t4 GND 0.13fF
C1108 x0_bar.t2 GND 0.19fF
C1109 x0_bar.n6 GND 0.23fF $ **FLOATING
C1110 CMOS_s1_0/CMOS_3in_AND_0/C GND 0.38fF $ **FLOATING
C1111 x0_bar.n7 GND 1.56fF $ **FLOATING
C1112 x0_bar.t6 GND 0.30fF
C1113 x0_bar.t7 GND 0.26fF
C1114 CMOS_s1_0/CMOS_XNOR_0/A_bar GND 0.64fF $ **FLOATING
C1115 x0_bar.n8 GND 1.94fF $ **FLOATING
C1116 CMOS_s1_0/x0_bar GND 1.34fF $ **FLOATING
C1117 x3.t10 GND 0.13fF
C1118 x3.t2 GND 0.20fF
C1119 x3.n0 GND 0.24fF $ **FLOATING
C1120 x3.t7 GND 0.76fF
C1121 x3.t12 GND 0.51fF
C1122 CMOS_s3_0/CMOS_XOR_0/B GND 0.49fF $ **FLOATING
C1123 x3.n1 GND 5.87fF $ **FLOATING
C1124 CMOS_s3_0/x3 GND 1.41fF $ **FLOATING
C1125 x3.t11 GND 0.26fF
C1126 x3.t13 GND 0.10fF
C1127 x3.n2 GND 0.30fF $ **FLOATING
C1128 CMOS_s2_0/CMOS_XNOR_0/A GND 0.25fF $ **FLOATING
C1129 x3.n3 GND 2.35fF $ **FLOATING
C1130 CMOS_s2_0/x3 GND 1.19fF $ **FLOATING
C1131 x3.t0 GND 0.14fF
C1132 x3.t8 GND 0.20fF
C1133 x3.n4 GND 0.28fF $ **FLOATING
C1134 CMOS_s1_0/CMOS_AND_1/B GND 0.04fF $ **FLOATING
C1135 x3.n5 GND 0.63fF $ **FLOATING
C1136 x3.n6 GND 2.95fF $ **FLOATING
C1137 x3.t6 GND 0.76fF
C1138 x3.t9 GND 0.51fF
C1139 CMOS_s1_0/CMOS_XOR_0/B GND 0.49fF $ **FLOATING
C1140 x3.n7 GND 3.12fF $ **FLOATING
C1141 CMOS_s1_0/x3 GND 0.76fF $ **FLOATING
C1142 x3.t1 GND 0.10fF
C1143 x3.t3 GND 0.26fF
C1144 x3.n8 GND 0.30fF $ **FLOATING
C1145 CMOS_s0_0/CMOS_XNOR_0/A GND 0.25fF $ **FLOATING
C1146 x3.n9 GND 2.30fF $ **FLOATING
C1147 x3.t4 GND 0.76fF
C1148 x3.t5 GND 0.51fF
C1149 CMOS_s0_0/CMOS_XOR_0/B GND 0.53fF $ **FLOATING
C1150 x3.n10 GND 1.76fF $ **FLOATING
C1151 CMOS_s0_0/x3 GND 0.08fF $ **FLOATING
C1152 VDD.t141 GND 0.05fF
C1153 VDD.t44 GND 0.05fF
C1154 VDD.n0 GND 0.22fF $ **FLOATING
C1155 CMOS_s3_0/CMOS_3in_AND_0/VDD GND 0.01fF $ **FLOATING
C1156 VDD.t57 GND 0.08fF
C1157 VDD.t73 GND 0.08fF
C1158 VDD.t55 GND 0.08fF
C1159 CMOS_s3_0/CMOS_AND_1/VDD GND 0.01fF $ **FLOATING
C1160 VDD.t69 GND 0.08fF
C1161 VDD.t67 GND 0.08fF
C1162 VDD.t111 GND 0.08fF
C1163 VDD.n1 GND 0.24fF $ **FLOATING
C1164 VDD.n2 GND 0.02fF $ **FLOATING
C1165 VDD.n3 GND 0.02fF $ **FLOATING
C1166 VDD.n4 GND 0.19fF $ **FLOATING
C1167 VDD.t110 GND 0.11fF
C1168 VDD.n5 GND 0.13fF $ **FLOATING
C1169 VDD.n6 GND 0.02fF $ **FLOATING
C1170 VDD.n7 GND 0.02fF $ **FLOATING
C1171 VDD.n8 GND 0.06fF $ **FLOATING
C1172 VDD.n9 GND 0.44fF $ **FLOATING
C1173 VDD.n10 GND 0.20fF $ **FLOATING
C1174 VDD.n11 GND 0.02fF $ **FLOATING
C1175 VDD.n12 GND 0.02fF $ **FLOATING
C1176 VDD.n13 GND 0.01fF $ **FLOATING
C1177 VDD.n14 GND 0.20fF $ **FLOATING
C1178 VDD.n15 GND 0.02fF $ **FLOATING
C1179 VDD.n16 GND 0.02fF $ **FLOATING
C1180 VDD.n17 GND 0.02fF $ **FLOATING
C1181 VDD.n18 GND 0.20fF $ **FLOATING
C1182 VDD.n19 GND 0.02fF $ **FLOATING
C1183 VDD.n20 GND 0.02fF $ **FLOATING
C1184 VDD.n21 GND 0.02fF $ **FLOATING
C1185 VDD.n22 GND 0.20fF $ **FLOATING
C1186 VDD.n23 GND 0.02fF $ **FLOATING
C1187 VDD.n24 GND 0.02fF $ **FLOATING
C1188 VDD.n25 GND 0.02fF $ **FLOATING
C1189 VDD.t0 GND 0.10fF
C1190 VDD.n26 GND 0.12fF $ **FLOATING
C1191 VDD.n27 GND 0.02fF $ **FLOATING
C1192 VDD.n28 GND 0.02fF $ **FLOATING
C1193 VDD.n29 GND 0.02fF $ **FLOATING
C1194 VDD.n30 GND 0.01fF $ **FLOATING
C1195 VDD.n31 GND 0.18fF $ **FLOATING
C1196 VDD.n32 GND 0.02fF $ **FLOATING
C1197 VDD.n33 GND 0.02fF $ **FLOATING
C1198 VDD.t133 GND 0.10fF
C1199 VDD.n34 GND 0.13fF $ **FLOATING
C1200 VDD.n35 GND 0.02fF $ **FLOATING
C1201 VDD.n36 GND 0.02fF $ **FLOATING
C1202 VDD.n37 GND 0.02fF $ **FLOATING
C1203 VDD.n38 GND 0.18fF $ **FLOATING
C1204 VDD.n39 GND 0.02fF $ **FLOATING
C1205 VDD.n40 GND 0.02fF $ **FLOATING
C1206 VDD.n41 GND 0.02fF $ **FLOATING
C1207 VDD.t66 GND 0.12fF
C1208 VDD.n42 GND 0.13fF $ **FLOATING
C1209 VDD.n43 GND 0.02fF $ **FLOATING
C1210 VDD.n44 GND 0.02fF $ **FLOATING
C1211 VDD.n45 GND 0.02fF $ **FLOATING
C1212 VDD.n46 GND 0.22fF $ **FLOATING
C1213 VDD.n47 GND 0.02fF $ **FLOATING
C1214 VDD.n48 GND 0.02fF $ **FLOATING
C1215 VDD.n49 GND 0.02fF $ **FLOATING
C1216 VDD.n50 GND 0.44fF $ **FLOATING
C1217 VDD.n51 GND 0.21fF $ **FLOATING
C1218 VDD.n52 GND 0.07fF $ **FLOATING
C1219 VDD.n53 GND 0.18fF $ **FLOATING
C1220 VDD.n54 GND 0.07fF $ **FLOATING
C1221 VDD.n55 GND 0.23fF $ **FLOATING
C1222 VDD.n56 GND 0.02fF $ **FLOATING
C1223 VDD.n57 GND 0.02fF $ **FLOATING
C1224 VDD.n58 GND 0.02fF $ **FLOATING
C1225 VDD.t68 GND 0.11fF
C1226 VDD.n59 GND 0.12fF $ **FLOATING
C1227 VDD.n60 GND 0.02fF $ **FLOATING
C1228 VDD.n61 GND 0.02fF $ **FLOATING
C1229 VDD.n62 GND 0.02fF $ **FLOATING
C1230 VDD.n63 GND 0.44fF $ **FLOATING
C1231 VDD.n64 GND 0.20fF $ **FLOATING
C1232 VDD.n65 GND 0.02fF $ **FLOATING
C1233 VDD.n66 GND 0.02fF $ **FLOATING
C1234 VDD.n67 GND 0.01fF $ **FLOATING
C1235 VDD.n68 GND 0.20fF $ **FLOATING
C1236 VDD.n69 GND 0.02fF $ **FLOATING
C1237 VDD.n70 GND 0.02fF $ **FLOATING
C1238 VDD.n71 GND 0.02fF $ **FLOATING
C1239 VDD.n72 GND 0.20fF $ **FLOATING
C1240 VDD.n73 GND 0.02fF $ **FLOATING
C1241 VDD.n74 GND 0.02fF $ **FLOATING
C1242 VDD.n75 GND 0.02fF $ **FLOATING
C1243 VDD.t71 GND 0.08fF
C1244 VDD.n76 GND 0.43fF $ **FLOATING
C1245 VDD.n77 GND 0.01fF $ **FLOATING
C1246 VDD.n78 GND 0.20fF $ **FLOATING
C1247 VDD.n79 GND 0.02fF $ **FLOATING
C1248 VDD.n80 GND 0.02fF $ **FLOATING
C1249 VDD.t70 GND 0.10fF
C1250 VDD.n81 GND 0.13fF $ **FLOATING
C1251 VDD.n82 GND 0.02fF $ **FLOATING
C1252 VDD.n83 GND 0.02fF $ **FLOATING
C1253 VDD.n84 GND 0.02fF $ **FLOATING
C1254 VDD.n85 GND 0.18fF $ **FLOATING
C1255 VDD.n86 GND 0.02fF $ **FLOATING
C1256 VDD.n87 GND 0.02fF $ **FLOATING
C1257 VDD.n88 GND 0.02fF $ **FLOATING
C1258 VDD.t54 GND 0.12fF
C1259 VDD.n89 GND 0.13fF $ **FLOATING
C1260 VDD.n90 GND 0.02fF $ **FLOATING
C1261 VDD.n91 GND 0.02fF $ **FLOATING
C1262 VDD.n92 GND 0.02fF $ **FLOATING
C1263 VDD.n93 GND 0.22fF $ **FLOATING
C1264 VDD.n94 GND 0.02fF $ **FLOATING
C1265 VDD.n95 GND 0.02fF $ **FLOATING
C1266 VDD.n96 GND 0.02fF $ **FLOATING
C1267 VDD.n97 GND 0.44fF $ **FLOATING
C1268 VDD.n98 GND 0.21fF $ **FLOATING
C1269 VDD.n99 GND 0.10fF $ **FLOATING
C1270 VDD.n100 GND 0.20fF $ **FLOATING
C1271 VDD.n101 GND 0.11fF $ **FLOATING
C1272 VDD.n102 GND 0.23fF $ **FLOATING
C1273 VDD.n103 GND 0.02fF $ **FLOATING
C1274 VDD.n104 GND 0.02fF $ **FLOATING
C1275 VDD.n105 GND 0.02fF $ **FLOATING
C1276 VDD.t72 GND 0.11fF
C1277 VDD.n106 GND 0.13fF $ **FLOATING
C1278 VDD.n107 GND 0.02fF $ **FLOATING
C1279 VDD.n108 GND 0.02fF $ **FLOATING
C1280 VDD.n109 GND 0.02fF $ **FLOATING
C1281 VDD.n110 GND 0.44fF $ **FLOATING
C1282 VDD.n111 GND 0.20fF $ **FLOATING
C1283 VDD.n112 GND 0.02fF $ **FLOATING
C1284 VDD.n113 GND 0.02fF $ **FLOATING
C1285 VDD.n114 GND 0.01fF $ **FLOATING
C1286 VDD.n115 GND 0.20fF $ **FLOATING
C1287 VDD.n116 GND 0.02fF $ **FLOATING
C1288 VDD.n117 GND 0.02fF $ **FLOATING
C1289 VDD.n118 GND 0.02fF $ **FLOATING
C1290 VDD.n119 GND 0.20fF $ **FLOATING
C1291 VDD.n120 GND 0.02fF $ **FLOATING
C1292 VDD.n121 GND 0.02fF $ **FLOATING
C1293 VDD.n122 GND 0.02fF $ **FLOATING
C1294 VDD.n123 GND 0.20fF $ **FLOATING
C1295 VDD.n124 GND 0.02fF $ **FLOATING
C1296 VDD.n125 GND 0.02fF $ **FLOATING
C1297 VDD.n126 GND 0.01fF $ **FLOATING
C1298 VDD.n127 GND 0.44fF $ **FLOATING
C1299 VDD.t56 GND 0.10fF
C1300 VDD.n128 GND 0.12fF $ **FLOATING
C1301 VDD.n129 GND 0.02fF $ **FLOATING
C1302 VDD.n130 GND 0.02fF $ **FLOATING
C1303 VDD.n131 GND 0.02fF $ **FLOATING
C1304 VDD.n132 GND 0.01fF $ **FLOATING
C1305 VDD.n133 GND 0.18fF $ **FLOATING
C1306 VDD.n134 GND 0.02fF $ **FLOATING
C1307 VDD.n135 GND 0.02fF $ **FLOATING
C1308 VDD.t140 GND 0.10fF
C1309 VDD.n136 GND 0.13fF $ **FLOATING
C1310 VDD.n137 GND 0.02fF $ **FLOATING
C1311 VDD.n138 GND 0.02fF $ **FLOATING
C1312 VDD.n139 GND 0.02fF $ **FLOATING
C1313 VDD.n140 GND 0.18fF $ **FLOATING
C1314 VDD.n141 GND 0.02fF $ **FLOATING
C1315 VDD.n142 GND 0.02fF $ **FLOATING
C1316 VDD.n143 GND 0.01fF $ **FLOATING
C1317 VDD.n144 GND 0.19fF $ **FLOATING
C1318 VDD.t43 GND 0.12fF
C1319 VDD.n145 GND 0.13fF $ **FLOATING
C1320 VDD.n146 GND 0.02fF $ **FLOATING
C1321 VDD.n147 GND 0.02fF $ **FLOATING
C1322 VDD.n148 GND 0.02fF $ **FLOATING
C1323 VDD.n149 GND 0.22fF $ **FLOATING
C1324 VDD.n150 GND 0.02fF $ **FLOATING
C1325 VDD.n151 GND 0.02fF $ **FLOATING
C1326 VDD.n152 GND 0.02fF $ **FLOATING
C1327 VDD.n153 GND 0.21fF $ **FLOATING
C1328 VDD.n154 GND 0.42fF $ **FLOATING
C1329 VDD.t115 GND 0.08fF
C1330 VDD.t145 GND 0.08fF
C1331 CMOS_s3_0/CMOS_XNOR_0/VDD GND 0.01fF $ **FLOATING
C1332 VDD.t88 GND 0.08fF
C1333 VDD.t126 GND 0.08fF
C1334 VDD.t6 GND 0.08fF
C1335 VDD.t13 GND 0.08fF
C1336 VDD.t128 GND 0.08fF
C1337 VDD.t139 GND 0.08fF
C1338 CMOS_s3_0/CMOS_XOR_0/VDD GND 0.02fF $ **FLOATING
C1339 VDD.t25 GND 0.08fF
C1340 VDD.t61 GND 0.08fF
C1341 VDD.t2 GND 0.08fF
C1342 VDD.t153 GND 0.08fF
C1343 CMOS_s3_0/CMOS_AND_0/VDD GND 0.02fF $ **FLOATING
C1344 VDD.t120 GND 0.08fF
C1345 VDD.t137 GND 0.08fF
C1346 VDD.n155 GND 0.30fF $ **FLOATING
C1347 VDD.n156 GND 0.02fF $ **FLOATING
C1348 VDD.n157 GND 0.02fF $ **FLOATING
C1349 VDD.n158 GND 0.11fF $ **FLOATING
C1350 VDD.t136 GND 0.17fF
C1351 VDD.n159 GND 0.14fF $ **FLOATING
C1352 VDD.n160 GND 0.04fF $ **FLOATING
C1353 VDD.n161 GND 0.03fF $ **FLOATING
C1354 VDD.n162 GND 0.08fF $ **FLOATING
C1355 VDD.n163 GND 0.44fF $ **FLOATING
C1356 VDD.n164 GND 0.23fF $ **FLOATING
C1357 VDD.n165 GND 0.04fF $ **FLOATING
C1358 VDD.n166 GND 0.03fF $ **FLOATING
C1359 VDD.n167 GND 0.02fF $ **FLOATING
C1360 VDD.n168 GND 0.23fF $ **FLOATING
C1361 VDD.n169 GND 0.04fF $ **FLOATING
C1362 VDD.n170 GND 0.03fF $ **FLOATING
C1363 VDD.n171 GND 0.04fF $ **FLOATING
C1364 VDD.n172 GND 0.44fF $ **FLOATING
C1365 VDD.n173 GND 0.23fF $ **FLOATING
C1366 VDD.n174 GND 0.04fF $ **FLOATING
C1367 VDD.n175 GND 0.03fF $ **FLOATING
C1368 VDD.n176 GND 0.02fF $ **FLOATING
C1369 VDD.n177 GND 0.23fF $ **FLOATING
C1370 VDD.n178 GND 0.04fF $ **FLOATING
C1371 VDD.n179 GND 0.03fF $ **FLOATING
C1372 VDD.n180 GND 0.04fF $ **FLOATING
C1373 VDD.t135 GND 0.07fF
C1374 VDD.n181 GND 0.13fF $ **FLOATING
C1375 VDD.n182 GND 0.04fF $ **FLOATING
C1376 VDD.n183 GND 0.03fF $ **FLOATING
C1377 VDD.n184 GND 0.04fF $ **FLOATING
C1378 VDD.t147 GND 0.08fF
C1379 VDD.n185 GND 0.43fF $ **FLOATING
C1380 VDD.n186 GND 0.02fF $ **FLOATING
C1381 VDD.t119 GND 0.65fF
C1382 VDD.t152 GND 0.52fF
C1383 VDD.t146 GND 0.28fF
C1384 VDD.n187 GND 0.50fF $ **FLOATING
C1385 VDD.n188 GND 0.16fF $ **FLOATING
C1386 VDD.n189 GND 0.04fF $ **FLOATING
C1387 VDD.n190 GND 0.03fF $ **FLOATING
C1388 VDD.t9 GND 0.11fF
C1389 VDD.n191 GND 0.14fF $ **FLOATING
C1390 VDD.n192 GND 0.04fF $ **FLOATING
C1391 VDD.n193 GND 0.03fF $ **FLOATING
C1392 VDD.n194 GND 0.03fF $ **FLOATING
C1393 VDD.n195 GND 0.20fF $ **FLOATING
C1394 VDD.n196 GND 0.04fF $ **FLOATING
C1395 VDD.n197 GND 0.03fF $ **FLOATING
C1396 VDD.n198 GND 0.04fF $ **FLOATING
C1397 VDD.t1 GND 0.13fF
C1398 VDD.n199 GND 0.15fF $ **FLOATING
C1399 VDD.n200 GND 0.04fF $ **FLOATING
C1400 VDD.n201 GND 0.03fF $ **FLOATING
C1401 VDD.n202 GND 0.04fF $ **FLOATING
C1402 VDD.n203 GND 0.24fF $ **FLOATING
C1403 VDD.n204 GND 0.04fF $ **FLOATING
C1404 VDD.n205 GND 0.03fF $ **FLOATING
C1405 VDD.n206 GND 0.03fF $ **FLOATING
C1406 VDD.n207 GND 0.87fF $ **FLOATING
C1407 VDD.n208 GND 0.29fF $ **FLOATING
C1408 VDD.n209 GND 0.12fF $ **FLOATING
C1409 VDD.n210 GND 0.24fF $ **FLOATING
C1410 VDD.n211 GND 0.13fF $ **FLOATING
C1411 VDD.n212 GND 0.25fF $ **FLOATING
C1412 VDD.n213 GND 0.04fF $ **FLOATING
C1413 VDD.n214 GND 0.03fF $ **FLOATING
C1414 VDD.n215 GND 0.02fF $ **FLOATING
C1415 VDD.n216 GND 0.44fF $ **FLOATING
C1416 VDD.t24 GND 0.12fF
C1417 VDD.n217 GND 0.13fF $ **FLOATING
C1418 VDD.n218 GND 0.04fF $ **FLOATING
C1419 VDD.n219 GND 0.03fF $ **FLOATING
C1420 VDD.n220 GND 0.03fF $ **FLOATING
C1421 VDD.n221 GND 0.44fF $ **FLOATING
C1422 VDD.n222 GND 0.23fF $ **FLOATING
C1423 VDD.n223 GND 0.04fF $ **FLOATING
C1424 VDD.n224 GND 0.03fF $ **FLOATING
C1425 VDD.n225 GND 0.02fF $ **FLOATING
C1426 VDD.n226 GND 0.23fF $ **FLOATING
C1427 VDD.n227 GND 0.04fF $ **FLOATING
C1428 VDD.n228 GND 0.03fF $ **FLOATING
C1429 VDD.n229 GND 0.04fF $ **FLOATING
C1430 VDD.t60 GND 0.59fF
C1431 VDD.t89 GND 0.23fF
C1432 VDD.t138 GND 0.57fF
C1433 VDD.t130 GND 0.24fF
C1434 VDD.n230 GND 0.27fF $ **FLOATING
C1435 VDD.n231 GND 0.16fF $ **FLOATING
C1436 VDD.n232 GND 0.04fF $ **FLOATING
C1437 VDD.n233 GND 0.03fF $ **FLOATING
C1438 VDD.n234 GND 0.04fF $ **FLOATING
C1439 VDD.t124 GND 0.08fF
C1440 VDD.n235 GND 0.43fF $ **FLOATING
C1441 VDD.n236 GND 0.02fF $ **FLOATING
C1442 VDD.n237 GND 0.19fF $ **FLOATING
C1443 VDD.n238 GND 0.04fF $ **FLOATING
C1444 VDD.n239 GND 0.03fF $ **FLOATING
C1445 VDD.t123 GND 0.11fF
C1446 VDD.n240 GND 0.14fF $ **FLOATING
C1447 VDD.n241 GND 0.04fF $ **FLOATING
C1448 VDD.n242 GND 0.03fF $ **FLOATING
C1449 VDD.n243 GND 0.03fF $ **FLOATING
C1450 VDD.n244 GND 0.20fF $ **FLOATING
C1451 VDD.n245 GND 0.04fF $ **FLOATING
C1452 VDD.n246 GND 0.03fF $ **FLOATING
C1453 VDD.n247 GND 0.04fF $ **FLOATING
C1454 VDD.t127 GND 0.13fF
C1455 VDD.n248 GND 0.15fF $ **FLOATING
C1456 VDD.n249 GND 0.04fF $ **FLOATING
C1457 VDD.n250 GND 0.03fF $ **FLOATING
C1458 VDD.n251 GND 0.03fF $ **FLOATING
C1459 VDD.n252 GND 0.44fF $ **FLOATING
C1460 VDD.n253 GND 0.24fF $ **FLOATING
C1461 VDD.n254 GND 0.04fF $ **FLOATING
C1462 VDD.n255 GND 0.03fF $ **FLOATING
C1463 VDD.n256 GND 0.01fF $ **FLOATING
C1464 VDD.n257 GND 0.44fF $ **FLOATING
C1465 VDD.n258 GND 0.29fF $ **FLOATING
C1466 VDD.n259 GND 0.12fF $ **FLOATING
C1467 VDD.n260 GND 0.05fF $ **FLOATING
C1468 VDD.n261 GND 0.02fF $ **FLOATING
C1469 VDD.n262 GND 0.02fF $ **FLOATING
C1470 VDD.n263 GND 0.13fF $ **FLOATING
C1471 VDD.n264 GND 0.30fF $ **FLOATING
C1472 VDD.n265 GND 0.04fF $ **FLOATING
C1473 VDD.n266 GND 0.03fF $ **FLOATING
C1474 VDD.n267 GND 0.04fF $ **FLOATING
C1475 VDD.n268 GND 0.19fF $ **FLOATING
C1476 VDD.n269 GND 0.04fF $ **FLOATING
C1477 VDD.n270 GND 0.03fF $ **FLOATING
C1478 VDD.n271 GND 0.03fF $ **FLOATING
C1479 VDD.n272 GND 0.44fF $ **FLOATING
C1480 VDD.t5 GND 0.11fF
C1481 VDD.n273 GND 0.15fF $ **FLOATING
C1482 VDD.n274 GND 0.04fF $ **FLOATING
C1483 VDD.n275 GND 0.03fF $ **FLOATING
C1484 VDD.n276 GND 0.02fF $ **FLOATING
C1485 VDD.n277 GND 0.44fF $ **FLOATING
C1486 VDD.n278 GND 0.23fF $ **FLOATING
C1487 VDD.n279 GND 0.04fF $ **FLOATING
C1488 VDD.n280 GND 0.03fF $ **FLOATING
C1489 VDD.n281 GND 0.02fF $ **FLOATING
C1490 VDD.n282 GND 0.23fF $ **FLOATING
C1491 VDD.n283 GND 0.04fF $ **FLOATING
C1492 VDD.n284 GND 0.03fF $ **FLOATING
C1493 VDD.n285 GND 0.04fF $ **FLOATING
C1494 VDD.n286 GND 0.23fF $ **FLOATING
C1495 VDD.n287 GND 0.04fF $ **FLOATING
C1496 VDD.n288 GND 0.03fF $ **FLOATING
C1497 VDD.n289 GND 0.02fF $ **FLOATING
C1498 VDD.n290 GND 0.44fF $ **FLOATING
C1499 VDD.n291 GND 0.23fF $ **FLOATING
C1500 VDD.n292 GND 0.04fF $ **FLOATING
C1501 VDD.n293 GND 0.03fF $ **FLOATING
C1502 VDD.n294 GND 0.01fF $ **FLOATING
C1503 VDD.n295 GND 0.44fF $ **FLOATING
C1504 VDD.t12 GND 0.77fF
C1505 VDD.t125 GND 0.49fF
C1506 VDD.t144 GND 0.57fF
C1507 VDD.t35 GND 0.31fF
C1508 VDD.t26 GND 0.24fF
C1509 VDD.n296 GND 0.26fF $ **FLOATING
C1510 VDD.t87 GND 0.03fF
C1511 VDD.n297 GND 0.12fF $ **FLOATING
C1512 VDD.n298 GND 0.04fF $ **FLOATING
C1513 VDD.n299 GND 0.03fF $ **FLOATING
C1514 VDD.n300 GND 0.04fF $ **FLOATING
C1515 VDD.n301 GND 0.20fF $ **FLOATING
C1516 VDD.n302 GND 0.04fF $ **FLOATING
C1517 VDD.n303 GND 0.03fF $ **FLOATING
C1518 VDD.n304 GND 0.04fF $ **FLOATING
C1519 VDD.t91 GND 0.11fF
C1520 VDD.n305 GND 0.13fF $ **FLOATING
C1521 VDD.n306 GND 0.04fF $ **FLOATING
C1522 VDD.n307 GND 0.03fF $ **FLOATING
C1523 VDD.n308 GND 0.04fF $ **FLOATING
C1524 VDD.t92 GND 0.05fF
C1525 VDD.t28 GND 0.05fF
C1526 VDD.n309 GND 0.22fF $ **FLOATING
C1527 VDD.n310 GND 0.18fF $ **FLOATING
C1528 VDD.n311 GND 0.02fF $ **FLOATING
C1529 VDD.n312 GND 0.21fF $ **FLOATING
C1530 VDD.n313 GND 0.04fF $ **FLOATING
C1531 VDD.n314 GND 0.03fF $ **FLOATING
C1532 VDD.t27 GND 0.11fF
C1533 VDD.n315 GND 0.14fF $ **FLOATING
C1534 VDD.n316 GND 0.04fF $ **FLOATING
C1535 VDD.n317 GND 0.03fF $ **FLOATING
C1536 VDD.n318 GND 0.03fF $ **FLOATING
C1537 VDD.n319 GND 0.20fF $ **FLOATING
C1538 VDD.n320 GND 0.04fF $ **FLOATING
C1539 VDD.n321 GND 0.03fF $ **FLOATING
C1540 VDD.n322 GND 0.04fF $ **FLOATING
C1541 VDD.t114 GND 0.13fF
C1542 VDD.n323 GND 0.15fF $ **FLOATING
C1543 VDD.n324 GND 0.04fF $ **FLOATING
C1544 VDD.n325 GND 0.03fF $ **FLOATING
C1545 VDD.n326 GND 0.03fF $ **FLOATING
C1546 VDD.n327 GND 0.44fF $ **FLOATING
C1547 VDD.n328 GND 0.24fF $ **FLOATING
C1548 VDD.n329 GND 0.04fF $ **FLOATING
C1549 VDD.n330 GND 0.03fF $ **FLOATING
C1550 VDD.n331 GND 0.01fF $ **FLOATING
C1551 VDD.n332 GND 0.44fF $ **FLOATING
C1552 VDD.n333 GND 0.29fF $ **FLOATING
C1553 VDD.n334 GND 0.04fF $ **FLOATING
C1554 CMOS_s3_0/VDD GND 0.02fF $ **FLOATING
C1555 VDD.n335 GND 0.79fF $ **FLOATING
C1556 VDD.t98 GND 0.08fF
C1557 VDD.t155 GND 0.05fF
C1558 VDD.t132 GND 0.05fF
C1559 VDD.n336 GND 0.22fF $ **FLOATING
C1560 CMOS_s2_0/CMOS_XNOR_0/VDD GND 0.02fF $ **FLOATING
C1561 VDD.t63 GND 0.08fF
C1562 VDD.t96 GND 0.08fF
C1563 VDD.t50 GND 0.08fF
C1564 VDD.t52 GND 0.08fF
C1565 VDD.t113 GND 0.08fF
C1566 VDD.t150 GND 0.08fF
C1567 CMOS_s2_0/CMOS_XOR_0/VDD GND 0.02fF $ **FLOATING
C1568 VDD.t84 GND 0.08fF
C1569 VDD.t38 GND 0.08fF
C1570 VDD.t80 GND 0.08fF
C1571 VDD.t15 GND 0.08fF
C1572 CMOS_s2_0/CMOS_AND_0/VDD GND 0.02fF $ **FLOATING
C1573 VDD.t109 GND 0.08fF
C1574 VDD.t59 GND 0.08fF
C1575 VDD.n337 GND 0.30fF $ **FLOATING
C1576 VDD.n338 GND 0.02fF $ **FLOATING
C1577 VDD.n339 GND 0.02fF $ **FLOATING
C1578 VDD.n340 GND 0.11fF $ **FLOATING
C1579 VDD.t58 GND 0.17fF
C1580 VDD.n341 GND 0.14fF $ **FLOATING
C1581 VDD.n342 GND 0.04fF $ **FLOATING
C1582 VDD.n343 GND 0.03fF $ **FLOATING
C1583 VDD.n344 GND 0.08fF $ **FLOATING
C1584 VDD.n345 GND 0.44fF $ **FLOATING
C1585 VDD.n346 GND 0.23fF $ **FLOATING
C1586 VDD.n347 GND 0.04fF $ **FLOATING
C1587 VDD.n348 GND 0.03fF $ **FLOATING
C1588 VDD.n349 GND 0.02fF $ **FLOATING
C1589 VDD.n350 GND 0.23fF $ **FLOATING
C1590 VDD.n351 GND 0.04fF $ **FLOATING
C1591 VDD.n352 GND 0.03fF $ **FLOATING
C1592 VDD.n353 GND 0.04fF $ **FLOATING
C1593 VDD.n354 GND 0.44fF $ **FLOATING
C1594 VDD.n355 GND 0.23fF $ **FLOATING
C1595 VDD.n356 GND 0.04fF $ **FLOATING
C1596 VDD.n357 GND 0.03fF $ **FLOATING
C1597 VDD.n358 GND 0.02fF $ **FLOATING
C1598 VDD.n359 GND 0.23fF $ **FLOATING
C1599 VDD.n360 GND 0.04fF $ **FLOATING
C1600 VDD.n361 GND 0.03fF $ **FLOATING
C1601 VDD.n362 GND 0.04fF $ **FLOATING
C1602 VDD.t129 GND 0.07fF
C1603 VDD.n363 GND 0.13fF $ **FLOATING
C1604 VDD.n364 GND 0.04fF $ **FLOATING
C1605 VDD.n365 GND 0.03fF $ **FLOATING
C1606 VDD.n366 GND 0.04fF $ **FLOATING
C1607 VDD.t65 GND 0.08fF
C1608 VDD.n367 GND 0.43fF $ **FLOATING
C1609 VDD.n368 GND 0.02fF $ **FLOATING
C1610 VDD.t108 GND 0.65fF
C1611 VDD.t14 GND 0.52fF
C1612 VDD.t64 GND 0.28fF
C1613 VDD.n369 GND 0.50fF $ **FLOATING
C1614 VDD.n370 GND 0.16fF $ **FLOATING
C1615 VDD.n371 GND 0.04fF $ **FLOATING
C1616 VDD.n372 GND 0.03fF $ **FLOATING
C1617 VDD.t134 GND 0.11fF
C1618 VDD.n373 GND 0.14fF $ **FLOATING
C1619 VDD.n374 GND 0.04fF $ **FLOATING
C1620 VDD.n375 GND 0.03fF $ **FLOATING
C1621 VDD.n376 GND 0.03fF $ **FLOATING
C1622 VDD.n377 GND 0.20fF $ **FLOATING
C1623 VDD.n378 GND 0.04fF $ **FLOATING
C1624 VDD.n379 GND 0.03fF $ **FLOATING
C1625 VDD.n380 GND 0.04fF $ **FLOATING
C1626 VDD.t79 GND 0.13fF
C1627 VDD.n381 GND 0.15fF $ **FLOATING
C1628 VDD.n382 GND 0.04fF $ **FLOATING
C1629 VDD.n383 GND 0.03fF $ **FLOATING
C1630 VDD.n384 GND 0.04fF $ **FLOATING
C1631 VDD.n385 GND 0.24fF $ **FLOATING
C1632 VDD.n386 GND 0.04fF $ **FLOATING
C1633 VDD.n387 GND 0.03fF $ **FLOATING
C1634 VDD.n388 GND 0.03fF $ **FLOATING
C1635 VDD.n389 GND 0.87fF $ **FLOATING
C1636 VDD.n390 GND 0.29fF $ **FLOATING
C1637 VDD.n391 GND 0.12fF $ **FLOATING
C1638 VDD.n392 GND 0.24fF $ **FLOATING
C1639 VDD.n393 GND 0.13fF $ **FLOATING
C1640 VDD.n394 GND 0.25fF $ **FLOATING
C1641 VDD.n395 GND 0.04fF $ **FLOATING
C1642 VDD.n396 GND 0.03fF $ **FLOATING
C1643 VDD.n397 GND 0.02fF $ **FLOATING
C1644 VDD.n398 GND 0.44fF $ **FLOATING
C1645 VDD.t83 GND 0.12fF
C1646 VDD.n399 GND 0.13fF $ **FLOATING
C1647 VDD.n400 GND 0.04fF $ **FLOATING
C1648 VDD.n401 GND 0.03fF $ **FLOATING
C1649 VDD.n402 GND 0.03fF $ **FLOATING
C1650 VDD.n403 GND 0.44fF $ **FLOATING
C1651 VDD.n404 GND 0.23fF $ **FLOATING
C1652 VDD.n405 GND 0.04fF $ **FLOATING
C1653 VDD.n406 GND 0.03fF $ **FLOATING
C1654 VDD.n407 GND 0.02fF $ **FLOATING
C1655 VDD.n408 GND 0.23fF $ **FLOATING
C1656 VDD.n409 GND 0.04fF $ **FLOATING
C1657 VDD.n410 GND 0.03fF $ **FLOATING
C1658 VDD.n411 GND 0.04fF $ **FLOATING
C1659 VDD.t37 GND 0.59fF
C1660 VDD.t29 GND 0.23fF
C1661 VDD.t149 GND 0.57fF
C1662 VDD.t151 GND 0.24fF
C1663 VDD.n412 GND 0.27fF $ **FLOATING
C1664 VDD.n413 GND 0.16fF $ **FLOATING
C1665 VDD.n414 GND 0.04fF $ **FLOATING
C1666 VDD.n415 GND 0.03fF $ **FLOATING
C1667 VDD.n416 GND 0.04fF $ **FLOATING
C1668 VDD.t77 GND 0.08fF
C1669 VDD.n417 GND 0.43fF $ **FLOATING
C1670 VDD.n418 GND 0.02fF $ **FLOATING
C1671 VDD.n419 GND 0.19fF $ **FLOATING
C1672 VDD.n420 GND 0.04fF $ **FLOATING
C1673 VDD.n421 GND 0.03fF $ **FLOATING
C1674 VDD.t76 GND 0.11fF
C1675 VDD.n422 GND 0.14fF $ **FLOATING
C1676 VDD.n423 GND 0.04fF $ **FLOATING
C1677 VDD.n424 GND 0.03fF $ **FLOATING
C1678 VDD.n425 GND 0.03fF $ **FLOATING
C1679 VDD.n426 GND 0.20fF $ **FLOATING
C1680 VDD.n427 GND 0.04fF $ **FLOATING
C1681 VDD.n428 GND 0.03fF $ **FLOATING
C1682 VDD.n429 GND 0.04fF $ **FLOATING
C1683 VDD.t112 GND 0.13fF
C1684 VDD.n430 GND 0.15fF $ **FLOATING
C1685 VDD.n431 GND 0.04fF $ **FLOATING
C1686 VDD.n432 GND 0.03fF $ **FLOATING
C1687 VDD.n433 GND 0.03fF $ **FLOATING
C1688 VDD.n434 GND 0.44fF $ **FLOATING
C1689 VDD.n435 GND 0.24fF $ **FLOATING
C1690 VDD.n436 GND 0.04fF $ **FLOATING
C1691 VDD.n437 GND 0.03fF $ **FLOATING
C1692 VDD.n438 GND 0.01fF $ **FLOATING
C1693 VDD.n439 GND 0.44fF $ **FLOATING
C1694 VDD.n440 GND 0.29fF $ **FLOATING
C1695 VDD.n441 GND 0.12fF $ **FLOATING
C1696 VDD.n442 GND 0.03fF $ **FLOATING
C1697 VDD.n443 GND 0.13fF $ **FLOATING
C1698 VDD.n444 GND 0.15fF $ **FLOATING
C1699 VDD.n445 GND 0.01fF $ **FLOATING
C1700 VDD.n446 GND 0.02fF $ **FLOATING
C1701 VDD.n447 GND 0.02fF $ **FLOATING
C1702 VDD.n448 GND 0.04fF $ **FLOATING
C1703 VDD.n449 GND 0.02fF $ **FLOATING
C1704 VDD.n450 GND 0.02fF $ **FLOATING
C1705 VDD.n451 GND 0.03fF $ **FLOATING
C1706 VDD.n452 GND 0.44fF $ **FLOATING
C1707 VDD.t51 GND 0.24fF
C1708 VDD.n453 GND 0.25fF $ **FLOATING
C1709 VDD.n454 GND 0.23fF $ **FLOATING
C1710 VDD.n455 GND 0.04fF $ **FLOATING
C1711 VDD.n456 GND 0.03fF $ **FLOATING
C1712 VDD.n457 GND 0.02fF $ **FLOATING
C1713 VDD.n458 GND 0.23fF $ **FLOATING
C1714 VDD.n459 GND 0.04fF $ **FLOATING
C1715 VDD.n460 GND 0.03fF $ **FLOATING
C1716 VDD.n461 GND 0.04fF $ **FLOATING
C1717 VDD.n462 GND 0.23fF $ **FLOATING
C1718 VDD.n463 GND 0.04fF $ **FLOATING
C1719 VDD.n464 GND 0.03fF $ **FLOATING
C1720 VDD.n465 GND 0.03fF $ **FLOATING
C1721 VDD.n466 GND 0.44fF $ **FLOATING
C1722 VDD.n467 GND 0.23fF $ **FLOATING
C1723 VDD.n468 GND 0.04fF $ **FLOATING
C1724 VDD.n469 GND 0.03fF $ **FLOATING
C1725 VDD.n470 GND 0.01fF $ **FLOATING
C1726 VDD.n471 GND 0.44fF $ **FLOATING
C1727 VDD.t95 GND 0.11fF
C1728 VDD.n472 GND 0.15fF $ **FLOATING
C1729 VDD.n473 GND 0.04fF $ **FLOATING
C1730 VDD.n474 GND 0.03fF $ **FLOATING
C1731 VDD.n475 GND 0.03fF $ **FLOATING
C1732 VDD.n476 GND 0.19fF $ **FLOATING
C1733 VDD.n477 GND 0.04fF $ **FLOATING
C1734 VDD.n478 GND 0.03fF $ **FLOATING
C1735 VDD.n479 GND 0.04fF $ **FLOATING
C1736 VDD.t49 GND 0.71fF
C1737 VDD.t131 GND 0.51fF
C1738 VDD.t154 GND 0.31fF
C1739 VDD.t62 GND 0.22fF
C1740 VDD.t45 GND 0.08fF
C1741 VDD.n480 GND 0.46fF $ **FLOATING
C1742 VDD.n481 GND 0.15fF $ **FLOATING
C1743 VDD.n482 GND 0.04fF $ **FLOATING
C1744 VDD.n483 GND 0.03fF $ **FLOATING
C1745 VDD.n484 GND 0.02fF $ **FLOATING
C1746 VDD.n485 GND 0.44fF $ **FLOATING
C1747 VDD.n486 GND 0.18fF $ **FLOATING
C1748 VDD.n487 GND 0.04fF $ **FLOATING
C1749 VDD.n488 GND 0.03fF $ **FLOATING
C1750 VDD.n489 GND 0.04fF $ **FLOATING
C1751 VDD.n490 GND 0.02fF $ **FLOATING
C1752 VDD.n491 GND 0.17fF $ **FLOATING
C1753 VDD.n492 GND 0.04fF $ **FLOATING
C1754 VDD.n493 GND 0.03fF $ **FLOATING
C1755 VDD.t53 GND 0.11fF
C1756 VDD.n494 GND 0.17fF $ **FLOATING
C1757 VDD.n495 GND 0.04fF $ **FLOATING
C1758 VDD.n496 GND 0.03fF $ **FLOATING
C1759 VDD.n497 GND 0.03fF $ **FLOATING
C1760 VDD.n498 GND 0.18fF $ **FLOATING
C1761 VDD.n499 GND 0.04fF $ **FLOATING
C1762 VDD.n500 GND 0.03fF $ **FLOATING
C1763 VDD.n501 GND 0.02fF $ **FLOATING
C1764 VDD.n502 GND 0.20fF $ **FLOATING
C1765 VDD.t97 GND 0.11fF
C1766 VDD.n503 GND 0.16fF $ **FLOATING
C1767 VDD.n504 GND 0.04fF $ **FLOATING
C1768 VDD.n505 GND 0.03fF $ **FLOATING
C1769 VDD.n506 GND 0.02fF $ **FLOATING
C1770 VDD.n507 GND 0.44fF $ **FLOATING
C1771 VDD.n508 GND 0.23fF $ **FLOATING
C1772 VDD.n509 GND 0.04fF $ **FLOATING
C1773 VDD.n510 GND 0.03fF $ **FLOATING
C1774 VDD.n511 GND 0.03fF $ **FLOATING
C1775 VDD.n512 GND 0.21fF $ **FLOATING
C1776 VDD.n513 GND 0.04fF $ **FLOATING
C1777 VDD.n514 GND 0.04fF $ **FLOATING
C1778 VDD.n515 GND 0.05fF $ **FLOATING
C1779 CMOS_s2_0/VDD GND 0.02fF $ **FLOATING
C1780 VDD.n516 GND 0.78fF $ **FLOATING
C1781 VDD.t23 GND 0.08fF
C1782 VDD.t90 GND 0.08fF
C1783 CMOS_s1_0/CMOS_XNOR_0/VDD GND 0.02fF $ **FLOATING
C1784 VDD.t148 GND 0.08fF
C1785 VDD.t117 GND 0.08fF
C1786 VDD.t46 GND 0.08fF
C1787 VDD.t20 GND 0.08fF
C1788 VDD.t103 GND 0.08fF
C1789 VDD.t32 GND 0.08fF
C1790 CMOS_s1_0/CMOS_XOR_0/VDD GND 0.02fF $ **FLOATING
C1791 VDD.t34 GND 0.08fF
C1792 VDD.t86 GND 0.08fF
C1793 VDD.t118 GND 0.08fF
C1794 VDD.t105 GND 0.08fF
C1795 CMOS_s1_0/CMOS_AND_0/VDD GND 0.02fF $ **FLOATING
C1796 VDD.t78 GND 0.08fF
C1797 VDD.t11 GND 0.08fF
C1798 VDD.n517 GND 0.44fF $ **FLOATING
C1799 VDD.n518 GND 0.04fF $ **FLOATING
C1800 VDD.n519 GND 0.03fF $ **FLOATING
C1801 VDD.n520 GND 0.35fF $ **FLOATING
C1802 VDD.t10 GND 0.21fF
C1803 VDD.n521 GND 0.22fF $ **FLOATING
C1804 VDD.n522 GND 0.04fF $ **FLOATING
C1805 VDD.n523 GND 0.03fF $ **FLOATING
C1806 VDD.n524 GND 0.11fF $ **FLOATING
C1807 VDD.n525 GND 0.87fF $ **FLOATING
C1808 VDD.n526 GND 0.38fF $ **FLOATING
C1809 VDD.n527 GND 0.04fF $ **FLOATING
C1810 VDD.n528 GND 0.03fF $ **FLOATING
C1811 VDD.n529 GND 0.02fF $ **FLOATING
C1812 VDD.n530 GND 0.38fF $ **FLOATING
C1813 VDD.n531 GND 0.04fF $ **FLOATING
C1814 VDD.n532 GND 0.03fF $ **FLOATING
C1815 VDD.n533 GND 0.04fF $ **FLOATING
C1816 VDD.n534 GND 0.38fF $ **FLOATING
C1817 VDD.n535 GND 0.04fF $ **FLOATING
C1818 VDD.n536 GND 0.03fF $ **FLOATING
C1819 VDD.n537 GND 0.04fF $ **FLOATING
C1820 VDD.t8 GND 0.08fF
C1821 VDD.t122 GND 0.08fF
C1822 VDD.n538 GND 0.86fF $ **FLOATING
C1823 VDD.n539 GND 0.02fF $ **FLOATING
C1824 VDD.n540 GND 0.38fF $ **FLOATING
C1825 VDD.n541 GND 0.04fF $ **FLOATING
C1826 VDD.n542 GND 0.03fF $ **FLOATING
C1827 VDD.t7 GND 0.19fF
C1828 VDD.n543 GND 0.24fF $ **FLOATING
C1829 VDD.n544 GND 0.04fF $ **FLOATING
C1830 VDD.n545 GND 0.03fF $ **FLOATING
C1831 VDD.n546 GND 0.03fF $ **FLOATING
C1832 VDD.n547 GND 0.33fF $ **FLOATING
C1833 VDD.n548 GND 0.04fF $ **FLOATING
C1834 VDD.n549 GND 0.03fF $ **FLOATING
C1835 VDD.n550 GND 0.04fF $ **FLOATING
C1836 VDD.t104 GND 0.22fF
C1837 VDD.n551 GND 0.25fF $ **FLOATING
C1838 VDD.n552 GND 0.04fF $ **FLOATING
C1839 VDD.n553 GND 0.03fF $ **FLOATING
C1840 VDD.n554 GND 0.04fF $ **FLOATING
C1841 VDD.n555 GND 0.41fF $ **FLOATING
C1842 VDD.n556 GND 0.04fF $ **FLOATING
C1843 VDD.n557 GND 0.03fF $ **FLOATING
C1844 VDD.n558 GND 0.03fF $ **FLOATING
C1845 VDD.n559 GND 0.87fF $ **FLOATING
C1846 VDD.n560 GND 0.41fF $ **FLOATING
C1847 VDD.n561 GND 0.12fF $ **FLOATING
C1848 VDD.n562 GND 0.24fF $ **FLOATING
C1849 VDD.n563 GND 0.13fF $ **FLOATING
C1850 VDD.n564 GND 0.25fF $ **FLOATING
C1851 VDD.n565 GND 0.04fF $ **FLOATING
C1852 VDD.n566 GND 0.03fF $ **FLOATING
C1853 VDD.n567 GND 0.02fF $ **FLOATING
C1854 VDD.n568 GND 0.44fF $ **FLOATING
C1855 VDD.t33 GND 0.12fF
C1856 VDD.n569 GND 0.13fF $ **FLOATING
C1857 VDD.n570 GND 0.04fF $ **FLOATING
C1858 VDD.n571 GND 0.03fF $ **FLOATING
C1859 VDD.n572 GND 0.03fF $ **FLOATING
C1860 VDD.n573 GND 0.44fF $ **FLOATING
C1861 VDD.n574 GND 0.23fF $ **FLOATING
C1862 VDD.n575 GND 0.04fF $ **FLOATING
C1863 VDD.n576 GND 0.03fF $ **FLOATING
C1864 VDD.n577 GND 0.02fF $ **FLOATING
C1865 VDD.n578 GND 0.23fF $ **FLOATING
C1866 VDD.n579 GND 0.04fF $ **FLOATING
C1867 VDD.n580 GND 0.03fF $ **FLOATING
C1868 VDD.n581 GND 0.04fF $ **FLOATING
C1869 VDD.t85 GND 0.59fF
C1870 VDD.t121 GND 0.23fF
C1871 VDD.t31 GND 0.57fF
C1872 VDD.t99 GND 0.24fF
C1873 VDD.n582 GND 0.27fF $ **FLOATING
C1874 VDD.n583 GND 0.16fF $ **FLOATING
C1875 VDD.n584 GND 0.04fF $ **FLOATING
C1876 VDD.n585 GND 0.03fF $ **FLOATING
C1877 VDD.n586 GND 0.04fF $ **FLOATING
C1878 VDD.t94 GND 0.08fF
C1879 VDD.n587 GND 0.43fF $ **FLOATING
C1880 VDD.n588 GND 0.02fF $ **FLOATING
C1881 VDD.n589 GND 0.19fF $ **FLOATING
C1882 VDD.n590 GND 0.04fF $ **FLOATING
C1883 VDD.n591 GND 0.03fF $ **FLOATING
C1884 VDD.t93 GND 0.11fF
C1885 VDD.n592 GND 0.14fF $ **FLOATING
C1886 VDD.n593 GND 0.04fF $ **FLOATING
C1887 VDD.n594 GND 0.03fF $ **FLOATING
C1888 VDD.n595 GND 0.03fF $ **FLOATING
C1889 VDD.n596 GND 0.20fF $ **FLOATING
C1890 VDD.n597 GND 0.04fF $ **FLOATING
C1891 VDD.n598 GND 0.03fF $ **FLOATING
C1892 VDD.n599 GND 0.04fF $ **FLOATING
C1893 VDD.t102 GND 0.13fF
C1894 VDD.n600 GND 0.15fF $ **FLOATING
C1895 VDD.n601 GND 0.04fF $ **FLOATING
C1896 VDD.n602 GND 0.03fF $ **FLOATING
C1897 VDD.n603 GND 0.03fF $ **FLOATING
C1898 VDD.n604 GND 0.44fF $ **FLOATING
C1899 VDD.n605 GND 0.24fF $ **FLOATING
C1900 VDD.n606 GND 0.04fF $ **FLOATING
C1901 VDD.n607 GND 0.03fF $ **FLOATING
C1902 VDD.n608 GND 0.01fF $ **FLOATING
C1903 VDD.n609 GND 0.44fF $ **FLOATING
C1904 VDD.n610 GND 0.29fF $ **FLOATING
C1905 VDD.n611 GND 0.12fF $ **FLOATING
C1906 VDD.n612 GND 0.38fF $ **FLOATING
C1907 VDD.n613 GND 0.13fF $ **FLOATING
C1908 VDD.n614 GND 0.42fF $ **FLOATING
C1909 VDD.n615 GND 0.04fF $ **FLOATING
C1910 VDD.n616 GND 0.03fF $ **FLOATING
C1911 VDD.n617 GND 0.04fF $ **FLOATING
C1912 VDD.t19 GND 0.21fF
C1913 VDD.n618 GND 0.24fF $ **FLOATING
C1914 VDD.n619 GND 0.04fF $ **FLOATING
C1915 VDD.n620 GND 0.03fF $ **FLOATING
C1916 VDD.n621 GND 0.03fF $ **FLOATING
C1917 VDD.n622 GND 0.87fF $ **FLOATING
C1918 VDD.n623 GND 0.38fF $ **FLOATING
C1919 VDD.n624 GND 0.04fF $ **FLOATING
C1920 VDD.n625 GND 0.03fF $ **FLOATING
C1921 VDD.n626 GND 0.02fF $ **FLOATING
C1922 VDD.n627 GND 0.38fF $ **FLOATING
C1923 VDD.n628 GND 0.04fF $ **FLOATING
C1924 VDD.n629 GND 0.03fF $ **FLOATING
C1925 VDD.n630 GND 0.04fF $ **FLOATING
C1926 VDD.n631 GND 0.38fF $ **FLOATING
C1927 VDD.n632 GND 0.04fF $ **FLOATING
C1928 VDD.n633 GND 0.03fF $ **FLOATING
C1929 VDD.n634 GND 0.04fF $ **FLOATING
C1930 VDD.n635 GND 0.38fF $ **FLOATING
C1931 VDD.n636 GND 0.04fF $ **FLOATING
C1932 VDD.n637 GND 0.03fF $ **FLOATING
C1933 VDD.n638 GND 0.02fF $ **FLOATING
C1934 VDD.n639 GND 0.87fF $ **FLOATING
C1935 VDD.t116 GND 0.19fF
C1936 VDD.n640 GND 0.25fF $ **FLOATING
C1937 VDD.n641 GND 0.04fF $ **FLOATING
C1938 VDD.n642 GND 0.03fF $ **FLOATING
C1939 VDD.n643 GND 0.03fF $ **FLOATING
C1940 VDD.n644 GND 0.32fF $ **FLOATING
C1941 VDD.n645 GND 0.04fF $ **FLOATING
C1942 VDD.n646 GND 0.03fF $ **FLOATING
C1943 VDD.n647 GND 0.04fF $ **FLOATING
C1944 VDD.t40 GND 0.19fF
C1945 VDD.n648 GND 0.27fF $ **FLOATING
C1946 VDD.n649 GND 0.04fF $ **FLOATING
C1947 VDD.n650 GND 0.03fF $ **FLOATING
C1948 VDD.n651 GND 0.04fF $ **FLOATING
C1949 VDD.n652 GND 0.30fF $ **FLOATING
C1950 VDD.n653 GND 0.04fF $ **FLOATING
C1951 VDD.n654 GND 0.03fF $ **FLOATING
C1952 VDD.n655 GND 0.04fF $ **FLOATING
C1953 VDD.n656 GND 0.02fF $ **FLOATING
C1954 VDD.n657 GND 0.28fF $ **FLOATING
C1955 VDD.n658 GND 0.04fF $ **FLOATING
C1956 VDD.n659 GND 0.03fF $ **FLOATING
C1957 VDD.t30 GND 0.19fF
C1958 VDD.n660 GND 0.29fF $ **FLOATING
C1959 VDD.n661 GND 0.04fF $ **FLOATING
C1960 VDD.n662 GND 0.03fF $ **FLOATING
C1961 VDD.n663 GND 0.03fF $ **FLOATING
C1962 VDD.n664 GND 0.30fF $ **FLOATING
C1963 VDD.n665 GND 0.04fF $ **FLOATING
C1964 VDD.n666 GND 0.03fF $ **FLOATING
C1965 VDD.n667 GND 0.04fF $ **FLOATING
C1966 VDD.t22 GND 0.19fF
C1967 VDD.n668 GND 0.29fF $ **FLOATING
C1968 VDD.n669 GND 0.04fF $ **FLOATING
C1969 VDD.n670 GND 0.03fF $ **FLOATING
C1970 VDD.n671 GND 0.03fF $ **FLOATING
C1971 VDD.n672 GND 0.87fF $ **FLOATING
C1972 VDD.n673 GND 0.43fF $ **FLOATING
C1973 VDD.n674 GND 0.04fF $ **FLOATING
C1974 VDD.n675 GND 0.03fF $ **FLOATING
C1975 VDD.n676 GND 0.03fF $ **FLOATING
C1976 VDD.n677 GND 0.24fF $ **FLOATING
C1977 VDD.n678 GND 0.05fF $ **FLOATING
C1978 CMOS_s1_0/VDD GND 0.02fF $ **FLOATING
C1979 VDD.n679 GND 0.78fF $ **FLOATING
C1980 VDD.t143 GND 0.08fF
C1981 CMOS_s0_0/CMOS_XOR_0/VDD GND 0.01fF $ **FLOATING
C1982 VDD.n680 GND 0.15fF $ **FLOATING
C1983 VDD.n681 GND 0.02fF $ **FLOATING
C1984 VDD.t17 GND 0.08fF
C1985 VDD.t101 GND 0.08fF
C1986 CMOS_s0_0/CMOS_OR_1/VDD GND 0.01fF $ **FLOATING
C1987 VDD.t48 GND 0.08fF
C1988 VDD.t42 GND 0.08fF
C1989 CMOS_s0_0/CMOS_AND_0/VDD GND 0.01fF $ **FLOATING
C1990 VDD.t82 GND 0.08fF
C1991 VDD.t75 GND 0.08fF
C1992 CMOS_s0_0/CMOS_OR_0/VDD GND 0.01fF $ **FLOATING
C1993 VDD.t4 GND 0.08fF
C1994 VDD.n682 GND 0.24fF $ **FLOATING
C1995 VDD.n683 GND 0.02fF $ **FLOATING
C1996 VDD.n684 GND 0.02fF $ **FLOATING
C1997 VDD.n685 GND 0.18fF $ **FLOATING
C1998 VDD.t3 GND 0.11fF
C1999 VDD.n686 GND 0.12fF $ **FLOATING
C2000 VDD.n687 GND 0.02fF $ **FLOATING
C2001 VDD.n688 GND 0.02fF $ **FLOATING
C2002 VDD.n689 GND 0.06fF $ **FLOATING
C2003 VDD.n690 GND 0.44fF $ **FLOATING
C2004 VDD.n691 GND 0.20fF $ **FLOATING
C2005 VDD.n692 GND 0.02fF $ **FLOATING
C2006 VDD.n693 GND 0.02fF $ **FLOATING
C2007 VDD.n694 GND 0.01fF $ **FLOATING
C2008 VDD.n695 GND 0.20fF $ **FLOATING
C2009 VDD.n696 GND 0.02fF $ **FLOATING
C2010 VDD.n697 GND 0.02fF $ **FLOATING
C2011 VDD.n698 GND 0.02fF $ **FLOATING
C2012 VDD.n699 GND 0.20fF $ **FLOATING
C2013 VDD.n700 GND 0.02fF $ **FLOATING
C2014 VDD.n701 GND 0.02fF $ **FLOATING
C2015 VDD.n702 GND 0.02fF $ **FLOATING
C2016 VDD.n703 GND 0.01fF $ **FLOATING
C2017 VDD.n704 GND 0.20fF $ **FLOATING
C2018 VDD.n705 GND 0.02fF $ **FLOATING
C2019 VDD.n706 GND 0.02fF $ **FLOATING
C2020 VDD.t36 GND 0.10fF
C2021 VDD.n707 GND 0.13fF $ **FLOATING
C2022 VDD.n708 GND 0.02fF $ **FLOATING
C2023 VDD.n709 GND 0.02fF $ **FLOATING
C2024 VDD.n710 GND 0.02fF $ **FLOATING
C2025 VDD.n711 GND 0.18fF $ **FLOATING
C2026 VDD.n712 GND 0.02fF $ **FLOATING
C2027 VDD.n713 GND 0.02fF $ **FLOATING
C2028 VDD.n714 GND 0.02fF $ **FLOATING
C2029 VDD.t74 GND 0.12fF
C2030 VDD.n715 GND 0.13fF $ **FLOATING
C2031 VDD.n716 GND 0.02fF $ **FLOATING
C2032 VDD.n717 GND 0.02fF $ **FLOATING
C2033 VDD.n718 GND 0.02fF $ **FLOATING
C2034 VDD.n719 GND 0.22fF $ **FLOATING
C2035 VDD.n720 GND 0.02fF $ **FLOATING
C2036 VDD.n721 GND 0.02fF $ **FLOATING
C2037 VDD.n722 GND 0.02fF $ **FLOATING
C2038 VDD.n723 GND 0.44fF $ **FLOATING
C2039 VDD.n724 GND 0.21fF $ **FLOATING
C2040 VDD.n725 GND 0.07fF $ **FLOATING
C2041 VDD.n726 GND 0.18fF $ **FLOATING
C2042 VDD.n727 GND 0.07fF $ **FLOATING
C2043 VDD.n728 GND 0.23fF $ **FLOATING
C2044 VDD.n729 GND 0.02fF $ **FLOATING
C2045 VDD.n730 GND 0.02fF $ **FLOATING
C2046 VDD.n731 GND 0.02fF $ **FLOATING
C2047 VDD.t81 GND 0.11fF
C2048 VDD.n732 GND 0.12fF $ **FLOATING
C2049 VDD.n733 GND 0.02fF $ **FLOATING
C2050 VDD.n734 GND 0.02fF $ **FLOATING
C2051 VDD.n735 GND 0.02fF $ **FLOATING
C2052 VDD.n736 GND 0.44fF $ **FLOATING
C2053 VDD.n737 GND 0.20fF $ **FLOATING
C2054 VDD.n738 GND 0.02fF $ **FLOATING
C2055 VDD.n739 GND 0.02fF $ **FLOATING
C2056 VDD.n740 GND 0.01fF $ **FLOATING
C2057 VDD.n741 GND 0.20fF $ **FLOATING
C2058 VDD.n742 GND 0.02fF $ **FLOATING
C2059 VDD.n743 GND 0.02fF $ **FLOATING
C2060 VDD.n744 GND 0.02fF $ **FLOATING
C2061 VDD.n745 GND 0.20fF $ **FLOATING
C2062 VDD.n746 GND 0.02fF $ **FLOATING
C2063 VDD.n747 GND 0.02fF $ **FLOATING
C2064 VDD.n748 GND 0.02fF $ **FLOATING
C2065 VDD.t107 GND 0.08fF
C2066 VDD.n749 GND 0.43fF $ **FLOATING
C2067 VDD.n750 GND 0.01fF $ **FLOATING
C2068 VDD.n751 GND 0.20fF $ **FLOATING
C2069 VDD.n752 GND 0.02fF $ **FLOATING
C2070 VDD.n753 GND 0.02fF $ **FLOATING
C2071 VDD.t106 GND 0.10fF
C2072 VDD.n754 GND 0.13fF $ **FLOATING
C2073 VDD.n755 GND 0.02fF $ **FLOATING
C2074 VDD.n756 GND 0.02fF $ **FLOATING
C2075 VDD.n757 GND 0.02fF $ **FLOATING
C2076 VDD.n758 GND 0.18fF $ **FLOATING
C2077 VDD.n759 GND 0.02fF $ **FLOATING
C2078 VDD.n760 GND 0.02fF $ **FLOATING
C2079 VDD.n761 GND 0.02fF $ **FLOATING
C2080 VDD.t41 GND 0.12fF
C2081 VDD.n762 GND 0.13fF $ **FLOATING
C2082 VDD.n763 GND 0.02fF $ **FLOATING
C2083 VDD.n764 GND 0.02fF $ **FLOATING
C2084 VDD.n765 GND 0.02fF $ **FLOATING
C2085 VDD.n766 GND 0.22fF $ **FLOATING
C2086 VDD.n767 GND 0.02fF $ **FLOATING
C2087 VDD.n768 GND 0.02fF $ **FLOATING
C2088 VDD.n769 GND 0.02fF $ **FLOATING
C2089 VDD.n770 GND 0.44fF $ **FLOATING
C2090 VDD.n771 GND 0.21fF $ **FLOATING
C2091 VDD.n772 GND 0.07fF $ **FLOATING
C2092 VDD.n773 GND 0.18fF $ **FLOATING
C2093 VDD.n774 GND 0.07fF $ **FLOATING
C2094 VDD.n775 GND 0.23fF $ **FLOATING
C2095 VDD.n776 GND 0.02fF $ **FLOATING
C2096 VDD.n777 GND 0.02fF $ **FLOATING
C2097 VDD.n778 GND 0.02fF $ **FLOATING
C2098 VDD.t47 GND 0.11fF
C2099 VDD.n779 GND 0.12fF $ **FLOATING
C2100 VDD.n780 GND 0.02fF $ **FLOATING
C2101 VDD.n781 GND 0.02fF $ **FLOATING
C2102 VDD.n782 GND 0.02fF $ **FLOATING
C2103 VDD.n783 GND 0.44fF $ **FLOATING
C2104 VDD.n784 GND 0.20fF $ **FLOATING
C2105 VDD.n785 GND 0.02fF $ **FLOATING
C2106 VDD.n786 GND 0.02fF $ **FLOATING
C2107 VDD.n787 GND 0.01fF $ **FLOATING
C2108 VDD.n788 GND 0.20fF $ **FLOATING
C2109 VDD.n789 GND 0.02fF $ **FLOATING
C2110 VDD.n790 GND 0.02fF $ **FLOATING
C2111 VDD.n791 GND 0.02fF $ **FLOATING
C2112 VDD.n792 GND 0.20fF $ **FLOATING
C2113 VDD.n793 GND 0.02fF $ **FLOATING
C2114 VDD.n794 GND 0.02fF $ **FLOATING
C2115 VDD.n795 GND 0.02fF $ **FLOATING
C2116 VDD.n796 GND 0.01fF $ **FLOATING
C2117 VDD.n797 GND 0.20fF $ **FLOATING
C2118 VDD.n798 GND 0.02fF $ **FLOATING
C2119 VDD.n799 GND 0.02fF $ **FLOATING
C2120 VDD.t18 GND 0.10fF
C2121 VDD.n800 GND 0.13fF $ **FLOATING
C2122 VDD.n801 GND 0.02fF $ **FLOATING
C2123 VDD.n802 GND 0.02fF $ **FLOATING
C2124 VDD.n803 GND 0.02fF $ **FLOATING
C2125 VDD.n804 GND 0.18fF $ **FLOATING
C2126 VDD.n805 GND 0.02fF $ **FLOATING
C2127 VDD.n806 GND 0.02fF $ **FLOATING
C2128 VDD.n807 GND 0.02fF $ **FLOATING
C2129 VDD.t100 GND 0.12fF
C2130 VDD.n808 GND 0.13fF $ **FLOATING
C2131 VDD.n809 GND 0.02fF $ **FLOATING
C2132 VDD.n810 GND 0.02fF $ **FLOATING
C2133 VDD.n811 GND 0.02fF $ **FLOATING
C2134 VDD.n812 GND 0.22fF $ **FLOATING
C2135 VDD.n813 GND 0.02fF $ **FLOATING
C2136 VDD.n814 GND 0.02fF $ **FLOATING
C2137 VDD.n815 GND 0.02fF $ **FLOATING
C2138 VDD.n816 GND 0.44fF $ **FLOATING
C2139 VDD.n817 GND 0.21fF $ **FLOATING
C2140 VDD.n818 GND 0.12fF $ **FLOATING
C2141 VDD.n819 GND 0.17fF $ **FLOATING
C2142 VDD.n820 GND 0.13fF $ **FLOATING
C2143 VDD.n821 GND 0.24fF $ **FLOATING
C2144 VDD.n822 GND 0.02fF $ **FLOATING
C2145 VDD.n823 GND 0.02fF $ **FLOATING
C2146 VDD.n824 GND 0.01fF $ **FLOATING
C2147 VDD.n825 GND 0.44fF $ **FLOATING
C2148 VDD.t16 GND 0.10fF
C2149 VDD.n826 GND 0.14fF $ **FLOATING
C2150 VDD.n827 GND 0.02fF $ **FLOATING
C2151 VDD.n828 GND 0.02fF $ **FLOATING
C2152 VDD.n829 GND 0.02fF $ **FLOATING
C2153 VDD.n830 GND 0.17fF $ **FLOATING
C2154 VDD.n831 GND 0.02fF $ **FLOATING
C2155 VDD.n832 GND 0.02fF $ **FLOATING
C2156 VDD.n833 GND 0.02fF $ **FLOATING
C2157 VDD.t21 GND 0.10fF
C2158 VDD.n834 GND 0.14fF $ **FLOATING
C2159 VDD.n835 GND 0.02fF $ **FLOATING
C2160 VDD.n836 GND 0.02fF $ **FLOATING
C2161 VDD.n837 GND 0.02fF $ **FLOATING
C2162 VDD.n838 GND 0.16fF $ **FLOATING
C2163 VDD.n839 GND 0.02fF $ **FLOATING
C2164 VDD.n840 GND 0.02fF $ **FLOATING
C2165 VDD.n841 GND 0.02fF $ **FLOATING
C2166 VDD.n842 GND 0.01fF $ **FLOATING
C2167 VDD.n843 GND 0.02fF $ **FLOATING
C2168 VDD.t39 GND 0.10fF
C2169 VDD.n844 GND 0.15fF $ **FLOATING
C2170 VDD.n845 GND 0.02fF $ **FLOATING
C2171 VDD.n846 GND 0.02fF $ **FLOATING
C2172 VDD.n847 GND 0.02fF $ **FLOATING
C2173 VDD.n848 GND 0.16fF $ **FLOATING
C2174 VDD.n849 GND 0.02fF $ **FLOATING
C2175 VDD.n850 GND 0.02fF $ **FLOATING
C2176 VDD.n851 GND 0.02fF $ **FLOATING
C2177 VDD.t142 GND 0.10fF
C2178 VDD.n852 GND 0.16fF $ **FLOATING
C2179 VDD.n853 GND 0.02fF $ **FLOATING
C2180 VDD.n854 GND 0.02fF $ **FLOATING
C2181 VDD.n855 GND 0.02fF $ **FLOATING
C2182 VDD.n856 GND 0.44fF $ **FLOATING
C2183 VDD.n857 GND 0.23fF $ **FLOATING
C2184 VDD.n858 GND 0.02fF $ **FLOATING
C2185 VDD.n859 GND 0.02fF $ **FLOATING
C2186 VDD.n860 GND 0.02fF $ **FLOATING
C2187 VDD.n861 GND 0.12fF $ **FLOATING
C2188 VDD.n862 GND 0.03fF $ **FLOATING
C2189 VDD.n863 GND 0.39fF $ **FLOATING
C2190 CMOS_s0_0/VDD GND 0.00fF $ **FLOATING
C2191 CMOS_s2_0/CMOS_4in_AND_0/OUT.t3 GND 0.11fF
C2192 CMOS_s2_0/CMOS_4in_AND_0/OUT.t2 GND 0.14fF
C2193 CMOS_s2_0/CMOS_4in_AND_0/OUT.t1 GND 0.37fF
C2194 CMOS_s2_0/CMOS_4in_AND_0/OUT.t0 GND 0.34fF
C2195 CMOS_s2_0/CMOS_4in_AND_0/OUT.n0 GND 0.81fF $ **FLOATING
C2196 CMOS_s2_0/CMOS_3in_OR_0/C GND 0.48fF $ **FLOATING
.ends

