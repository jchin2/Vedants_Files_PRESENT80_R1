magic
tech sky130A
timestamp 1679780349
<< metal2 >>
rect 0 0 30 30
rect 0 50 30 80
rect 0 100 30 130
rect 0 150 30 180
rect 0 200 30 230
rect 0 250 30 280
rect 0 300 30 330
rect 0 350 30 380
rect 0 400 30 430
rect 0 450 30 480
rect 0 500 30 530
rect 0 550 30 580
rect 0 600 30 630
rect 0 650 30 680
rect 0 700 30 730
rect 0 750 30 780
rect 0 800 30 830
rect 0 850 30 880
rect 0 900 30 930
rect 0 950 30 980
rect 0 1000 30 1030
rect 0 1050 30 1080
rect 0 1100 30 1130
rect 0 1150 30 1180
rect 0 1200 30 1230
rect 0 1250 30 1280
rect 0 1300 30 1330
rect 0 1350 30 1380
rect 0 1400 30 1430
rect 0 1450 30 1480
rect 0 1500 30 1530
rect 0 1550 30 1580
rect 0 1600 30 1630
rect 0 1650 30 1680
rect 0 1700 30 1730
rect 0 1750 30 1780
rect 0 1800 30 1830
rect 0 1850 30 1880
rect 0 1900 30 1930
rect 0 1950 30 1980
rect 0 2000 30 2030
rect 0 2050 30 2080
rect 0 2100 30 2130
rect 0 2150 30 2180
rect 0 2200 30 2230
rect 0 2250 30 2280
rect 0 2300 30 2330
rect 0 2350 30 2380
rect 0 2400 30 2430
rect 0 2450 30 2480
rect 0 2500 30 2530
rect 0 2550 30 2580
rect 0 2600 30 2630
rect 0 2650 30 2680
rect 0 2700 30 2730
rect 0 2750 30 2780
rect 0 2800 30 2830
rect 0 2850 30 2880
rect 0 2900 30 2930
rect 0 2950 30 2980
rect 0 3000 30 3030
rect 0 3050 30 3080
rect 0 3100 30 3130
rect 0 3150 30 3180
<< labels >>
rlabel metal2 0 0 30 30 1 s0
port 0 n
rlabel metal2 0 50 30 80 1 s1
port 1 n
rlabel metal2 0 100 30 130 1 s2
port 2 n
rlabel metal2 0 150 30 180 1 s3
port 3 n
rlabel metal2 0 200 30 230 1 s4
port 4 n
rlabel metal2 0 250 30 280 1 s5
port 5 n
rlabel metal2 0 300 30 330 1 s6
port 6 n
rlabel metal2 0 350 30 380 1 s7
port 7 n
rlabel metal2 0 400 30 430 1 s8
port 8 n
rlabel metal2 0 450 30 480 1 s9
port 9 n
rlabel metal2 0 500 30 530 1 s10
port 10 n
rlabel metal2 0 550 30 580 1 s11
port 11 n
rlabel metal2 0 600 30 630 1 s12
port 12 n
rlabel metal2 0 650 30 680 1 s13
port 13 n
rlabel metal2 0 700 30 730 1 s14
port 14 n
rlabel metal2 0 750 30 780 1 s15
port 15 n
rlabel metal2 0 800 30 830 1 s16
port 16 n
rlabel metal2 0 850 30 880 1 s17
port 17 n
rlabel metal2 0 900 30 930 1 s18
port 18 n
rlabel metal2 0 950 30 980 1 s19
port 19 n
rlabel metal2 0 1000 30 1030 1 s20
port 20 n
rlabel metal2 0 1050 30 1080 1 s21
port 21 n
rlabel metal2 0 1100 30 1130 1 s22
port 22 n
rlabel metal2 0 1150 30 1180 1 s23
port 23 n
rlabel metal2 0 1200 30 1230 1 s24
port 24 n
rlabel metal2 0 1250 30 1280 1 s25
port 25 n
rlabel metal2 0 1300 30 1330 1 s26
port 26 n
rlabel metal2 0 1350 30 1380 1 s27
port 27 n
rlabel metal2 0 1400 30 1430 1 s28
port 28 n
rlabel metal2 0 1450 30 1480 1 s29
port 29 n
rlabel metal2 0 1500 30 1530 1 s30
port 30 n
rlabel metal2 0 1550 30 1580 1 s31
port 31 n
rlabel metal2 0 1600 30 1630 1 s32
port 32 n
rlabel metal2 0 1650 30 1680 1 s33
port 33 n
rlabel metal2 0 1700 30 1730 1 s34
port 34 n
rlabel metal2 0 1750 30 1780 1 s35
port 35 n
rlabel metal2 0 1800 30 1830 1 s36
port 36 n
rlabel metal2 0 1850 30 1880 1 s37
port 37 n
rlabel metal2 0 1900 30 1930 1 s38
port 38 n
rlabel metal2 0 1950 30 1980 1 s39
port 39 n
rlabel metal2 0 2000 30 2030 1 s40
port 40 n
rlabel metal2 0 2050 30 2080 1 s41
port 41 n
rlabel metal2 0 2100 30 2130 1 s42
port 42 n
rlabel metal2 0 2150 30 2180 1 s43
port 43 n
rlabel metal2 0 2200 30 2230 1 s44
port 44 n
rlabel metal2 0 2250 30 2280 1 s45
port 45 n
rlabel metal2 0 2300 30 2330 1 s46
port 46 n
rlabel metal2 0 2350 30 2380 1 s47
port 47 n
rlabel metal2 0 2400 30 2430 1 s48
port 48 n
rlabel metal2 0 2450 30 2480 1 s49
port 49 n
rlabel metal2 0 2500 30 2530 1 s50
port 50 n
rlabel metal2 0 2550 30 2580 1 s51
port 51 n
rlabel metal2 0 2600 30 2630 1 s52
port 52 n
rlabel metal2 0 2650 30 2680 1 s53
port 53 n
rlabel metal2 0 2700 30 2730 1 s54
port 54 n
rlabel metal2 0 2750 30 2780 1 s55
port 55 n
rlabel metal2 0 2800 30 2830 1 s56
port 56 n
rlabel metal2 0 2850 30 2880 1 s57
port 57 n
rlabel metal2 0 2900 30 2930 1 s58
port 58 n
rlabel metal2 0 2950 30 2980 1 s59
port 59 n
rlabel metal2 0 3000 30 3030 1 s60
port 60 n
rlabel metal2 0 3050 30 3080 1 s61
port 61 n
rlabel metal2 0 3100 30 3130 1 s62
port 62 n
rlabel metal2 0 3150 30 3180 1 s63
port 63 n
<< end >>
