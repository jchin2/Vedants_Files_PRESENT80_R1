magic
tech sky130A
magscale 1 2
timestamp 1675786016
<< nwell >>
rect -2340 1470 -260 1660
rect -1710 1080 -890 1470
<< pwell >>
rect -2316 456 -284 896
rect -2326 304 -274 456
<< nmos >>
rect -2170 570 -2140 870
rect -2020 570 -1990 870
rect -1870 570 -1840 870
rect -1540 570 -1510 870
rect -1390 570 -1360 870
rect -1240 570 -1210 870
rect -1090 570 -1060 870
rect -760 570 -730 870
rect -610 570 -580 870
rect -460 570 -430 870
<< pmos >>
rect -1540 1130 -1510 1430
rect -1390 1130 -1360 1430
rect -1240 1130 -1210 1430
rect -1090 1130 -1060 1430
<< ndiff >>
rect -2290 797 -2170 870
rect -2290 763 -2247 797
rect -2213 763 -2170 797
rect -2290 717 -2170 763
rect -2290 683 -2247 717
rect -2213 683 -2170 717
rect -2290 637 -2170 683
rect -2290 603 -2247 637
rect -2213 603 -2170 637
rect -2290 570 -2170 603
rect -2140 570 -2020 870
rect -1990 570 -1870 870
rect -1840 797 -1720 870
rect -1840 763 -1797 797
rect -1763 763 -1720 797
rect -1840 717 -1720 763
rect -1840 683 -1797 717
rect -1763 683 -1720 717
rect -1840 637 -1720 683
rect -1840 603 -1797 637
rect -1763 603 -1720 637
rect -1840 570 -1720 603
rect -1660 797 -1540 870
rect -1660 763 -1617 797
rect -1583 763 -1540 797
rect -1660 717 -1540 763
rect -1660 683 -1617 717
rect -1583 683 -1540 717
rect -1660 637 -1540 683
rect -1660 603 -1617 637
rect -1583 603 -1540 637
rect -1660 570 -1540 603
rect -1510 797 -1390 870
rect -1510 763 -1467 797
rect -1433 763 -1390 797
rect -1510 717 -1390 763
rect -1510 683 -1467 717
rect -1433 683 -1390 717
rect -1510 637 -1390 683
rect -1510 603 -1467 637
rect -1433 603 -1390 637
rect -1510 570 -1390 603
rect -1360 797 -1240 870
rect -1360 763 -1317 797
rect -1283 763 -1240 797
rect -1360 717 -1240 763
rect -1360 683 -1317 717
rect -1283 683 -1240 717
rect -1360 637 -1240 683
rect -1360 603 -1317 637
rect -1283 603 -1240 637
rect -1360 570 -1240 603
rect -1210 797 -1090 870
rect -1210 763 -1167 797
rect -1133 763 -1090 797
rect -1210 717 -1090 763
rect -1210 683 -1167 717
rect -1133 683 -1090 717
rect -1210 637 -1090 683
rect -1210 603 -1167 637
rect -1133 603 -1090 637
rect -1210 570 -1090 603
rect -1060 797 -940 870
rect -1060 763 -1017 797
rect -983 763 -940 797
rect -1060 717 -940 763
rect -1060 683 -1017 717
rect -983 683 -940 717
rect -1060 637 -940 683
rect -1060 603 -1017 637
rect -983 603 -940 637
rect -1060 570 -940 603
rect -880 797 -760 870
rect -880 763 -837 797
rect -803 763 -760 797
rect -880 717 -760 763
rect -880 683 -837 717
rect -803 683 -760 717
rect -880 637 -760 683
rect -880 603 -837 637
rect -803 603 -760 637
rect -880 570 -760 603
rect -730 797 -610 870
rect -730 763 -687 797
rect -653 763 -610 797
rect -730 717 -610 763
rect -730 683 -687 717
rect -653 683 -610 717
rect -730 637 -610 683
rect -730 603 -687 637
rect -653 603 -610 637
rect -730 570 -610 603
rect -580 797 -460 870
rect -580 763 -537 797
rect -503 763 -460 797
rect -580 717 -460 763
rect -580 683 -537 717
rect -503 683 -460 717
rect -580 637 -460 683
rect -580 603 -537 637
rect -503 603 -460 637
rect -580 570 -460 603
rect -430 797 -310 870
rect -430 763 -387 797
rect -353 763 -310 797
rect -430 717 -310 763
rect -430 683 -387 717
rect -353 683 -310 717
rect -430 637 -310 683
rect -430 603 -387 637
rect -353 603 -310 637
rect -430 570 -310 603
<< pdiff >>
rect -1660 1357 -1540 1430
rect -1660 1323 -1617 1357
rect -1583 1323 -1540 1357
rect -1660 1277 -1540 1323
rect -1660 1243 -1617 1277
rect -1583 1243 -1540 1277
rect -1660 1197 -1540 1243
rect -1660 1163 -1617 1197
rect -1583 1163 -1540 1197
rect -1660 1130 -1540 1163
rect -1510 1357 -1390 1430
rect -1510 1323 -1467 1357
rect -1433 1323 -1390 1357
rect -1510 1277 -1390 1323
rect -1510 1243 -1467 1277
rect -1433 1243 -1390 1277
rect -1510 1197 -1390 1243
rect -1510 1163 -1467 1197
rect -1433 1163 -1390 1197
rect -1510 1130 -1390 1163
rect -1360 1357 -1240 1430
rect -1360 1323 -1317 1357
rect -1283 1323 -1240 1357
rect -1360 1277 -1240 1323
rect -1360 1243 -1317 1277
rect -1283 1243 -1240 1277
rect -1360 1197 -1240 1243
rect -1360 1163 -1317 1197
rect -1283 1163 -1240 1197
rect -1360 1130 -1240 1163
rect -1210 1357 -1090 1430
rect -1210 1323 -1167 1357
rect -1133 1323 -1090 1357
rect -1210 1277 -1090 1323
rect -1210 1243 -1167 1277
rect -1133 1243 -1090 1277
rect -1210 1197 -1090 1243
rect -1210 1163 -1167 1197
rect -1133 1163 -1090 1197
rect -1210 1130 -1090 1163
rect -1060 1357 -940 1430
rect -1060 1323 -1017 1357
rect -983 1323 -940 1357
rect -1060 1277 -940 1323
rect -1060 1243 -1017 1277
rect -983 1243 -940 1277
rect -1060 1197 -940 1243
rect -1060 1163 -1017 1197
rect -983 1163 -940 1197
rect -1060 1130 -940 1163
<< ndiffc >>
rect -2247 763 -2213 797
rect -2247 683 -2213 717
rect -2247 603 -2213 637
rect -1797 763 -1763 797
rect -1797 683 -1763 717
rect -1797 603 -1763 637
rect -1617 763 -1583 797
rect -1617 683 -1583 717
rect -1617 603 -1583 637
rect -1467 763 -1433 797
rect -1467 683 -1433 717
rect -1467 603 -1433 637
rect -1317 763 -1283 797
rect -1317 683 -1283 717
rect -1317 603 -1283 637
rect -1167 763 -1133 797
rect -1167 683 -1133 717
rect -1167 603 -1133 637
rect -1017 763 -983 797
rect -1017 683 -983 717
rect -1017 603 -983 637
rect -837 763 -803 797
rect -837 683 -803 717
rect -837 603 -803 637
rect -687 763 -653 797
rect -687 683 -653 717
rect -687 603 -653 637
rect -537 763 -503 797
rect -537 683 -503 717
rect -537 603 -503 637
rect -387 763 -353 797
rect -387 683 -353 717
rect -387 603 -353 637
<< pdiffc >>
rect -1617 1323 -1583 1357
rect -1617 1243 -1583 1277
rect -1617 1163 -1583 1197
rect -1467 1323 -1433 1357
rect -1467 1243 -1433 1277
rect -1467 1163 -1433 1197
rect -1317 1323 -1283 1357
rect -1317 1243 -1283 1277
rect -1317 1163 -1283 1197
rect -1167 1323 -1133 1357
rect -1167 1243 -1133 1277
rect -1167 1163 -1133 1197
rect -1017 1323 -983 1357
rect -1017 1243 -983 1277
rect -1017 1163 -983 1197
<< psubdiff >>
rect -2300 397 -300 430
rect -2300 363 -2277 397
rect -2243 363 -2197 397
rect -2163 363 -2117 397
rect -2083 363 -2037 397
rect -2003 363 -1957 397
rect -1923 363 -1877 397
rect -1843 363 -1797 397
rect -1763 363 -1717 397
rect -1683 363 -1637 397
rect -1603 363 -1557 397
rect -1523 363 -1477 397
rect -1443 363 -1397 397
rect -1363 363 -1317 397
rect -1283 363 -1237 397
rect -1203 363 -1157 397
rect -1123 363 -1077 397
rect -1043 363 -997 397
rect -963 363 -917 397
rect -883 363 -837 397
rect -803 363 -757 397
rect -723 363 -677 397
rect -643 363 -597 397
rect -563 363 -517 397
rect -483 363 -437 397
rect -403 363 -357 397
rect -323 363 -300 397
rect -2300 330 -300 363
<< nsubdiff >>
rect -2300 1577 -300 1610
rect -2300 1543 -2277 1577
rect -2243 1543 -2197 1577
rect -2163 1543 -2117 1577
rect -2083 1543 -2037 1577
rect -2003 1543 -1957 1577
rect -1923 1543 -1877 1577
rect -1843 1543 -1797 1577
rect -1763 1543 -1717 1577
rect -1683 1543 -1637 1577
rect -1603 1543 -1557 1577
rect -1523 1543 -1477 1577
rect -1443 1543 -1397 1577
rect -1363 1543 -1317 1577
rect -1283 1543 -1237 1577
rect -1203 1543 -1157 1577
rect -1123 1543 -1077 1577
rect -1043 1543 -997 1577
rect -963 1543 -917 1577
rect -883 1543 -837 1577
rect -803 1543 -757 1577
rect -723 1543 -677 1577
rect -643 1543 -597 1577
rect -563 1543 -517 1577
rect -483 1543 -437 1577
rect -403 1543 -357 1577
rect -323 1543 -300 1577
rect -2300 1510 -300 1543
<< psubdiffcont >>
rect -2277 363 -2243 397
rect -2197 363 -2163 397
rect -2117 363 -2083 397
rect -2037 363 -2003 397
rect -1957 363 -1923 397
rect -1877 363 -1843 397
rect -1797 363 -1763 397
rect -1717 363 -1683 397
rect -1637 363 -1603 397
rect -1557 363 -1523 397
rect -1477 363 -1443 397
rect -1397 363 -1363 397
rect -1317 363 -1283 397
rect -1237 363 -1203 397
rect -1157 363 -1123 397
rect -1077 363 -1043 397
rect -997 363 -963 397
rect -917 363 -883 397
rect -837 363 -803 397
rect -757 363 -723 397
rect -677 363 -643 397
rect -597 363 -563 397
rect -517 363 -483 397
rect -437 363 -403 397
rect -357 363 -323 397
<< nsubdiffcont >>
rect -2277 1543 -2243 1577
rect -2197 1543 -2163 1577
rect -2117 1543 -2083 1577
rect -2037 1543 -2003 1577
rect -1957 1543 -1923 1577
rect -1877 1543 -1843 1577
rect -1797 1543 -1763 1577
rect -1717 1543 -1683 1577
rect -1637 1543 -1603 1577
rect -1557 1543 -1523 1577
rect -1477 1543 -1443 1577
rect -1397 1543 -1363 1577
rect -1317 1543 -1283 1577
rect -1237 1543 -1203 1577
rect -1157 1543 -1123 1577
rect -1077 1543 -1043 1577
rect -997 1543 -963 1577
rect -917 1543 -883 1577
rect -837 1543 -803 1577
rect -757 1543 -723 1577
rect -677 1543 -643 1577
rect -597 1543 -563 1577
rect -517 1543 -483 1577
rect -437 1543 -403 1577
rect -357 1543 -323 1577
<< poly >>
rect -1540 1460 -1360 1490
rect -1540 1430 -1510 1460
rect -1390 1430 -1360 1460
rect -1240 1460 -1060 1490
rect -1240 1430 -1210 1460
rect -1090 1430 -1060 1460
rect -510 1452 -430 1475
rect -2210 1127 -2130 1150
rect -510 1418 -487 1452
rect -453 1418 -430 1452
rect -510 1395 -430 1418
rect -610 1327 -530 1350
rect -610 1293 -587 1327
rect -553 1293 -530 1327
rect -610 1270 -530 1293
rect -810 1237 -730 1260
rect -810 1203 -787 1237
rect -753 1203 -730 1237
rect -810 1180 -730 1203
rect -2210 1093 -2187 1127
rect -2153 1093 -2130 1127
rect -1540 1100 -1510 1130
rect -2210 1070 -2130 1093
rect -2170 870 -2140 1070
rect -2070 1027 -1990 1050
rect -2070 993 -2047 1027
rect -2013 993 -1990 1027
rect -2070 970 -1990 993
rect -1390 975 -1360 1130
rect -1240 1100 -1210 1130
rect -1090 1100 -1060 1130
rect -1290 1077 -1210 1100
rect -1290 1043 -1267 1077
rect -1233 1043 -1210 1077
rect -1290 1020 -1210 1043
rect -2020 870 -1990 970
rect -1920 947 -1840 970
rect -1920 913 -1897 947
rect -1863 913 -1840 947
rect -1920 890 -1840 913
rect -1390 952 -1310 975
rect -1390 918 -1367 952
rect -1333 918 -1310 952
rect -1870 870 -1840 890
rect -1540 870 -1510 900
rect -1390 895 -1310 918
rect -1390 870 -1360 895
rect -1240 870 -1210 1020
rect -1090 870 -1060 900
rect -760 870 -730 1180
rect -610 870 -580 1270
rect -460 870 -430 1395
rect -2170 540 -2140 570
rect -2020 540 -1990 570
rect -1870 540 -1840 570
rect -1540 540 -1510 570
rect -1390 540 -1360 570
rect -1240 540 -1210 570
rect -1090 540 -1060 570
rect -760 540 -730 570
rect -610 540 -580 570
rect -460 540 -430 570
rect -1540 517 -1460 540
rect -1540 483 -1517 517
rect -1483 483 -1460 517
rect -1540 460 -1460 483
rect -1140 517 -1060 540
rect -1140 483 -1117 517
rect -1083 483 -1060 517
rect -1140 460 -1060 483
<< polycont >>
rect -487 1418 -453 1452
rect -587 1293 -553 1327
rect -787 1203 -753 1237
rect -2187 1093 -2153 1127
rect -2047 993 -2013 1027
rect -1267 1043 -1233 1077
rect -1897 913 -1863 947
rect -1367 918 -1333 952
rect -1517 483 -1483 517
rect -1117 483 -1083 517
<< locali >>
rect -2300 1577 -300 1600
rect -2300 1543 -2277 1577
rect -2243 1543 -2197 1577
rect -2163 1543 -2117 1577
rect -2083 1543 -2037 1577
rect -2003 1543 -1957 1577
rect -1923 1543 -1877 1577
rect -1843 1543 -1797 1577
rect -1763 1543 -1717 1577
rect -1683 1543 -1637 1577
rect -1603 1543 -1557 1577
rect -1523 1543 -1477 1577
rect -1443 1543 -1397 1577
rect -1363 1543 -1317 1577
rect -1283 1543 -1237 1577
rect -1203 1543 -1157 1577
rect -1123 1543 -1077 1577
rect -1043 1543 -997 1577
rect -963 1543 -917 1577
rect -883 1543 -837 1577
rect -803 1543 -757 1577
rect -723 1543 -677 1577
rect -643 1543 -597 1577
rect -563 1543 -517 1577
rect -483 1543 -437 1577
rect -403 1543 -357 1577
rect -323 1543 -300 1577
rect -2300 1520 -300 1543
rect -1790 1450 -1710 1470
rect -2290 1447 -1710 1450
rect -2290 1413 -1767 1447
rect -1733 1413 -1710 1447
rect -2290 1410 -1710 1413
rect -1790 1390 -1710 1410
rect -510 1452 -430 1475
rect -510 1418 -487 1452
rect -453 1418 -430 1452
rect -510 1395 -430 1418
rect -1910 1340 -1830 1360
rect -2290 1337 -1830 1340
rect -2290 1303 -1887 1337
rect -1853 1303 -1830 1337
rect -2290 1300 -1830 1303
rect -1910 1280 -1830 1300
rect -1640 1357 -1560 1390
rect -1640 1323 -1617 1357
rect -1583 1323 -1560 1357
rect -1640 1277 -1560 1323
rect -1790 1240 -1710 1260
rect -2290 1237 -1710 1240
rect -2290 1203 -1767 1237
rect -1733 1203 -1710 1237
rect -2290 1200 -1710 1203
rect -1790 1180 -1710 1200
rect -1640 1243 -1617 1277
rect -1583 1243 -1560 1277
rect -1640 1197 -1560 1243
rect -1640 1163 -1617 1197
rect -1583 1163 -1560 1197
rect -2290 1127 -2130 1150
rect -1640 1140 -1560 1163
rect -1490 1357 -1410 1390
rect -1490 1323 -1467 1357
rect -1433 1323 -1410 1357
rect -1490 1277 -1410 1323
rect -1490 1243 -1467 1277
rect -1433 1243 -1410 1277
rect -1490 1197 -1410 1243
rect -1490 1163 -1467 1197
rect -1433 1163 -1410 1197
rect -1490 1130 -1410 1163
rect -1340 1357 -1260 1390
rect -1340 1323 -1317 1357
rect -1283 1323 -1260 1357
rect -1340 1277 -1260 1323
rect -1340 1243 -1317 1277
rect -1283 1243 -1260 1277
rect -1340 1197 -1260 1243
rect -1340 1163 -1317 1197
rect -1283 1163 -1260 1197
rect -1340 1140 -1260 1163
rect -1190 1357 -1110 1390
rect -1190 1323 -1167 1357
rect -1133 1323 -1110 1357
rect -1190 1277 -1110 1323
rect -1190 1243 -1167 1277
rect -1133 1243 -1110 1277
rect -1190 1197 -1110 1243
rect -1190 1163 -1167 1197
rect -1133 1163 -1110 1197
rect -1190 1130 -1110 1163
rect -1040 1357 -960 1390
rect -1040 1323 -1017 1357
rect -983 1323 -960 1357
rect -1040 1277 -960 1323
rect -1040 1243 -1017 1277
rect -983 1243 -960 1277
rect -610 1327 -530 1350
rect -610 1293 -587 1327
rect -553 1293 -530 1327
rect -610 1270 -530 1293
rect -1040 1197 -960 1243
rect -1040 1163 -1017 1197
rect -983 1163 -960 1197
rect -810 1237 -730 1260
rect -810 1203 -787 1237
rect -753 1203 -730 1237
rect -810 1180 -730 1203
rect -1040 1140 -960 1163
rect -2290 1110 -2187 1127
rect -2210 1093 -2187 1110
rect -2153 1093 -2130 1127
rect -2210 1070 -2130 1093
rect -1470 1080 -1430 1130
rect -1290 1080 -1210 1100
rect -1470 1077 -1210 1080
rect -2070 1030 -1990 1050
rect -2290 1027 -1990 1030
rect -2290 993 -2047 1027
rect -2013 993 -1990 1027
rect -2290 990 -1990 993
rect -2070 970 -1990 990
rect -1470 1043 -1267 1077
rect -1233 1043 -1210 1077
rect -1470 1040 -1210 1043
rect -1920 947 -1840 970
rect -1920 930 -1897 947
rect -2290 913 -1897 930
rect -1863 913 -1840 947
rect -2290 890 -1840 913
rect -1470 910 -1430 1040
rect -1290 1020 -1210 1040
rect -1780 870 -1430 910
rect -1390 960 -1310 975
rect -1170 960 -1130 1130
rect -890 1080 -810 1100
rect -890 1077 -310 1080
rect -890 1043 -867 1077
rect -833 1043 -310 1077
rect -890 1040 -310 1043
rect -890 1020 -810 1040
rect -1390 952 -310 960
rect -1390 918 -1367 952
rect -1333 920 -310 952
rect -1333 918 -1310 920
rect -1390 895 -1310 918
rect -1780 830 -1740 870
rect -1470 830 -1430 870
rect -1170 830 -1130 920
rect -840 830 -800 920
rect -540 830 -500 920
rect -2270 797 -2190 830
rect -2270 763 -2247 797
rect -2213 763 -2190 797
rect -2270 717 -2190 763
rect -2270 683 -2247 717
rect -2213 683 -2190 717
rect -2270 637 -2190 683
rect -2270 603 -2247 637
rect -2213 603 -2190 637
rect -2270 580 -2190 603
rect -1820 797 -1740 830
rect -1820 763 -1797 797
rect -1763 763 -1740 797
rect -1820 717 -1740 763
rect -1820 683 -1797 717
rect -1763 683 -1740 717
rect -1820 637 -1740 683
rect -1820 603 -1797 637
rect -1763 603 -1740 637
rect -1820 580 -1740 603
rect -1640 797 -1560 830
rect -1640 763 -1617 797
rect -1583 763 -1560 797
rect -1640 717 -1560 763
rect -1640 683 -1617 717
rect -1583 683 -1560 717
rect -1640 637 -1560 683
rect -1640 603 -1617 637
rect -1583 603 -1560 637
rect -1640 580 -1560 603
rect -1490 797 -1410 830
rect -1490 763 -1467 797
rect -1433 763 -1410 797
rect -1490 717 -1410 763
rect -1490 683 -1467 717
rect -1433 683 -1410 717
rect -1490 637 -1410 683
rect -1490 603 -1467 637
rect -1433 603 -1410 637
rect -1490 580 -1410 603
rect -1340 797 -1260 830
rect -1340 763 -1317 797
rect -1283 763 -1260 797
rect -1340 717 -1260 763
rect -1340 683 -1317 717
rect -1283 683 -1260 717
rect -1340 637 -1260 683
rect -1340 603 -1317 637
rect -1283 603 -1260 637
rect -1340 580 -1260 603
rect -1190 797 -1110 830
rect -1190 763 -1167 797
rect -1133 763 -1110 797
rect -1190 717 -1110 763
rect -1190 683 -1167 717
rect -1133 683 -1110 717
rect -1190 637 -1110 683
rect -1190 603 -1167 637
rect -1133 603 -1110 637
rect -1190 580 -1110 603
rect -1040 797 -960 830
rect -1040 763 -1017 797
rect -983 763 -960 797
rect -1040 717 -960 763
rect -1040 683 -1017 717
rect -983 683 -960 717
rect -1040 637 -960 683
rect -1040 603 -1017 637
rect -983 603 -960 637
rect -1040 580 -960 603
rect -860 797 -780 830
rect -860 763 -837 797
rect -803 763 -780 797
rect -860 717 -780 763
rect -860 683 -837 717
rect -803 683 -780 717
rect -860 637 -780 683
rect -860 603 -837 637
rect -803 603 -780 637
rect -860 580 -780 603
rect -710 797 -630 830
rect -710 763 -687 797
rect -653 763 -630 797
rect -710 717 -630 763
rect -710 683 -687 717
rect -653 683 -630 717
rect -710 637 -630 683
rect -710 603 -687 637
rect -653 603 -630 637
rect -710 580 -630 603
rect -560 797 -480 830
rect -560 763 -537 797
rect -503 763 -480 797
rect -560 717 -480 763
rect -560 683 -537 717
rect -503 683 -480 717
rect -560 637 -480 683
rect -560 603 -537 637
rect -503 603 -480 637
rect -560 580 -480 603
rect -410 797 -330 830
rect -410 763 -387 797
rect -353 763 -330 797
rect -410 717 -330 763
rect -410 683 -387 717
rect -353 683 -330 717
rect -410 637 -330 683
rect -410 603 -387 637
rect -353 603 -330 637
rect -410 580 -330 603
rect -1540 520 -1460 540
rect -1140 520 -1060 540
rect -2290 517 -1060 520
rect -2290 483 -1517 517
rect -1483 483 -1117 517
rect -1083 483 -1060 517
rect -2290 480 -1060 483
rect -1540 460 -1460 480
rect -1140 460 -1060 480
rect -2300 397 -300 420
rect -2300 363 -2277 397
rect -2243 363 -2197 397
rect -2163 363 -2117 397
rect -2083 363 -2037 397
rect -2003 363 -1957 397
rect -1923 363 -1877 397
rect -1843 363 -1797 397
rect -1763 363 -1717 397
rect -1683 363 -1637 397
rect -1603 363 -1557 397
rect -1523 363 -1477 397
rect -1443 363 -1397 397
rect -1363 363 -1317 397
rect -1283 363 -1237 397
rect -1203 363 -1157 397
rect -1123 363 -1077 397
rect -1043 363 -997 397
rect -963 363 -917 397
rect -883 363 -837 397
rect -803 363 -757 397
rect -723 363 -677 397
rect -643 363 -597 397
rect -563 363 -517 397
rect -483 363 -437 397
rect -403 363 -357 397
rect -323 363 -300 397
rect -2300 340 -300 363
<< viali >>
rect -2277 1543 -2243 1577
rect -2197 1543 -2163 1577
rect -2117 1543 -2083 1577
rect -2037 1543 -2003 1577
rect -1957 1543 -1923 1577
rect -1877 1543 -1843 1577
rect -1797 1543 -1763 1577
rect -1717 1543 -1683 1577
rect -1637 1543 -1603 1577
rect -1557 1543 -1523 1577
rect -1477 1543 -1443 1577
rect -1397 1543 -1363 1577
rect -1317 1543 -1283 1577
rect -1237 1543 -1203 1577
rect -1157 1543 -1123 1577
rect -1077 1543 -1043 1577
rect -997 1543 -963 1577
rect -917 1543 -883 1577
rect -837 1543 -803 1577
rect -757 1543 -723 1577
rect -677 1543 -643 1577
rect -597 1543 -563 1577
rect -517 1543 -483 1577
rect -437 1543 -403 1577
rect -357 1543 -323 1577
rect -1767 1413 -1733 1447
rect -487 1418 -453 1452
rect -1887 1303 -1853 1337
rect -1617 1323 -1583 1357
rect -1767 1203 -1733 1237
rect -1617 1243 -1583 1277
rect -1617 1163 -1583 1197
rect -1317 1323 -1283 1357
rect -1317 1243 -1283 1277
rect -1317 1163 -1283 1197
rect -1017 1323 -983 1357
rect -1017 1243 -983 1277
rect -587 1293 -553 1327
rect -1017 1163 -983 1197
rect -787 1203 -753 1237
rect -1267 1043 -1233 1077
rect -867 1043 -833 1077
rect -2247 763 -2213 797
rect -2247 683 -2213 717
rect -2247 603 -2213 637
rect -1617 763 -1583 797
rect -1617 683 -1583 717
rect -1617 603 -1583 637
rect -1317 763 -1283 797
rect -1317 683 -1283 717
rect -1317 603 -1283 637
rect -1017 763 -983 797
rect -1017 683 -983 717
rect -1017 603 -983 637
rect -687 763 -653 797
rect -687 683 -653 717
rect -687 603 -653 637
rect -387 763 -353 797
rect -387 683 -353 717
rect -387 603 -353 637
rect -2277 363 -2243 397
rect -2197 363 -2163 397
rect -2117 363 -2083 397
rect -2037 363 -2003 397
rect -1957 363 -1923 397
rect -1877 363 -1843 397
rect -1797 363 -1763 397
rect -1717 363 -1683 397
rect -1637 363 -1603 397
rect -1557 363 -1523 397
rect -1477 363 -1443 397
rect -1397 363 -1363 397
rect -1317 363 -1283 397
rect -1237 363 -1203 397
rect -1157 363 -1123 397
rect -1077 363 -1043 397
rect -997 363 -963 397
rect -917 363 -883 397
rect -837 363 -803 397
rect -757 363 -723 397
rect -677 363 -643 397
rect -597 363 -563 397
rect -517 363 -483 397
rect -437 363 -403 397
rect -357 363 -323 397
<< metal1 >>
rect -2300 1577 -300 1610
rect -2300 1543 -2277 1577
rect -2243 1543 -2197 1577
rect -2163 1543 -2117 1577
rect -2083 1543 -2037 1577
rect -2003 1543 -1957 1577
rect -1923 1543 -1877 1577
rect -1843 1543 -1797 1577
rect -1763 1543 -1717 1577
rect -1683 1543 -1637 1577
rect -1603 1543 -1557 1577
rect -1523 1543 -1477 1577
rect -1443 1543 -1397 1577
rect -1363 1543 -1317 1577
rect -1283 1543 -1237 1577
rect -1203 1543 -1157 1577
rect -1123 1543 -1077 1577
rect -1043 1543 -997 1577
rect -963 1543 -917 1577
rect -883 1543 -837 1577
rect -803 1543 -757 1577
rect -723 1543 -677 1577
rect -643 1543 -597 1577
rect -563 1543 -517 1577
rect -483 1543 -437 1577
rect -403 1543 -357 1577
rect -323 1543 -300 1577
rect -2300 1510 -300 1543
rect -2250 830 -2210 1510
rect -1790 1456 -1710 1470
rect -1790 1404 -1776 1456
rect -1724 1404 -1710 1456
rect -1790 1390 -1710 1404
rect -1910 1346 -1830 1360
rect -1910 1294 -1896 1346
rect -1844 1294 -1830 1346
rect -1910 1280 -1830 1294
rect -1640 1357 -1560 1510
rect -1640 1323 -1617 1357
rect -1583 1323 -1560 1357
rect -1640 1277 -1560 1323
rect -1790 1246 -1710 1260
rect -1790 1194 -1776 1246
rect -1724 1194 -1710 1246
rect -1790 1180 -1710 1194
rect -1640 1243 -1617 1277
rect -1583 1243 -1560 1277
rect -1640 1197 -1560 1243
rect -1640 1163 -1617 1197
rect -1583 1163 -1560 1197
rect -1640 1140 -1560 1163
rect -1340 1357 -1260 1510
rect -1340 1323 -1317 1357
rect -1283 1323 -1260 1357
rect -1340 1277 -1260 1323
rect -1340 1243 -1317 1277
rect -1283 1243 -1260 1277
rect -1340 1197 -1260 1243
rect -1340 1163 -1317 1197
rect -1283 1163 -1260 1197
rect -1340 1140 -1260 1163
rect -1040 1357 -960 1510
rect -1040 1323 -1017 1357
rect -983 1323 -960 1357
rect -1040 1277 -960 1323
rect -1040 1243 -1017 1277
rect -983 1243 -960 1277
rect -1040 1197 -960 1243
rect -1040 1163 -1017 1197
rect -983 1163 -960 1197
rect -810 1246 -730 1260
rect -810 1194 -796 1246
rect -744 1194 -730 1246
rect -810 1180 -730 1194
rect -1040 1140 -960 1163
rect -1290 1080 -1210 1100
rect -890 1080 -810 1100
rect -1290 1077 -810 1080
rect -1290 1043 -1267 1077
rect -1233 1043 -867 1077
rect -833 1043 -810 1077
rect -1290 1040 -810 1043
rect -1290 1020 -1210 1040
rect -890 1020 -810 1040
rect -690 830 -650 1510
rect -510 1461 -430 1475
rect -510 1409 -496 1461
rect -444 1409 -430 1461
rect -510 1395 -430 1409
rect -610 1336 -530 1350
rect -610 1284 -596 1336
rect -544 1284 -530 1336
rect -610 1270 -530 1284
rect -390 830 -350 1510
rect -2270 797 -2190 830
rect -2270 763 -2247 797
rect -2213 763 -2190 797
rect -2270 717 -2190 763
rect -2270 683 -2247 717
rect -2213 683 -2190 717
rect -2270 637 -2190 683
rect -2270 603 -2247 637
rect -2213 603 -2190 637
rect -2270 580 -2190 603
rect -1640 797 -1560 830
rect -1640 763 -1617 797
rect -1583 763 -1560 797
rect -1640 717 -1560 763
rect -1640 683 -1617 717
rect -1583 683 -1560 717
rect -1640 637 -1560 683
rect -1640 603 -1617 637
rect -1583 603 -1560 637
rect -1640 580 -1560 603
rect -1340 797 -1260 830
rect -1340 763 -1317 797
rect -1283 763 -1260 797
rect -1340 717 -1260 763
rect -1340 683 -1317 717
rect -1283 683 -1260 717
rect -1340 637 -1260 683
rect -1340 603 -1317 637
rect -1283 603 -1260 637
rect -1340 580 -1260 603
rect -1040 797 -960 830
rect -1040 763 -1017 797
rect -983 763 -960 797
rect -1040 717 -960 763
rect -1040 683 -1017 717
rect -983 683 -960 717
rect -1040 637 -960 683
rect -1040 603 -1017 637
rect -983 603 -960 637
rect -1040 580 -960 603
rect -710 797 -630 830
rect -710 763 -687 797
rect -653 763 -630 797
rect -710 717 -630 763
rect -710 683 -687 717
rect -653 683 -630 717
rect -710 637 -630 683
rect -710 603 -687 637
rect -653 603 -630 637
rect -710 580 -630 603
rect -410 797 -330 830
rect -410 763 -387 797
rect -353 763 -330 797
rect -410 717 -330 763
rect -410 683 -387 717
rect -353 683 -330 717
rect -410 637 -330 683
rect -410 603 -387 637
rect -353 603 -330 637
rect -410 580 -330 603
rect -1620 430 -1580 580
rect -1320 430 -1280 580
rect -1020 430 -980 580
rect -2300 397 -300 430
rect -2300 363 -2277 397
rect -2243 363 -2197 397
rect -2163 363 -2117 397
rect -2083 363 -2037 397
rect -2003 363 -1957 397
rect -1923 363 -1877 397
rect -1843 363 -1797 397
rect -1763 363 -1717 397
rect -1683 363 -1637 397
rect -1603 363 -1557 397
rect -1523 363 -1477 397
rect -1443 363 -1397 397
rect -1363 363 -1317 397
rect -1283 363 -1237 397
rect -1203 363 -1157 397
rect -1123 363 -1077 397
rect -1043 363 -997 397
rect -963 363 -917 397
rect -883 363 -837 397
rect -803 363 -757 397
rect -723 363 -677 397
rect -643 363 -597 397
rect -563 363 -517 397
rect -483 363 -437 397
rect -403 363 -357 397
rect -323 363 -300 397
rect -2300 330 -300 363
<< via1 >>
rect -1776 1447 -1724 1456
rect -1776 1413 -1767 1447
rect -1767 1413 -1733 1447
rect -1733 1413 -1724 1447
rect -1776 1404 -1724 1413
rect -1896 1337 -1844 1346
rect -1896 1303 -1887 1337
rect -1887 1303 -1853 1337
rect -1853 1303 -1844 1337
rect -1896 1294 -1844 1303
rect -1776 1237 -1724 1246
rect -1776 1203 -1767 1237
rect -1767 1203 -1733 1237
rect -1733 1203 -1724 1237
rect -1776 1194 -1724 1203
rect -796 1237 -744 1246
rect -796 1203 -787 1237
rect -787 1203 -753 1237
rect -753 1203 -744 1237
rect -796 1194 -744 1203
rect -496 1452 -444 1461
rect -496 1418 -487 1452
rect -487 1418 -453 1452
rect -453 1418 -444 1452
rect -496 1409 -444 1418
rect -596 1327 -544 1336
rect -596 1293 -587 1327
rect -587 1293 -553 1327
rect -553 1293 -544 1327
rect -596 1284 -544 1293
<< metal2 >>
rect -1790 1456 -1710 1470
rect -1790 1404 -1776 1456
rect -1724 1450 -1710 1456
rect -510 1461 -430 1475
rect -510 1450 -496 1461
rect -1724 1410 -496 1450
rect -1724 1404 -1710 1410
rect -1790 1390 -1710 1404
rect -510 1409 -496 1410
rect -444 1409 -430 1461
rect -510 1395 -430 1409
rect -1910 1346 -1830 1360
rect -1910 1294 -1896 1346
rect -1844 1340 -1830 1346
rect -610 1340 -530 1350
rect -1844 1336 -530 1340
rect -1844 1300 -596 1336
rect -1844 1294 -1830 1300
rect -1910 1280 -1830 1294
rect -610 1284 -596 1300
rect -544 1284 -530 1336
rect -610 1270 -530 1284
rect -1790 1246 -1710 1260
rect -1790 1194 -1776 1246
rect -1724 1240 -1710 1246
rect -810 1246 -730 1260
rect -810 1240 -796 1246
rect -1724 1200 -796 1240
rect -1724 1194 -1710 1200
rect -1790 1180 -1710 1194
rect -810 1194 -796 1200
rect -744 1194 -730 1246
rect -810 1180 -730 1194
<< labels >>
rlabel metal1 s -1270 1040 -1230 1080 4 OUT_bar
port 1 nsew
rlabel metal1 s -1320 360 -1280 400 4 GND!
port 2 nsew
rlabel metal1 s -1320 1540 -1280 1580 4 CLK
port 3 nsew
rlabel locali s -1370 915 -1330 955 4 OUT
port 4 nsew
rlabel locali s -2280 1420 -2260 1440 4 A
port 5 nsew
rlabel locali s -2280 1120 -2260 1140 4 A_bar
port 6 nsew
rlabel locali s -2280 1310 -2260 1330 4 B
port 7 nsew
rlabel locali s -2280 1000 -2260 1020 4 B_bar
port 8 nsew
rlabel locali s -2280 1210 -2260 1230 4 C
port 9 nsew
rlabel locali s -2280 900 -2260 920 4 C_bar
port 10 nsew
rlabel locali s -1520 480 -1480 520 4 Dis
port 11 nsew
<< end >>
