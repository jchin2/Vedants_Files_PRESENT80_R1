magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -568 -20 -183 550
<< l67d20 >>
rect -460 520 -290 540
rect -460 500 -440 520
rect -310 500 -290 520
rect -545 20 -505 500
rect -470 20 -430 500
rect -395 20 -355 500
rect -320 20 -280 500
rect -245 20 -205 500
rect -535 0 -515 20
rect -385 0 -365 20
rect -235 0 -215 20
rect -535 -20 -215 0
<< l66d20 >>
rect -495 535 -255 550
rect -495 -5 -480 535
rect -420 -5 -405 535
rect -345 -5 -330 535
rect -270 -5 -255 535
<< l66d44 >>
rect -534 464 -517 481
rect -459 464 -442 481
rect -384 464 -367 481
rect -309 464 -292 481
rect -234 464 -217 481
rect -534 414 -517 431
rect -459 409 -442 426
rect -384 414 -367 431
rect -309 414 -292 431
rect -234 414 -217 431
rect -534 380 -517 397
rect -459 375 -442 392
rect -384 380 -367 397
rect -309 380 -292 397
rect -234 380 -217 397
rect -534 346 -517 363
rect -459 341 -442 358
rect -384 346 -367 363
rect -309 346 -292 363
rect -234 346 -217 363
rect -534 312 -517 329
rect -459 307 -442 324
rect -384 312 -367 329
rect -309 312 -292 329
rect -234 312 -217 329
rect -534 278 -517 295
rect -459 273 -442 290
rect -384 278 -367 295
rect -309 278 -292 295
rect -234 278 -217 295
rect -534 244 -517 261
rect -459 239 -442 256
rect -384 244 -367 261
rect -309 244 -292 261
rect -234 244 -217 261
rect -534 210 -517 227
rect -459 205 -442 222
rect -384 210 -367 227
rect -309 210 -292 227
rect -234 210 -217 227
rect -534 176 -517 193
rect -459 171 -442 188
rect -384 176 -367 193
rect -309 176 -292 193
rect -234 176 -217 193
rect -534 142 -517 159
rect -459 137 -442 154
rect -384 142 -367 159
rect -309 142 -292 159
rect -234 142 -217 159
rect -534 108 -517 125
rect -459 103 -442 120
rect -384 108 -367 125
rect -309 108 -292 125
rect -234 108 -217 125
rect -534 74 -517 91
rect -459 69 -442 86
rect -384 74 -367 91
rect -309 74 -292 91
rect -234 74 -217 91
rect -534 40 -517 57
rect -459 35 -442 52
rect -384 40 -367 57
rect -309 40 -292 57
rect -234 40 -217 57
<< l65d20 >>
rect -555 10 -195 510
<< l93d44 >>
rect -568 -3 -183 523
<< l125d44 >>
rect -513 -8 -237 528
<< end >>
