magic
tech sky130A
magscale 1 2
timestamp 1671041739
<< pwell >>
rect -2136 -6 -964 996
<< nmoslvt >>
rect -1870 20 -1770 970
rect -1650 20 -1550 970
rect -1430 20 -1330 970
rect -1210 20 -1110 970
<< ndiff >>
rect -1990 920 -1870 970
rect -1990 886 -1947 920
rect -1913 886 -1870 920
rect -1990 852 -1870 886
rect -1990 818 -1947 852
rect -1913 818 -1870 852
rect -1990 784 -1870 818
rect -1990 750 -1947 784
rect -1913 750 -1870 784
rect -1990 716 -1870 750
rect -1990 682 -1947 716
rect -1913 682 -1870 716
rect -1990 648 -1870 682
rect -1990 614 -1947 648
rect -1913 614 -1870 648
rect -1990 580 -1870 614
rect -1990 546 -1947 580
rect -1913 546 -1870 580
rect -1990 512 -1870 546
rect -1990 478 -1947 512
rect -1913 478 -1870 512
rect -1990 444 -1870 478
rect -1990 410 -1947 444
rect -1913 410 -1870 444
rect -1990 376 -1870 410
rect -1990 342 -1947 376
rect -1913 342 -1870 376
rect -1990 308 -1870 342
rect -1990 274 -1947 308
rect -1913 274 -1870 308
rect -1990 240 -1870 274
rect -1990 206 -1947 240
rect -1913 206 -1870 240
rect -1990 172 -1870 206
rect -1990 138 -1947 172
rect -1913 138 -1870 172
rect -1990 104 -1870 138
rect -1990 70 -1947 104
rect -1913 70 -1870 104
rect -1990 20 -1870 70
rect -1770 920 -1650 970
rect -1770 886 -1727 920
rect -1693 886 -1650 920
rect -1770 852 -1650 886
rect -1770 818 -1727 852
rect -1693 818 -1650 852
rect -1770 784 -1650 818
rect -1770 750 -1727 784
rect -1693 750 -1650 784
rect -1770 716 -1650 750
rect -1770 682 -1727 716
rect -1693 682 -1650 716
rect -1770 648 -1650 682
rect -1770 614 -1727 648
rect -1693 614 -1650 648
rect -1770 580 -1650 614
rect -1770 546 -1727 580
rect -1693 546 -1650 580
rect -1770 512 -1650 546
rect -1770 478 -1727 512
rect -1693 478 -1650 512
rect -1770 444 -1650 478
rect -1770 410 -1727 444
rect -1693 410 -1650 444
rect -1770 376 -1650 410
rect -1770 342 -1727 376
rect -1693 342 -1650 376
rect -1770 308 -1650 342
rect -1770 274 -1727 308
rect -1693 274 -1650 308
rect -1770 240 -1650 274
rect -1770 206 -1727 240
rect -1693 206 -1650 240
rect -1770 172 -1650 206
rect -1770 138 -1727 172
rect -1693 138 -1650 172
rect -1770 104 -1650 138
rect -1770 70 -1727 104
rect -1693 70 -1650 104
rect -1770 20 -1650 70
rect -1550 920 -1430 970
rect -1550 886 -1507 920
rect -1473 886 -1430 920
rect -1550 852 -1430 886
rect -1550 818 -1507 852
rect -1473 818 -1430 852
rect -1550 784 -1430 818
rect -1550 750 -1507 784
rect -1473 750 -1430 784
rect -1550 716 -1430 750
rect -1550 682 -1507 716
rect -1473 682 -1430 716
rect -1550 648 -1430 682
rect -1550 614 -1507 648
rect -1473 614 -1430 648
rect -1550 580 -1430 614
rect -1550 546 -1507 580
rect -1473 546 -1430 580
rect -1550 512 -1430 546
rect -1550 478 -1507 512
rect -1473 478 -1430 512
rect -1550 444 -1430 478
rect -1550 410 -1507 444
rect -1473 410 -1430 444
rect -1550 376 -1430 410
rect -1550 342 -1507 376
rect -1473 342 -1430 376
rect -1550 308 -1430 342
rect -1550 274 -1507 308
rect -1473 274 -1430 308
rect -1550 240 -1430 274
rect -1550 206 -1507 240
rect -1473 206 -1430 240
rect -1550 172 -1430 206
rect -1550 138 -1507 172
rect -1473 138 -1430 172
rect -1550 104 -1430 138
rect -1550 70 -1507 104
rect -1473 70 -1430 104
rect -1550 20 -1430 70
rect -1330 920 -1210 970
rect -1330 886 -1287 920
rect -1253 886 -1210 920
rect -1330 852 -1210 886
rect -1330 818 -1287 852
rect -1253 818 -1210 852
rect -1330 784 -1210 818
rect -1330 750 -1287 784
rect -1253 750 -1210 784
rect -1330 716 -1210 750
rect -1330 682 -1287 716
rect -1253 682 -1210 716
rect -1330 648 -1210 682
rect -1330 614 -1287 648
rect -1253 614 -1210 648
rect -1330 580 -1210 614
rect -1330 546 -1287 580
rect -1253 546 -1210 580
rect -1330 512 -1210 546
rect -1330 478 -1287 512
rect -1253 478 -1210 512
rect -1330 444 -1210 478
rect -1330 410 -1287 444
rect -1253 410 -1210 444
rect -1330 376 -1210 410
rect -1330 342 -1287 376
rect -1253 342 -1210 376
rect -1330 308 -1210 342
rect -1330 274 -1287 308
rect -1253 274 -1210 308
rect -1330 240 -1210 274
rect -1330 206 -1287 240
rect -1253 206 -1210 240
rect -1330 172 -1210 206
rect -1330 138 -1287 172
rect -1253 138 -1210 172
rect -1330 104 -1210 138
rect -1330 70 -1287 104
rect -1253 70 -1210 104
rect -1330 20 -1210 70
rect -1110 920 -990 970
rect -1110 886 -1067 920
rect -1033 886 -990 920
rect -1110 852 -990 886
rect -1110 818 -1067 852
rect -1033 818 -990 852
rect -1110 784 -990 818
rect -1110 750 -1067 784
rect -1033 750 -990 784
rect -1110 716 -990 750
rect -1110 682 -1067 716
rect -1033 682 -990 716
rect -1110 648 -990 682
rect -1110 614 -1067 648
rect -1033 614 -990 648
rect -1110 580 -990 614
rect -1110 546 -1067 580
rect -1033 546 -990 580
rect -1110 512 -990 546
rect -1110 478 -1067 512
rect -1033 478 -990 512
rect -1110 444 -990 478
rect -1110 410 -1067 444
rect -1033 410 -990 444
rect -1110 376 -990 410
rect -1110 342 -1067 376
rect -1033 342 -990 376
rect -1110 308 -990 342
rect -1110 274 -1067 308
rect -1033 274 -990 308
rect -1110 240 -990 274
rect -1110 206 -1067 240
rect -1033 206 -990 240
rect -1110 172 -990 206
rect -1110 138 -1067 172
rect -1033 138 -990 172
rect -1110 104 -990 138
rect -1110 70 -1067 104
rect -1033 70 -990 104
rect -1110 20 -990 70
<< ndiffc >>
rect -1947 886 -1913 920
rect -1947 818 -1913 852
rect -1947 750 -1913 784
rect -1947 682 -1913 716
rect -1947 614 -1913 648
rect -1947 546 -1913 580
rect -1947 478 -1913 512
rect -1947 410 -1913 444
rect -1947 342 -1913 376
rect -1947 274 -1913 308
rect -1947 206 -1913 240
rect -1947 138 -1913 172
rect -1947 70 -1913 104
rect -1727 886 -1693 920
rect -1727 818 -1693 852
rect -1727 750 -1693 784
rect -1727 682 -1693 716
rect -1727 614 -1693 648
rect -1727 546 -1693 580
rect -1727 478 -1693 512
rect -1727 410 -1693 444
rect -1727 342 -1693 376
rect -1727 274 -1693 308
rect -1727 206 -1693 240
rect -1727 138 -1693 172
rect -1727 70 -1693 104
rect -1507 886 -1473 920
rect -1507 818 -1473 852
rect -1507 750 -1473 784
rect -1507 682 -1473 716
rect -1507 614 -1473 648
rect -1507 546 -1473 580
rect -1507 478 -1473 512
rect -1507 410 -1473 444
rect -1507 342 -1473 376
rect -1507 274 -1473 308
rect -1507 206 -1473 240
rect -1507 138 -1473 172
rect -1507 70 -1473 104
rect -1287 886 -1253 920
rect -1287 818 -1253 852
rect -1287 750 -1253 784
rect -1287 682 -1253 716
rect -1287 614 -1253 648
rect -1287 546 -1253 580
rect -1287 478 -1253 512
rect -1287 410 -1253 444
rect -1287 342 -1253 376
rect -1287 274 -1253 308
rect -1287 206 -1253 240
rect -1287 138 -1253 172
rect -1287 70 -1253 104
rect -1067 886 -1033 920
rect -1067 818 -1033 852
rect -1067 750 -1033 784
rect -1067 682 -1033 716
rect -1067 614 -1033 648
rect -1067 546 -1033 580
rect -1067 478 -1033 512
rect -1067 410 -1033 444
rect -1067 342 -1033 376
rect -1067 274 -1033 308
rect -1067 206 -1033 240
rect -1067 138 -1033 172
rect -1067 70 -1033 104
<< psubdiff >>
rect -2110 920 -1990 970
rect -2110 886 -2067 920
rect -2033 886 -1990 920
rect -2110 852 -1990 886
rect -2110 818 -2067 852
rect -2033 818 -1990 852
rect -2110 784 -1990 818
rect -2110 750 -2067 784
rect -2033 750 -1990 784
rect -2110 716 -1990 750
rect -2110 682 -2067 716
rect -2033 682 -1990 716
rect -2110 648 -1990 682
rect -2110 614 -2067 648
rect -2033 614 -1990 648
rect -2110 580 -1990 614
rect -2110 546 -2067 580
rect -2033 546 -1990 580
rect -2110 512 -1990 546
rect -2110 478 -2067 512
rect -2033 478 -1990 512
rect -2110 444 -1990 478
rect -2110 410 -2067 444
rect -2033 410 -1990 444
rect -2110 376 -1990 410
rect -2110 342 -2067 376
rect -2033 342 -1990 376
rect -2110 308 -1990 342
rect -2110 274 -2067 308
rect -2033 274 -1990 308
rect -2110 240 -1990 274
rect -2110 206 -2067 240
rect -2033 206 -1990 240
rect -2110 172 -1990 206
rect -2110 138 -2067 172
rect -2033 138 -1990 172
rect -2110 104 -1990 138
rect -2110 70 -2067 104
rect -2033 70 -1990 104
rect -2110 20 -1990 70
<< psubdiffcont >>
rect -2067 886 -2033 920
rect -2067 818 -2033 852
rect -2067 750 -2033 784
rect -2067 682 -2033 716
rect -2067 614 -2033 648
rect -2067 546 -2033 580
rect -2067 478 -2033 512
rect -2067 410 -2033 444
rect -2067 342 -2033 376
rect -2067 274 -2033 308
rect -2067 206 -2033 240
rect -2067 138 -2033 172
rect -2067 70 -2033 104
<< poly >>
rect -1870 1020 -1110 1050
rect -1870 970 -1770 1020
rect -1650 970 -1550 1020
rect -1430 970 -1330 1020
rect -1210 970 -1110 1020
rect -1870 -10 -1770 20
rect -1650 -10 -1550 20
rect -1430 -10 -1330 20
rect -1210 -10 -1110 20
<< locali >>
rect -1730 990 -1250 1030
rect -1730 950 -1690 990
rect -1290 950 -1250 990
rect -2090 920 -2010 950
rect -2090 886 -2067 920
rect -2033 886 -2010 920
rect -2090 852 -2010 886
rect -2090 818 -2067 852
rect -2033 818 -2010 852
rect -2090 784 -2010 818
rect -2090 750 -2067 784
rect -2033 750 -2010 784
rect -2090 716 -2010 750
rect -2090 682 -2067 716
rect -2033 682 -2010 716
rect -2090 648 -2010 682
rect -2090 614 -2067 648
rect -2033 614 -2010 648
rect -2090 580 -2010 614
rect -2090 546 -2067 580
rect -2033 546 -2010 580
rect -2090 512 -2010 546
rect -2090 478 -2067 512
rect -2033 478 -2010 512
rect -2090 444 -2010 478
rect -2090 410 -2067 444
rect -2033 410 -2010 444
rect -2090 376 -2010 410
rect -2090 342 -2067 376
rect -2033 342 -2010 376
rect -2090 308 -2010 342
rect -2090 274 -2067 308
rect -2033 274 -2010 308
rect -2090 240 -2010 274
rect -2090 206 -2067 240
rect -2033 206 -2010 240
rect -2090 172 -2010 206
rect -2090 138 -2067 172
rect -2033 138 -2010 172
rect -2090 104 -2010 138
rect -2090 70 -2067 104
rect -2033 70 -2010 104
rect -2090 40 -2010 70
rect -1970 920 -1890 950
rect -1970 886 -1947 920
rect -1913 886 -1890 920
rect -1970 852 -1890 886
rect -1970 818 -1947 852
rect -1913 818 -1890 852
rect -1970 784 -1890 818
rect -1970 750 -1947 784
rect -1913 750 -1890 784
rect -1970 716 -1890 750
rect -1970 682 -1947 716
rect -1913 682 -1890 716
rect -1970 648 -1890 682
rect -1970 614 -1947 648
rect -1913 614 -1890 648
rect -1970 580 -1890 614
rect -1970 546 -1947 580
rect -1913 546 -1890 580
rect -1970 512 -1890 546
rect -1970 478 -1947 512
rect -1913 478 -1890 512
rect -1970 444 -1890 478
rect -1970 410 -1947 444
rect -1913 410 -1890 444
rect -1970 376 -1890 410
rect -1970 342 -1947 376
rect -1913 342 -1890 376
rect -1970 308 -1890 342
rect -1970 274 -1947 308
rect -1913 274 -1890 308
rect -1970 240 -1890 274
rect -1970 206 -1947 240
rect -1913 206 -1890 240
rect -1970 172 -1890 206
rect -1970 138 -1947 172
rect -1913 138 -1890 172
rect -1970 104 -1890 138
rect -1970 70 -1947 104
rect -1913 70 -1890 104
rect -1970 40 -1890 70
rect -1750 920 -1670 950
rect -1750 886 -1727 920
rect -1693 886 -1670 920
rect -1750 852 -1670 886
rect -1750 818 -1727 852
rect -1693 818 -1670 852
rect -1750 784 -1670 818
rect -1750 750 -1727 784
rect -1693 750 -1670 784
rect -1750 716 -1670 750
rect -1750 682 -1727 716
rect -1693 682 -1670 716
rect -1750 648 -1670 682
rect -1750 614 -1727 648
rect -1693 614 -1670 648
rect -1750 580 -1670 614
rect -1750 546 -1727 580
rect -1693 546 -1670 580
rect -1750 512 -1670 546
rect -1750 478 -1727 512
rect -1693 478 -1670 512
rect -1750 444 -1670 478
rect -1750 410 -1727 444
rect -1693 410 -1670 444
rect -1750 376 -1670 410
rect -1750 342 -1727 376
rect -1693 342 -1670 376
rect -1750 308 -1670 342
rect -1750 274 -1727 308
rect -1693 274 -1670 308
rect -1750 240 -1670 274
rect -1750 206 -1727 240
rect -1693 206 -1670 240
rect -1750 172 -1670 206
rect -1750 138 -1727 172
rect -1693 138 -1670 172
rect -1750 104 -1670 138
rect -1750 70 -1727 104
rect -1693 70 -1670 104
rect -1750 40 -1670 70
rect -1530 920 -1450 950
rect -1530 886 -1507 920
rect -1473 886 -1450 920
rect -1530 852 -1450 886
rect -1530 818 -1507 852
rect -1473 818 -1450 852
rect -1530 784 -1450 818
rect -1530 750 -1507 784
rect -1473 750 -1450 784
rect -1530 716 -1450 750
rect -1530 682 -1507 716
rect -1473 682 -1450 716
rect -1530 648 -1450 682
rect -1530 614 -1507 648
rect -1473 614 -1450 648
rect -1530 580 -1450 614
rect -1530 546 -1507 580
rect -1473 546 -1450 580
rect -1530 512 -1450 546
rect -1530 478 -1507 512
rect -1473 478 -1450 512
rect -1530 444 -1450 478
rect -1530 410 -1507 444
rect -1473 410 -1450 444
rect -1530 376 -1450 410
rect -1530 342 -1507 376
rect -1473 342 -1450 376
rect -1530 308 -1450 342
rect -1530 274 -1507 308
rect -1473 274 -1450 308
rect -1530 240 -1450 274
rect -1530 206 -1507 240
rect -1473 206 -1450 240
rect -1530 172 -1450 206
rect -1530 138 -1507 172
rect -1473 138 -1450 172
rect -1530 104 -1450 138
rect -1530 70 -1507 104
rect -1473 70 -1450 104
rect -1530 40 -1450 70
rect -1310 920 -1230 950
rect -1310 886 -1287 920
rect -1253 886 -1230 920
rect -1310 852 -1230 886
rect -1310 818 -1287 852
rect -1253 818 -1230 852
rect -1310 784 -1230 818
rect -1310 750 -1287 784
rect -1253 750 -1230 784
rect -1310 716 -1230 750
rect -1310 682 -1287 716
rect -1253 682 -1230 716
rect -1310 648 -1230 682
rect -1310 614 -1287 648
rect -1253 614 -1230 648
rect -1310 580 -1230 614
rect -1310 546 -1287 580
rect -1253 546 -1230 580
rect -1310 512 -1230 546
rect -1310 478 -1287 512
rect -1253 478 -1230 512
rect -1310 444 -1230 478
rect -1310 410 -1287 444
rect -1253 410 -1230 444
rect -1310 376 -1230 410
rect -1310 342 -1287 376
rect -1253 342 -1230 376
rect -1310 308 -1230 342
rect -1310 274 -1287 308
rect -1253 274 -1230 308
rect -1310 240 -1230 274
rect -1310 206 -1287 240
rect -1253 206 -1230 240
rect -1310 172 -1230 206
rect -1310 138 -1287 172
rect -1253 138 -1230 172
rect -1310 104 -1230 138
rect -1310 70 -1287 104
rect -1253 70 -1230 104
rect -1310 40 -1230 70
rect -1090 920 -1010 950
rect -1090 886 -1067 920
rect -1033 886 -1010 920
rect -1090 852 -1010 886
rect -1090 818 -1067 852
rect -1033 818 -1010 852
rect -1090 784 -1010 818
rect -1090 750 -1067 784
rect -1033 750 -1010 784
rect -1090 716 -1010 750
rect -1090 682 -1067 716
rect -1033 682 -1010 716
rect -1090 648 -1010 682
rect -1090 614 -1067 648
rect -1033 614 -1010 648
rect -1090 580 -1010 614
rect -1090 546 -1067 580
rect -1033 546 -1010 580
rect -1090 512 -1010 546
rect -1090 478 -1067 512
rect -1033 478 -1010 512
rect -1090 444 -1010 478
rect -1090 410 -1067 444
rect -1033 410 -1010 444
rect -1090 376 -1010 410
rect -1090 342 -1067 376
rect -1033 342 -1010 376
rect -1090 308 -1010 342
rect -1090 274 -1067 308
rect -1033 274 -1010 308
rect -1090 240 -1010 274
rect -1090 206 -1067 240
rect -1033 206 -1010 240
rect -1090 172 -1010 206
rect -1090 138 -1067 172
rect -1033 138 -1010 172
rect -1090 104 -1010 138
rect -1090 70 -1067 104
rect -1033 70 -1010 104
rect -1090 40 -1010 70
rect -1950 0 -1910 40
rect -1510 0 -1470 40
rect -1070 0 -1030 40
rect -1950 -40 -1030 0
<< end >>
