magic
tech sky130A
timestamp 1676416811
<< nwell >>
rect -680 655 -160 1000
<< nmos >>
rect -600 450 -585 600
rect -525 450 -510 600
rect -450 450 -435 600
rect -255 450 -240 600
<< pmos >>
rect -600 680 -585 980
rect -525 680 -510 980
rect -450 680 -435 980
rect -255 680 -240 980
<< ndiff >>
rect -660 585 -600 600
rect -660 465 -640 585
rect -620 465 -600 585
rect -660 450 -600 465
rect -585 585 -525 600
rect -585 465 -565 585
rect -545 465 -525 585
rect -585 450 -525 465
rect -510 585 -450 600
rect -510 465 -490 585
rect -470 465 -450 585
rect -510 450 -450 465
rect -435 585 -375 600
rect -435 465 -415 585
rect -395 465 -375 585
rect -435 450 -375 465
rect -315 585 -255 600
rect -315 465 -295 585
rect -275 465 -255 585
rect -315 450 -255 465
rect -240 585 -180 600
rect -240 465 -220 585
rect -200 465 -180 585
rect -240 450 -180 465
<< pdiff >>
rect -660 965 -600 980
rect -660 695 -640 965
rect -620 695 -600 965
rect -660 680 -600 695
rect -585 680 -525 980
rect -510 680 -450 980
rect -435 965 -375 980
rect -435 695 -415 965
rect -395 695 -375 965
rect -435 680 -375 695
rect -315 965 -255 980
rect -315 695 -295 965
rect -275 695 -255 965
rect -315 680 -255 695
rect -240 960 -180 980
rect -240 700 -220 960
rect -200 700 -180 960
rect -240 680 -180 700
<< ndiffc >>
rect -640 465 -620 585
rect -565 465 -545 585
rect -490 465 -470 585
rect -415 465 -395 585
rect -295 465 -275 585
rect -220 465 -200 585
<< pdiffc >>
rect -640 695 -620 965
rect -415 695 -395 965
rect -295 695 -275 965
rect -220 700 -200 960
<< poly >>
rect -600 980 -585 995
rect -525 980 -510 995
rect -450 980 -435 995
rect -255 980 -240 995
rect -600 660 -585 680
rect -625 650 -585 660
rect -625 630 -615 650
rect -595 630 -585 650
rect -625 620 -585 630
rect -600 600 -585 620
rect -525 600 -510 680
rect -450 600 -435 680
rect -255 665 -240 680
rect -295 655 -240 665
rect -295 635 -285 655
rect -265 635 -240 655
rect -295 625 -240 635
rect -255 600 -240 625
rect -600 435 -585 450
rect -525 400 -510 450
rect -450 400 -435 450
rect -255 435 -240 450
rect -550 390 -510 400
rect -550 370 -540 390
rect -520 370 -510 390
rect -550 360 -510 370
rect -465 390 -425 400
rect -465 370 -455 390
rect -435 370 -425 390
rect -465 360 -425 370
<< polycont >>
rect -615 630 -595 650
rect -285 635 -265 655
rect -540 370 -520 390
rect -455 370 -435 390
<< locali >>
rect -650 965 -610 970
rect -650 695 -640 965
rect -620 695 -610 965
rect -650 690 -610 695
rect -425 965 -385 970
rect -425 695 -415 965
rect -395 695 -385 965
rect -425 690 -385 695
rect -305 965 -265 970
rect -305 695 -295 965
rect -275 695 -265 965
rect -305 690 -265 695
rect -230 960 -190 970
rect -230 700 -220 960
rect -200 700 -190 960
rect -230 690 -190 700
rect -625 650 -585 660
rect -415 655 -395 690
rect -295 655 -255 665
rect -625 630 -615 650
rect -595 630 -585 650
rect -625 620 -585 630
rect -490 635 -285 655
rect -265 635 -255 655
rect -490 590 -470 635
rect -295 625 -255 635
rect -220 590 -200 690
rect -650 585 -610 590
rect -650 465 -640 585
rect -620 465 -610 585
rect -650 460 -610 465
rect -575 585 -535 590
rect -575 465 -565 585
rect -545 465 -535 585
rect -575 460 -535 465
rect -500 585 -460 590
rect -500 465 -490 585
rect -470 465 -460 585
rect -500 460 -460 465
rect -425 585 -385 590
rect -425 465 -415 585
rect -395 465 -385 585
rect -425 460 -385 465
rect -305 585 -265 590
rect -305 465 -295 585
rect -275 465 -265 585
rect -305 460 -265 465
rect -230 585 -190 590
rect -230 465 -220 585
rect -200 465 -190 585
rect -230 460 -190 465
rect -640 440 -620 460
rect -490 440 -470 460
rect -640 420 -470 440
rect -550 390 -510 400
rect -550 370 -540 390
rect -520 370 -510 390
rect -550 360 -510 370
rect -465 390 -425 400
rect -465 370 -455 390
rect -435 370 -425 390
rect -465 360 -425 370
<< viali >>
rect -640 695 -620 965
rect -295 695 -275 965
rect -565 465 -545 585
rect -415 465 -395 585
rect -295 465 -275 585
<< metal1 >>
rect -650 965 -610 970
rect -650 695 -640 965
rect -620 695 -610 965
rect -650 690 -610 695
rect -305 965 -265 970
rect -305 695 -295 965
rect -275 695 -265 965
rect -305 690 -265 695
rect -575 585 -535 590
rect -575 465 -565 585
rect -545 465 -535 585
rect -575 460 -535 465
rect -425 585 -385 590
rect -425 465 -415 585
rect -395 465 -385 585
rect -425 460 -385 465
rect -305 585 -265 590
rect -305 465 -295 585
rect -275 465 -265 585
rect -305 460 -265 465
<< end >>
