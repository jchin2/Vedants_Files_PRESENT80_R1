magic
tech sky130A
magscale 1 2
timestamp 1675786016
<< nwell >>
rect -2010 1450 -250 1640
rect -1540 1060 -720 1450
<< pwell >>
rect -1996 284 -264 876
<< nmos >>
rect -1850 550 -1820 850
rect -1700 550 -1670 850
rect -1370 550 -1340 850
rect -1220 550 -1190 850
rect -1070 550 -1040 850
rect -920 550 -890 850
rect -590 550 -560 850
rect -440 550 -410 850
<< pmos >>
rect -1370 1110 -1340 1410
rect -1220 1110 -1190 1410
rect -1070 1110 -1040 1410
rect -920 1110 -890 1410
<< ndiff >>
rect -1970 777 -1850 850
rect -1970 743 -1927 777
rect -1893 743 -1850 777
rect -1970 697 -1850 743
rect -1970 663 -1927 697
rect -1893 663 -1850 697
rect -1970 617 -1850 663
rect -1970 583 -1927 617
rect -1893 583 -1850 617
rect -1970 550 -1850 583
rect -1820 550 -1700 850
rect -1670 777 -1550 850
rect -1670 743 -1627 777
rect -1593 743 -1550 777
rect -1670 697 -1550 743
rect -1670 663 -1627 697
rect -1593 663 -1550 697
rect -1670 617 -1550 663
rect -1670 583 -1627 617
rect -1593 583 -1550 617
rect -1670 550 -1550 583
rect -1490 777 -1370 850
rect -1490 743 -1447 777
rect -1413 743 -1370 777
rect -1490 697 -1370 743
rect -1490 663 -1447 697
rect -1413 663 -1370 697
rect -1490 617 -1370 663
rect -1490 583 -1447 617
rect -1413 583 -1370 617
rect -1490 550 -1370 583
rect -1340 777 -1220 850
rect -1340 743 -1297 777
rect -1263 743 -1220 777
rect -1340 697 -1220 743
rect -1340 663 -1297 697
rect -1263 663 -1220 697
rect -1340 617 -1220 663
rect -1340 583 -1297 617
rect -1263 583 -1220 617
rect -1340 550 -1220 583
rect -1190 777 -1070 850
rect -1190 743 -1147 777
rect -1113 743 -1070 777
rect -1190 697 -1070 743
rect -1190 663 -1147 697
rect -1113 663 -1070 697
rect -1190 617 -1070 663
rect -1190 583 -1147 617
rect -1113 583 -1070 617
rect -1190 550 -1070 583
rect -1040 777 -920 850
rect -1040 743 -997 777
rect -963 743 -920 777
rect -1040 697 -920 743
rect -1040 663 -997 697
rect -963 663 -920 697
rect -1040 617 -920 663
rect -1040 583 -997 617
rect -963 583 -920 617
rect -1040 550 -920 583
rect -890 777 -770 850
rect -890 743 -847 777
rect -813 743 -770 777
rect -890 697 -770 743
rect -890 663 -847 697
rect -813 663 -770 697
rect -890 617 -770 663
rect -890 583 -847 617
rect -813 583 -770 617
rect -890 550 -770 583
rect -710 777 -590 850
rect -710 743 -667 777
rect -633 743 -590 777
rect -710 697 -590 743
rect -710 663 -667 697
rect -633 663 -590 697
rect -710 617 -590 663
rect -710 583 -667 617
rect -633 583 -590 617
rect -710 550 -590 583
rect -560 777 -440 850
rect -560 743 -517 777
rect -483 743 -440 777
rect -560 697 -440 743
rect -560 663 -517 697
rect -483 663 -440 697
rect -560 617 -440 663
rect -560 583 -517 617
rect -483 583 -440 617
rect -560 550 -440 583
rect -410 777 -290 850
rect -410 743 -367 777
rect -333 743 -290 777
rect -410 697 -290 743
rect -410 663 -367 697
rect -333 663 -290 697
rect -410 617 -290 663
rect -410 583 -367 617
rect -333 583 -290 617
rect -410 550 -290 583
<< pdiff >>
rect -1490 1337 -1370 1410
rect -1490 1303 -1447 1337
rect -1413 1303 -1370 1337
rect -1490 1257 -1370 1303
rect -1490 1223 -1447 1257
rect -1413 1223 -1370 1257
rect -1490 1177 -1370 1223
rect -1490 1143 -1447 1177
rect -1413 1143 -1370 1177
rect -1490 1110 -1370 1143
rect -1340 1337 -1220 1410
rect -1340 1303 -1297 1337
rect -1263 1303 -1220 1337
rect -1340 1257 -1220 1303
rect -1340 1223 -1297 1257
rect -1263 1223 -1220 1257
rect -1340 1177 -1220 1223
rect -1340 1143 -1297 1177
rect -1263 1143 -1220 1177
rect -1340 1110 -1220 1143
rect -1190 1337 -1070 1410
rect -1190 1303 -1147 1337
rect -1113 1303 -1070 1337
rect -1190 1257 -1070 1303
rect -1190 1223 -1147 1257
rect -1113 1223 -1070 1257
rect -1190 1177 -1070 1223
rect -1190 1143 -1147 1177
rect -1113 1143 -1070 1177
rect -1190 1110 -1070 1143
rect -1040 1337 -920 1410
rect -1040 1303 -997 1337
rect -963 1303 -920 1337
rect -1040 1257 -920 1303
rect -1040 1223 -997 1257
rect -963 1223 -920 1257
rect -1040 1177 -920 1223
rect -1040 1143 -997 1177
rect -963 1143 -920 1177
rect -1040 1110 -920 1143
rect -890 1337 -770 1410
rect -890 1303 -847 1337
rect -813 1303 -770 1337
rect -890 1257 -770 1303
rect -890 1223 -847 1257
rect -813 1223 -770 1257
rect -890 1177 -770 1223
rect -890 1143 -847 1177
rect -813 1143 -770 1177
rect -890 1110 -770 1143
<< ndiffc >>
rect -1927 743 -1893 777
rect -1927 663 -1893 697
rect -1927 583 -1893 617
rect -1627 743 -1593 777
rect -1627 663 -1593 697
rect -1627 583 -1593 617
rect -1447 743 -1413 777
rect -1447 663 -1413 697
rect -1447 583 -1413 617
rect -1297 743 -1263 777
rect -1297 663 -1263 697
rect -1297 583 -1263 617
rect -1147 743 -1113 777
rect -1147 663 -1113 697
rect -1147 583 -1113 617
rect -997 743 -963 777
rect -997 663 -963 697
rect -997 583 -963 617
rect -847 743 -813 777
rect -847 663 -813 697
rect -847 583 -813 617
rect -667 743 -633 777
rect -667 663 -633 697
rect -667 583 -633 617
rect -517 743 -483 777
rect -517 663 -483 697
rect -517 583 -483 617
rect -367 743 -333 777
rect -367 663 -333 697
rect -367 583 -333 617
<< pdiffc >>
rect -1447 1303 -1413 1337
rect -1447 1223 -1413 1257
rect -1447 1143 -1413 1177
rect -1297 1303 -1263 1337
rect -1297 1223 -1263 1257
rect -1297 1143 -1263 1177
rect -1147 1303 -1113 1337
rect -1147 1223 -1113 1257
rect -1147 1143 -1113 1177
rect -997 1303 -963 1337
rect -997 1223 -963 1257
rect -997 1143 -963 1177
rect -847 1303 -813 1337
rect -847 1223 -813 1257
rect -847 1143 -813 1177
<< psubdiff >>
rect -1970 377 -290 410
rect -1970 343 -1947 377
rect -1913 343 -1867 377
rect -1833 343 -1787 377
rect -1753 343 -1707 377
rect -1673 343 -1627 377
rect -1593 343 -1547 377
rect -1513 343 -1467 377
rect -1433 343 -1387 377
rect -1353 343 -1307 377
rect -1273 343 -1227 377
rect -1193 343 -1147 377
rect -1113 343 -1067 377
rect -1033 343 -987 377
rect -953 343 -907 377
rect -873 343 -827 377
rect -793 343 -747 377
rect -713 343 -667 377
rect -633 343 -587 377
rect -553 343 -507 377
rect -473 343 -427 377
rect -393 343 -347 377
rect -313 343 -290 377
rect -1970 310 -290 343
<< nsubdiff >>
rect -1970 1557 -290 1590
rect -1970 1523 -1947 1557
rect -1913 1523 -1867 1557
rect -1833 1523 -1787 1557
rect -1753 1523 -1707 1557
rect -1673 1523 -1627 1557
rect -1593 1523 -1547 1557
rect -1513 1523 -1467 1557
rect -1433 1523 -1387 1557
rect -1353 1523 -1307 1557
rect -1273 1523 -1227 1557
rect -1193 1523 -1147 1557
rect -1113 1523 -1067 1557
rect -1033 1523 -987 1557
rect -953 1523 -907 1557
rect -873 1523 -827 1557
rect -793 1523 -747 1557
rect -713 1523 -667 1557
rect -633 1523 -587 1557
rect -553 1523 -507 1557
rect -473 1523 -427 1557
rect -393 1523 -347 1557
rect -313 1523 -290 1557
rect -1970 1490 -290 1523
<< psubdiffcont >>
rect -1947 343 -1913 377
rect -1867 343 -1833 377
rect -1787 343 -1753 377
rect -1707 343 -1673 377
rect -1627 343 -1593 377
rect -1547 343 -1513 377
rect -1467 343 -1433 377
rect -1387 343 -1353 377
rect -1307 343 -1273 377
rect -1227 343 -1193 377
rect -1147 343 -1113 377
rect -1067 343 -1033 377
rect -987 343 -953 377
rect -907 343 -873 377
rect -827 343 -793 377
rect -747 343 -713 377
rect -667 343 -633 377
rect -587 343 -553 377
rect -507 343 -473 377
rect -427 343 -393 377
rect -347 343 -313 377
<< nsubdiffcont >>
rect -1947 1523 -1913 1557
rect -1867 1523 -1833 1557
rect -1787 1523 -1753 1557
rect -1707 1523 -1673 1557
rect -1627 1523 -1593 1557
rect -1547 1523 -1513 1557
rect -1467 1523 -1433 1557
rect -1387 1523 -1353 1557
rect -1307 1523 -1273 1557
rect -1227 1523 -1193 1557
rect -1147 1523 -1113 1557
rect -1067 1523 -1033 1557
rect -987 1523 -953 1557
rect -907 1523 -873 1557
rect -827 1523 -793 1557
rect -747 1523 -713 1557
rect -667 1523 -633 1557
rect -587 1523 -553 1557
rect -507 1523 -473 1557
rect -427 1523 -393 1557
rect -347 1523 -313 1557
<< poly >>
rect -1370 1440 -1190 1470
rect -1370 1410 -1340 1440
rect -1220 1410 -1190 1440
rect -1070 1440 -890 1470
rect -1070 1410 -1040 1440
rect -920 1410 -890 1440
rect -440 1297 -360 1320
rect -440 1263 -417 1297
rect -383 1263 -360 1297
rect -440 1240 -360 1263
rect -640 1177 -560 1200
rect -640 1143 -617 1177
rect -583 1143 -560 1177
rect -640 1120 -560 1143
rect -1750 1077 -1670 1100
rect -1370 1080 -1340 1110
rect -1750 1043 -1727 1077
rect -1693 1043 -1670 1077
rect -1750 1020 -1670 1043
rect -1900 977 -1820 1000
rect -1900 943 -1877 977
rect -1843 943 -1820 977
rect -1900 920 -1820 943
rect -1850 850 -1820 920
rect -1700 850 -1670 1020
rect -1220 955 -1190 1110
rect -1070 1080 -1040 1110
rect -920 1080 -890 1110
rect -1120 1057 -1040 1080
rect -1120 1023 -1097 1057
rect -1063 1023 -1040 1057
rect -1120 1000 -1040 1023
rect -1220 932 -1140 955
rect -1220 898 -1197 932
rect -1163 898 -1140 932
rect -1370 850 -1340 880
rect -1220 875 -1140 898
rect -1220 850 -1190 875
rect -1070 850 -1040 1000
rect -920 850 -890 880
rect -590 850 -560 1120
rect -440 850 -410 1240
rect -1850 520 -1820 550
rect -1700 520 -1670 550
rect -1370 520 -1340 550
rect -1220 520 -1190 550
rect -1070 520 -1040 550
rect -920 520 -890 550
rect -590 520 -560 550
rect -440 520 -410 550
rect -1370 497 -1290 520
rect -1370 463 -1347 497
rect -1313 463 -1290 497
rect -1370 440 -1290 463
rect -970 497 -890 520
rect -970 463 -947 497
rect -913 463 -890 497
rect -970 440 -890 463
<< polycont >>
rect -417 1263 -383 1297
rect -617 1143 -583 1177
rect -1727 1043 -1693 1077
rect -1877 943 -1843 977
rect -1097 1023 -1063 1057
rect -1197 898 -1163 932
rect -1347 463 -1313 497
rect -947 463 -913 497
<< locali >>
rect -1970 1557 -290 1580
rect -1970 1523 -1947 1557
rect -1913 1523 -1867 1557
rect -1833 1523 -1787 1557
rect -1753 1523 -1707 1557
rect -1673 1523 -1627 1557
rect -1593 1523 -1547 1557
rect -1513 1523 -1467 1557
rect -1433 1523 -1387 1557
rect -1353 1523 -1307 1557
rect -1273 1523 -1227 1557
rect -1193 1523 -1147 1557
rect -1113 1523 -1067 1557
rect -1033 1523 -987 1557
rect -953 1523 -907 1557
rect -873 1523 -827 1557
rect -793 1523 -747 1557
rect -713 1523 -667 1557
rect -633 1523 -587 1557
rect -553 1523 -507 1557
rect -473 1523 -427 1557
rect -393 1523 -347 1557
rect -313 1523 -290 1557
rect -1970 1500 -290 1523
rect -1470 1337 -1390 1370
rect -1620 1300 -1540 1320
rect -1970 1297 -1540 1300
rect -1970 1263 -1597 1297
rect -1563 1263 -1540 1297
rect -1970 1260 -1540 1263
rect -1620 1240 -1540 1260
rect -1470 1303 -1447 1337
rect -1413 1303 -1390 1337
rect -1470 1257 -1390 1303
rect -1470 1223 -1447 1257
rect -1413 1223 -1390 1257
rect -1620 1180 -1540 1200
rect -1970 1177 -1540 1180
rect -1970 1143 -1597 1177
rect -1563 1143 -1540 1177
rect -1970 1140 -1540 1143
rect -1620 1120 -1540 1140
rect -1470 1177 -1390 1223
rect -1470 1143 -1447 1177
rect -1413 1143 -1390 1177
rect -1470 1120 -1390 1143
rect -1320 1337 -1240 1370
rect -1320 1303 -1297 1337
rect -1263 1303 -1240 1337
rect -1320 1257 -1240 1303
rect -1320 1223 -1297 1257
rect -1263 1223 -1240 1257
rect -1320 1177 -1240 1223
rect -1320 1143 -1297 1177
rect -1263 1143 -1240 1177
rect -1320 1110 -1240 1143
rect -1170 1337 -1090 1370
rect -1170 1303 -1147 1337
rect -1113 1303 -1090 1337
rect -1170 1257 -1090 1303
rect -1170 1223 -1147 1257
rect -1113 1223 -1090 1257
rect -1170 1177 -1090 1223
rect -1170 1143 -1147 1177
rect -1113 1143 -1090 1177
rect -1170 1120 -1090 1143
rect -1020 1337 -940 1370
rect -1020 1303 -997 1337
rect -963 1303 -940 1337
rect -1020 1257 -940 1303
rect -1020 1223 -997 1257
rect -963 1223 -940 1257
rect -1020 1177 -940 1223
rect -1020 1143 -997 1177
rect -963 1143 -940 1177
rect -1020 1110 -940 1143
rect -870 1337 -790 1370
rect -870 1303 -847 1337
rect -813 1303 -790 1337
rect -870 1257 -790 1303
rect -870 1223 -847 1257
rect -813 1223 -790 1257
rect -440 1297 -360 1320
rect -440 1263 -417 1297
rect -383 1263 -360 1297
rect -440 1240 -360 1263
rect -870 1177 -790 1223
rect -870 1143 -847 1177
rect -813 1143 -790 1177
rect -870 1120 -790 1143
rect -640 1177 -560 1200
rect -640 1143 -617 1177
rect -583 1143 -560 1177
rect -640 1120 -560 1143
rect -1750 1080 -1670 1100
rect -1970 1077 -1670 1080
rect -1970 1043 -1727 1077
rect -1693 1043 -1670 1077
rect -1970 1040 -1670 1043
rect -1750 1020 -1670 1040
rect -1300 1060 -1260 1110
rect -1120 1060 -1040 1080
rect -1300 1057 -1040 1060
rect -1300 1023 -1097 1057
rect -1063 1023 -1040 1057
rect -1300 1020 -1040 1023
rect -1900 980 -1820 1000
rect -1970 977 -1820 980
rect -1970 943 -1877 977
rect -1843 943 -1820 977
rect -1970 940 -1820 943
rect -1900 920 -1820 940
rect -1300 890 -1260 1020
rect -1120 1000 -1040 1020
rect -1630 850 -1260 890
rect -1220 940 -1140 955
rect -1000 940 -960 1110
rect -720 1060 -640 1080
rect -720 1057 -290 1060
rect -720 1023 -697 1057
rect -663 1023 -290 1057
rect -720 1020 -290 1023
rect -720 1000 -640 1020
rect -1220 932 -290 940
rect -1220 898 -1197 932
rect -1163 900 -290 932
rect -1163 898 -1140 900
rect -1220 875 -1140 898
rect -1630 810 -1590 850
rect -1300 810 -1260 850
rect -1000 810 -960 900
rect -690 810 -650 900
rect -370 810 -330 900
rect -1950 777 -1870 810
rect -1950 743 -1927 777
rect -1893 743 -1870 777
rect -1950 697 -1870 743
rect -1950 663 -1927 697
rect -1893 663 -1870 697
rect -1950 617 -1870 663
rect -1950 583 -1927 617
rect -1893 583 -1870 617
rect -1950 560 -1870 583
rect -1650 777 -1570 810
rect -1650 743 -1627 777
rect -1593 743 -1570 777
rect -1650 697 -1570 743
rect -1650 663 -1627 697
rect -1593 663 -1570 697
rect -1650 617 -1570 663
rect -1650 583 -1627 617
rect -1593 583 -1570 617
rect -1650 560 -1570 583
rect -1470 777 -1390 810
rect -1470 743 -1447 777
rect -1413 743 -1390 777
rect -1470 697 -1390 743
rect -1470 663 -1447 697
rect -1413 663 -1390 697
rect -1470 617 -1390 663
rect -1470 583 -1447 617
rect -1413 583 -1390 617
rect -1470 560 -1390 583
rect -1320 777 -1240 810
rect -1320 743 -1297 777
rect -1263 743 -1240 777
rect -1320 697 -1240 743
rect -1320 663 -1297 697
rect -1263 663 -1240 697
rect -1320 617 -1240 663
rect -1320 583 -1297 617
rect -1263 583 -1240 617
rect -1320 560 -1240 583
rect -1170 777 -1090 810
rect -1170 743 -1147 777
rect -1113 743 -1090 777
rect -1170 697 -1090 743
rect -1170 663 -1147 697
rect -1113 663 -1090 697
rect -1170 617 -1090 663
rect -1170 583 -1147 617
rect -1113 583 -1090 617
rect -1170 560 -1090 583
rect -1020 777 -940 810
rect -1020 743 -997 777
rect -963 743 -940 777
rect -1020 697 -940 743
rect -1020 663 -997 697
rect -963 663 -940 697
rect -1020 617 -940 663
rect -1020 583 -997 617
rect -963 583 -940 617
rect -1020 560 -940 583
rect -870 777 -790 810
rect -870 743 -847 777
rect -813 743 -790 777
rect -870 697 -790 743
rect -870 663 -847 697
rect -813 663 -790 697
rect -870 617 -790 663
rect -870 583 -847 617
rect -813 583 -790 617
rect -870 560 -790 583
rect -690 777 -610 810
rect -690 743 -667 777
rect -633 743 -610 777
rect -690 697 -610 743
rect -690 663 -667 697
rect -633 663 -610 697
rect -690 617 -610 663
rect -690 583 -667 617
rect -633 583 -610 617
rect -690 560 -610 583
rect -540 777 -460 810
rect -540 743 -517 777
rect -483 743 -460 777
rect -540 697 -460 743
rect -540 663 -517 697
rect -483 663 -460 697
rect -540 617 -460 663
rect -540 583 -517 617
rect -483 583 -460 617
rect -540 560 -460 583
rect -390 777 -310 810
rect -390 743 -367 777
rect -333 743 -310 777
rect -390 697 -310 743
rect -390 663 -367 697
rect -333 663 -310 697
rect -390 617 -310 663
rect -390 583 -367 617
rect -333 583 -310 617
rect -390 560 -310 583
rect -1370 500 -1290 520
rect -970 500 -890 520
rect -1970 497 -890 500
rect -1970 463 -1347 497
rect -1313 463 -947 497
rect -913 463 -890 497
rect -1970 460 -890 463
rect -1370 440 -1290 460
rect -970 440 -890 460
rect -1970 377 -290 400
rect -1970 343 -1947 377
rect -1913 343 -1867 377
rect -1833 343 -1787 377
rect -1753 343 -1707 377
rect -1673 343 -1627 377
rect -1593 343 -1547 377
rect -1513 343 -1467 377
rect -1433 343 -1387 377
rect -1353 343 -1307 377
rect -1273 343 -1227 377
rect -1193 343 -1147 377
rect -1113 343 -1067 377
rect -1033 343 -987 377
rect -953 343 -907 377
rect -873 343 -827 377
rect -793 343 -747 377
rect -713 343 -667 377
rect -633 343 -587 377
rect -553 343 -507 377
rect -473 343 -427 377
rect -393 343 -347 377
rect -313 343 -290 377
rect -1970 320 -290 343
<< viali >>
rect -1947 1523 -1913 1557
rect -1867 1523 -1833 1557
rect -1787 1523 -1753 1557
rect -1707 1523 -1673 1557
rect -1627 1523 -1593 1557
rect -1547 1523 -1513 1557
rect -1467 1523 -1433 1557
rect -1387 1523 -1353 1557
rect -1307 1523 -1273 1557
rect -1227 1523 -1193 1557
rect -1147 1523 -1113 1557
rect -1067 1523 -1033 1557
rect -987 1523 -953 1557
rect -907 1523 -873 1557
rect -827 1523 -793 1557
rect -747 1523 -713 1557
rect -667 1523 -633 1557
rect -587 1523 -553 1557
rect -507 1523 -473 1557
rect -427 1523 -393 1557
rect -347 1523 -313 1557
rect -1597 1263 -1563 1297
rect -1447 1303 -1413 1337
rect -1447 1223 -1413 1257
rect -1597 1143 -1563 1177
rect -1447 1143 -1413 1177
rect -1147 1303 -1113 1337
rect -1147 1223 -1113 1257
rect -1147 1143 -1113 1177
rect -847 1303 -813 1337
rect -847 1223 -813 1257
rect -417 1263 -383 1297
rect -847 1143 -813 1177
rect -617 1143 -583 1177
rect -1097 1023 -1063 1057
rect -697 1023 -663 1057
rect -1927 743 -1893 777
rect -1927 663 -1893 697
rect -1927 583 -1893 617
rect -1447 743 -1413 777
rect -1447 663 -1413 697
rect -1447 583 -1413 617
rect -1147 743 -1113 777
rect -1147 663 -1113 697
rect -1147 583 -1113 617
rect -847 743 -813 777
rect -847 663 -813 697
rect -847 583 -813 617
rect -517 743 -483 777
rect -517 663 -483 697
rect -517 583 -483 617
rect -1947 343 -1913 377
rect -1867 343 -1833 377
rect -1787 343 -1753 377
rect -1707 343 -1673 377
rect -1627 343 -1593 377
rect -1547 343 -1513 377
rect -1467 343 -1433 377
rect -1387 343 -1353 377
rect -1307 343 -1273 377
rect -1227 343 -1193 377
rect -1147 343 -1113 377
rect -1067 343 -1033 377
rect -987 343 -953 377
rect -907 343 -873 377
rect -827 343 -793 377
rect -747 343 -713 377
rect -667 343 -633 377
rect -587 343 -553 377
rect -507 343 -473 377
rect -427 343 -393 377
rect -347 343 -313 377
<< metal1 >>
rect -1970 1557 -290 1590
rect -1970 1523 -1947 1557
rect -1913 1523 -1867 1557
rect -1833 1523 -1787 1557
rect -1753 1523 -1707 1557
rect -1673 1523 -1627 1557
rect -1593 1523 -1547 1557
rect -1513 1523 -1467 1557
rect -1433 1523 -1387 1557
rect -1353 1523 -1307 1557
rect -1273 1523 -1227 1557
rect -1193 1523 -1147 1557
rect -1113 1523 -1067 1557
rect -1033 1523 -987 1557
rect -953 1523 -907 1557
rect -873 1523 -827 1557
rect -793 1523 -747 1557
rect -713 1523 -667 1557
rect -633 1523 -587 1557
rect -553 1523 -507 1557
rect -473 1523 -427 1557
rect -393 1523 -347 1557
rect -313 1523 -290 1557
rect -1970 1490 -290 1523
rect -1930 810 -1890 1490
rect -1470 1337 -1390 1490
rect -1620 1306 -1540 1320
rect -1620 1254 -1606 1306
rect -1554 1254 -1540 1306
rect -1620 1240 -1540 1254
rect -1470 1303 -1447 1337
rect -1413 1303 -1390 1337
rect -1470 1257 -1390 1303
rect -1470 1223 -1447 1257
rect -1413 1223 -1390 1257
rect -1620 1186 -1540 1200
rect -1620 1134 -1606 1186
rect -1554 1134 -1540 1186
rect -1620 1120 -1540 1134
rect -1470 1177 -1390 1223
rect -1470 1143 -1447 1177
rect -1413 1143 -1390 1177
rect -1470 1120 -1390 1143
rect -1170 1337 -1090 1490
rect -1170 1303 -1147 1337
rect -1113 1303 -1090 1337
rect -1170 1257 -1090 1303
rect -1170 1223 -1147 1257
rect -1113 1223 -1090 1257
rect -1170 1177 -1090 1223
rect -1170 1143 -1147 1177
rect -1113 1143 -1090 1177
rect -1170 1120 -1090 1143
rect -870 1337 -790 1490
rect -870 1303 -847 1337
rect -813 1303 -790 1337
rect -870 1257 -790 1303
rect -870 1223 -847 1257
rect -813 1223 -790 1257
rect -870 1177 -790 1223
rect -870 1143 -847 1177
rect -813 1143 -790 1177
rect -870 1120 -790 1143
rect -640 1186 -560 1200
rect -640 1134 -626 1186
rect -574 1134 -560 1186
rect -640 1120 -560 1134
rect -1120 1060 -1040 1080
rect -720 1060 -640 1080
rect -1120 1057 -640 1060
rect -1120 1023 -1097 1057
rect -1063 1023 -697 1057
rect -663 1023 -640 1057
rect -1120 1020 -640 1023
rect -1120 1000 -1040 1020
rect -720 1000 -640 1020
rect -520 810 -480 1490
rect -440 1306 -360 1320
rect -440 1254 -426 1306
rect -374 1254 -360 1306
rect -440 1240 -360 1254
rect -1950 777 -1870 810
rect -1950 743 -1927 777
rect -1893 743 -1870 777
rect -1950 697 -1870 743
rect -1950 663 -1927 697
rect -1893 663 -1870 697
rect -1950 617 -1870 663
rect -1950 583 -1927 617
rect -1893 583 -1870 617
rect -1950 560 -1870 583
rect -1470 777 -1390 810
rect -1470 743 -1447 777
rect -1413 743 -1390 777
rect -1470 697 -1390 743
rect -1470 663 -1447 697
rect -1413 663 -1390 697
rect -1470 617 -1390 663
rect -1470 583 -1447 617
rect -1413 583 -1390 617
rect -1470 560 -1390 583
rect -1170 777 -1090 810
rect -1170 743 -1147 777
rect -1113 743 -1090 777
rect -1170 697 -1090 743
rect -1170 663 -1147 697
rect -1113 663 -1090 697
rect -1170 617 -1090 663
rect -1170 583 -1147 617
rect -1113 583 -1090 617
rect -1170 560 -1090 583
rect -870 777 -790 810
rect -870 743 -847 777
rect -813 743 -790 777
rect -870 697 -790 743
rect -870 663 -847 697
rect -813 663 -790 697
rect -870 617 -790 663
rect -870 583 -847 617
rect -813 583 -790 617
rect -870 560 -790 583
rect -540 777 -460 810
rect -540 743 -517 777
rect -483 743 -460 777
rect -540 697 -460 743
rect -540 663 -517 697
rect -483 663 -460 697
rect -540 617 -460 663
rect -540 583 -517 617
rect -483 583 -460 617
rect -540 560 -460 583
rect -1450 410 -1410 560
rect -1150 410 -1110 560
rect -850 410 -810 560
rect -1970 377 -290 410
rect -1970 343 -1947 377
rect -1913 343 -1867 377
rect -1833 343 -1787 377
rect -1753 343 -1707 377
rect -1673 343 -1627 377
rect -1593 343 -1547 377
rect -1513 343 -1467 377
rect -1433 343 -1387 377
rect -1353 343 -1307 377
rect -1273 343 -1227 377
rect -1193 343 -1147 377
rect -1113 343 -1067 377
rect -1033 343 -987 377
rect -953 343 -907 377
rect -873 343 -827 377
rect -793 343 -747 377
rect -713 343 -667 377
rect -633 343 -587 377
rect -553 343 -507 377
rect -473 343 -427 377
rect -393 343 -347 377
rect -313 343 -290 377
rect -1970 310 -290 343
<< via1 >>
rect -1606 1297 -1554 1306
rect -1606 1263 -1597 1297
rect -1597 1263 -1563 1297
rect -1563 1263 -1554 1297
rect -1606 1254 -1554 1263
rect -1606 1177 -1554 1186
rect -1606 1143 -1597 1177
rect -1597 1143 -1563 1177
rect -1563 1143 -1554 1177
rect -1606 1134 -1554 1143
rect -626 1177 -574 1186
rect -626 1143 -617 1177
rect -617 1143 -583 1177
rect -583 1143 -574 1177
rect -626 1134 -574 1143
rect -426 1297 -374 1306
rect -426 1263 -417 1297
rect -417 1263 -383 1297
rect -383 1263 -374 1297
rect -426 1254 -374 1263
<< metal2 >>
rect -1620 1306 -1540 1320
rect -1620 1254 -1606 1306
rect -1554 1300 -1540 1306
rect -440 1306 -360 1320
rect -440 1300 -426 1306
rect -1554 1260 -426 1300
rect -1554 1254 -1540 1260
rect -1620 1240 -1540 1254
rect -440 1254 -426 1260
rect -374 1254 -360 1306
rect -440 1240 -360 1254
rect -1620 1186 -1540 1200
rect -1620 1134 -1606 1186
rect -1554 1180 -1540 1186
rect -640 1186 -560 1200
rect -640 1180 -626 1186
rect -1554 1140 -626 1180
rect -1554 1134 -1540 1140
rect -1620 1120 -1540 1134
rect -640 1134 -626 1140
rect -574 1134 -560 1186
rect -640 1120 -560 1134
<< labels >>
rlabel metal1 s -1100 1020 -1060 1060 4 OUT_bar
port 1 nsew
rlabel metal1 s -1150 340 -1110 380 4 GND!
port 2 nsew
rlabel metal1 s -1150 1520 -1110 1560 4 CLK
port 3 nsew
rlabel locali s -1200 895 -1160 935 4 OUT
port 4 nsew
rlabel locali s -1960 1270 -1940 1290 4 A
port 5 nsew
rlabel locali s -1960 950 -1940 970 4 A_bar
port 6 nsew
rlabel locali s -1960 1150 -1940 1170 4 B
port 7 nsew
rlabel locali s -1960 1050 -1940 1070 4 B_bar
port 8 nsew
rlabel locali s -1350 460 -1310 500 4 Dis
port 9 nsew
<< end >>
