magic
tech sky130A
timestamp 1679781200
<< metal2 >>
rect 0 0 30 30
rect 0 50 30 80
rect 0 100 30 130
rect 0 150 30 180
rect 0 200 30 230
rect 0 250 30 280
rect 0 300 30 330
rect 0 350 30 380
rect 0 400 30 430
rect 0 450 30 480
rect 0 500 30 530
rect 0 550 30 580
rect 0 600 30 630
rect 0 650 30 680
rect 0 700 30 730
rect 0 750 30 780
rect 0 800 30 830
rect 0 850 30 880
rect 0 900 30 930
rect 0 950 30 980
rect 0 1000 30 1030
rect 0 1050 30 1080
rect 0 1100 30 1130
rect 0 1150 30 1180
rect 0 1200 30 1230
rect 0 1250 30 1280
rect 0 1300 30 1330
rect 0 1350 30 1380
rect 0 1400 30 1430
rect 0 1450 30 1480
rect 0 1500 30 1530
rect 0 1550 30 1580
rect 0 1600 30 1630
rect 0 1650 30 1680
rect 0 1700 30 1730
rect 0 1750 30 1780
rect 0 1800 30 1830
rect 0 1850 30 1880
rect 0 1900 30 1930
rect 0 1950 30 1980
rect 0 2000 30 2030
rect 0 2050 30 2080
rect 0 2100 30 2130
rect 0 2150 30 2180
rect 0 2200 30 2230
rect 0 2250 30 2280
rect 0 2300 30 2330
rect 0 2350 30 2380
rect 0 2400 30 2430
rect 0 2450 30 2480
rect 0 2500 30 2530
rect 0 2550 30 2580
rect 0 2600 30 2630
rect 0 2650 30 2680
rect 0 2700 30 2730
rect 0 2750 30 2780
rect 0 2800 30 2830
rect 0 2850 30 2880
rect 0 2900 30 2930
rect 0 2950 30 2980
rect 0 3000 30 3030
rect 0 3050 30 3080
rect 0 3100 30 3130
rect 0 3150 30 3180
<< labels >>
rlabel metal2 0 0 30 30 1 s0_bar
port 0 n
rlabel metal2 0 50 30 80 1 s1_bar
port 1 n
rlabel metal2 0 100 30 130 1 s2_bar
port 2 n
rlabel metal2 0 150 30 180 1 s3_bar
port 3 n
rlabel metal2 0 200 30 230 1 s4_bar
port 4 n
rlabel metal2 0 250 30 280 1 s5_bar
port 5 n
rlabel metal2 0 300 30 330 1 s6_bar
port 6 n
rlabel metal2 0 350 30 380 1 s7_bar
port 7 n
rlabel metal2 0 400 30 430 1 s8_bar
port 8 n
rlabel metal2 0 450 30 480 1 s9_bar
port 9 n
rlabel metal2 0 500 30 530 1 s10_bar
port 10 n
rlabel metal2 0 550 30 580 1 s11_bar
port 11 n
rlabel metal2 0 600 30 630 1 s12_bar
port 12 n
rlabel metal2 0 650 30 680 1 s13_bar
port 13 n
rlabel metal2 0 700 30 730 1 s14_bar
port 14 n
rlabel metal2 0 750 30 780 1 s15_bar
port 15 n
rlabel metal2 0 800 30 830 1 s16_bar
port 16 n
rlabel metal2 0 850 30 880 1 s17_bar
port 17 n
rlabel metal2 0 900 30 930 1 s18_bar
port 18 n
rlabel metal2 0 950 30 980 1 s19_bar
port 19 n
rlabel metal2 0 1000 30 1030 1 s20_bar
port 20 n
rlabel metal2 0 1050 30 1080 1 s21_bar
port 21 n
rlabel metal2 0 1100 30 1130 1 s22_bar
port 22 n
rlabel metal2 0 1150 30 1180 1 s23_bar
port 23 n
rlabel metal2 0 1200 30 1230 1 s24_bar
port 24 n
rlabel metal2 0 1250 30 1280 1 s25_bar
port 25 n
rlabel metal2 0 1300 30 1330 1 s26_bar
port 26 n
rlabel metal2 0 1350 30 1380 1 s27_bar
port 27 n
rlabel metal2 0 1400 30 1430 1 s28_bar
port 28 n
rlabel metal2 0 1450 30 1480 1 s29_bar
port 29 n
rlabel metal2 0 1500 30 1530 1 s30_bar
port 30 n
rlabel metal2 0 1550 30 1580 1 s31_bar
port 31 n
rlabel metal2 0 1600 30 1630 1 s32_bar
port 32 n
rlabel metal2 0 1650 30 1680 1 s33_bar
port 33 n
rlabel metal2 0 1700 30 1730 1 s34_bar
port 34 n
rlabel metal2 0 1750 30 1780 1 s35_bar
port 35 n
rlabel metal2 0 1800 30 1830 1 s36_bar
port 36 n
rlabel metal2 0 1850 30 1880 1 s37_bar
port 37 n
rlabel metal2 0 1900 30 1930 1 s38_bar
port 38 n
rlabel metal2 0 1950 30 1980 1 s39_bar
port 39 n
rlabel metal2 0 2000 30 2030 1 s40_bar
port 40 n
rlabel metal2 0 2050 30 2080 1 s41_bar
port 41 n
rlabel metal2 0 2100 30 2130 1 s42_bar
port 42 n
rlabel metal2 0 2150 30 2180 1 s43_bar
port 43 n
rlabel metal2 0 2200 30 2230 1 s44_bar
port 44 n
rlabel metal2 0 2250 30 2280 1 s45_bar
port 45 n
rlabel metal2 0 2300 30 2330 1 s46_bar
port 46 n
rlabel metal2 0 2350 30 2380 1 s47_bar
port 47 n
rlabel metal2 0 2400 30 2430 1 s48_bar
port 48 n
rlabel metal2 0 2450 30 2480 1 s49_bar
port 49 n
rlabel metal2 0 2500 30 2530 1 s50_bar
port 50 n
rlabel metal2 0 2550 30 2580 1 s51_bar
port 51 n
rlabel metal2 0 2600 30 2630 1 s52_bar
port 52 n
rlabel metal2 0 2650 30 2680 1 s53_bar
port 53 n
rlabel metal2 0 2700 30 2730 1 s54_bar
port 54 n
rlabel metal2 0 2750 30 2780 1 s55_bar
port 55 n
rlabel metal2 0 2800 30 2830 1 s56_bar
port 56 n
rlabel metal2 0 2850 30 2880 1 s57_bar
port 57 n
rlabel metal2 0 2900 30 2930 1 s58_bar
port 58 n
rlabel metal2 0 2950 30 2980 1 s59_bar
port 59 n
rlabel metal2 0 3000 30 3030 1 s60_bar
port 60 n
rlabel metal2 0 3050 30 3080 1 s61_bar
port 61 n
rlabel metal2 0 3100 30 3130 1 s62_bar
port 62 n
rlabel metal2 0 3150 30 3180 1 s63_bar
port 63 n
<< end >>
