magic
tech sky130A
magscale 1 2
timestamp 1671080676
<< poly >>
rect -421 1107 1219 1157
<< locali >>
rect -561 127 -521 1037
rect 1319 127 1359 1037
use pmos_1v8_lvt_4p75_Lbody_4finger  pmos_1v8_lvt_4p75_Lbody_4finger_0
timestamp 1671080676
transform 1 0 -511 0 1 -273
box -242 245 1178 1505
use pmos_1v8_lvt_4p75_Rbody_4finger  pmos_1v8_lvt_4p75_Rbody_4finger_0
timestamp 1671080676
transform 1 0 369 0 1 -273
box -240 245 1180 1505
<< properties >>
string path -2.105 5.660 6.095 5.660 
<< end >>
