magic
tech sky130A
magscale 1 2
timestamp 1675193052
<< nwell >>
rect -3910 967 -1550 1157
rect -1290 967 200 1157
rect 460 967 2220 1157
rect -3140 577 -2320 967
rect -950 577 -130 967
rect 930 577 1750 967
rect -3140 -1213 -2320 -823
rect -950 -1213 -130 -823
rect 930 -1213 1750 -823
rect -3910 -1403 -1550 -1213
rect -1290 -1403 200 -1213
rect 460 -1403 2220 -1213
rect -3769 -1853 -1689 -1663
rect -1429 -1853 61 -1663
rect -3139 -2243 -2319 -1853
rect -1089 -2243 -269 -1853
rect 321 -1854 2401 -1664
rect 951 -2244 1771 -1854
<< pwell >>
rect -3896 -639 -1564 393
rect -1256 -639 176 393
rect 474 -639 2206 393
rect -3745 -2867 -1713 -2427
rect -3755 -3019 -1703 -2867
rect -1395 -3019 37 -2427
rect 345 -2868 2377 -2428
rect 335 -3020 2387 -2868
<< nmos >>
rect -3750 67 -3720 367
rect -3600 67 -3570 367
rect -3450 67 -3420 367
rect -3300 67 -3270 367
rect -2970 67 -2940 367
rect -2820 67 -2790 367
rect -2670 67 -2640 367
rect -2520 67 -2490 367
rect -2190 67 -2160 367
rect -2040 67 -2010 367
rect -1890 67 -1860 367
rect -1740 67 -1710 367
rect -1110 67 -1080 367
rect -780 67 -750 367
rect -630 67 -600 367
rect -480 67 -450 367
rect -330 67 -300 367
rect 0 67 30 367
rect 620 67 650 367
rect 770 67 800 367
rect 1100 67 1130 367
rect 1250 67 1280 367
rect 1400 67 1430 367
rect 1550 67 1580 367
rect 1880 67 1910 367
rect 2030 67 2060 367
rect -3750 -613 -3720 -313
rect -3600 -613 -3570 -313
rect -3450 -613 -3420 -313
rect -3300 -613 -3270 -313
rect -2970 -613 -2940 -313
rect -2820 -613 -2790 -313
rect -2670 -613 -2640 -313
rect -2520 -613 -2490 -313
rect -2190 -613 -2160 -313
rect -2040 -613 -2010 -313
rect -1890 -613 -1860 -313
rect -1740 -613 -1710 -313
rect -1110 -613 -1080 -313
rect -780 -613 -750 -313
rect -630 -613 -600 -313
rect -480 -613 -450 -313
rect -330 -613 -300 -313
rect 0 -613 30 -313
rect 620 -613 650 -313
rect 770 -613 800 -313
rect 1100 -613 1130 -313
rect 1250 -613 1280 -313
rect 1400 -613 1430 -313
rect 1550 -613 1580 -313
rect 1880 -613 1910 -313
rect 2030 -613 2060 -313
rect -3599 -2753 -3569 -2453
rect -3449 -2753 -3419 -2453
rect -3299 -2753 -3269 -2453
rect -2969 -2753 -2939 -2453
rect -2819 -2753 -2789 -2453
rect -2669 -2753 -2639 -2453
rect -2519 -2753 -2489 -2453
rect -2189 -2753 -2159 -2453
rect -2039 -2753 -2009 -2453
rect -1889 -2753 -1859 -2453
rect -1249 -2753 -1219 -2453
rect -919 -2753 -889 -2453
rect -769 -2753 -739 -2453
rect -619 -2753 -589 -2453
rect -469 -2753 -439 -2453
rect -139 -2753 -109 -2453
rect 491 -2754 521 -2454
rect 641 -2754 671 -2454
rect 791 -2754 821 -2454
rect 1121 -2754 1151 -2454
rect 1271 -2754 1301 -2454
rect 1421 -2754 1451 -2454
rect 1571 -2754 1601 -2454
rect 1901 -2754 1931 -2454
rect 2051 -2754 2081 -2454
rect 2201 -2754 2231 -2454
<< pmos >>
rect -2970 627 -2940 927
rect -2820 627 -2790 927
rect -2670 627 -2640 927
rect -2520 627 -2490 927
rect -780 627 -750 927
rect -630 627 -600 927
rect -480 627 -450 927
rect -330 627 -300 927
rect 1100 627 1130 927
rect 1250 627 1280 927
rect 1400 627 1430 927
rect 1550 627 1580 927
rect -2970 -1173 -2940 -873
rect -2820 -1173 -2790 -873
rect -2670 -1173 -2640 -873
rect -2520 -1173 -2490 -873
rect -780 -1173 -750 -873
rect -630 -1173 -600 -873
rect -480 -1173 -450 -873
rect -330 -1173 -300 -873
rect 1100 -1173 1130 -873
rect 1250 -1173 1280 -873
rect 1400 -1173 1430 -873
rect 1550 -1173 1580 -873
rect -2969 -2193 -2939 -1893
rect -2819 -2193 -2789 -1893
rect -2669 -2193 -2639 -1893
rect -2519 -2193 -2489 -1893
rect -919 -2193 -889 -1893
rect -769 -2193 -739 -1893
rect -619 -2193 -589 -1893
rect -469 -2193 -439 -1893
rect 1121 -2194 1151 -1894
rect 1271 -2194 1301 -1894
rect 1421 -2194 1451 -1894
rect 1571 -2194 1601 -1894
<< ndiff >>
rect -3870 294 -3750 367
rect -3870 260 -3827 294
rect -3793 260 -3750 294
rect -3870 214 -3750 260
rect -3870 180 -3827 214
rect -3793 180 -3750 214
rect -3870 134 -3750 180
rect -3870 100 -3827 134
rect -3793 100 -3750 134
rect -3870 67 -3750 100
rect -3720 67 -3600 367
rect -3570 294 -3450 367
rect -3570 260 -3527 294
rect -3493 260 -3450 294
rect -3570 214 -3450 260
rect -3570 180 -3527 214
rect -3493 180 -3450 214
rect -3570 134 -3450 180
rect -3570 100 -3527 134
rect -3493 100 -3450 134
rect -3570 67 -3450 100
rect -3420 67 -3300 367
rect -3270 294 -3150 367
rect -3270 260 -3227 294
rect -3193 260 -3150 294
rect -3270 214 -3150 260
rect -3270 180 -3227 214
rect -3193 180 -3150 214
rect -3270 134 -3150 180
rect -3270 100 -3227 134
rect -3193 100 -3150 134
rect -3270 67 -3150 100
rect -3090 294 -2970 367
rect -3090 260 -3047 294
rect -3013 260 -2970 294
rect -3090 214 -2970 260
rect -3090 180 -3047 214
rect -3013 180 -2970 214
rect -3090 134 -2970 180
rect -3090 100 -3047 134
rect -3013 100 -2970 134
rect -3090 67 -2970 100
rect -2940 294 -2820 367
rect -2940 260 -2897 294
rect -2863 260 -2820 294
rect -2940 214 -2820 260
rect -2940 180 -2897 214
rect -2863 180 -2820 214
rect -2940 134 -2820 180
rect -2940 100 -2897 134
rect -2863 100 -2820 134
rect -2940 67 -2820 100
rect -2790 294 -2670 367
rect -2790 260 -2747 294
rect -2713 260 -2670 294
rect -2790 214 -2670 260
rect -2790 180 -2747 214
rect -2713 180 -2670 214
rect -2790 134 -2670 180
rect -2790 100 -2747 134
rect -2713 100 -2670 134
rect -2790 67 -2670 100
rect -2640 294 -2520 367
rect -2640 260 -2597 294
rect -2563 260 -2520 294
rect -2640 214 -2520 260
rect -2640 180 -2597 214
rect -2563 180 -2520 214
rect -2640 134 -2520 180
rect -2640 100 -2597 134
rect -2563 100 -2520 134
rect -2640 67 -2520 100
rect -2490 294 -2370 367
rect -2490 260 -2447 294
rect -2413 260 -2370 294
rect -2490 214 -2370 260
rect -2490 180 -2447 214
rect -2413 180 -2370 214
rect -2490 134 -2370 180
rect -2490 100 -2447 134
rect -2413 100 -2370 134
rect -2490 67 -2370 100
rect -2310 294 -2190 367
rect -2310 260 -2267 294
rect -2233 260 -2190 294
rect -2310 214 -2190 260
rect -2310 180 -2267 214
rect -2233 180 -2190 214
rect -2310 134 -2190 180
rect -2310 100 -2267 134
rect -2233 100 -2190 134
rect -2310 67 -2190 100
rect -2160 67 -2040 367
rect -2010 294 -1890 367
rect -2010 260 -1967 294
rect -1933 260 -1890 294
rect -2010 214 -1890 260
rect -2010 180 -1967 214
rect -1933 180 -1890 214
rect -2010 134 -1890 180
rect -2010 100 -1967 134
rect -1933 100 -1890 134
rect -2010 67 -1890 100
rect -1860 67 -1740 367
rect -1710 294 -1590 367
rect -1710 260 -1667 294
rect -1633 260 -1590 294
rect -1710 214 -1590 260
rect -1710 180 -1667 214
rect -1633 180 -1590 214
rect -1710 134 -1590 180
rect -1710 100 -1667 134
rect -1633 100 -1590 134
rect -1710 67 -1590 100
rect -1230 294 -1110 367
rect -1230 260 -1187 294
rect -1153 260 -1110 294
rect -1230 214 -1110 260
rect -1230 180 -1187 214
rect -1153 180 -1110 214
rect -1230 134 -1110 180
rect -1230 100 -1187 134
rect -1153 100 -1110 134
rect -1230 67 -1110 100
rect -1080 294 -960 367
rect -1080 260 -1037 294
rect -1003 260 -960 294
rect -1080 214 -960 260
rect -1080 180 -1037 214
rect -1003 180 -960 214
rect -1080 134 -960 180
rect -1080 100 -1037 134
rect -1003 100 -960 134
rect -1080 67 -960 100
rect -900 294 -780 367
rect -900 260 -857 294
rect -823 260 -780 294
rect -900 214 -780 260
rect -900 180 -857 214
rect -823 180 -780 214
rect -900 134 -780 180
rect -900 100 -857 134
rect -823 100 -780 134
rect -900 67 -780 100
rect -750 294 -630 367
rect -750 260 -707 294
rect -673 260 -630 294
rect -750 214 -630 260
rect -750 180 -707 214
rect -673 180 -630 214
rect -750 134 -630 180
rect -750 100 -707 134
rect -673 100 -630 134
rect -750 67 -630 100
rect -600 294 -480 367
rect -600 260 -557 294
rect -523 260 -480 294
rect -600 214 -480 260
rect -600 180 -557 214
rect -523 180 -480 214
rect -600 134 -480 180
rect -600 100 -557 134
rect -523 100 -480 134
rect -600 67 -480 100
rect -450 294 -330 367
rect -450 260 -407 294
rect -373 260 -330 294
rect -450 214 -330 260
rect -450 180 -407 214
rect -373 180 -330 214
rect -450 134 -330 180
rect -450 100 -407 134
rect -373 100 -330 134
rect -450 67 -330 100
rect -300 294 -180 367
rect -300 260 -257 294
rect -223 260 -180 294
rect -300 214 -180 260
rect -300 180 -257 214
rect -223 180 -180 214
rect -300 134 -180 180
rect -300 100 -257 134
rect -223 100 -180 134
rect -300 67 -180 100
rect -120 294 0 367
rect -120 260 -77 294
rect -43 260 0 294
rect -120 214 0 260
rect -120 180 -77 214
rect -43 180 0 214
rect -120 134 0 180
rect -120 100 -77 134
rect -43 100 0 134
rect -120 67 0 100
rect 30 294 150 367
rect 30 260 73 294
rect 107 260 150 294
rect 30 214 150 260
rect 30 180 73 214
rect 107 180 150 214
rect 30 134 150 180
rect 30 100 73 134
rect 107 100 150 134
rect 30 67 150 100
rect 500 294 620 367
rect 500 260 543 294
rect 577 260 620 294
rect 500 214 620 260
rect 500 180 543 214
rect 577 180 620 214
rect 500 134 620 180
rect 500 100 543 134
rect 577 100 620 134
rect 500 67 620 100
rect 650 294 770 367
rect 650 260 693 294
rect 727 260 770 294
rect 650 214 770 260
rect 650 180 693 214
rect 727 180 770 214
rect 650 134 770 180
rect 650 100 693 134
rect 727 100 770 134
rect 650 67 770 100
rect 800 294 920 367
rect 800 260 843 294
rect 877 260 920 294
rect 800 214 920 260
rect 800 180 843 214
rect 877 180 920 214
rect 800 134 920 180
rect 800 100 843 134
rect 877 100 920 134
rect 800 67 920 100
rect 980 294 1100 367
rect 980 260 1023 294
rect 1057 260 1100 294
rect 980 214 1100 260
rect 980 180 1023 214
rect 1057 180 1100 214
rect 980 134 1100 180
rect 980 100 1023 134
rect 1057 100 1100 134
rect 980 67 1100 100
rect 1130 294 1250 367
rect 1130 260 1173 294
rect 1207 260 1250 294
rect 1130 214 1250 260
rect 1130 180 1173 214
rect 1207 180 1250 214
rect 1130 134 1250 180
rect 1130 100 1173 134
rect 1207 100 1250 134
rect 1130 67 1250 100
rect 1280 294 1400 367
rect 1280 260 1323 294
rect 1357 260 1400 294
rect 1280 214 1400 260
rect 1280 180 1323 214
rect 1357 180 1400 214
rect 1280 134 1400 180
rect 1280 100 1323 134
rect 1357 100 1400 134
rect 1280 67 1400 100
rect 1430 294 1550 367
rect 1430 260 1473 294
rect 1507 260 1550 294
rect 1430 214 1550 260
rect 1430 180 1473 214
rect 1507 180 1550 214
rect 1430 134 1550 180
rect 1430 100 1473 134
rect 1507 100 1550 134
rect 1430 67 1550 100
rect 1580 294 1700 367
rect 1580 260 1623 294
rect 1657 260 1700 294
rect 1580 214 1700 260
rect 1580 180 1623 214
rect 1657 180 1700 214
rect 1580 134 1700 180
rect 1580 100 1623 134
rect 1657 100 1700 134
rect 1580 67 1700 100
rect 1760 294 1880 367
rect 1760 260 1803 294
rect 1837 260 1880 294
rect 1760 214 1880 260
rect 1760 180 1803 214
rect 1837 180 1880 214
rect 1760 134 1880 180
rect 1760 100 1803 134
rect 1837 100 1880 134
rect 1760 67 1880 100
rect 1910 67 2030 367
rect 2060 294 2180 367
rect 2060 260 2103 294
rect 2137 260 2180 294
rect 2060 214 2180 260
rect 2060 180 2103 214
rect 2137 180 2180 214
rect 2060 134 2180 180
rect 2060 100 2103 134
rect 2137 100 2180 134
rect 2060 67 2180 100
rect -3870 -346 -3750 -313
rect -3870 -380 -3827 -346
rect -3793 -380 -3750 -346
rect -3870 -426 -3750 -380
rect -3870 -460 -3827 -426
rect -3793 -460 -3750 -426
rect -3870 -506 -3750 -460
rect -3870 -540 -3827 -506
rect -3793 -540 -3750 -506
rect -3870 -613 -3750 -540
rect -3720 -613 -3600 -313
rect -3570 -346 -3450 -313
rect -3570 -380 -3527 -346
rect -3493 -380 -3450 -346
rect -3570 -426 -3450 -380
rect -3570 -460 -3527 -426
rect -3493 -460 -3450 -426
rect -3570 -506 -3450 -460
rect -3570 -540 -3527 -506
rect -3493 -540 -3450 -506
rect -3570 -613 -3450 -540
rect -3420 -613 -3300 -313
rect -3270 -346 -3150 -313
rect -3270 -380 -3227 -346
rect -3193 -380 -3150 -346
rect -3270 -426 -3150 -380
rect -3270 -460 -3227 -426
rect -3193 -460 -3150 -426
rect -3270 -506 -3150 -460
rect -3270 -540 -3227 -506
rect -3193 -540 -3150 -506
rect -3270 -613 -3150 -540
rect -3090 -346 -2970 -313
rect -3090 -380 -3047 -346
rect -3013 -380 -2970 -346
rect -3090 -426 -2970 -380
rect -3090 -460 -3047 -426
rect -3013 -460 -2970 -426
rect -3090 -506 -2970 -460
rect -3090 -540 -3047 -506
rect -3013 -540 -2970 -506
rect -3090 -613 -2970 -540
rect -2940 -346 -2820 -313
rect -2940 -380 -2897 -346
rect -2863 -380 -2820 -346
rect -2940 -426 -2820 -380
rect -2940 -460 -2897 -426
rect -2863 -460 -2820 -426
rect -2940 -506 -2820 -460
rect -2940 -540 -2897 -506
rect -2863 -540 -2820 -506
rect -2940 -613 -2820 -540
rect -2790 -346 -2670 -313
rect -2790 -380 -2747 -346
rect -2713 -380 -2670 -346
rect -2790 -426 -2670 -380
rect -2790 -460 -2747 -426
rect -2713 -460 -2670 -426
rect -2790 -506 -2670 -460
rect -2790 -540 -2747 -506
rect -2713 -540 -2670 -506
rect -2790 -613 -2670 -540
rect -2640 -346 -2520 -313
rect -2640 -380 -2597 -346
rect -2563 -380 -2520 -346
rect -2640 -426 -2520 -380
rect -2640 -460 -2597 -426
rect -2563 -460 -2520 -426
rect -2640 -506 -2520 -460
rect -2640 -540 -2597 -506
rect -2563 -540 -2520 -506
rect -2640 -613 -2520 -540
rect -2490 -346 -2370 -313
rect -2490 -380 -2447 -346
rect -2413 -380 -2370 -346
rect -2490 -426 -2370 -380
rect -2490 -460 -2447 -426
rect -2413 -460 -2370 -426
rect -2490 -506 -2370 -460
rect -2490 -540 -2447 -506
rect -2413 -540 -2370 -506
rect -2490 -613 -2370 -540
rect -2310 -346 -2190 -313
rect -2310 -380 -2267 -346
rect -2233 -380 -2190 -346
rect -2310 -426 -2190 -380
rect -2310 -460 -2267 -426
rect -2233 -460 -2190 -426
rect -2310 -506 -2190 -460
rect -2310 -540 -2267 -506
rect -2233 -540 -2190 -506
rect -2310 -613 -2190 -540
rect -2160 -613 -2040 -313
rect -2010 -346 -1890 -313
rect -2010 -380 -1967 -346
rect -1933 -380 -1890 -346
rect -2010 -426 -1890 -380
rect -2010 -460 -1967 -426
rect -1933 -460 -1890 -426
rect -2010 -506 -1890 -460
rect -2010 -540 -1967 -506
rect -1933 -540 -1890 -506
rect -2010 -613 -1890 -540
rect -1860 -613 -1740 -313
rect -1710 -346 -1590 -313
rect -1710 -380 -1667 -346
rect -1633 -380 -1590 -346
rect -1710 -426 -1590 -380
rect -1710 -460 -1667 -426
rect -1633 -460 -1590 -426
rect -1710 -506 -1590 -460
rect -1710 -540 -1667 -506
rect -1633 -540 -1590 -506
rect -1710 -613 -1590 -540
rect -1230 -346 -1110 -313
rect -1230 -380 -1187 -346
rect -1153 -380 -1110 -346
rect -1230 -426 -1110 -380
rect -1230 -460 -1187 -426
rect -1153 -460 -1110 -426
rect -1230 -506 -1110 -460
rect -1230 -540 -1187 -506
rect -1153 -540 -1110 -506
rect -1230 -613 -1110 -540
rect -1080 -346 -960 -313
rect -1080 -380 -1037 -346
rect -1003 -380 -960 -346
rect -1080 -426 -960 -380
rect -1080 -460 -1037 -426
rect -1003 -460 -960 -426
rect -1080 -506 -960 -460
rect -1080 -540 -1037 -506
rect -1003 -540 -960 -506
rect -1080 -613 -960 -540
rect -900 -346 -780 -313
rect -900 -380 -857 -346
rect -823 -380 -780 -346
rect -900 -426 -780 -380
rect -900 -460 -857 -426
rect -823 -460 -780 -426
rect -900 -506 -780 -460
rect -900 -540 -857 -506
rect -823 -540 -780 -506
rect -900 -613 -780 -540
rect -750 -346 -630 -313
rect -750 -380 -707 -346
rect -673 -380 -630 -346
rect -750 -426 -630 -380
rect -750 -460 -707 -426
rect -673 -460 -630 -426
rect -750 -506 -630 -460
rect -750 -540 -707 -506
rect -673 -540 -630 -506
rect -750 -613 -630 -540
rect -600 -346 -480 -313
rect -600 -380 -557 -346
rect -523 -380 -480 -346
rect -600 -426 -480 -380
rect -600 -460 -557 -426
rect -523 -460 -480 -426
rect -600 -506 -480 -460
rect -600 -540 -557 -506
rect -523 -540 -480 -506
rect -600 -613 -480 -540
rect -450 -346 -330 -313
rect -450 -380 -407 -346
rect -373 -380 -330 -346
rect -450 -426 -330 -380
rect -450 -460 -407 -426
rect -373 -460 -330 -426
rect -450 -506 -330 -460
rect -450 -540 -407 -506
rect -373 -540 -330 -506
rect -450 -613 -330 -540
rect -300 -346 -180 -313
rect -300 -380 -257 -346
rect -223 -380 -180 -346
rect -300 -426 -180 -380
rect -300 -460 -257 -426
rect -223 -460 -180 -426
rect -300 -506 -180 -460
rect -300 -540 -257 -506
rect -223 -540 -180 -506
rect -300 -613 -180 -540
rect -120 -346 0 -313
rect -120 -380 -77 -346
rect -43 -380 0 -346
rect -120 -426 0 -380
rect -120 -460 -77 -426
rect -43 -460 0 -426
rect -120 -506 0 -460
rect -120 -540 -77 -506
rect -43 -540 0 -506
rect -120 -613 0 -540
rect 30 -346 150 -313
rect 30 -380 73 -346
rect 107 -380 150 -346
rect 30 -426 150 -380
rect 30 -460 73 -426
rect 107 -460 150 -426
rect 30 -506 150 -460
rect 30 -540 73 -506
rect 107 -540 150 -506
rect 30 -613 150 -540
rect 500 -346 620 -313
rect 500 -380 543 -346
rect 577 -380 620 -346
rect 500 -426 620 -380
rect 500 -460 543 -426
rect 577 -460 620 -426
rect 500 -506 620 -460
rect 500 -540 543 -506
rect 577 -540 620 -506
rect 500 -613 620 -540
rect 650 -346 770 -313
rect 650 -380 693 -346
rect 727 -380 770 -346
rect 650 -426 770 -380
rect 650 -460 693 -426
rect 727 -460 770 -426
rect 650 -506 770 -460
rect 650 -540 693 -506
rect 727 -540 770 -506
rect 650 -613 770 -540
rect 800 -346 920 -313
rect 800 -380 843 -346
rect 877 -380 920 -346
rect 800 -426 920 -380
rect 800 -460 843 -426
rect 877 -460 920 -426
rect 800 -506 920 -460
rect 800 -540 843 -506
rect 877 -540 920 -506
rect 800 -613 920 -540
rect 980 -346 1100 -313
rect 980 -380 1023 -346
rect 1057 -380 1100 -346
rect 980 -426 1100 -380
rect 980 -460 1023 -426
rect 1057 -460 1100 -426
rect 980 -506 1100 -460
rect 980 -540 1023 -506
rect 1057 -540 1100 -506
rect 980 -613 1100 -540
rect 1130 -346 1250 -313
rect 1130 -380 1173 -346
rect 1207 -380 1250 -346
rect 1130 -426 1250 -380
rect 1130 -460 1173 -426
rect 1207 -460 1250 -426
rect 1130 -506 1250 -460
rect 1130 -540 1173 -506
rect 1207 -540 1250 -506
rect 1130 -613 1250 -540
rect 1280 -346 1400 -313
rect 1280 -380 1323 -346
rect 1357 -380 1400 -346
rect 1280 -426 1400 -380
rect 1280 -460 1323 -426
rect 1357 -460 1400 -426
rect 1280 -506 1400 -460
rect 1280 -540 1323 -506
rect 1357 -540 1400 -506
rect 1280 -613 1400 -540
rect 1430 -346 1550 -313
rect 1430 -380 1473 -346
rect 1507 -380 1550 -346
rect 1430 -426 1550 -380
rect 1430 -460 1473 -426
rect 1507 -460 1550 -426
rect 1430 -506 1550 -460
rect 1430 -540 1473 -506
rect 1507 -540 1550 -506
rect 1430 -613 1550 -540
rect 1580 -346 1700 -313
rect 1580 -380 1623 -346
rect 1657 -380 1700 -346
rect 1580 -426 1700 -380
rect 1580 -460 1623 -426
rect 1657 -460 1700 -426
rect 1580 -506 1700 -460
rect 1580 -540 1623 -506
rect 1657 -540 1700 -506
rect 1580 -613 1700 -540
rect 1760 -346 1880 -313
rect 1760 -380 1803 -346
rect 1837 -380 1880 -346
rect 1760 -426 1880 -380
rect 1760 -460 1803 -426
rect 1837 -460 1880 -426
rect 1760 -506 1880 -460
rect 1760 -540 1803 -506
rect 1837 -540 1880 -506
rect 1760 -613 1880 -540
rect 1910 -613 2030 -313
rect 2060 -346 2180 -313
rect 2060 -380 2103 -346
rect 2137 -380 2180 -346
rect 2060 -426 2180 -380
rect 2060 -460 2103 -426
rect 2137 -460 2180 -426
rect 2060 -506 2180 -460
rect 2060 -540 2103 -506
rect 2137 -540 2180 -506
rect 2060 -613 2180 -540
rect -3719 -2526 -3599 -2453
rect -3719 -2560 -3676 -2526
rect -3642 -2560 -3599 -2526
rect -3719 -2606 -3599 -2560
rect -3719 -2640 -3676 -2606
rect -3642 -2640 -3599 -2606
rect -3719 -2686 -3599 -2640
rect -3719 -2720 -3676 -2686
rect -3642 -2720 -3599 -2686
rect -3719 -2753 -3599 -2720
rect -3569 -2526 -3449 -2453
rect -3569 -2560 -3526 -2526
rect -3492 -2560 -3449 -2526
rect -3569 -2606 -3449 -2560
rect -3569 -2640 -3526 -2606
rect -3492 -2640 -3449 -2606
rect -3569 -2686 -3449 -2640
rect -3569 -2720 -3526 -2686
rect -3492 -2720 -3449 -2686
rect -3569 -2753 -3449 -2720
rect -3419 -2526 -3299 -2453
rect -3419 -2560 -3376 -2526
rect -3342 -2560 -3299 -2526
rect -3419 -2606 -3299 -2560
rect -3419 -2640 -3376 -2606
rect -3342 -2640 -3299 -2606
rect -3419 -2686 -3299 -2640
rect -3419 -2720 -3376 -2686
rect -3342 -2720 -3299 -2686
rect -3419 -2753 -3299 -2720
rect -3269 -2526 -3149 -2453
rect -3269 -2560 -3226 -2526
rect -3192 -2560 -3149 -2526
rect -3269 -2606 -3149 -2560
rect -3269 -2640 -3226 -2606
rect -3192 -2640 -3149 -2606
rect -3269 -2686 -3149 -2640
rect -3269 -2720 -3226 -2686
rect -3192 -2720 -3149 -2686
rect -3269 -2753 -3149 -2720
rect -3089 -2526 -2969 -2453
rect -3089 -2560 -3046 -2526
rect -3012 -2560 -2969 -2526
rect -3089 -2606 -2969 -2560
rect -3089 -2640 -3046 -2606
rect -3012 -2640 -2969 -2606
rect -3089 -2686 -2969 -2640
rect -3089 -2720 -3046 -2686
rect -3012 -2720 -2969 -2686
rect -3089 -2753 -2969 -2720
rect -2939 -2526 -2819 -2453
rect -2939 -2560 -2896 -2526
rect -2862 -2560 -2819 -2526
rect -2939 -2606 -2819 -2560
rect -2939 -2640 -2896 -2606
rect -2862 -2640 -2819 -2606
rect -2939 -2686 -2819 -2640
rect -2939 -2720 -2896 -2686
rect -2862 -2720 -2819 -2686
rect -2939 -2753 -2819 -2720
rect -2789 -2526 -2669 -2453
rect -2789 -2560 -2746 -2526
rect -2712 -2560 -2669 -2526
rect -2789 -2606 -2669 -2560
rect -2789 -2640 -2746 -2606
rect -2712 -2640 -2669 -2606
rect -2789 -2686 -2669 -2640
rect -2789 -2720 -2746 -2686
rect -2712 -2720 -2669 -2686
rect -2789 -2753 -2669 -2720
rect -2639 -2526 -2519 -2453
rect -2639 -2560 -2596 -2526
rect -2562 -2560 -2519 -2526
rect -2639 -2606 -2519 -2560
rect -2639 -2640 -2596 -2606
rect -2562 -2640 -2519 -2606
rect -2639 -2686 -2519 -2640
rect -2639 -2720 -2596 -2686
rect -2562 -2720 -2519 -2686
rect -2639 -2753 -2519 -2720
rect -2489 -2526 -2369 -2453
rect -2489 -2560 -2446 -2526
rect -2412 -2560 -2369 -2526
rect -2489 -2606 -2369 -2560
rect -2489 -2640 -2446 -2606
rect -2412 -2640 -2369 -2606
rect -2489 -2686 -2369 -2640
rect -2489 -2720 -2446 -2686
rect -2412 -2720 -2369 -2686
rect -2489 -2753 -2369 -2720
rect -2309 -2526 -2189 -2453
rect -2309 -2560 -2266 -2526
rect -2232 -2560 -2189 -2526
rect -2309 -2606 -2189 -2560
rect -2309 -2640 -2266 -2606
rect -2232 -2640 -2189 -2606
rect -2309 -2686 -2189 -2640
rect -2309 -2720 -2266 -2686
rect -2232 -2720 -2189 -2686
rect -2309 -2753 -2189 -2720
rect -2159 -2753 -2039 -2453
rect -2009 -2753 -1889 -2453
rect -1859 -2526 -1739 -2453
rect -1859 -2560 -1816 -2526
rect -1782 -2560 -1739 -2526
rect -1859 -2606 -1739 -2560
rect -1859 -2640 -1816 -2606
rect -1782 -2640 -1739 -2606
rect -1859 -2686 -1739 -2640
rect -1859 -2720 -1816 -2686
rect -1782 -2720 -1739 -2686
rect -1859 -2753 -1739 -2720
rect -1369 -2526 -1249 -2453
rect -1369 -2560 -1326 -2526
rect -1292 -2560 -1249 -2526
rect -1369 -2606 -1249 -2560
rect -1369 -2640 -1326 -2606
rect -1292 -2640 -1249 -2606
rect -1369 -2686 -1249 -2640
rect -1369 -2720 -1326 -2686
rect -1292 -2720 -1249 -2686
rect -1369 -2753 -1249 -2720
rect -1219 -2526 -1099 -2453
rect -1219 -2560 -1176 -2526
rect -1142 -2560 -1099 -2526
rect -1219 -2606 -1099 -2560
rect -1219 -2640 -1176 -2606
rect -1142 -2640 -1099 -2606
rect -1219 -2686 -1099 -2640
rect -1219 -2720 -1176 -2686
rect -1142 -2720 -1099 -2686
rect -1219 -2753 -1099 -2720
rect -1039 -2526 -919 -2453
rect -1039 -2560 -996 -2526
rect -962 -2560 -919 -2526
rect -1039 -2606 -919 -2560
rect -1039 -2640 -996 -2606
rect -962 -2640 -919 -2606
rect -1039 -2686 -919 -2640
rect -1039 -2720 -996 -2686
rect -962 -2720 -919 -2686
rect -1039 -2753 -919 -2720
rect -889 -2526 -769 -2453
rect -889 -2560 -846 -2526
rect -812 -2560 -769 -2526
rect -889 -2606 -769 -2560
rect -889 -2640 -846 -2606
rect -812 -2640 -769 -2606
rect -889 -2686 -769 -2640
rect -889 -2720 -846 -2686
rect -812 -2720 -769 -2686
rect -889 -2753 -769 -2720
rect -739 -2526 -619 -2453
rect -739 -2560 -696 -2526
rect -662 -2560 -619 -2526
rect -739 -2606 -619 -2560
rect -739 -2640 -696 -2606
rect -662 -2640 -619 -2606
rect -739 -2686 -619 -2640
rect -739 -2720 -696 -2686
rect -662 -2720 -619 -2686
rect -739 -2753 -619 -2720
rect -589 -2526 -469 -2453
rect -589 -2560 -546 -2526
rect -512 -2560 -469 -2526
rect -589 -2606 -469 -2560
rect -589 -2640 -546 -2606
rect -512 -2640 -469 -2606
rect -589 -2686 -469 -2640
rect -589 -2720 -546 -2686
rect -512 -2720 -469 -2686
rect -589 -2753 -469 -2720
rect -439 -2526 -319 -2453
rect -439 -2560 -396 -2526
rect -362 -2560 -319 -2526
rect -439 -2606 -319 -2560
rect -439 -2640 -396 -2606
rect -362 -2640 -319 -2606
rect -439 -2686 -319 -2640
rect -439 -2720 -396 -2686
rect -362 -2720 -319 -2686
rect -439 -2753 -319 -2720
rect -259 -2526 -139 -2453
rect -259 -2560 -216 -2526
rect -182 -2560 -139 -2526
rect -259 -2606 -139 -2560
rect -259 -2640 -216 -2606
rect -182 -2640 -139 -2606
rect -259 -2686 -139 -2640
rect -259 -2720 -216 -2686
rect -182 -2720 -139 -2686
rect -259 -2753 -139 -2720
rect -109 -2526 11 -2453
rect -109 -2560 -66 -2526
rect -32 -2560 11 -2526
rect -109 -2606 11 -2560
rect -109 -2640 -66 -2606
rect -32 -2640 11 -2606
rect -109 -2686 11 -2640
rect -109 -2720 -66 -2686
rect -32 -2720 11 -2686
rect -109 -2753 11 -2720
rect 371 -2527 491 -2454
rect 371 -2561 414 -2527
rect 448 -2561 491 -2527
rect 371 -2607 491 -2561
rect 371 -2641 414 -2607
rect 448 -2641 491 -2607
rect 371 -2687 491 -2641
rect 371 -2721 414 -2687
rect 448 -2721 491 -2687
rect 371 -2754 491 -2721
rect 521 -2527 641 -2454
rect 521 -2561 564 -2527
rect 598 -2561 641 -2527
rect 521 -2607 641 -2561
rect 521 -2641 564 -2607
rect 598 -2641 641 -2607
rect 521 -2687 641 -2641
rect 521 -2721 564 -2687
rect 598 -2721 641 -2687
rect 521 -2754 641 -2721
rect 671 -2527 791 -2454
rect 671 -2561 714 -2527
rect 748 -2561 791 -2527
rect 671 -2607 791 -2561
rect 671 -2641 714 -2607
rect 748 -2641 791 -2607
rect 671 -2687 791 -2641
rect 671 -2721 714 -2687
rect 748 -2721 791 -2687
rect 671 -2754 791 -2721
rect 821 -2527 941 -2454
rect 821 -2561 864 -2527
rect 898 -2561 941 -2527
rect 821 -2607 941 -2561
rect 821 -2641 864 -2607
rect 898 -2641 941 -2607
rect 821 -2687 941 -2641
rect 821 -2721 864 -2687
rect 898 -2721 941 -2687
rect 821 -2754 941 -2721
rect 1001 -2527 1121 -2454
rect 1001 -2561 1044 -2527
rect 1078 -2561 1121 -2527
rect 1001 -2607 1121 -2561
rect 1001 -2641 1044 -2607
rect 1078 -2641 1121 -2607
rect 1001 -2687 1121 -2641
rect 1001 -2721 1044 -2687
rect 1078 -2721 1121 -2687
rect 1001 -2754 1121 -2721
rect 1151 -2527 1271 -2454
rect 1151 -2561 1194 -2527
rect 1228 -2561 1271 -2527
rect 1151 -2607 1271 -2561
rect 1151 -2641 1194 -2607
rect 1228 -2641 1271 -2607
rect 1151 -2687 1271 -2641
rect 1151 -2721 1194 -2687
rect 1228 -2721 1271 -2687
rect 1151 -2754 1271 -2721
rect 1301 -2527 1421 -2454
rect 1301 -2561 1344 -2527
rect 1378 -2561 1421 -2527
rect 1301 -2607 1421 -2561
rect 1301 -2641 1344 -2607
rect 1378 -2641 1421 -2607
rect 1301 -2687 1421 -2641
rect 1301 -2721 1344 -2687
rect 1378 -2721 1421 -2687
rect 1301 -2754 1421 -2721
rect 1451 -2527 1571 -2454
rect 1451 -2561 1494 -2527
rect 1528 -2561 1571 -2527
rect 1451 -2607 1571 -2561
rect 1451 -2641 1494 -2607
rect 1528 -2641 1571 -2607
rect 1451 -2687 1571 -2641
rect 1451 -2721 1494 -2687
rect 1528 -2721 1571 -2687
rect 1451 -2754 1571 -2721
rect 1601 -2527 1721 -2454
rect 1601 -2561 1644 -2527
rect 1678 -2561 1721 -2527
rect 1601 -2607 1721 -2561
rect 1601 -2641 1644 -2607
rect 1678 -2641 1721 -2607
rect 1601 -2687 1721 -2641
rect 1601 -2721 1644 -2687
rect 1678 -2721 1721 -2687
rect 1601 -2754 1721 -2721
rect 1781 -2527 1901 -2454
rect 1781 -2561 1824 -2527
rect 1858 -2561 1901 -2527
rect 1781 -2607 1901 -2561
rect 1781 -2641 1824 -2607
rect 1858 -2641 1901 -2607
rect 1781 -2687 1901 -2641
rect 1781 -2721 1824 -2687
rect 1858 -2721 1901 -2687
rect 1781 -2754 1901 -2721
rect 1931 -2754 2051 -2454
rect 2081 -2754 2201 -2454
rect 2231 -2527 2351 -2454
rect 2231 -2561 2274 -2527
rect 2308 -2561 2351 -2527
rect 2231 -2607 2351 -2561
rect 2231 -2641 2274 -2607
rect 2308 -2641 2351 -2607
rect 2231 -2687 2351 -2641
rect 2231 -2721 2274 -2687
rect 2308 -2721 2351 -2687
rect 2231 -2754 2351 -2721
<< pdiff >>
rect -3090 854 -2970 927
rect -3090 820 -3047 854
rect -3013 820 -2970 854
rect -3090 774 -2970 820
rect -3090 740 -3047 774
rect -3013 740 -2970 774
rect -3090 694 -2970 740
rect -3090 660 -3047 694
rect -3013 660 -2970 694
rect -3090 627 -2970 660
rect -2940 854 -2820 927
rect -2940 820 -2897 854
rect -2863 820 -2820 854
rect -2940 774 -2820 820
rect -2940 740 -2897 774
rect -2863 740 -2820 774
rect -2940 694 -2820 740
rect -2940 660 -2897 694
rect -2863 660 -2820 694
rect -2940 627 -2820 660
rect -2790 854 -2670 927
rect -2790 820 -2747 854
rect -2713 820 -2670 854
rect -2790 774 -2670 820
rect -2790 740 -2747 774
rect -2713 740 -2670 774
rect -2790 694 -2670 740
rect -2790 660 -2747 694
rect -2713 660 -2670 694
rect -2790 627 -2670 660
rect -2640 854 -2520 927
rect -2640 820 -2597 854
rect -2563 820 -2520 854
rect -2640 774 -2520 820
rect -2640 740 -2597 774
rect -2563 740 -2520 774
rect -2640 694 -2520 740
rect -2640 660 -2597 694
rect -2563 660 -2520 694
rect -2640 627 -2520 660
rect -2490 854 -2370 927
rect -2490 820 -2447 854
rect -2413 820 -2370 854
rect -2490 774 -2370 820
rect -2490 740 -2447 774
rect -2413 740 -2370 774
rect -2490 694 -2370 740
rect -2490 660 -2447 694
rect -2413 660 -2370 694
rect -2490 627 -2370 660
rect -900 854 -780 927
rect -900 820 -857 854
rect -823 820 -780 854
rect -900 774 -780 820
rect -900 740 -857 774
rect -823 740 -780 774
rect -900 694 -780 740
rect -900 660 -857 694
rect -823 660 -780 694
rect -900 627 -780 660
rect -750 854 -630 927
rect -750 820 -707 854
rect -673 820 -630 854
rect -750 774 -630 820
rect -750 740 -707 774
rect -673 740 -630 774
rect -750 694 -630 740
rect -750 660 -707 694
rect -673 660 -630 694
rect -750 627 -630 660
rect -600 854 -480 927
rect -600 820 -557 854
rect -523 820 -480 854
rect -600 774 -480 820
rect -600 740 -557 774
rect -523 740 -480 774
rect -600 694 -480 740
rect -600 660 -557 694
rect -523 660 -480 694
rect -600 627 -480 660
rect -450 854 -330 927
rect -450 820 -407 854
rect -373 820 -330 854
rect -450 774 -330 820
rect -450 740 -407 774
rect -373 740 -330 774
rect -450 694 -330 740
rect -450 660 -407 694
rect -373 660 -330 694
rect -450 627 -330 660
rect -300 854 -180 927
rect -300 820 -257 854
rect -223 820 -180 854
rect -300 774 -180 820
rect -300 740 -257 774
rect -223 740 -180 774
rect -300 694 -180 740
rect 980 854 1100 927
rect 980 820 1023 854
rect 1057 820 1100 854
rect 980 774 1100 820
rect 980 740 1023 774
rect 1057 740 1100 774
rect -300 660 -257 694
rect -223 660 -180 694
rect -300 627 -180 660
rect 980 694 1100 740
rect 980 660 1023 694
rect 1057 660 1100 694
rect 980 627 1100 660
rect 1130 854 1250 927
rect 1130 820 1173 854
rect 1207 820 1250 854
rect 1130 774 1250 820
rect 1130 740 1173 774
rect 1207 740 1250 774
rect 1130 694 1250 740
rect 1130 660 1173 694
rect 1207 660 1250 694
rect 1130 627 1250 660
rect 1280 854 1400 927
rect 1280 820 1323 854
rect 1357 820 1400 854
rect 1280 774 1400 820
rect 1280 740 1323 774
rect 1357 740 1400 774
rect 1280 694 1400 740
rect 1280 660 1323 694
rect 1357 660 1400 694
rect 1280 627 1400 660
rect 1430 854 1550 927
rect 1430 820 1473 854
rect 1507 820 1550 854
rect 1430 774 1550 820
rect 1430 740 1473 774
rect 1507 740 1550 774
rect 1430 694 1550 740
rect 1430 660 1473 694
rect 1507 660 1550 694
rect 1430 627 1550 660
rect 1580 854 1700 927
rect 1580 820 1623 854
rect 1657 820 1700 854
rect 1580 774 1700 820
rect 1580 740 1623 774
rect 1657 740 1700 774
rect 1580 694 1700 740
rect 1580 660 1623 694
rect 1657 660 1700 694
rect 1580 627 1700 660
rect -3090 -906 -2970 -873
rect -3090 -940 -3047 -906
rect -3013 -940 -2970 -906
rect -3090 -986 -2970 -940
rect -3090 -1020 -3047 -986
rect -3013 -1020 -2970 -986
rect -3090 -1066 -2970 -1020
rect -3090 -1100 -3047 -1066
rect -3013 -1100 -2970 -1066
rect -3090 -1173 -2970 -1100
rect -2940 -906 -2820 -873
rect -2940 -940 -2897 -906
rect -2863 -940 -2820 -906
rect -2940 -986 -2820 -940
rect -2940 -1020 -2897 -986
rect -2863 -1020 -2820 -986
rect -2940 -1066 -2820 -1020
rect -2940 -1100 -2897 -1066
rect -2863 -1100 -2820 -1066
rect -2940 -1173 -2820 -1100
rect -2790 -906 -2670 -873
rect -2790 -940 -2747 -906
rect -2713 -940 -2670 -906
rect -2790 -986 -2670 -940
rect -2790 -1020 -2747 -986
rect -2713 -1020 -2670 -986
rect -2790 -1066 -2670 -1020
rect -2790 -1100 -2747 -1066
rect -2713 -1100 -2670 -1066
rect -2790 -1173 -2670 -1100
rect -2640 -906 -2520 -873
rect -2640 -940 -2597 -906
rect -2563 -940 -2520 -906
rect -2640 -986 -2520 -940
rect -2640 -1020 -2597 -986
rect -2563 -1020 -2520 -986
rect -2640 -1066 -2520 -1020
rect -2640 -1100 -2597 -1066
rect -2563 -1100 -2520 -1066
rect -2640 -1173 -2520 -1100
rect -2490 -906 -2370 -873
rect -2490 -940 -2447 -906
rect -2413 -940 -2370 -906
rect -2490 -986 -2370 -940
rect -2490 -1020 -2447 -986
rect -2413 -1020 -2370 -986
rect -2490 -1066 -2370 -1020
rect -2490 -1100 -2447 -1066
rect -2413 -1100 -2370 -1066
rect -2490 -1173 -2370 -1100
rect -900 -906 -780 -873
rect -900 -940 -857 -906
rect -823 -940 -780 -906
rect -900 -986 -780 -940
rect -900 -1020 -857 -986
rect -823 -1020 -780 -986
rect -900 -1066 -780 -1020
rect -900 -1100 -857 -1066
rect -823 -1100 -780 -1066
rect -900 -1173 -780 -1100
rect -750 -906 -630 -873
rect -750 -940 -707 -906
rect -673 -940 -630 -906
rect -750 -986 -630 -940
rect -750 -1020 -707 -986
rect -673 -1020 -630 -986
rect -750 -1066 -630 -1020
rect -750 -1100 -707 -1066
rect -673 -1100 -630 -1066
rect -750 -1173 -630 -1100
rect -600 -906 -480 -873
rect -600 -940 -557 -906
rect -523 -940 -480 -906
rect -600 -986 -480 -940
rect -600 -1020 -557 -986
rect -523 -1020 -480 -986
rect -600 -1066 -480 -1020
rect -600 -1100 -557 -1066
rect -523 -1100 -480 -1066
rect -600 -1173 -480 -1100
rect -450 -906 -330 -873
rect -450 -940 -407 -906
rect -373 -940 -330 -906
rect -450 -986 -330 -940
rect -450 -1020 -407 -986
rect -373 -1020 -330 -986
rect -450 -1066 -330 -1020
rect -450 -1100 -407 -1066
rect -373 -1100 -330 -1066
rect -450 -1173 -330 -1100
rect -300 -906 -180 -873
rect -300 -940 -257 -906
rect -223 -940 -180 -906
rect -300 -986 -180 -940
rect 980 -906 1100 -873
rect 980 -940 1023 -906
rect 1057 -940 1100 -906
rect -300 -1020 -257 -986
rect -223 -1020 -180 -986
rect -300 -1066 -180 -1020
rect -300 -1100 -257 -1066
rect -223 -1100 -180 -1066
rect -300 -1173 -180 -1100
rect 980 -986 1100 -940
rect 980 -1020 1023 -986
rect 1057 -1020 1100 -986
rect 980 -1066 1100 -1020
rect 980 -1100 1023 -1066
rect 1057 -1100 1100 -1066
rect 980 -1173 1100 -1100
rect 1130 -906 1250 -873
rect 1130 -940 1173 -906
rect 1207 -940 1250 -906
rect 1130 -986 1250 -940
rect 1130 -1020 1173 -986
rect 1207 -1020 1250 -986
rect 1130 -1066 1250 -1020
rect 1130 -1100 1173 -1066
rect 1207 -1100 1250 -1066
rect 1130 -1173 1250 -1100
rect 1280 -906 1400 -873
rect 1280 -940 1323 -906
rect 1357 -940 1400 -906
rect 1280 -986 1400 -940
rect 1280 -1020 1323 -986
rect 1357 -1020 1400 -986
rect 1280 -1066 1400 -1020
rect 1280 -1100 1323 -1066
rect 1357 -1100 1400 -1066
rect 1280 -1173 1400 -1100
rect 1430 -906 1550 -873
rect 1430 -940 1473 -906
rect 1507 -940 1550 -906
rect 1430 -986 1550 -940
rect 1430 -1020 1473 -986
rect 1507 -1020 1550 -986
rect 1430 -1066 1550 -1020
rect 1430 -1100 1473 -1066
rect 1507 -1100 1550 -1066
rect 1430 -1173 1550 -1100
rect 1580 -906 1700 -873
rect 1580 -940 1623 -906
rect 1657 -940 1700 -906
rect 1580 -986 1700 -940
rect 1580 -1020 1623 -986
rect 1657 -1020 1700 -986
rect 1580 -1066 1700 -1020
rect 1580 -1100 1623 -1066
rect 1657 -1100 1700 -1066
rect 1580 -1173 1700 -1100
rect -3089 -1966 -2969 -1893
rect -3089 -2000 -3046 -1966
rect -3012 -2000 -2969 -1966
rect -3089 -2046 -2969 -2000
rect -3089 -2080 -3046 -2046
rect -3012 -2080 -2969 -2046
rect -3089 -2126 -2969 -2080
rect -3089 -2160 -3046 -2126
rect -3012 -2160 -2969 -2126
rect -3089 -2193 -2969 -2160
rect -2939 -1966 -2819 -1893
rect -2939 -2000 -2896 -1966
rect -2862 -2000 -2819 -1966
rect -2939 -2046 -2819 -2000
rect -2939 -2080 -2896 -2046
rect -2862 -2080 -2819 -2046
rect -2939 -2126 -2819 -2080
rect -2939 -2160 -2896 -2126
rect -2862 -2160 -2819 -2126
rect -2939 -2193 -2819 -2160
rect -2789 -1966 -2669 -1893
rect -2789 -2000 -2746 -1966
rect -2712 -2000 -2669 -1966
rect -2789 -2046 -2669 -2000
rect -2789 -2080 -2746 -2046
rect -2712 -2080 -2669 -2046
rect -2789 -2126 -2669 -2080
rect -2789 -2160 -2746 -2126
rect -2712 -2160 -2669 -2126
rect -2789 -2193 -2669 -2160
rect -2639 -1966 -2519 -1893
rect -2639 -2000 -2596 -1966
rect -2562 -2000 -2519 -1966
rect -2639 -2046 -2519 -2000
rect -2639 -2080 -2596 -2046
rect -2562 -2080 -2519 -2046
rect -2639 -2126 -2519 -2080
rect -2639 -2160 -2596 -2126
rect -2562 -2160 -2519 -2126
rect -2639 -2193 -2519 -2160
rect -2489 -1966 -2369 -1893
rect -2489 -2000 -2446 -1966
rect -2412 -2000 -2369 -1966
rect -2489 -2046 -2369 -2000
rect -2489 -2080 -2446 -2046
rect -2412 -2080 -2369 -2046
rect -2489 -2126 -2369 -2080
rect -2489 -2160 -2446 -2126
rect -2412 -2160 -2369 -2126
rect -2489 -2193 -2369 -2160
rect -1039 -1966 -919 -1893
rect -1039 -2000 -996 -1966
rect -962 -2000 -919 -1966
rect -1039 -2046 -919 -2000
rect -1039 -2080 -996 -2046
rect -962 -2080 -919 -2046
rect -1039 -2126 -919 -2080
rect -1039 -2160 -996 -2126
rect -962 -2160 -919 -2126
rect -1039 -2193 -919 -2160
rect -889 -1966 -769 -1893
rect -889 -2000 -846 -1966
rect -812 -2000 -769 -1966
rect -889 -2046 -769 -2000
rect -889 -2080 -846 -2046
rect -812 -2080 -769 -2046
rect -889 -2126 -769 -2080
rect -889 -2160 -846 -2126
rect -812 -2160 -769 -2126
rect -889 -2193 -769 -2160
rect -739 -1966 -619 -1893
rect -739 -2000 -696 -1966
rect -662 -2000 -619 -1966
rect -739 -2046 -619 -2000
rect -739 -2080 -696 -2046
rect -662 -2080 -619 -2046
rect -739 -2126 -619 -2080
rect -739 -2160 -696 -2126
rect -662 -2160 -619 -2126
rect -739 -2193 -619 -2160
rect -589 -1966 -469 -1893
rect -589 -2000 -546 -1966
rect -512 -2000 -469 -1966
rect -589 -2046 -469 -2000
rect -589 -2080 -546 -2046
rect -512 -2080 -469 -2046
rect -589 -2126 -469 -2080
rect -589 -2160 -546 -2126
rect -512 -2160 -469 -2126
rect -589 -2193 -469 -2160
rect -439 -1966 -319 -1893
rect -439 -2000 -396 -1966
rect -362 -2000 -319 -1966
rect -439 -2046 -319 -2000
rect -439 -2080 -396 -2046
rect -362 -2080 -319 -2046
rect -439 -2126 -319 -2080
rect -439 -2160 -396 -2126
rect -362 -2160 -319 -2126
rect -439 -2193 -319 -2160
rect 1001 -1967 1121 -1894
rect 1001 -2001 1044 -1967
rect 1078 -2001 1121 -1967
rect 1001 -2047 1121 -2001
rect 1001 -2081 1044 -2047
rect 1078 -2081 1121 -2047
rect 1001 -2127 1121 -2081
rect 1001 -2161 1044 -2127
rect 1078 -2161 1121 -2127
rect 1001 -2194 1121 -2161
rect 1151 -1967 1271 -1894
rect 1151 -2001 1194 -1967
rect 1228 -2001 1271 -1967
rect 1151 -2047 1271 -2001
rect 1151 -2081 1194 -2047
rect 1228 -2081 1271 -2047
rect 1151 -2127 1271 -2081
rect 1151 -2161 1194 -2127
rect 1228 -2161 1271 -2127
rect 1151 -2194 1271 -2161
rect 1301 -1967 1421 -1894
rect 1301 -2001 1344 -1967
rect 1378 -2001 1421 -1967
rect 1301 -2047 1421 -2001
rect 1301 -2081 1344 -2047
rect 1378 -2081 1421 -2047
rect 1301 -2127 1421 -2081
rect 1301 -2161 1344 -2127
rect 1378 -2161 1421 -2127
rect 1301 -2194 1421 -2161
rect 1451 -1967 1571 -1894
rect 1451 -2001 1494 -1967
rect 1528 -2001 1571 -1967
rect 1451 -2047 1571 -2001
rect 1451 -2081 1494 -2047
rect 1528 -2081 1571 -2047
rect 1451 -2127 1571 -2081
rect 1451 -2161 1494 -2127
rect 1528 -2161 1571 -2127
rect 1451 -2194 1571 -2161
rect 1601 -1967 1721 -1894
rect 1601 -2001 1644 -1967
rect 1678 -2001 1721 -1967
rect 1601 -2047 1721 -2001
rect 1601 -2081 1644 -2047
rect 1678 -2081 1721 -2047
rect 1601 -2127 1721 -2081
rect 1601 -2161 1644 -2127
rect 1678 -2161 1721 -2127
rect 1601 -2194 1721 -2161
<< ndiffc >>
rect -3827 260 -3793 294
rect -3827 180 -3793 214
rect -3827 100 -3793 134
rect -3527 260 -3493 294
rect -3527 180 -3493 214
rect -3527 100 -3493 134
rect -3227 260 -3193 294
rect -3227 180 -3193 214
rect -3227 100 -3193 134
rect -3047 260 -3013 294
rect -3047 180 -3013 214
rect -3047 100 -3013 134
rect -2897 260 -2863 294
rect -2897 180 -2863 214
rect -2897 100 -2863 134
rect -2747 260 -2713 294
rect -2747 180 -2713 214
rect -2747 100 -2713 134
rect -2597 260 -2563 294
rect -2597 180 -2563 214
rect -2597 100 -2563 134
rect -2447 260 -2413 294
rect -2447 180 -2413 214
rect -2447 100 -2413 134
rect -2267 260 -2233 294
rect -2267 180 -2233 214
rect -2267 100 -2233 134
rect -1967 260 -1933 294
rect -1967 180 -1933 214
rect -1967 100 -1933 134
rect -1667 260 -1633 294
rect -1667 180 -1633 214
rect -1667 100 -1633 134
rect -1187 260 -1153 294
rect -1187 180 -1153 214
rect -1187 100 -1153 134
rect -1037 260 -1003 294
rect -1037 180 -1003 214
rect -1037 100 -1003 134
rect -857 260 -823 294
rect -857 180 -823 214
rect -857 100 -823 134
rect -707 260 -673 294
rect -707 180 -673 214
rect -707 100 -673 134
rect -557 260 -523 294
rect -557 180 -523 214
rect -557 100 -523 134
rect -407 260 -373 294
rect -407 180 -373 214
rect -407 100 -373 134
rect -257 260 -223 294
rect -257 180 -223 214
rect -257 100 -223 134
rect -77 260 -43 294
rect -77 180 -43 214
rect -77 100 -43 134
rect 73 260 107 294
rect 73 180 107 214
rect 73 100 107 134
rect 543 260 577 294
rect 543 180 577 214
rect 543 100 577 134
rect 693 260 727 294
rect 693 180 727 214
rect 693 100 727 134
rect 843 260 877 294
rect 843 180 877 214
rect 843 100 877 134
rect 1023 260 1057 294
rect 1023 180 1057 214
rect 1023 100 1057 134
rect 1173 260 1207 294
rect 1173 180 1207 214
rect 1173 100 1207 134
rect 1323 260 1357 294
rect 1323 180 1357 214
rect 1323 100 1357 134
rect 1473 260 1507 294
rect 1473 180 1507 214
rect 1473 100 1507 134
rect 1623 260 1657 294
rect 1623 180 1657 214
rect 1623 100 1657 134
rect 1803 260 1837 294
rect 1803 180 1837 214
rect 1803 100 1837 134
rect 2103 260 2137 294
rect 2103 180 2137 214
rect 2103 100 2137 134
rect -3827 -380 -3793 -346
rect -3827 -460 -3793 -426
rect -3827 -540 -3793 -506
rect -3527 -380 -3493 -346
rect -3527 -460 -3493 -426
rect -3527 -540 -3493 -506
rect -3227 -380 -3193 -346
rect -3227 -460 -3193 -426
rect -3227 -540 -3193 -506
rect -3047 -380 -3013 -346
rect -3047 -460 -3013 -426
rect -3047 -540 -3013 -506
rect -2897 -380 -2863 -346
rect -2897 -460 -2863 -426
rect -2897 -540 -2863 -506
rect -2747 -380 -2713 -346
rect -2747 -460 -2713 -426
rect -2747 -540 -2713 -506
rect -2597 -380 -2563 -346
rect -2597 -460 -2563 -426
rect -2597 -540 -2563 -506
rect -2447 -380 -2413 -346
rect -2447 -460 -2413 -426
rect -2447 -540 -2413 -506
rect -2267 -380 -2233 -346
rect -2267 -460 -2233 -426
rect -2267 -540 -2233 -506
rect -1967 -380 -1933 -346
rect -1967 -460 -1933 -426
rect -1967 -540 -1933 -506
rect -1667 -380 -1633 -346
rect -1667 -460 -1633 -426
rect -1667 -540 -1633 -506
rect -1187 -380 -1153 -346
rect -1187 -460 -1153 -426
rect -1187 -540 -1153 -506
rect -1037 -380 -1003 -346
rect -1037 -460 -1003 -426
rect -1037 -540 -1003 -506
rect -857 -380 -823 -346
rect -857 -460 -823 -426
rect -857 -540 -823 -506
rect -707 -380 -673 -346
rect -707 -460 -673 -426
rect -707 -540 -673 -506
rect -557 -380 -523 -346
rect -557 -460 -523 -426
rect -557 -540 -523 -506
rect -407 -380 -373 -346
rect -407 -460 -373 -426
rect -407 -540 -373 -506
rect -257 -380 -223 -346
rect -257 -460 -223 -426
rect -257 -540 -223 -506
rect -77 -380 -43 -346
rect -77 -460 -43 -426
rect -77 -540 -43 -506
rect 73 -380 107 -346
rect 73 -460 107 -426
rect 73 -540 107 -506
rect 543 -380 577 -346
rect 543 -460 577 -426
rect 543 -540 577 -506
rect 693 -380 727 -346
rect 693 -460 727 -426
rect 693 -540 727 -506
rect 843 -380 877 -346
rect 843 -460 877 -426
rect 843 -540 877 -506
rect 1023 -380 1057 -346
rect 1023 -460 1057 -426
rect 1023 -540 1057 -506
rect 1173 -380 1207 -346
rect 1173 -460 1207 -426
rect 1173 -540 1207 -506
rect 1323 -380 1357 -346
rect 1323 -460 1357 -426
rect 1323 -540 1357 -506
rect 1473 -380 1507 -346
rect 1473 -460 1507 -426
rect 1473 -540 1507 -506
rect 1623 -380 1657 -346
rect 1623 -460 1657 -426
rect 1623 -540 1657 -506
rect 1803 -380 1837 -346
rect 1803 -460 1837 -426
rect 1803 -540 1837 -506
rect 2103 -380 2137 -346
rect 2103 -460 2137 -426
rect 2103 -540 2137 -506
rect -3676 -2560 -3642 -2526
rect -3676 -2640 -3642 -2606
rect -3676 -2720 -3642 -2686
rect -3526 -2560 -3492 -2526
rect -3526 -2640 -3492 -2606
rect -3526 -2720 -3492 -2686
rect -3376 -2560 -3342 -2526
rect -3376 -2640 -3342 -2606
rect -3376 -2720 -3342 -2686
rect -3226 -2560 -3192 -2526
rect -3226 -2640 -3192 -2606
rect -3226 -2720 -3192 -2686
rect -3046 -2560 -3012 -2526
rect -3046 -2640 -3012 -2606
rect -3046 -2720 -3012 -2686
rect -2896 -2560 -2862 -2526
rect -2896 -2640 -2862 -2606
rect -2896 -2720 -2862 -2686
rect -2746 -2560 -2712 -2526
rect -2746 -2640 -2712 -2606
rect -2746 -2720 -2712 -2686
rect -2596 -2560 -2562 -2526
rect -2596 -2640 -2562 -2606
rect -2596 -2720 -2562 -2686
rect -2446 -2560 -2412 -2526
rect -2446 -2640 -2412 -2606
rect -2446 -2720 -2412 -2686
rect -2266 -2560 -2232 -2526
rect -2266 -2640 -2232 -2606
rect -2266 -2720 -2232 -2686
rect -1816 -2560 -1782 -2526
rect -1816 -2640 -1782 -2606
rect -1816 -2720 -1782 -2686
rect -1326 -2560 -1292 -2526
rect -1326 -2640 -1292 -2606
rect -1326 -2720 -1292 -2686
rect -1176 -2560 -1142 -2526
rect -1176 -2640 -1142 -2606
rect -1176 -2720 -1142 -2686
rect -996 -2560 -962 -2526
rect -996 -2640 -962 -2606
rect -996 -2720 -962 -2686
rect -846 -2560 -812 -2526
rect -846 -2640 -812 -2606
rect -846 -2720 -812 -2686
rect -696 -2560 -662 -2526
rect -696 -2640 -662 -2606
rect -696 -2720 -662 -2686
rect -546 -2560 -512 -2526
rect -546 -2640 -512 -2606
rect -546 -2720 -512 -2686
rect -396 -2560 -362 -2526
rect -396 -2640 -362 -2606
rect -396 -2720 -362 -2686
rect -216 -2560 -182 -2526
rect -216 -2640 -182 -2606
rect -216 -2720 -182 -2686
rect -66 -2560 -32 -2526
rect -66 -2640 -32 -2606
rect -66 -2720 -32 -2686
rect 414 -2561 448 -2527
rect 414 -2641 448 -2607
rect 414 -2721 448 -2687
rect 564 -2561 598 -2527
rect 564 -2641 598 -2607
rect 564 -2721 598 -2687
rect 714 -2561 748 -2527
rect 714 -2641 748 -2607
rect 714 -2721 748 -2687
rect 864 -2561 898 -2527
rect 864 -2641 898 -2607
rect 864 -2721 898 -2687
rect 1044 -2561 1078 -2527
rect 1044 -2641 1078 -2607
rect 1044 -2721 1078 -2687
rect 1194 -2561 1228 -2527
rect 1194 -2641 1228 -2607
rect 1194 -2721 1228 -2687
rect 1344 -2561 1378 -2527
rect 1344 -2641 1378 -2607
rect 1344 -2721 1378 -2687
rect 1494 -2561 1528 -2527
rect 1494 -2641 1528 -2607
rect 1494 -2721 1528 -2687
rect 1644 -2561 1678 -2527
rect 1644 -2641 1678 -2607
rect 1644 -2721 1678 -2687
rect 1824 -2561 1858 -2527
rect 1824 -2641 1858 -2607
rect 1824 -2721 1858 -2687
rect 2274 -2561 2308 -2527
rect 2274 -2641 2308 -2607
rect 2274 -2721 2308 -2687
<< pdiffc >>
rect -3047 820 -3013 854
rect -3047 740 -3013 774
rect -3047 660 -3013 694
rect -2897 820 -2863 854
rect -2897 740 -2863 774
rect -2897 660 -2863 694
rect -2747 820 -2713 854
rect -2747 740 -2713 774
rect -2747 660 -2713 694
rect -2597 820 -2563 854
rect -2597 740 -2563 774
rect -2597 660 -2563 694
rect -2447 820 -2413 854
rect -2447 740 -2413 774
rect -2447 660 -2413 694
rect -857 820 -823 854
rect -857 740 -823 774
rect -857 660 -823 694
rect -707 820 -673 854
rect -707 740 -673 774
rect -707 660 -673 694
rect -557 820 -523 854
rect -557 740 -523 774
rect -557 660 -523 694
rect -407 820 -373 854
rect -407 740 -373 774
rect -407 660 -373 694
rect -257 820 -223 854
rect -257 740 -223 774
rect 1023 820 1057 854
rect 1023 740 1057 774
rect -257 660 -223 694
rect 1023 660 1057 694
rect 1173 820 1207 854
rect 1173 740 1207 774
rect 1173 660 1207 694
rect 1323 820 1357 854
rect 1323 740 1357 774
rect 1323 660 1357 694
rect 1473 820 1507 854
rect 1473 740 1507 774
rect 1473 660 1507 694
rect 1623 820 1657 854
rect 1623 740 1657 774
rect 1623 660 1657 694
rect -3047 -940 -3013 -906
rect -3047 -1020 -3013 -986
rect -3047 -1100 -3013 -1066
rect -2897 -940 -2863 -906
rect -2897 -1020 -2863 -986
rect -2897 -1100 -2863 -1066
rect -2747 -940 -2713 -906
rect -2747 -1020 -2713 -986
rect -2747 -1100 -2713 -1066
rect -2597 -940 -2563 -906
rect -2597 -1020 -2563 -986
rect -2597 -1100 -2563 -1066
rect -2447 -940 -2413 -906
rect -2447 -1020 -2413 -986
rect -2447 -1100 -2413 -1066
rect -857 -940 -823 -906
rect -857 -1020 -823 -986
rect -857 -1100 -823 -1066
rect -707 -940 -673 -906
rect -707 -1020 -673 -986
rect -707 -1100 -673 -1066
rect -557 -940 -523 -906
rect -557 -1020 -523 -986
rect -557 -1100 -523 -1066
rect -407 -940 -373 -906
rect -407 -1020 -373 -986
rect -407 -1100 -373 -1066
rect -257 -940 -223 -906
rect 1023 -940 1057 -906
rect -257 -1020 -223 -986
rect -257 -1100 -223 -1066
rect 1023 -1020 1057 -986
rect 1023 -1100 1057 -1066
rect 1173 -940 1207 -906
rect 1173 -1020 1207 -986
rect 1173 -1100 1207 -1066
rect 1323 -940 1357 -906
rect 1323 -1020 1357 -986
rect 1323 -1100 1357 -1066
rect 1473 -940 1507 -906
rect 1473 -1020 1507 -986
rect 1473 -1100 1507 -1066
rect 1623 -940 1657 -906
rect 1623 -1020 1657 -986
rect 1623 -1100 1657 -1066
rect -3046 -2000 -3012 -1966
rect -3046 -2080 -3012 -2046
rect -3046 -2160 -3012 -2126
rect -2896 -2000 -2862 -1966
rect -2896 -2080 -2862 -2046
rect -2896 -2160 -2862 -2126
rect -2746 -2000 -2712 -1966
rect -2746 -2080 -2712 -2046
rect -2746 -2160 -2712 -2126
rect -2596 -2000 -2562 -1966
rect -2596 -2080 -2562 -2046
rect -2596 -2160 -2562 -2126
rect -2446 -2000 -2412 -1966
rect -2446 -2080 -2412 -2046
rect -2446 -2160 -2412 -2126
rect -996 -2000 -962 -1966
rect -996 -2080 -962 -2046
rect -996 -2160 -962 -2126
rect -846 -2000 -812 -1966
rect -846 -2080 -812 -2046
rect -846 -2160 -812 -2126
rect -696 -2000 -662 -1966
rect -696 -2080 -662 -2046
rect -696 -2160 -662 -2126
rect -546 -2000 -512 -1966
rect -546 -2080 -512 -2046
rect -546 -2160 -512 -2126
rect -396 -2000 -362 -1966
rect -396 -2080 -362 -2046
rect -396 -2160 -362 -2126
rect 1044 -2001 1078 -1967
rect 1044 -2081 1078 -2047
rect 1044 -2161 1078 -2127
rect 1194 -2001 1228 -1967
rect 1194 -2081 1228 -2047
rect 1194 -2161 1228 -2127
rect 1344 -2001 1378 -1967
rect 1344 -2081 1378 -2047
rect 1344 -2161 1378 -2127
rect 1494 -2001 1528 -1967
rect 1494 -2081 1528 -2047
rect 1494 -2161 1528 -2127
rect 1644 -2001 1678 -1967
rect 1644 -2081 1678 -2047
rect 1644 -2161 1678 -2127
<< psubdiff >>
rect -3870 -106 -1590 -73
rect -3870 -140 -3787 -106
rect -3753 -140 -3707 -106
rect -3673 -140 -3627 -106
rect -3593 -140 -3547 -106
rect -3513 -140 -3467 -106
rect -3433 -140 -3387 -106
rect -3353 -140 -3307 -106
rect -3273 -140 -3227 -106
rect -3193 -140 -3147 -106
rect -3113 -140 -3067 -106
rect -3033 -140 -2987 -106
rect -2953 -140 -2907 -106
rect -2873 -140 -2827 -106
rect -2793 -140 -2747 -106
rect -2713 -140 -2667 -106
rect -2633 -140 -2587 -106
rect -2553 -140 -2507 -106
rect -2473 -140 -2427 -106
rect -2393 -140 -2347 -106
rect -2313 -140 -2267 -106
rect -2233 -140 -2187 -106
rect -2153 -140 -2107 -106
rect -2073 -140 -2027 -106
rect -1993 -140 -1947 -106
rect -1913 -140 -1867 -106
rect -1833 -140 -1787 -106
rect -1753 -140 -1707 -106
rect -1673 -140 -1590 -106
rect -3870 -173 -1590 -140
rect -1230 -106 150 -73
rect -1230 -140 -1197 -106
rect -1163 -140 -1117 -106
rect -1083 -140 -1037 -106
rect -1003 -140 -957 -106
rect -923 -140 -877 -106
rect -843 -140 -797 -106
rect -763 -140 -717 -106
rect -683 -140 -637 -106
rect -603 -140 -557 -106
rect -523 -140 -477 -106
rect -443 -140 -397 -106
rect -363 -140 -317 -106
rect -283 -140 -237 -106
rect -203 -140 -157 -106
rect -123 -140 -77 -106
rect -43 -140 3 -106
rect 37 -140 83 -106
rect 117 -140 150 -106
rect -1230 -173 150 -140
rect 500 -106 2180 -73
rect 500 -140 523 -106
rect 557 -140 603 -106
rect 637 -140 683 -106
rect 717 -140 763 -106
rect 797 -140 843 -106
rect 877 -140 923 -106
rect 957 -140 1003 -106
rect 1037 -140 1083 -106
rect 1117 -140 1163 -106
rect 1197 -140 1243 -106
rect 1277 -140 1323 -106
rect 1357 -140 1403 -106
rect 1437 -140 1483 -106
rect 1517 -140 1563 -106
rect 1597 -140 1643 -106
rect 1677 -140 1723 -106
rect 1757 -140 1803 -106
rect 1837 -140 1883 -106
rect 1917 -140 1963 -106
rect 1997 -140 2043 -106
rect 2077 -140 2123 -106
rect 2157 -140 2180 -106
rect 500 -173 2180 -140
rect -3729 -2926 -1729 -2893
rect -3729 -2960 -3706 -2926
rect -3672 -2960 -3626 -2926
rect -3592 -2960 -3546 -2926
rect -3512 -2960 -3466 -2926
rect -3432 -2960 -3386 -2926
rect -3352 -2960 -3306 -2926
rect -3272 -2960 -3226 -2926
rect -3192 -2960 -3146 -2926
rect -3112 -2960 -3066 -2926
rect -3032 -2960 -2986 -2926
rect -2952 -2960 -2906 -2926
rect -2872 -2960 -2826 -2926
rect -2792 -2960 -2746 -2926
rect -2712 -2960 -2666 -2926
rect -2632 -2960 -2586 -2926
rect -2552 -2960 -2506 -2926
rect -2472 -2960 -2426 -2926
rect -2392 -2960 -2346 -2926
rect -2312 -2960 -2266 -2926
rect -2232 -2960 -2186 -2926
rect -2152 -2960 -2106 -2926
rect -2072 -2960 -2026 -2926
rect -1992 -2960 -1946 -2926
rect -1912 -2960 -1866 -2926
rect -1832 -2960 -1786 -2926
rect -1752 -2960 -1729 -2926
rect -3729 -2993 -1729 -2960
rect -1369 -2926 11 -2893
rect -1369 -2960 -1336 -2926
rect -1302 -2960 -1256 -2926
rect -1222 -2960 -1176 -2926
rect -1142 -2960 -1096 -2926
rect -1062 -2960 -1016 -2926
rect -982 -2960 -936 -2926
rect -902 -2960 -856 -2926
rect -822 -2960 -776 -2926
rect -742 -2960 -696 -2926
rect -662 -2960 -616 -2926
rect -582 -2960 -536 -2926
rect -502 -2960 -456 -2926
rect -422 -2960 -376 -2926
rect -342 -2960 -296 -2926
rect -262 -2960 -216 -2926
rect -182 -2960 -136 -2926
rect -102 -2960 -56 -2926
rect -22 -2960 11 -2926
rect -1369 -2993 11 -2960
rect 361 -2927 2361 -2894
rect 361 -2961 384 -2927
rect 418 -2961 464 -2927
rect 498 -2961 544 -2927
rect 578 -2961 624 -2927
rect 658 -2961 704 -2927
rect 738 -2961 784 -2927
rect 818 -2961 864 -2927
rect 898 -2961 944 -2927
rect 978 -2961 1024 -2927
rect 1058 -2961 1104 -2927
rect 1138 -2961 1184 -2927
rect 1218 -2961 1264 -2927
rect 1298 -2961 1344 -2927
rect 1378 -2961 1424 -2927
rect 1458 -2961 1504 -2927
rect 1538 -2961 1584 -2927
rect 1618 -2961 1664 -2927
rect 1698 -2961 1744 -2927
rect 1778 -2961 1824 -2927
rect 1858 -2961 1904 -2927
rect 1938 -2961 1984 -2927
rect 2018 -2961 2064 -2927
rect 2098 -2961 2144 -2927
rect 2178 -2961 2224 -2927
rect 2258 -2961 2304 -2927
rect 2338 -2961 2361 -2927
rect 361 -2994 2361 -2961
<< nsubdiff >>
rect -3870 1074 -1590 1107
rect -3870 1040 -3787 1074
rect -3753 1040 -3707 1074
rect -3673 1040 -3627 1074
rect -3593 1040 -3547 1074
rect -3513 1040 -3467 1074
rect -3433 1040 -3387 1074
rect -3353 1040 -3307 1074
rect -3273 1040 -3227 1074
rect -3193 1040 -3147 1074
rect -3113 1040 -3067 1074
rect -3033 1040 -2987 1074
rect -2953 1040 -2907 1074
rect -2873 1040 -2827 1074
rect -2793 1040 -2747 1074
rect -2713 1040 -2667 1074
rect -2633 1040 -2587 1074
rect -2553 1040 -2507 1074
rect -2473 1040 -2427 1074
rect -2393 1040 -2347 1074
rect -2313 1040 -2267 1074
rect -2233 1040 -2187 1074
rect -2153 1040 -2107 1074
rect -2073 1040 -2027 1074
rect -1993 1040 -1947 1074
rect -1913 1040 -1867 1074
rect -1833 1040 -1787 1074
rect -1753 1040 -1707 1074
rect -1673 1040 -1590 1074
rect -3870 1007 -1590 1040
rect -1230 1074 150 1107
rect -1230 1040 -1197 1074
rect -1163 1040 -1117 1074
rect -1083 1040 -1037 1074
rect -1003 1040 -957 1074
rect -923 1040 -877 1074
rect -843 1040 -797 1074
rect -763 1040 -717 1074
rect -683 1040 -637 1074
rect -603 1040 -557 1074
rect -523 1040 -477 1074
rect -443 1040 -397 1074
rect -363 1040 -317 1074
rect -283 1040 -237 1074
rect -203 1040 -157 1074
rect -123 1040 -77 1074
rect -43 1040 3 1074
rect 37 1040 83 1074
rect 117 1040 150 1074
rect -1230 1007 150 1040
rect 500 1074 2180 1107
rect 500 1040 523 1074
rect 557 1040 603 1074
rect 637 1040 683 1074
rect 717 1040 763 1074
rect 797 1040 843 1074
rect 877 1040 923 1074
rect 957 1040 1003 1074
rect 1037 1040 1083 1074
rect 1117 1040 1163 1074
rect 1197 1040 1243 1074
rect 1277 1040 1323 1074
rect 1357 1040 1403 1074
rect 1437 1040 1483 1074
rect 1517 1040 1563 1074
rect 1597 1040 1643 1074
rect 1677 1040 1723 1074
rect 1757 1040 1803 1074
rect 1837 1040 1883 1074
rect 1917 1040 1963 1074
rect 1997 1040 2043 1074
rect 2077 1040 2123 1074
rect 2157 1040 2180 1074
rect 500 1007 2180 1040
rect -3870 -1286 -1590 -1253
rect -3870 -1320 -3787 -1286
rect -3753 -1320 -3707 -1286
rect -3673 -1320 -3627 -1286
rect -3593 -1320 -3547 -1286
rect -3513 -1320 -3467 -1286
rect -3433 -1320 -3387 -1286
rect -3353 -1320 -3307 -1286
rect -3273 -1320 -3227 -1286
rect -3193 -1320 -3147 -1286
rect -3113 -1320 -3067 -1286
rect -3033 -1320 -2987 -1286
rect -2953 -1320 -2907 -1286
rect -2873 -1320 -2827 -1286
rect -2793 -1320 -2747 -1286
rect -2713 -1320 -2667 -1286
rect -2633 -1320 -2587 -1286
rect -2553 -1320 -2507 -1286
rect -2473 -1320 -2427 -1286
rect -2393 -1320 -2347 -1286
rect -2313 -1320 -2267 -1286
rect -2233 -1320 -2187 -1286
rect -2153 -1320 -2107 -1286
rect -2073 -1320 -2027 -1286
rect -1993 -1320 -1947 -1286
rect -1913 -1320 -1867 -1286
rect -1833 -1320 -1787 -1286
rect -1753 -1320 -1707 -1286
rect -1673 -1320 -1590 -1286
rect -3870 -1353 -1590 -1320
rect -1230 -1286 150 -1253
rect -1230 -1320 -1197 -1286
rect -1163 -1320 -1117 -1286
rect -1083 -1320 -1037 -1286
rect -1003 -1320 -957 -1286
rect -923 -1320 -877 -1286
rect -843 -1320 -797 -1286
rect -763 -1320 -717 -1286
rect -683 -1320 -637 -1286
rect -603 -1320 -557 -1286
rect -523 -1320 -477 -1286
rect -443 -1320 -397 -1286
rect -363 -1320 -317 -1286
rect -283 -1320 -237 -1286
rect -203 -1320 -157 -1286
rect -123 -1320 -77 -1286
rect -43 -1320 3 -1286
rect 37 -1320 83 -1286
rect 117 -1320 150 -1286
rect -1230 -1353 150 -1320
rect 500 -1286 2180 -1253
rect 500 -1320 523 -1286
rect 557 -1320 603 -1286
rect 637 -1320 683 -1286
rect 717 -1320 763 -1286
rect 797 -1320 843 -1286
rect 877 -1320 923 -1286
rect 957 -1320 1003 -1286
rect 1037 -1320 1083 -1286
rect 1117 -1320 1163 -1286
rect 1197 -1320 1243 -1286
rect 1277 -1320 1323 -1286
rect 1357 -1320 1403 -1286
rect 1437 -1320 1483 -1286
rect 1517 -1320 1563 -1286
rect 1597 -1320 1643 -1286
rect 1677 -1320 1723 -1286
rect 1757 -1320 1803 -1286
rect 1837 -1320 1883 -1286
rect 1917 -1320 1963 -1286
rect 1997 -1320 2043 -1286
rect 2077 -1320 2123 -1286
rect 2157 -1320 2180 -1286
rect 500 -1353 2180 -1320
rect -3729 -1746 -1729 -1713
rect -3729 -1780 -3706 -1746
rect -3672 -1780 -3626 -1746
rect -3592 -1780 -3546 -1746
rect -3512 -1780 -3466 -1746
rect -3432 -1780 -3386 -1746
rect -3352 -1780 -3306 -1746
rect -3272 -1780 -3226 -1746
rect -3192 -1780 -3146 -1746
rect -3112 -1780 -3066 -1746
rect -3032 -1780 -2986 -1746
rect -2952 -1780 -2906 -1746
rect -2872 -1780 -2826 -1746
rect -2792 -1780 -2746 -1746
rect -2712 -1780 -2666 -1746
rect -2632 -1780 -2586 -1746
rect -2552 -1780 -2506 -1746
rect -2472 -1780 -2426 -1746
rect -2392 -1780 -2346 -1746
rect -2312 -1780 -2266 -1746
rect -2232 -1780 -2186 -1746
rect -2152 -1780 -2106 -1746
rect -2072 -1780 -2026 -1746
rect -1992 -1780 -1946 -1746
rect -1912 -1780 -1866 -1746
rect -1832 -1780 -1786 -1746
rect -1752 -1780 -1729 -1746
rect -3729 -1813 -1729 -1780
rect -1369 -1746 11 -1713
rect -1369 -1780 -1336 -1746
rect -1302 -1780 -1256 -1746
rect -1222 -1780 -1176 -1746
rect -1142 -1780 -1096 -1746
rect -1062 -1780 -1016 -1746
rect -982 -1780 -936 -1746
rect -902 -1780 -856 -1746
rect -822 -1780 -776 -1746
rect -742 -1780 -696 -1746
rect -662 -1780 -616 -1746
rect -582 -1780 -536 -1746
rect -502 -1780 -456 -1746
rect -422 -1780 -376 -1746
rect -342 -1780 -296 -1746
rect -262 -1780 -216 -1746
rect -182 -1780 -136 -1746
rect -102 -1780 -56 -1746
rect -22 -1780 11 -1746
rect -1369 -1813 11 -1780
rect 361 -1747 2361 -1714
rect 361 -1781 384 -1747
rect 418 -1781 464 -1747
rect 498 -1781 544 -1747
rect 578 -1781 624 -1747
rect 658 -1781 704 -1747
rect 738 -1781 784 -1747
rect 818 -1781 864 -1747
rect 898 -1781 944 -1747
rect 978 -1781 1024 -1747
rect 1058 -1781 1104 -1747
rect 1138 -1781 1184 -1747
rect 1218 -1781 1264 -1747
rect 1298 -1781 1344 -1747
rect 1378 -1781 1424 -1747
rect 1458 -1781 1504 -1747
rect 1538 -1781 1584 -1747
rect 1618 -1781 1664 -1747
rect 1698 -1781 1744 -1747
rect 1778 -1781 1824 -1747
rect 1858 -1781 1904 -1747
rect 1938 -1781 1984 -1747
rect 2018 -1781 2064 -1747
rect 2098 -1781 2144 -1747
rect 2178 -1781 2224 -1747
rect 2258 -1781 2304 -1747
rect 2338 -1781 2361 -1747
rect 361 -1814 2361 -1781
<< psubdiffcont >>
rect -3787 -140 -3753 -106
rect -3707 -140 -3673 -106
rect -3627 -140 -3593 -106
rect -3547 -140 -3513 -106
rect -3467 -140 -3433 -106
rect -3387 -140 -3353 -106
rect -3307 -140 -3273 -106
rect -3227 -140 -3193 -106
rect -3147 -140 -3113 -106
rect -3067 -140 -3033 -106
rect -2987 -140 -2953 -106
rect -2907 -140 -2873 -106
rect -2827 -140 -2793 -106
rect -2747 -140 -2713 -106
rect -2667 -140 -2633 -106
rect -2587 -140 -2553 -106
rect -2507 -140 -2473 -106
rect -2427 -140 -2393 -106
rect -2347 -140 -2313 -106
rect -2267 -140 -2233 -106
rect -2187 -140 -2153 -106
rect -2107 -140 -2073 -106
rect -2027 -140 -1993 -106
rect -1947 -140 -1913 -106
rect -1867 -140 -1833 -106
rect -1787 -140 -1753 -106
rect -1707 -140 -1673 -106
rect -1197 -140 -1163 -106
rect -1117 -140 -1083 -106
rect -1037 -140 -1003 -106
rect -957 -140 -923 -106
rect -877 -140 -843 -106
rect -797 -140 -763 -106
rect -717 -140 -683 -106
rect -637 -140 -603 -106
rect -557 -140 -523 -106
rect -477 -140 -443 -106
rect -397 -140 -363 -106
rect -317 -140 -283 -106
rect -237 -140 -203 -106
rect -157 -140 -123 -106
rect -77 -140 -43 -106
rect 3 -140 37 -106
rect 83 -140 117 -106
rect 523 -140 557 -106
rect 603 -140 637 -106
rect 683 -140 717 -106
rect 763 -140 797 -106
rect 843 -140 877 -106
rect 923 -140 957 -106
rect 1003 -140 1037 -106
rect 1083 -140 1117 -106
rect 1163 -140 1197 -106
rect 1243 -140 1277 -106
rect 1323 -140 1357 -106
rect 1403 -140 1437 -106
rect 1483 -140 1517 -106
rect 1563 -140 1597 -106
rect 1643 -140 1677 -106
rect 1723 -140 1757 -106
rect 1803 -140 1837 -106
rect 1883 -140 1917 -106
rect 1963 -140 1997 -106
rect 2043 -140 2077 -106
rect 2123 -140 2157 -106
rect -3706 -2960 -3672 -2926
rect -3626 -2960 -3592 -2926
rect -3546 -2960 -3512 -2926
rect -3466 -2960 -3432 -2926
rect -3386 -2960 -3352 -2926
rect -3306 -2960 -3272 -2926
rect -3226 -2960 -3192 -2926
rect -3146 -2960 -3112 -2926
rect -3066 -2960 -3032 -2926
rect -2986 -2960 -2952 -2926
rect -2906 -2960 -2872 -2926
rect -2826 -2960 -2792 -2926
rect -2746 -2960 -2712 -2926
rect -2666 -2960 -2632 -2926
rect -2586 -2960 -2552 -2926
rect -2506 -2960 -2472 -2926
rect -2426 -2960 -2392 -2926
rect -2346 -2960 -2312 -2926
rect -2266 -2960 -2232 -2926
rect -2186 -2960 -2152 -2926
rect -2106 -2960 -2072 -2926
rect -2026 -2960 -1992 -2926
rect -1946 -2960 -1912 -2926
rect -1866 -2960 -1832 -2926
rect -1786 -2960 -1752 -2926
rect -1336 -2960 -1302 -2926
rect -1256 -2960 -1222 -2926
rect -1176 -2960 -1142 -2926
rect -1096 -2960 -1062 -2926
rect -1016 -2960 -982 -2926
rect -936 -2960 -902 -2926
rect -856 -2960 -822 -2926
rect -776 -2960 -742 -2926
rect -696 -2960 -662 -2926
rect -616 -2960 -582 -2926
rect -536 -2960 -502 -2926
rect -456 -2960 -422 -2926
rect -376 -2960 -342 -2926
rect -296 -2960 -262 -2926
rect -216 -2960 -182 -2926
rect -136 -2960 -102 -2926
rect -56 -2960 -22 -2926
rect 384 -2961 418 -2927
rect 464 -2961 498 -2927
rect 544 -2961 578 -2927
rect 624 -2961 658 -2927
rect 704 -2961 738 -2927
rect 784 -2961 818 -2927
rect 864 -2961 898 -2927
rect 944 -2961 978 -2927
rect 1024 -2961 1058 -2927
rect 1104 -2961 1138 -2927
rect 1184 -2961 1218 -2927
rect 1264 -2961 1298 -2927
rect 1344 -2961 1378 -2927
rect 1424 -2961 1458 -2927
rect 1504 -2961 1538 -2927
rect 1584 -2961 1618 -2927
rect 1664 -2961 1698 -2927
rect 1744 -2961 1778 -2927
rect 1824 -2961 1858 -2927
rect 1904 -2961 1938 -2927
rect 1984 -2961 2018 -2927
rect 2064 -2961 2098 -2927
rect 2144 -2961 2178 -2927
rect 2224 -2961 2258 -2927
rect 2304 -2961 2338 -2927
<< nsubdiffcont >>
rect -3787 1040 -3753 1074
rect -3707 1040 -3673 1074
rect -3627 1040 -3593 1074
rect -3547 1040 -3513 1074
rect -3467 1040 -3433 1074
rect -3387 1040 -3353 1074
rect -3307 1040 -3273 1074
rect -3227 1040 -3193 1074
rect -3147 1040 -3113 1074
rect -3067 1040 -3033 1074
rect -2987 1040 -2953 1074
rect -2907 1040 -2873 1074
rect -2827 1040 -2793 1074
rect -2747 1040 -2713 1074
rect -2667 1040 -2633 1074
rect -2587 1040 -2553 1074
rect -2507 1040 -2473 1074
rect -2427 1040 -2393 1074
rect -2347 1040 -2313 1074
rect -2267 1040 -2233 1074
rect -2187 1040 -2153 1074
rect -2107 1040 -2073 1074
rect -2027 1040 -1993 1074
rect -1947 1040 -1913 1074
rect -1867 1040 -1833 1074
rect -1787 1040 -1753 1074
rect -1707 1040 -1673 1074
rect -1197 1040 -1163 1074
rect -1117 1040 -1083 1074
rect -1037 1040 -1003 1074
rect -957 1040 -923 1074
rect -877 1040 -843 1074
rect -797 1040 -763 1074
rect -717 1040 -683 1074
rect -637 1040 -603 1074
rect -557 1040 -523 1074
rect -477 1040 -443 1074
rect -397 1040 -363 1074
rect -317 1040 -283 1074
rect -237 1040 -203 1074
rect -157 1040 -123 1074
rect -77 1040 -43 1074
rect 3 1040 37 1074
rect 83 1040 117 1074
rect 523 1040 557 1074
rect 603 1040 637 1074
rect 683 1040 717 1074
rect 763 1040 797 1074
rect 843 1040 877 1074
rect 923 1040 957 1074
rect 1003 1040 1037 1074
rect 1083 1040 1117 1074
rect 1163 1040 1197 1074
rect 1243 1040 1277 1074
rect 1323 1040 1357 1074
rect 1403 1040 1437 1074
rect 1483 1040 1517 1074
rect 1563 1040 1597 1074
rect 1643 1040 1677 1074
rect 1723 1040 1757 1074
rect 1803 1040 1837 1074
rect 1883 1040 1917 1074
rect 1963 1040 1997 1074
rect 2043 1040 2077 1074
rect 2123 1040 2157 1074
rect -3787 -1320 -3753 -1286
rect -3707 -1320 -3673 -1286
rect -3627 -1320 -3593 -1286
rect -3547 -1320 -3513 -1286
rect -3467 -1320 -3433 -1286
rect -3387 -1320 -3353 -1286
rect -3307 -1320 -3273 -1286
rect -3227 -1320 -3193 -1286
rect -3147 -1320 -3113 -1286
rect -3067 -1320 -3033 -1286
rect -2987 -1320 -2953 -1286
rect -2907 -1320 -2873 -1286
rect -2827 -1320 -2793 -1286
rect -2747 -1320 -2713 -1286
rect -2667 -1320 -2633 -1286
rect -2587 -1320 -2553 -1286
rect -2507 -1320 -2473 -1286
rect -2427 -1320 -2393 -1286
rect -2347 -1320 -2313 -1286
rect -2267 -1320 -2233 -1286
rect -2187 -1320 -2153 -1286
rect -2107 -1320 -2073 -1286
rect -2027 -1320 -1993 -1286
rect -1947 -1320 -1913 -1286
rect -1867 -1320 -1833 -1286
rect -1787 -1320 -1753 -1286
rect -1707 -1320 -1673 -1286
rect -1197 -1320 -1163 -1286
rect -1117 -1320 -1083 -1286
rect -1037 -1320 -1003 -1286
rect -957 -1320 -923 -1286
rect -877 -1320 -843 -1286
rect -797 -1320 -763 -1286
rect -717 -1320 -683 -1286
rect -637 -1320 -603 -1286
rect -557 -1320 -523 -1286
rect -477 -1320 -443 -1286
rect -397 -1320 -363 -1286
rect -317 -1320 -283 -1286
rect -237 -1320 -203 -1286
rect -157 -1320 -123 -1286
rect -77 -1320 -43 -1286
rect 3 -1320 37 -1286
rect 83 -1320 117 -1286
rect 523 -1320 557 -1286
rect 603 -1320 637 -1286
rect 683 -1320 717 -1286
rect 763 -1320 797 -1286
rect 843 -1320 877 -1286
rect 923 -1320 957 -1286
rect 1003 -1320 1037 -1286
rect 1083 -1320 1117 -1286
rect 1163 -1320 1197 -1286
rect 1243 -1320 1277 -1286
rect 1323 -1320 1357 -1286
rect 1403 -1320 1437 -1286
rect 1483 -1320 1517 -1286
rect 1563 -1320 1597 -1286
rect 1643 -1320 1677 -1286
rect 1723 -1320 1757 -1286
rect 1803 -1320 1837 -1286
rect 1883 -1320 1917 -1286
rect 1963 -1320 1997 -1286
rect 2043 -1320 2077 -1286
rect 2123 -1320 2157 -1286
rect -3706 -1780 -3672 -1746
rect -3626 -1780 -3592 -1746
rect -3546 -1780 -3512 -1746
rect -3466 -1780 -3432 -1746
rect -3386 -1780 -3352 -1746
rect -3306 -1780 -3272 -1746
rect -3226 -1780 -3192 -1746
rect -3146 -1780 -3112 -1746
rect -3066 -1780 -3032 -1746
rect -2986 -1780 -2952 -1746
rect -2906 -1780 -2872 -1746
rect -2826 -1780 -2792 -1746
rect -2746 -1780 -2712 -1746
rect -2666 -1780 -2632 -1746
rect -2586 -1780 -2552 -1746
rect -2506 -1780 -2472 -1746
rect -2426 -1780 -2392 -1746
rect -2346 -1780 -2312 -1746
rect -2266 -1780 -2232 -1746
rect -2186 -1780 -2152 -1746
rect -2106 -1780 -2072 -1746
rect -2026 -1780 -1992 -1746
rect -1946 -1780 -1912 -1746
rect -1866 -1780 -1832 -1746
rect -1786 -1780 -1752 -1746
rect -1336 -1780 -1302 -1746
rect -1256 -1780 -1222 -1746
rect -1176 -1780 -1142 -1746
rect -1096 -1780 -1062 -1746
rect -1016 -1780 -982 -1746
rect -936 -1780 -902 -1746
rect -856 -1780 -822 -1746
rect -776 -1780 -742 -1746
rect -696 -1780 -662 -1746
rect -616 -1780 -582 -1746
rect -536 -1780 -502 -1746
rect -456 -1780 -422 -1746
rect -376 -1780 -342 -1746
rect -296 -1780 -262 -1746
rect -216 -1780 -182 -1746
rect -136 -1780 -102 -1746
rect -56 -1780 -22 -1746
rect 384 -1781 418 -1747
rect 464 -1781 498 -1747
rect 544 -1781 578 -1747
rect 624 -1781 658 -1747
rect 704 -1781 738 -1747
rect 784 -1781 818 -1747
rect 864 -1781 898 -1747
rect 944 -1781 978 -1747
rect 1024 -1781 1058 -1747
rect 1104 -1781 1138 -1747
rect 1184 -1781 1218 -1747
rect 1264 -1781 1298 -1747
rect 1344 -1781 1378 -1747
rect 1424 -1781 1458 -1747
rect 1504 -1781 1538 -1747
rect 1584 -1781 1618 -1747
rect 1664 -1781 1698 -1747
rect 1744 -1781 1778 -1747
rect 1824 -1781 1858 -1747
rect 1904 -1781 1938 -1747
rect 1984 -1781 2018 -1747
rect 2064 -1781 2098 -1747
rect 2144 -1781 2178 -1747
rect 2224 -1781 2258 -1747
rect 2304 -1781 2338 -1747
<< poly >>
rect -3480 944 -3400 967
rect -3480 910 -3457 944
rect -3423 910 -3400 944
rect -2970 957 -2790 987
rect -2970 927 -2940 957
rect -2820 927 -2790 957
rect -2670 957 -2490 987
rect -2670 927 -2640 957
rect -2520 927 -2490 957
rect -2090 944 -2010 967
rect -3480 887 -3400 910
rect -3600 844 -3520 867
rect -3600 810 -3577 844
rect -3543 810 -3520 844
rect -3600 787 -3520 810
rect -3800 644 -3720 667
rect -3800 610 -3777 644
rect -3743 610 -3720 644
rect -3800 587 -3720 610
rect -3750 367 -3720 587
rect -3600 367 -3570 787
rect -3450 367 -3420 887
rect -3350 744 -3270 767
rect -3350 710 -3327 744
rect -3293 710 -3270 744
rect -3350 687 -3270 710
rect -3300 367 -3270 687
rect -2090 910 -2067 944
rect -2033 910 -2010 944
rect -780 957 -600 987
rect -780 927 -750 957
rect -630 927 -600 957
rect -480 957 -300 987
rect -480 927 -450 957
rect -330 927 -300 957
rect 1100 957 1280 987
rect 1100 927 1130 957
rect 1250 927 1280 957
rect 1400 957 1580 987
rect 1400 927 1430 957
rect 1550 927 1580 957
rect -2090 887 -2010 910
rect -2190 644 -2110 667
rect -2970 597 -2940 627
rect -2820 472 -2790 627
rect -2670 597 -2640 627
rect -2520 597 -2490 627
rect -2190 610 -2167 644
rect -2133 610 -2110 644
rect -2720 574 -2640 597
rect -2720 540 -2697 574
rect -2663 540 -2640 574
rect -2720 517 -2640 540
rect -2820 449 -2740 472
rect -2820 415 -2797 449
rect -2763 415 -2740 449
rect -2970 367 -2940 397
rect -2820 392 -2740 415
rect -2820 367 -2790 392
rect -2670 367 -2640 517
rect -2190 587 -2110 610
rect -2520 367 -2490 397
rect -2190 367 -2160 587
rect -2040 367 -2010 887
rect -1890 844 -1810 867
rect -1890 810 -1867 844
rect -1833 810 -1810 844
rect -1890 787 -1810 810
rect -1890 367 -1860 787
rect -1740 744 -1660 767
rect -1740 710 -1717 744
rect -1683 710 -1660 744
rect -1740 687 -1660 710
rect -1740 367 -1710 687
rect 0 694 80 717
rect 0 660 23 694
rect 57 660 80 694
rect 0 637 80 660
rect -780 597 -750 627
rect -1160 454 -1080 477
rect -1160 420 -1137 454
rect -1103 420 -1080 454
rect -1160 397 -1080 420
rect -630 472 -600 627
rect -480 597 -450 627
rect -330 597 -300 627
rect -530 574 -450 597
rect -530 540 -507 574
rect -473 540 -450 574
rect -530 517 -450 540
rect -630 449 -550 472
rect -630 415 -607 449
rect -573 415 -550 449
rect -1110 367 -1080 397
rect -780 367 -750 397
rect -630 392 -550 415
rect -630 367 -600 392
rect -480 367 -450 517
rect -330 367 -300 397
rect 0 367 30 637
rect 720 624 800 647
rect 1980 844 2060 867
rect 1980 810 2003 844
rect 2037 810 2060 844
rect 1980 787 2060 810
rect 1830 724 1910 747
rect 1830 690 1853 724
rect 1887 690 1910 724
rect 1830 667 1910 690
rect 720 590 743 624
rect 777 590 800 624
rect 1100 597 1130 627
rect 720 567 800 590
rect 570 524 650 547
rect 570 490 593 524
rect 627 490 650 524
rect 570 467 650 490
rect 620 367 650 467
rect 770 367 800 567
rect 1250 472 1280 627
rect 1400 597 1430 627
rect 1550 597 1580 627
rect 1350 574 1430 597
rect 1350 540 1373 574
rect 1407 540 1430 574
rect 1350 517 1430 540
rect 1250 449 1330 472
rect 1250 415 1273 449
rect 1307 415 1330 449
rect 1100 367 1130 397
rect 1250 392 1330 415
rect 1250 367 1280 392
rect 1400 367 1430 517
rect 1550 367 1580 397
rect 1880 367 1910 667
rect 2030 367 2060 787
rect -3750 37 -3720 67
rect -3600 37 -3570 67
rect -3450 37 -3420 67
rect -3300 37 -3270 67
rect -2970 37 -2940 67
rect -2820 37 -2790 67
rect -2670 37 -2640 67
rect -2520 37 -2490 67
rect -2190 37 -2160 67
rect -2970 14 -2890 37
rect -2970 -20 -2947 14
rect -2913 -20 -2890 14
rect -2970 -43 -2890 -20
rect -2570 14 -2490 37
rect -2040 27 -2010 67
rect -1890 27 -1860 67
rect -1740 27 -1710 67
rect -1110 37 -1080 67
rect -780 37 -750 67
rect -630 37 -600 67
rect -480 37 -450 67
rect -330 37 -300 67
rect 0 37 30 67
rect 620 37 650 67
rect 770 37 800 67
rect 1100 37 1130 67
rect 1250 37 1280 67
rect 1400 37 1430 67
rect 1550 37 1580 67
rect 1880 37 1910 67
rect 2030 37 2060 67
rect -2570 -20 -2547 14
rect -2513 -20 -2490 14
rect -2570 -43 -2490 -20
rect -780 14 -700 37
rect -780 -20 -757 14
rect -723 -20 -700 14
rect -780 -43 -700 -20
rect -380 14 -300 37
rect -380 -20 -357 14
rect -323 -20 -300 14
rect -380 -43 -300 -20
rect 1100 14 1180 37
rect 1100 -20 1123 14
rect 1157 -20 1180 14
rect 1100 -43 1180 -20
rect 1500 14 1580 37
rect 1500 -20 1523 14
rect 1557 -20 1580 14
rect 1500 -43 1580 -20
rect -2970 -226 -2890 -203
rect -2970 -260 -2947 -226
rect -2913 -260 -2890 -226
rect -2970 -283 -2890 -260
rect -2570 -226 -2490 -203
rect -2570 -260 -2547 -226
rect -2513 -260 -2490 -226
rect -2570 -283 -2490 -260
rect -780 -226 -700 -203
rect -780 -260 -757 -226
rect -723 -260 -700 -226
rect -3750 -313 -3720 -283
rect -3600 -313 -3570 -283
rect -3450 -313 -3420 -283
rect -3300 -313 -3270 -283
rect -2970 -313 -2940 -283
rect -2820 -313 -2790 -283
rect -2670 -313 -2640 -283
rect -2520 -313 -2490 -283
rect -2190 -313 -2160 -283
rect -2040 -313 -2010 -273
rect -1890 -313 -1860 -273
rect -1740 -313 -1710 -273
rect -780 -283 -700 -260
rect -380 -226 -300 -203
rect -380 -260 -357 -226
rect -323 -260 -300 -226
rect -380 -283 -300 -260
rect 1100 -226 1180 -203
rect 1100 -260 1123 -226
rect 1157 -260 1180 -226
rect 1100 -283 1180 -260
rect 1500 -226 1580 -203
rect 1500 -260 1523 -226
rect 1557 -260 1580 -226
rect 1500 -283 1580 -260
rect -1110 -313 -1080 -283
rect -780 -313 -750 -283
rect -630 -313 -600 -283
rect -480 -313 -450 -283
rect -330 -313 -300 -283
rect 0 -313 30 -283
rect 620 -313 650 -283
rect 770 -313 800 -283
rect 1100 -313 1130 -283
rect 1250 -313 1280 -283
rect 1400 -313 1430 -283
rect 1550 -313 1580 -283
rect 1880 -313 1910 -283
rect 2030 -313 2060 -283
rect -3750 -833 -3720 -613
rect -3800 -856 -3720 -833
rect -3800 -890 -3777 -856
rect -3743 -890 -3720 -856
rect -3800 -913 -3720 -890
rect -3600 -1033 -3570 -613
rect -3600 -1056 -3520 -1033
rect -3600 -1090 -3577 -1056
rect -3543 -1090 -3520 -1056
rect -3600 -1113 -3520 -1090
rect -3450 -1133 -3420 -613
rect -3300 -933 -3270 -613
rect -2970 -643 -2940 -613
rect -2820 -638 -2790 -613
rect -2820 -661 -2740 -638
rect -2820 -695 -2797 -661
rect -2763 -695 -2740 -661
rect -2820 -718 -2740 -695
rect -2970 -873 -2940 -843
rect -2820 -873 -2790 -718
rect -2670 -763 -2640 -613
rect -2520 -643 -2490 -613
rect -2720 -786 -2640 -763
rect -2720 -820 -2697 -786
rect -2663 -820 -2640 -786
rect -2720 -843 -2640 -820
rect -2190 -833 -2160 -613
rect -2670 -873 -2640 -843
rect -2520 -873 -2490 -843
rect -2190 -856 -2110 -833
rect -3350 -956 -3270 -933
rect -3350 -990 -3327 -956
rect -3293 -990 -3270 -956
rect -3350 -1013 -3270 -990
rect -3480 -1156 -3400 -1133
rect -3480 -1190 -3457 -1156
rect -3423 -1190 -3400 -1156
rect -2190 -890 -2167 -856
rect -2133 -890 -2110 -856
rect -2190 -913 -2110 -890
rect -2040 -1133 -2010 -613
rect -1890 -1033 -1860 -613
rect -1740 -933 -1710 -613
rect -1110 -643 -1080 -613
rect -780 -643 -750 -613
rect -630 -638 -600 -613
rect -1160 -666 -1080 -643
rect -1160 -700 -1137 -666
rect -1103 -700 -1080 -666
rect -1160 -723 -1080 -700
rect -630 -661 -550 -638
rect -630 -695 -607 -661
rect -573 -695 -550 -661
rect -630 -718 -550 -695
rect -780 -873 -750 -843
rect -630 -873 -600 -718
rect -480 -763 -450 -613
rect -330 -643 -300 -613
rect -530 -786 -450 -763
rect -530 -820 -507 -786
rect -473 -820 -450 -786
rect -530 -843 -450 -820
rect -480 -873 -450 -843
rect -330 -873 -300 -843
rect -1740 -956 -1660 -933
rect -1740 -990 -1717 -956
rect -1683 -990 -1660 -956
rect -1740 -1013 -1660 -990
rect -1890 -1056 -1810 -1033
rect -1890 -1090 -1867 -1056
rect -1833 -1090 -1810 -1056
rect -1890 -1113 -1810 -1090
rect -2090 -1156 -2010 -1133
rect -3480 -1213 -3400 -1190
rect -2970 -1203 -2940 -1173
rect -2820 -1203 -2790 -1173
rect -2970 -1233 -2790 -1203
rect -2670 -1203 -2640 -1173
rect -2520 -1203 -2490 -1173
rect -2670 -1233 -2490 -1203
rect -2090 -1190 -2067 -1156
rect -2033 -1190 -2010 -1156
rect 0 -883 30 -613
rect 620 -713 650 -613
rect 570 -736 650 -713
rect 570 -770 593 -736
rect 627 -770 650 -736
rect 570 -793 650 -770
rect 770 -813 800 -613
rect 1100 -643 1130 -613
rect 1250 -638 1280 -613
rect 720 -836 800 -813
rect 720 -870 743 -836
rect 777 -870 800 -836
rect 1250 -661 1330 -638
rect 1250 -695 1273 -661
rect 1307 -695 1330 -661
rect 1250 -718 1330 -695
rect 0 -906 80 -883
rect 720 -893 800 -870
rect 1100 -873 1130 -843
rect 1250 -873 1280 -718
rect 1400 -763 1430 -613
rect 1550 -643 1580 -613
rect 1350 -786 1430 -763
rect 1350 -820 1373 -786
rect 1407 -820 1430 -786
rect 1350 -843 1430 -820
rect 1400 -873 1430 -843
rect 1550 -873 1580 -843
rect 0 -940 23 -906
rect 57 -940 80 -906
rect 0 -963 80 -940
rect 1880 -913 1910 -613
rect 1830 -936 1910 -913
rect 1830 -970 1853 -936
rect 1887 -970 1910 -936
rect 1830 -993 1910 -970
rect 2030 -1033 2060 -613
rect 1980 -1056 2060 -1033
rect 1980 -1090 2003 -1056
rect 2037 -1090 2060 -1056
rect 1980 -1113 2060 -1090
rect -2090 -1213 -2010 -1190
rect -780 -1203 -750 -1173
rect -630 -1203 -600 -1173
rect -780 -1233 -600 -1203
rect -480 -1203 -450 -1173
rect -330 -1203 -300 -1173
rect -480 -1233 -300 -1203
rect 1100 -1203 1130 -1173
rect 1250 -1203 1280 -1173
rect 1100 -1233 1280 -1203
rect 1400 -1203 1430 -1173
rect 1550 -1203 1580 -1173
rect 1400 -1233 1580 -1203
rect -2969 -1863 -2789 -1833
rect -2969 -1893 -2939 -1863
rect -2819 -1893 -2789 -1863
rect -2669 -1863 -2489 -1833
rect -2669 -1893 -2639 -1863
rect -2519 -1893 -2489 -1863
rect -1939 -1866 -1859 -1843
rect -1939 -1900 -1916 -1866
rect -1882 -1900 -1859 -1866
rect -919 -1863 -739 -1833
rect -919 -1893 -889 -1863
rect -769 -1893 -739 -1863
rect -619 -1863 -439 -1833
rect -619 -1893 -589 -1863
rect -469 -1893 -439 -1863
rect 491 -1872 571 -1849
rect -1939 -1923 -1859 -1900
rect -2089 -1986 -2009 -1963
rect -2089 -2020 -2066 -1986
rect -2032 -2020 -2009 -1986
rect -2089 -2043 -2009 -2020
rect -2219 -2106 -2139 -2083
rect -2219 -2140 -2196 -2106
rect -2162 -2140 -2139 -2106
rect -2219 -2163 -2139 -2140
rect -2969 -2223 -2939 -2193
rect -3519 -2276 -3419 -2253
rect -3519 -2310 -3496 -2276
rect -3462 -2310 -3419 -2276
rect -3519 -2333 -3419 -2310
rect -3349 -2256 -3269 -2233
rect -3349 -2290 -3326 -2256
rect -3292 -2290 -3269 -2256
rect -3349 -2313 -3269 -2290
rect -3649 -2356 -3569 -2333
rect -3649 -2390 -3626 -2356
rect -3592 -2390 -3569 -2356
rect -3649 -2413 -3569 -2390
rect -3599 -2453 -3569 -2413
rect -3449 -2453 -3419 -2333
rect -3299 -2453 -3269 -2313
rect -2819 -2348 -2789 -2193
rect -2669 -2223 -2639 -2193
rect -2519 -2223 -2489 -2193
rect -2719 -2246 -2639 -2223
rect -2719 -2280 -2696 -2246
rect -2662 -2280 -2639 -2246
rect -2719 -2303 -2639 -2280
rect -2819 -2371 -2739 -2348
rect -2819 -2405 -2796 -2371
rect -2762 -2405 -2739 -2371
rect -2969 -2453 -2939 -2423
rect -2819 -2428 -2739 -2405
rect -2819 -2453 -2789 -2428
rect -2669 -2453 -2639 -2303
rect -2519 -2453 -2489 -2423
rect -2189 -2453 -2159 -2163
rect -2039 -2453 -2009 -2043
rect -1889 -2453 -1859 -1923
rect 491 -1906 514 -1872
rect 548 -1906 571 -1872
rect 1121 -1864 1301 -1834
rect 1121 -1894 1151 -1864
rect 1271 -1894 1301 -1864
rect 1421 -1864 1601 -1834
rect 1421 -1894 1451 -1864
rect 1571 -1894 1601 -1864
rect 491 -1929 571 -1906
rect -139 -2126 -59 -2103
rect -139 -2160 -116 -2126
rect -82 -2160 -59 -2126
rect -139 -2183 -59 -2160
rect -919 -2223 -889 -2193
rect -1299 -2366 -1219 -2343
rect -1299 -2400 -1276 -2366
rect -1242 -2400 -1219 -2366
rect -1299 -2423 -1219 -2400
rect -769 -2348 -739 -2193
rect -619 -2223 -589 -2193
rect -469 -2223 -439 -2193
rect -669 -2246 -589 -2223
rect -669 -2280 -646 -2246
rect -612 -2280 -589 -2246
rect -669 -2303 -589 -2280
rect -769 -2371 -689 -2348
rect -769 -2405 -746 -2371
rect -712 -2405 -689 -2371
rect -1249 -2453 -1219 -2423
rect -919 -2453 -889 -2423
rect -769 -2428 -689 -2405
rect -769 -2453 -739 -2428
rect -619 -2453 -589 -2303
rect -469 -2453 -439 -2423
rect -139 -2453 -109 -2183
rect 491 -2454 521 -1929
rect 591 -1997 671 -1974
rect 591 -2031 614 -1997
rect 648 -2031 671 -1997
rect 591 -2054 671 -2031
rect 641 -2454 671 -2054
rect 791 -2087 871 -2064
rect 791 -2121 814 -2087
rect 848 -2121 871 -2087
rect 791 -2144 871 -2121
rect 791 -2454 821 -2144
rect 1121 -2224 1151 -2194
rect 1271 -2224 1301 -2194
rect 1271 -2247 1351 -2224
rect 1271 -2281 1294 -2247
rect 1328 -2281 1351 -2247
rect 1271 -2304 1351 -2281
rect 1121 -2454 1151 -2424
rect 1271 -2454 1301 -2304
rect 1421 -2349 1451 -2194
rect 1571 -2224 1601 -2194
rect 2191 -2197 2271 -2174
rect 2191 -2231 2214 -2197
rect 2248 -2231 2271 -2197
rect 2191 -2254 2271 -2231
rect 1371 -2372 1451 -2349
rect 2051 -2297 2131 -2274
rect 2051 -2331 2074 -2297
rect 2108 -2331 2131 -2297
rect 2051 -2354 2131 -2331
rect 1371 -2406 1394 -2372
rect 1428 -2406 1451 -2372
rect 1371 -2429 1451 -2406
rect 1901 -2377 1981 -2354
rect 1901 -2411 1924 -2377
rect 1958 -2411 1981 -2377
rect 1421 -2454 1451 -2429
rect 1571 -2454 1601 -2424
rect 1901 -2434 1981 -2411
rect 1901 -2454 1931 -2434
rect 2051 -2454 2081 -2354
rect 2201 -2454 2231 -2254
rect -3599 -2783 -3569 -2753
rect -3449 -2783 -3419 -2753
rect -3299 -2783 -3269 -2753
rect -2969 -2783 -2939 -2753
rect -2819 -2783 -2789 -2753
rect -2669 -2783 -2639 -2753
rect -2519 -2783 -2489 -2753
rect -2189 -2783 -2159 -2753
rect -2039 -2783 -2009 -2753
rect -1889 -2783 -1859 -2753
rect -1249 -2783 -1219 -2753
rect -919 -2783 -889 -2753
rect -769 -2783 -739 -2753
rect -619 -2783 -589 -2753
rect -469 -2783 -439 -2753
rect -139 -2783 -109 -2753
rect -2969 -2806 -2889 -2783
rect -2969 -2840 -2946 -2806
rect -2912 -2840 -2889 -2806
rect -2969 -2863 -2889 -2840
rect -2569 -2806 -2489 -2783
rect -2569 -2840 -2546 -2806
rect -2512 -2840 -2489 -2806
rect -2569 -2863 -2489 -2840
rect -919 -2806 -839 -2783
rect -919 -2840 -896 -2806
rect -862 -2840 -839 -2806
rect -919 -2863 -839 -2840
rect -519 -2806 -439 -2783
rect 491 -2784 521 -2754
rect 641 -2784 671 -2754
rect 791 -2784 821 -2754
rect 1121 -2784 1151 -2754
rect 1271 -2784 1301 -2754
rect 1421 -2784 1451 -2754
rect 1571 -2784 1601 -2754
rect 1901 -2784 1931 -2754
rect 2051 -2784 2081 -2754
rect 2201 -2784 2231 -2754
rect -519 -2840 -496 -2806
rect -462 -2840 -439 -2806
rect -519 -2863 -439 -2840
rect 1121 -2807 1201 -2784
rect 1121 -2841 1144 -2807
rect 1178 -2841 1201 -2807
rect 1121 -2864 1201 -2841
rect 1521 -2807 1601 -2784
rect 1521 -2841 1544 -2807
rect 1578 -2841 1601 -2807
rect 1521 -2864 1601 -2841
<< polycont >>
rect -3457 910 -3423 944
rect -3577 810 -3543 844
rect -3777 610 -3743 644
rect -3327 710 -3293 744
rect -2067 910 -2033 944
rect -2167 610 -2133 644
rect -2697 540 -2663 574
rect -2797 415 -2763 449
rect -1867 810 -1833 844
rect -1717 710 -1683 744
rect 23 660 57 694
rect -1137 420 -1103 454
rect -507 540 -473 574
rect -607 415 -573 449
rect 2003 810 2037 844
rect 1853 690 1887 724
rect 743 590 777 624
rect 593 490 627 524
rect 1373 540 1407 574
rect 1273 415 1307 449
rect -2947 -20 -2913 14
rect -2547 -20 -2513 14
rect -757 -20 -723 14
rect -357 -20 -323 14
rect 1123 -20 1157 14
rect 1523 -20 1557 14
rect -2947 -260 -2913 -226
rect -2547 -260 -2513 -226
rect -757 -260 -723 -226
rect -357 -260 -323 -226
rect 1123 -260 1157 -226
rect 1523 -260 1557 -226
rect -3777 -890 -3743 -856
rect -3577 -1090 -3543 -1056
rect -2797 -695 -2763 -661
rect -2697 -820 -2663 -786
rect -3327 -990 -3293 -956
rect -3457 -1190 -3423 -1156
rect -2167 -890 -2133 -856
rect -1137 -700 -1103 -666
rect -607 -695 -573 -661
rect -507 -820 -473 -786
rect -1717 -990 -1683 -956
rect -1867 -1090 -1833 -1056
rect -2067 -1190 -2033 -1156
rect 593 -770 627 -736
rect 743 -870 777 -836
rect 1273 -695 1307 -661
rect 1373 -820 1407 -786
rect 23 -940 57 -906
rect 1853 -970 1887 -936
rect 2003 -1090 2037 -1056
rect -1916 -1900 -1882 -1866
rect -2066 -2020 -2032 -1986
rect -2196 -2140 -2162 -2106
rect -3496 -2310 -3462 -2276
rect -3326 -2290 -3292 -2256
rect -3626 -2390 -3592 -2356
rect -2696 -2280 -2662 -2246
rect -2796 -2405 -2762 -2371
rect 514 -1906 548 -1872
rect -116 -2160 -82 -2126
rect -1276 -2400 -1242 -2366
rect -646 -2280 -612 -2246
rect -746 -2405 -712 -2371
rect 614 -2031 648 -1997
rect 814 -2121 848 -2087
rect 1294 -2281 1328 -2247
rect 2214 -2231 2248 -2197
rect 2074 -2331 2108 -2297
rect 1394 -2406 1428 -2372
rect 1924 -2411 1958 -2377
rect -2946 -2840 -2912 -2806
rect -2546 -2840 -2512 -2806
rect -896 -2840 -862 -2806
rect -496 -2840 -462 -2806
rect 1144 -2841 1178 -2807
rect 1544 -2841 1578 -2807
<< locali >>
rect -3870 1074 -1590 1097
rect -3870 1040 -3787 1074
rect -3753 1040 -3707 1074
rect -3673 1040 -3627 1074
rect -3593 1040 -3547 1074
rect -3513 1040 -3467 1074
rect -3433 1040 -3387 1074
rect -3353 1040 -3307 1074
rect -3273 1040 -3227 1074
rect -3193 1040 -3147 1074
rect -3113 1040 -3067 1074
rect -3033 1040 -2987 1074
rect -2953 1040 -2907 1074
rect -2873 1040 -2827 1074
rect -2793 1040 -2747 1074
rect -2713 1040 -2667 1074
rect -2633 1040 -2587 1074
rect -2553 1040 -2507 1074
rect -2473 1040 -2427 1074
rect -2393 1040 -2347 1074
rect -2313 1040 -2267 1074
rect -2233 1040 -2187 1074
rect -2153 1040 -2107 1074
rect -2073 1040 -2027 1074
rect -1993 1040 -1947 1074
rect -1913 1040 -1867 1074
rect -1833 1040 -1787 1074
rect -1753 1040 -1707 1074
rect -1673 1040 -1590 1074
rect -3870 1017 -1590 1040
rect -1230 1074 150 1097
rect -1230 1040 -1197 1074
rect -1163 1040 -1117 1074
rect -1083 1040 -1037 1074
rect -1003 1040 -957 1074
rect -923 1040 -877 1074
rect -843 1040 -797 1074
rect -763 1040 -717 1074
rect -683 1040 -637 1074
rect -603 1040 -557 1074
rect -523 1040 -477 1074
rect -443 1040 -397 1074
rect -363 1040 -317 1074
rect -283 1040 -237 1074
rect -203 1040 -157 1074
rect -123 1040 -77 1074
rect -43 1040 3 1074
rect 37 1040 83 1074
rect 117 1040 150 1074
rect -1230 1017 150 1040
rect 500 1074 2180 1097
rect 500 1040 523 1074
rect 557 1040 603 1074
rect 637 1040 683 1074
rect 717 1040 763 1074
rect 797 1040 843 1074
rect 877 1040 923 1074
rect 957 1040 1003 1074
rect 1037 1040 1083 1074
rect 1117 1040 1163 1074
rect 1197 1040 1243 1074
rect 1277 1040 1323 1074
rect 1357 1040 1403 1074
rect 1437 1040 1483 1074
rect 1517 1040 1563 1074
rect 1597 1040 1643 1074
rect 1677 1040 1723 1074
rect 1757 1040 1803 1074
rect 1837 1040 1883 1074
rect 1917 1040 1963 1074
rect 1997 1040 2043 1074
rect 2077 1040 2123 1074
rect 2157 1040 2180 1074
rect 500 1017 2180 1040
rect -4662 947 -4582 967
rect -3480 947 -3400 967
rect -3350 947 -3270 967
rect -4662 944 -3270 947
rect -4662 910 -4639 944
rect -4605 910 -3457 944
rect -3423 910 -3327 944
rect -3293 910 -3270 944
rect -4662 907 -3270 910
rect -4662 887 -4582 907
rect -3480 887 -3400 907
rect -3350 887 -3270 907
rect -2090 944 -2010 967
rect -2090 910 -2067 944
rect -2033 910 -2010 944
rect -2090 887 -2010 910
rect -4548 847 -4468 867
rect -3600 847 -3520 867
rect -3220 847 -3140 867
rect -4548 844 -3140 847
rect -4548 810 -4525 844
rect -4491 810 -3577 844
rect -3543 810 -3197 844
rect -3163 810 -3140 844
rect -4548 807 -3140 810
rect -4548 787 -4468 807
rect -3600 787 -3520 807
rect -3220 787 -3140 807
rect -3070 854 -2990 887
rect -3070 820 -3047 854
rect -3013 820 -2990 854
rect -3070 774 -2990 820
rect -4890 747 -4810 767
rect -3350 747 -3270 767
rect -4890 744 -3270 747
rect -4890 710 -4867 744
rect -4833 710 -3327 744
rect -3293 710 -3270 744
rect -4890 707 -3270 710
rect -4890 687 -4810 707
rect -3350 687 -3270 707
rect -3070 740 -3047 774
rect -3013 740 -2990 774
rect -3070 694 -2990 740
rect -4776 647 -4696 667
rect -3800 647 -3720 667
rect -3220 647 -3140 667
rect -4776 644 -3140 647
rect -4776 610 -4753 644
rect -4719 610 -3777 644
rect -3743 610 -3197 644
rect -3163 610 -3140 644
rect -3070 660 -3047 694
rect -3013 660 -2990 694
rect -3070 637 -2990 660
rect -2920 854 -2840 887
rect -2920 820 -2897 854
rect -2863 820 -2840 854
rect -2920 774 -2840 820
rect -2920 740 -2897 774
rect -2863 740 -2840 774
rect -2920 694 -2840 740
rect -2920 660 -2897 694
rect -2863 660 -2840 694
rect -2920 627 -2840 660
rect -2770 854 -2690 887
rect -2770 820 -2747 854
rect -2713 820 -2690 854
rect -2770 774 -2690 820
rect -2770 740 -2747 774
rect -2713 740 -2690 774
rect -2770 694 -2690 740
rect -2770 660 -2747 694
rect -2713 660 -2690 694
rect -2770 637 -2690 660
rect -2620 854 -2540 887
rect -2620 820 -2597 854
rect -2563 820 -2540 854
rect -2620 774 -2540 820
rect -2620 740 -2597 774
rect -2563 740 -2540 774
rect -2620 694 -2540 740
rect -2620 660 -2597 694
rect -2563 660 -2540 694
rect -2620 627 -2540 660
rect -2470 854 -2390 887
rect -1318 879 -1238 901
rect -1591 878 -1238 879
rect -2470 820 -2447 854
rect -2413 820 -2390 854
rect -2470 774 -2390 820
rect -1890 844 -1810 867
rect -1890 810 -1867 844
rect -1833 810 -1810 844
rect -1890 787 -1810 810
rect -1591 844 -1295 878
rect -1261 844 -1238 878
rect -1591 839 -1238 844
rect -2470 740 -2447 774
rect -2413 740 -2390 774
rect -2470 694 -2390 740
rect -2470 660 -2447 694
rect -2413 660 -2390 694
rect -1740 744 -1660 767
rect -1740 710 -1717 744
rect -1683 710 -1660 744
rect -1740 687 -1660 710
rect -2470 637 -2390 660
rect -2190 644 -2110 667
rect -4776 607 -3140 610
rect -4776 587 -4696 607
rect -3800 587 -3720 607
rect -3220 587 -3140 607
rect -2900 577 -2860 627
rect -2720 577 -2640 597
rect -2900 574 -2640 577
rect -2900 540 -2697 574
rect -2663 540 -2640 574
rect -2900 537 -2640 540
rect -2900 407 -2860 537
rect -2720 517 -2640 537
rect -3830 367 -2860 407
rect -2820 457 -2740 472
rect -2600 457 -2560 627
rect -2190 610 -2167 644
rect -2133 610 -2110 644
rect -2190 587 -2110 610
rect -2350 564 -2270 587
rect -2350 530 -2327 564
rect -2293 547 -2270 564
rect -1591 547 -1551 839
rect -1318 821 -1238 839
rect -880 854 -800 887
rect -880 820 -857 854
rect -823 820 -800 854
rect -880 774 -800 820
rect -880 740 -857 774
rect -823 740 -800 774
rect -1030 697 -950 717
rect -1230 694 -950 697
rect -1230 660 -1007 694
rect -973 660 -950 694
rect -1230 657 -950 660
rect -1030 637 -950 657
rect -880 694 -800 740
rect -880 660 -857 694
rect -823 660 -800 694
rect -880 637 -800 660
rect -730 854 -650 887
rect -730 820 -707 854
rect -673 820 -650 854
rect -730 774 -650 820
rect -730 740 -707 774
rect -673 740 -650 774
rect -730 694 -650 740
rect -730 660 -707 694
rect -673 660 -650 694
rect -730 627 -650 660
rect -580 854 -500 887
rect -580 820 -557 854
rect -523 820 -500 854
rect -580 774 -500 820
rect -580 740 -557 774
rect -523 740 -500 774
rect -580 694 -500 740
rect -580 660 -557 694
rect -523 660 -500 694
rect -580 637 -500 660
rect -430 854 -350 887
rect -430 820 -407 854
rect -373 820 -350 854
rect -430 774 -350 820
rect -430 740 -407 774
rect -373 740 -350 774
rect -430 694 -350 740
rect -430 660 -407 694
rect -373 660 -350 694
rect -430 627 -350 660
rect -280 854 -200 887
rect -280 820 -257 854
rect -223 820 -200 854
rect -280 774 -200 820
rect 420 847 500 867
rect 850 847 930 867
rect 420 844 930 847
rect 420 810 443 844
rect 477 810 873 844
rect 907 810 930 844
rect 420 807 930 810
rect 420 787 500 807
rect 850 787 930 807
rect 1000 854 1080 887
rect 1000 820 1023 854
rect 1057 820 1080 854
rect -280 740 -257 774
rect -223 740 -200 774
rect 1000 774 1080 820
rect -280 694 -200 740
rect 272 727 661 732
rect 850 727 930 747
rect 272 724 930 727
rect -280 660 -257 694
rect -223 660 -200 694
rect -280 637 -200 660
rect -130 697 -50 717
rect 0 697 80 717
rect -130 694 80 697
rect -130 660 -107 694
rect -73 660 23 694
rect 57 660 80 694
rect -130 657 80 660
rect -130 637 -50 657
rect 0 637 80 657
rect 272 692 873 724
rect -2293 530 -1551 547
rect -2350 507 -1551 530
rect -710 577 -670 627
rect -530 577 -450 597
rect -710 574 -450 577
rect -710 540 -507 574
rect -473 540 -450 574
rect -710 537 -450 540
rect -1590 457 -1510 473
rect -1160 457 -1080 477
rect -2820 450 -1510 457
rect -2820 449 -1567 450
rect -2820 415 -2797 449
rect -2763 417 -1567 449
rect -2763 415 -2740 417
rect -2820 392 -2740 415
rect -3830 327 -3790 367
rect -3230 327 -3190 367
rect -2900 327 -2860 367
rect -2600 327 -2560 417
rect -2270 327 -2230 417
rect -1670 327 -1630 417
rect -1590 416 -1567 417
rect -1533 416 -1510 450
rect -1590 393 -1510 416
rect -1284 454 -1080 457
rect -1284 420 -1137 454
rect -1103 420 -1080 454
rect -1284 417 -1080 420
rect -3850 294 -3770 327
rect -3850 260 -3827 294
rect -3793 260 -3770 294
rect -3850 214 -3770 260
rect -3850 180 -3827 214
rect -3793 180 -3770 214
rect -3850 134 -3770 180
rect -3850 100 -3827 134
rect -3793 100 -3770 134
rect -3850 77 -3770 100
rect -3550 294 -3470 327
rect -3550 260 -3527 294
rect -3493 260 -3470 294
rect -3550 214 -3470 260
rect -3550 180 -3527 214
rect -3493 180 -3470 214
rect -3550 134 -3470 180
rect -3550 100 -3527 134
rect -3493 100 -3470 134
rect -3550 77 -3470 100
rect -3250 294 -3170 327
rect -3250 260 -3227 294
rect -3193 260 -3170 294
rect -3250 214 -3170 260
rect -3250 180 -3227 214
rect -3193 180 -3170 214
rect -3250 134 -3170 180
rect -3250 100 -3227 134
rect -3193 100 -3170 134
rect -3250 77 -3170 100
rect -3070 294 -2990 327
rect -3070 260 -3047 294
rect -3013 260 -2990 294
rect -3070 214 -2990 260
rect -3070 180 -3047 214
rect -3013 180 -2990 214
rect -3070 134 -2990 180
rect -3070 100 -3047 134
rect -3013 100 -2990 134
rect -3070 77 -2990 100
rect -2920 294 -2840 327
rect -2920 260 -2897 294
rect -2863 260 -2840 294
rect -2920 214 -2840 260
rect -2920 180 -2897 214
rect -2863 180 -2840 214
rect -2920 134 -2840 180
rect -2920 100 -2897 134
rect -2863 100 -2840 134
rect -2920 77 -2840 100
rect -2770 294 -2690 327
rect -2770 260 -2747 294
rect -2713 260 -2690 294
rect -2770 214 -2690 260
rect -2770 180 -2747 214
rect -2713 180 -2690 214
rect -2770 134 -2690 180
rect -2770 100 -2747 134
rect -2713 100 -2690 134
rect -2770 77 -2690 100
rect -2620 294 -2540 327
rect -2620 260 -2597 294
rect -2563 260 -2540 294
rect -2620 214 -2540 260
rect -2620 180 -2597 214
rect -2563 180 -2540 214
rect -2620 134 -2540 180
rect -2620 100 -2597 134
rect -2563 100 -2540 134
rect -2620 77 -2540 100
rect -2470 294 -2390 327
rect -2470 260 -2447 294
rect -2413 260 -2390 294
rect -2470 214 -2390 260
rect -2470 180 -2447 214
rect -2413 180 -2390 214
rect -2470 134 -2390 180
rect -2470 100 -2447 134
rect -2413 100 -2390 134
rect -2470 77 -2390 100
rect -2290 294 -2210 327
rect -2290 260 -2267 294
rect -2233 260 -2210 294
rect -2290 214 -2210 260
rect -2290 180 -2267 214
rect -2233 180 -2210 214
rect -2290 134 -2210 180
rect -2290 100 -2267 134
rect -2233 100 -2210 134
rect -2290 77 -2210 100
rect -1990 294 -1910 327
rect -1990 260 -1967 294
rect -1933 260 -1910 294
rect -1990 214 -1910 260
rect -1990 180 -1967 214
rect -1933 180 -1910 214
rect -1990 134 -1910 180
rect -1990 100 -1967 134
rect -1933 100 -1910 134
rect -1990 77 -1910 100
rect -1690 294 -1610 327
rect -1690 260 -1667 294
rect -1633 260 -1610 294
rect -1690 214 -1610 260
rect -1690 180 -1667 214
rect -1633 180 -1610 214
rect -1576 249 -1496 268
rect -1284 249 -1244 417
rect -1160 397 -1080 417
rect -710 407 -670 537
rect -530 517 -450 537
rect -1040 367 -670 407
rect -630 457 -550 472
rect -410 457 -370 627
rect -130 577 -50 597
rect 158 577 238 591
rect -130 574 238 577
rect -130 540 -107 574
rect -73 568 238 574
rect -73 540 181 568
rect -130 537 181 540
rect -130 517 -50 537
rect 158 534 181 537
rect 215 534 238 568
rect 158 511 238 534
rect -630 449 -370 457
rect -630 415 -607 449
rect -573 417 -370 449
rect -573 415 -550 417
rect -630 392 -550 415
rect -410 407 -370 417
rect 272 407 312 692
rect 500 690 873 692
rect 907 690 930 724
rect 500 687 930 690
rect 850 667 930 687
rect 1000 740 1023 774
rect 1057 740 1080 774
rect 1000 694 1080 740
rect 1000 660 1023 694
rect 1057 660 1080 694
rect 420 627 500 647
rect 720 627 800 647
rect 1000 637 1080 660
rect 1150 854 1230 887
rect 1150 820 1173 854
rect 1207 820 1230 854
rect 1150 774 1230 820
rect 1150 740 1173 774
rect 1207 740 1230 774
rect 1150 694 1230 740
rect 1150 660 1173 694
rect 1207 660 1230 694
rect 1150 627 1230 660
rect 1300 854 1380 887
rect 1300 820 1323 854
rect 1357 820 1380 854
rect 1300 774 1380 820
rect 1300 740 1323 774
rect 1357 740 1380 774
rect 1300 694 1380 740
rect 1300 660 1323 694
rect 1357 660 1380 694
rect 1300 637 1380 660
rect 1450 854 1530 887
rect 1450 820 1473 854
rect 1507 820 1530 854
rect 1450 774 1530 820
rect 1450 740 1473 774
rect 1507 740 1530 774
rect 1450 694 1530 740
rect 1450 660 1473 694
rect 1507 660 1530 694
rect 1450 627 1530 660
rect 1600 854 1680 887
rect 1600 820 1623 854
rect 1657 820 1680 854
rect 1600 774 1680 820
rect 1980 844 2060 867
rect 1980 810 2003 844
rect 2037 810 2060 844
rect 1980 787 2060 810
rect 1600 740 1623 774
rect 1657 740 1680 774
rect 1600 694 1680 740
rect 1600 660 1623 694
rect 1657 660 1680 694
rect 1830 724 1910 747
rect 1830 690 1853 724
rect 1887 690 1910 724
rect 1830 667 1910 690
rect 1600 637 1680 660
rect 420 624 800 627
rect 420 590 443 624
rect 477 590 743 624
rect 777 590 800 624
rect 420 587 800 590
rect 420 567 500 587
rect 720 567 800 587
rect 1170 577 1210 627
rect 1350 577 1430 597
rect 1170 574 1430 577
rect 570 527 650 547
rect 420 524 650 527
rect 420 504 593 524
rect 420 470 443 504
rect 477 490 593 504
rect 627 490 650 524
rect 477 487 650 490
rect 477 470 500 487
rect 420 447 500 470
rect 570 467 650 487
rect 1170 540 1373 574
rect 1407 540 1430 574
rect 1170 537 1430 540
rect 1170 407 1210 537
rect 1350 517 1430 537
rect -410 367 312 407
rect 540 367 1210 407
rect 1250 457 1330 472
rect 1470 457 1510 627
rect 1750 577 1830 597
rect 1750 574 2337 577
rect 1750 540 1773 574
rect 1807 540 2337 574
rect 1750 537 2337 540
rect 1750 517 1830 537
rect 2183 457 2263 477
rect 1250 454 2263 457
rect 1250 449 2206 454
rect 1250 415 1273 449
rect 1307 420 2206 449
rect 2240 420 2263 454
rect 1307 417 2263 420
rect 1307 415 1330 417
rect 1250 392 1330 415
rect -1040 327 -1000 367
rect -710 327 -670 367
rect -1576 246 -1244 249
rect -1576 212 -1553 246
rect -1519 212 -1244 246
rect -1576 209 -1244 212
rect -1210 294 -1130 327
rect -1210 260 -1187 294
rect -1153 260 -1130 294
rect -1210 214 -1130 260
rect -1576 188 -1496 209
rect -1690 134 -1610 180
rect -1690 100 -1667 134
rect -1633 100 -1610 134
rect -1690 77 -1610 100
rect -1210 180 -1187 214
rect -1153 180 -1130 214
rect -1210 134 -1130 180
rect -1210 100 -1187 134
rect -1153 100 -1130 134
rect -1210 77 -1130 100
rect -1060 294 -980 327
rect -1060 260 -1037 294
rect -1003 260 -980 294
rect -1060 214 -980 260
rect -1060 180 -1037 214
rect -1003 180 -980 214
rect -1060 134 -980 180
rect -1060 100 -1037 134
rect -1003 100 -980 134
rect -1060 77 -980 100
rect -880 294 -800 327
rect -880 260 -857 294
rect -823 260 -800 294
rect -880 214 -800 260
rect -880 180 -857 214
rect -823 180 -800 214
rect -880 134 -800 180
rect -880 100 -857 134
rect -823 100 -800 134
rect -880 77 -800 100
rect -730 294 -650 327
rect -730 260 -707 294
rect -673 260 -650 294
rect -730 214 -650 260
rect -730 180 -707 214
rect -673 180 -650 214
rect -730 134 -650 180
rect -730 100 -707 134
rect -673 100 -650 134
rect -730 77 -650 100
rect -580 294 -500 327
rect -580 260 -557 294
rect -523 260 -500 294
rect -580 214 -500 260
rect -580 180 -557 214
rect -523 180 -500 214
rect -580 134 -500 180
rect -580 100 -557 134
rect -523 100 -500 134
rect -580 77 -500 100
rect -430 294 -350 367
rect -80 327 -40 367
rect 540 327 580 367
rect 840 327 880 367
rect 1171 327 1210 367
rect 1470 327 1510 417
rect 1800 327 1840 417
rect 2183 397 2263 417
rect -430 260 -407 294
rect -373 260 -350 294
rect -430 214 -350 260
rect -430 180 -407 214
rect -373 180 -350 214
rect -430 134 -350 180
rect -430 100 -407 134
rect -373 100 -350 134
rect -430 77 -350 100
rect -280 294 -200 327
rect -280 260 -257 294
rect -223 260 -200 294
rect -280 214 -200 260
rect -280 180 -257 214
rect -223 180 -200 214
rect -280 134 -200 180
rect -280 100 -257 134
rect -223 100 -200 134
rect -280 77 -200 100
rect -100 294 -20 327
rect -100 260 -77 294
rect -43 260 -20 294
rect -100 214 -20 260
rect -100 180 -77 214
rect -43 180 -20 214
rect -100 134 -20 180
rect -100 100 -77 134
rect -43 100 -20 134
rect -100 77 -20 100
rect 50 294 130 327
rect 50 260 73 294
rect 107 260 130 294
rect 50 214 130 260
rect 50 180 73 214
rect 107 180 130 214
rect 50 134 130 180
rect 50 100 73 134
rect 107 100 130 134
rect 50 77 130 100
rect 520 294 600 327
rect 520 260 543 294
rect 577 260 600 294
rect 520 214 600 260
rect 520 180 543 214
rect 577 180 600 214
rect 520 134 600 180
rect 520 100 543 134
rect 577 100 600 134
rect 520 77 600 100
rect 670 294 750 327
rect 670 260 693 294
rect 727 260 750 294
rect 670 214 750 260
rect 670 180 693 214
rect 727 180 750 214
rect 670 134 750 180
rect 670 100 693 134
rect 727 100 750 134
rect 670 77 750 100
rect 820 294 900 327
rect 820 260 843 294
rect 877 260 900 294
rect 820 214 900 260
rect 820 180 843 214
rect 877 180 900 214
rect 820 134 900 180
rect 820 100 843 134
rect 877 100 900 134
rect 820 77 900 100
rect 1000 294 1080 327
rect 1000 260 1023 294
rect 1057 260 1080 294
rect 1000 214 1080 260
rect 1000 180 1023 214
rect 1057 180 1080 214
rect 1000 134 1080 180
rect 1000 100 1023 134
rect 1057 100 1080 134
rect 1000 77 1080 100
rect 1150 294 1230 327
rect 1150 260 1173 294
rect 1207 260 1230 294
rect 1150 214 1230 260
rect 1150 180 1173 214
rect 1207 180 1230 214
rect 1150 134 1230 180
rect 1150 100 1173 134
rect 1207 100 1230 134
rect 1150 77 1230 100
rect 1300 294 1380 327
rect 1300 260 1323 294
rect 1357 260 1380 294
rect 1300 214 1380 260
rect 1300 180 1323 214
rect 1357 180 1380 214
rect 1300 134 1380 180
rect 1300 100 1323 134
rect 1357 100 1380 134
rect 1300 77 1380 100
rect 1450 294 1530 327
rect 1450 260 1473 294
rect 1507 260 1530 294
rect 1450 214 1530 260
rect 1450 180 1473 214
rect 1507 180 1530 214
rect 1450 134 1530 180
rect 1450 100 1473 134
rect 1507 100 1530 134
rect 1450 77 1530 100
rect 1600 294 1680 327
rect 1600 260 1623 294
rect 1657 260 1680 294
rect 1600 214 1680 260
rect 1600 180 1623 214
rect 1657 180 1680 214
rect 1600 134 1680 180
rect 1600 100 1623 134
rect 1657 100 1680 134
rect 1600 77 1680 100
rect 1780 294 1860 327
rect 1780 260 1803 294
rect 1837 260 1860 294
rect 1780 214 1860 260
rect 1780 180 1803 214
rect 1837 180 1860 214
rect 1780 134 1860 180
rect 1780 100 1803 134
rect 1837 100 1860 134
rect 1780 77 1860 100
rect 2080 294 2160 327
rect 2080 260 2103 294
rect 2137 260 2160 294
rect 2080 214 2160 260
rect 2080 180 2103 214
rect 2137 180 2160 214
rect 2080 134 2160 180
rect 2080 100 2103 134
rect 2137 100 2160 134
rect 2080 77 2160 100
rect -3719 17 -3639 37
rect -2970 17 -2890 37
rect -2570 17 -2490 37
rect -780 17 -700 37
rect -380 17 -300 37
rect 508 17 588 37
rect 1100 17 1180 37
rect 1500 17 1580 37
rect -3870 14 -300 17
rect -3870 -20 -3696 14
rect -3662 -20 -2947 14
rect -2913 -20 -2547 14
rect -2513 -20 -757 14
rect -723 -20 -357 14
rect -323 -20 -300 14
rect -3870 -23 -300 -20
rect 500 14 1580 17
rect 500 -20 531 14
rect 565 -20 1123 14
rect 1157 -20 1523 14
rect 1557 -20 1580 14
rect 500 -23 1580 -20
rect -3719 -43 -3639 -23
rect -2970 -43 -2890 -23
rect -2570 -43 -2490 -23
rect -780 -43 -700 -23
rect -380 -43 -300 -23
rect 508 -43 588 -23
rect 1100 -43 1180 -23
rect 1500 -43 1580 -23
rect -3978 -106 -1590 -83
rect -3978 -140 -3955 -106
rect -3921 -140 -3787 -106
rect -3753 -140 -3707 -106
rect -3673 -140 -3627 -106
rect -3593 -140 -3547 -106
rect -3513 -140 -3467 -106
rect -3433 -140 -3387 -106
rect -3353 -140 -3307 -106
rect -3273 -140 -3227 -106
rect -3193 -140 -3147 -106
rect -3113 -140 -3067 -106
rect -3033 -140 -2987 -106
rect -2953 -140 -2907 -106
rect -2873 -140 -2827 -106
rect -2793 -140 -2747 -106
rect -2713 -140 -2667 -106
rect -2633 -140 -2587 -106
rect -2553 -140 -2507 -106
rect -2473 -140 -2427 -106
rect -2393 -140 -2347 -106
rect -2313 -140 -2267 -106
rect -2233 -140 -2187 -106
rect -2153 -140 -2107 -106
rect -2073 -140 -2027 -106
rect -1993 -140 -1947 -106
rect -1913 -140 -1867 -106
rect -1833 -140 -1787 -106
rect -1753 -140 -1707 -106
rect -1673 -140 -1590 -106
rect -3978 -163 -1590 -140
rect -1230 -106 150 -83
rect -1230 -140 -1197 -106
rect -1163 -140 -1117 -106
rect -1083 -140 -1037 -106
rect -1003 -140 -957 -106
rect -923 -140 -877 -106
rect -843 -140 -797 -106
rect -763 -140 -717 -106
rect -683 -140 -637 -106
rect -603 -140 -557 -106
rect -523 -140 -477 -106
rect -443 -140 -397 -106
rect -363 -140 -317 -106
rect -283 -140 -237 -106
rect -203 -140 -157 -106
rect -123 -140 -77 -106
rect -43 -140 3 -106
rect 37 -140 83 -106
rect 117 -140 150 -106
rect -1230 -163 150 -140
rect 500 -106 2180 -83
rect 500 -140 523 -106
rect 557 -140 603 -106
rect 637 -140 683 -106
rect 717 -140 763 -106
rect 797 -140 843 -106
rect 877 -140 923 -106
rect 957 -140 1003 -106
rect 1037 -140 1083 -106
rect 1117 -140 1163 -106
rect 1197 -140 1243 -106
rect 1277 -140 1323 -106
rect 1357 -140 1403 -106
rect 1437 -140 1483 -106
rect 1517 -140 1563 -106
rect 1597 -140 1643 -106
rect 1677 -140 1723 -106
rect 1757 -140 1803 -106
rect 1837 -140 1883 -106
rect 1917 -140 1963 -106
rect 1997 -140 2043 -106
rect 2077 -140 2123 -106
rect 2157 -140 2180 -106
rect 500 -163 2180 -140
rect -3719 -223 -3639 -203
rect -2970 -223 -2890 -203
rect -2570 -223 -2490 -203
rect -780 -223 -700 -203
rect -380 -223 -300 -203
rect 508 -223 588 -202
rect 1100 -223 1180 -203
rect 1500 -223 1580 -203
rect -3870 -226 -300 -223
rect -3870 -260 -3696 -226
rect -3662 -260 -2947 -226
rect -2913 -260 -2547 -226
rect -2513 -260 -757 -226
rect -723 -260 -357 -226
rect -323 -260 -300 -226
rect -3870 -263 -300 -260
rect 500 -225 1580 -223
rect 500 -259 531 -225
rect 565 -226 1580 -225
rect 565 -259 1123 -226
rect 500 -260 1123 -259
rect 1157 -260 1523 -226
rect 1557 -260 1580 -226
rect 500 -263 1580 -260
rect -3719 -283 -3639 -263
rect -2970 -283 -2890 -263
rect -2570 -283 -2490 -263
rect -780 -283 -700 -263
rect -380 -283 -300 -263
rect 508 -282 588 -263
rect 1100 -283 1180 -263
rect 1500 -283 1580 -263
rect -3850 -346 -3770 -323
rect -3850 -380 -3827 -346
rect -3793 -380 -3770 -346
rect -3850 -426 -3770 -380
rect -3850 -460 -3827 -426
rect -3793 -460 -3770 -426
rect -3850 -506 -3770 -460
rect -3850 -540 -3827 -506
rect -3793 -540 -3770 -506
rect -3850 -573 -3770 -540
rect -3550 -346 -3470 -323
rect -3550 -380 -3527 -346
rect -3493 -380 -3470 -346
rect -3550 -426 -3470 -380
rect -3550 -460 -3527 -426
rect -3493 -460 -3470 -426
rect -3550 -506 -3470 -460
rect -3550 -540 -3527 -506
rect -3493 -540 -3470 -506
rect -3550 -573 -3470 -540
rect -3250 -346 -3170 -323
rect -3250 -380 -3227 -346
rect -3193 -380 -3170 -346
rect -3250 -426 -3170 -380
rect -3250 -460 -3227 -426
rect -3193 -460 -3170 -426
rect -3250 -506 -3170 -460
rect -3250 -540 -3227 -506
rect -3193 -540 -3170 -506
rect -3250 -573 -3170 -540
rect -3070 -346 -2990 -323
rect -3070 -380 -3047 -346
rect -3013 -380 -2990 -346
rect -3070 -426 -2990 -380
rect -3070 -460 -3047 -426
rect -3013 -460 -2990 -426
rect -3070 -506 -2990 -460
rect -3070 -540 -3047 -506
rect -3013 -540 -2990 -506
rect -3070 -573 -2990 -540
rect -2920 -346 -2840 -323
rect -2920 -380 -2897 -346
rect -2863 -380 -2840 -346
rect -2920 -426 -2840 -380
rect -2920 -460 -2897 -426
rect -2863 -460 -2840 -426
rect -2920 -506 -2840 -460
rect -2920 -540 -2897 -506
rect -2863 -540 -2840 -506
rect -2920 -573 -2840 -540
rect -2770 -346 -2690 -323
rect -2770 -380 -2747 -346
rect -2713 -380 -2690 -346
rect -2770 -426 -2690 -380
rect -2770 -460 -2747 -426
rect -2713 -460 -2690 -426
rect -2770 -506 -2690 -460
rect -2770 -540 -2747 -506
rect -2713 -540 -2690 -506
rect -2770 -573 -2690 -540
rect -2620 -346 -2540 -323
rect -2620 -380 -2597 -346
rect -2563 -380 -2540 -346
rect -2620 -426 -2540 -380
rect -2620 -460 -2597 -426
rect -2563 -460 -2540 -426
rect -2620 -506 -2540 -460
rect -2620 -540 -2597 -506
rect -2563 -540 -2540 -506
rect -2620 -573 -2540 -540
rect -2470 -346 -2390 -323
rect -2470 -380 -2447 -346
rect -2413 -380 -2390 -346
rect -2470 -426 -2390 -380
rect -2470 -460 -2447 -426
rect -2413 -460 -2390 -426
rect -2470 -506 -2390 -460
rect -2470 -540 -2447 -506
rect -2413 -540 -2390 -506
rect -2470 -573 -2390 -540
rect -2290 -346 -2210 -323
rect -2290 -380 -2267 -346
rect -2233 -380 -2210 -346
rect -2290 -426 -2210 -380
rect -2290 -460 -2267 -426
rect -2233 -460 -2210 -426
rect -2290 -506 -2210 -460
rect -2290 -540 -2267 -506
rect -2233 -540 -2210 -506
rect -2290 -573 -2210 -540
rect -1990 -346 -1910 -323
rect -1990 -380 -1967 -346
rect -1933 -380 -1910 -346
rect -1990 -426 -1910 -380
rect -1990 -460 -1967 -426
rect -1933 -460 -1910 -426
rect -1990 -506 -1910 -460
rect -1990 -540 -1967 -506
rect -1933 -540 -1910 -506
rect -1990 -573 -1910 -540
rect -1690 -346 -1610 -323
rect -1690 -380 -1667 -346
rect -1633 -380 -1610 -346
rect -1690 -426 -1610 -380
rect -1690 -460 -1667 -426
rect -1633 -460 -1610 -426
rect -1210 -346 -1130 -323
rect -1210 -380 -1187 -346
rect -1153 -380 -1130 -346
rect -1210 -426 -1130 -380
rect -1690 -506 -1610 -460
rect -1690 -540 -1667 -506
rect -1633 -540 -1610 -506
rect -1576 -446 -1496 -427
rect -1576 -449 -1244 -446
rect -1576 -483 -1553 -449
rect -1519 -483 -1244 -449
rect -1576 -486 -1244 -483
rect -1576 -507 -1496 -486
rect -1690 -573 -1610 -540
rect -3830 -613 -3790 -573
rect -3230 -613 -3190 -573
rect -2900 -613 -2860 -573
rect -3830 -653 -2860 -613
rect -2900 -783 -2860 -653
rect -2820 -661 -2740 -638
rect -2820 -695 -2797 -661
rect -2763 -663 -2740 -661
rect -2600 -663 -2560 -573
rect -2270 -663 -2230 -573
rect -1670 -663 -1630 -573
rect -1284 -663 -1244 -486
rect -1210 -460 -1187 -426
rect -1153 -460 -1130 -426
rect -1210 -506 -1130 -460
rect -1210 -540 -1187 -506
rect -1153 -540 -1130 -506
rect -1210 -573 -1130 -540
rect -1060 -346 -980 -323
rect -1060 -380 -1037 -346
rect -1003 -380 -980 -346
rect -1060 -426 -980 -380
rect -1060 -460 -1037 -426
rect -1003 -460 -980 -426
rect -1060 -506 -980 -460
rect -1060 -540 -1037 -506
rect -1003 -540 -980 -506
rect -1060 -573 -980 -540
rect -880 -346 -800 -323
rect -880 -380 -857 -346
rect -823 -380 -800 -346
rect -880 -426 -800 -380
rect -880 -460 -857 -426
rect -823 -460 -800 -426
rect -880 -506 -800 -460
rect -880 -540 -857 -506
rect -823 -540 -800 -506
rect -880 -573 -800 -540
rect -730 -346 -650 -323
rect -730 -380 -707 -346
rect -673 -380 -650 -346
rect -730 -426 -650 -380
rect -730 -460 -707 -426
rect -673 -460 -650 -426
rect -730 -506 -650 -460
rect -730 -540 -707 -506
rect -673 -540 -650 -506
rect -730 -573 -650 -540
rect -580 -346 -500 -323
rect -580 -380 -557 -346
rect -523 -380 -500 -346
rect -580 -426 -500 -380
rect -580 -460 -557 -426
rect -523 -460 -500 -426
rect -580 -506 -500 -460
rect -580 -540 -557 -506
rect -523 -540 -500 -506
rect -580 -573 -500 -540
rect -430 -346 -350 -323
rect -430 -380 -407 -346
rect -373 -380 -350 -346
rect -430 -426 -350 -380
rect -430 -460 -407 -426
rect -373 -460 -350 -426
rect -430 -506 -350 -460
rect -430 -540 -407 -506
rect -373 -540 -350 -506
rect -1040 -613 -1000 -573
rect -710 -613 -670 -573
rect -430 -613 -350 -540
rect -280 -346 -200 -323
rect -280 -380 -257 -346
rect -223 -380 -200 -346
rect -280 -426 -200 -380
rect -280 -460 -257 -426
rect -223 -460 -200 -426
rect -280 -506 -200 -460
rect -280 -540 -257 -506
rect -223 -540 -200 -506
rect -280 -573 -200 -540
rect -100 -346 -20 -323
rect -100 -380 -77 -346
rect -43 -380 -20 -346
rect -100 -426 -20 -380
rect -100 -460 -77 -426
rect -43 -460 -20 -426
rect -100 -506 -20 -460
rect -100 -540 -77 -506
rect -43 -540 -20 -506
rect -100 -573 -20 -540
rect 50 -346 130 -323
rect 50 -380 73 -346
rect 107 -380 130 -346
rect 50 -426 130 -380
rect 50 -460 73 -426
rect 107 -460 130 -426
rect 50 -506 130 -460
rect 50 -540 73 -506
rect 107 -540 130 -506
rect 50 -573 130 -540
rect 520 -346 600 -323
rect 520 -380 543 -346
rect 577 -380 600 -346
rect 520 -426 600 -380
rect 520 -460 543 -426
rect 577 -460 600 -426
rect 520 -506 600 -460
rect 520 -540 543 -506
rect 577 -540 600 -506
rect 520 -573 600 -540
rect 670 -346 750 -323
rect 670 -380 693 -346
rect 727 -380 750 -346
rect 670 -426 750 -380
rect 670 -460 693 -426
rect 727 -460 750 -426
rect 670 -506 750 -460
rect 670 -540 693 -506
rect 727 -540 750 -506
rect 670 -573 750 -540
rect 820 -346 900 -323
rect 820 -380 843 -346
rect 877 -380 900 -346
rect 820 -426 900 -380
rect 820 -460 843 -426
rect 877 -460 900 -426
rect 820 -506 900 -460
rect 820 -540 843 -506
rect 877 -540 900 -506
rect 820 -573 900 -540
rect 1000 -346 1080 -323
rect 1000 -380 1023 -346
rect 1057 -380 1080 -346
rect 1000 -426 1080 -380
rect 1000 -460 1023 -426
rect 1057 -460 1080 -426
rect 1000 -506 1080 -460
rect 1000 -540 1023 -506
rect 1057 -540 1080 -506
rect 1000 -573 1080 -540
rect 1150 -346 1230 -323
rect 1150 -380 1173 -346
rect 1207 -380 1230 -346
rect 1150 -426 1230 -380
rect 1150 -460 1173 -426
rect 1207 -460 1230 -426
rect 1150 -506 1230 -460
rect 1150 -540 1173 -506
rect 1207 -540 1230 -506
rect 1150 -573 1230 -540
rect 1300 -346 1380 -323
rect 1300 -380 1323 -346
rect 1357 -380 1380 -346
rect 1300 -426 1380 -380
rect 1300 -460 1323 -426
rect 1357 -460 1380 -426
rect 1300 -506 1380 -460
rect 1300 -540 1323 -506
rect 1357 -540 1380 -506
rect 1300 -573 1380 -540
rect 1450 -346 1530 -323
rect 1450 -380 1473 -346
rect 1507 -380 1530 -346
rect 1450 -426 1530 -380
rect 1450 -460 1473 -426
rect 1507 -460 1530 -426
rect 1450 -506 1530 -460
rect 1450 -540 1473 -506
rect 1507 -540 1530 -506
rect 1450 -573 1530 -540
rect 1600 -346 1680 -323
rect 1600 -380 1623 -346
rect 1657 -380 1680 -346
rect 1600 -426 1680 -380
rect 1600 -460 1623 -426
rect 1657 -460 1680 -426
rect 1600 -506 1680 -460
rect 1600 -540 1623 -506
rect 1657 -540 1680 -506
rect 1600 -573 1680 -540
rect 1780 -346 1860 -323
rect 1780 -380 1803 -346
rect 1837 -380 1860 -346
rect 1780 -426 1860 -380
rect 1780 -460 1803 -426
rect 1837 -460 1860 -426
rect 1780 -506 1860 -460
rect 1780 -540 1803 -506
rect 1837 -540 1860 -506
rect 1780 -573 1860 -540
rect 2080 -346 2160 -323
rect 2080 -380 2103 -346
rect 2137 -380 2160 -346
rect 2080 -426 2160 -380
rect 2080 -460 2103 -426
rect 2137 -460 2160 -426
rect 2080 -506 2160 -460
rect 2080 -540 2103 -506
rect 2137 -540 2160 -506
rect 2080 -573 2160 -540
rect -80 -613 -40 -573
rect 158 -613 238 -593
rect -1160 -663 -1080 -643
rect -1040 -653 -670 -613
rect -410 -616 238 -613
rect -2763 -695 -1385 -663
rect -2820 -703 -1385 -695
rect -1284 -666 -1080 -663
rect -1284 -700 -1137 -666
rect -1103 -700 -1080 -666
rect -1284 -703 -1080 -700
rect -2820 -718 -2740 -703
rect -2720 -783 -2640 -763
rect -2900 -786 -2640 -783
rect -2900 -820 -2697 -786
rect -2663 -820 -2640 -786
rect -2900 -823 -2640 -820
rect -4092 -853 -4012 -833
rect -3800 -853 -3720 -833
rect -3220 -853 -3140 -833
rect -4092 -856 -3140 -853
rect -4092 -890 -4069 -856
rect -4035 -890 -3777 -856
rect -3743 -890 -3197 -856
rect -3163 -890 -3140 -856
rect -2900 -873 -2860 -823
rect -2720 -843 -2640 -823
rect -2600 -873 -2560 -703
rect -2350 -776 -1510 -753
rect -2350 -810 -2327 -776
rect -2293 -793 -1567 -776
rect -2293 -810 -2270 -793
rect -2350 -833 -2270 -810
rect -1590 -810 -1567 -793
rect -1533 -810 -1510 -776
rect -1590 -833 -1510 -810
rect -2190 -856 -2110 -833
rect -4092 -893 -3140 -890
rect -4092 -913 -4012 -893
rect -3800 -913 -3720 -893
rect -3220 -913 -3140 -893
rect -3070 -906 -2990 -883
rect -4206 -953 -4126 -933
rect -3350 -953 -3270 -933
rect -4206 -956 -3270 -953
rect -4206 -990 -4183 -956
rect -4149 -990 -3327 -956
rect -3293 -990 -3270 -956
rect -4206 -993 -3270 -990
rect -4206 -1013 -4126 -993
rect -3350 -1013 -3270 -993
rect -3070 -940 -3047 -906
rect -3013 -940 -2990 -906
rect -3070 -986 -2990 -940
rect -3070 -1020 -3047 -986
rect -3013 -1020 -2990 -986
rect -4320 -1053 -4240 -1033
rect -3600 -1053 -3520 -1033
rect -3220 -1053 -3140 -1033
rect -4320 -1056 -3140 -1053
rect -4320 -1090 -4297 -1056
rect -4263 -1090 -3577 -1056
rect -3543 -1090 -3197 -1056
rect -3163 -1090 -3140 -1056
rect -4320 -1093 -3140 -1090
rect -4320 -1113 -4240 -1093
rect -3600 -1113 -3520 -1093
rect -3220 -1113 -3140 -1093
rect -3070 -1066 -2990 -1020
rect -3070 -1100 -3047 -1066
rect -3013 -1100 -2990 -1066
rect -3070 -1133 -2990 -1100
rect -2920 -906 -2840 -873
rect -2920 -940 -2897 -906
rect -2863 -940 -2840 -906
rect -2920 -986 -2840 -940
rect -2920 -1020 -2897 -986
rect -2863 -1020 -2840 -986
rect -2920 -1066 -2840 -1020
rect -2920 -1100 -2897 -1066
rect -2863 -1100 -2840 -1066
rect -2920 -1133 -2840 -1100
rect -2770 -906 -2690 -883
rect -2770 -940 -2747 -906
rect -2713 -940 -2690 -906
rect -2770 -986 -2690 -940
rect -2770 -1020 -2747 -986
rect -2713 -1020 -2690 -986
rect -2770 -1066 -2690 -1020
rect -2770 -1100 -2747 -1066
rect -2713 -1100 -2690 -1066
rect -2770 -1133 -2690 -1100
rect -2620 -906 -2540 -873
rect -2620 -940 -2597 -906
rect -2563 -940 -2540 -906
rect -2620 -986 -2540 -940
rect -2620 -1020 -2597 -986
rect -2563 -1020 -2540 -986
rect -2620 -1066 -2540 -1020
rect -2620 -1100 -2597 -1066
rect -2563 -1100 -2540 -1066
rect -2620 -1133 -2540 -1100
rect -2470 -906 -2390 -883
rect -2470 -940 -2447 -906
rect -2413 -940 -2390 -906
rect -2190 -890 -2167 -856
rect -2133 -890 -2110 -856
rect -2190 -913 -2110 -890
rect -2470 -986 -2390 -940
rect -2470 -1020 -2447 -986
rect -2413 -1020 -2390 -986
rect -1740 -956 -1660 -933
rect -1740 -990 -1717 -956
rect -1683 -990 -1660 -956
rect -1740 -1013 -1660 -990
rect -2470 -1066 -2390 -1020
rect -2470 -1100 -2447 -1066
rect -2413 -1100 -2390 -1066
rect -2470 -1133 -2390 -1100
rect -1890 -1056 -1810 -1033
rect -1890 -1090 -1867 -1056
rect -1833 -1090 -1810 -1056
rect -1890 -1113 -1810 -1090
rect -1425 -1085 -1385 -703
rect -1160 -723 -1080 -703
rect -710 -783 -670 -653
rect -630 -661 -550 -638
rect -630 -695 -607 -661
rect -573 -663 -550 -661
rect -410 -650 181 -616
rect 215 -650 238 -616
rect -410 -653 238 -650
rect 540 -613 580 -573
rect 840 -613 880 -573
rect 1171 -613 1210 -573
rect 540 -653 1210 -613
rect -410 -663 -370 -653
rect -573 -695 -370 -663
rect 158 -673 238 -653
rect -630 -703 -370 -695
rect -630 -718 -550 -703
rect -530 -783 -450 -763
rect -710 -786 -450 -783
rect -710 -820 -507 -786
rect -473 -820 -450 -786
rect -710 -823 -450 -820
rect -710 -873 -670 -823
rect -530 -843 -450 -823
rect -410 -873 -370 -703
rect 570 -733 650 -713
rect 130 -736 650 -733
rect -130 -783 -50 -763
rect 130 -770 593 -736
rect 627 -770 650 -736
rect 130 -773 650 -770
rect 130 -783 170 -773
rect -130 -786 170 -783
rect -130 -820 -107 -786
rect -73 -820 170 -786
rect 570 -793 650 -773
rect 1170 -783 1210 -653
rect 1250 -661 1330 -638
rect 1250 -695 1273 -661
rect 1307 -663 1330 -661
rect 1470 -663 1510 -573
rect 1800 -663 1840 -573
rect 2183 -663 2263 -643
rect 1307 -666 2263 -663
rect 1307 -695 2206 -666
rect 1250 -700 2206 -695
rect 2240 -700 2263 -666
rect 1250 -703 2263 -700
rect 1250 -718 1330 -703
rect 1350 -783 1430 -763
rect 1170 -786 1430 -783
rect -130 -823 170 -820
rect -130 -843 -50 -823
rect 720 -833 800 -813
rect 272 -836 800 -833
rect 272 -870 743 -836
rect 777 -870 800 -836
rect 272 -873 800 -870
rect 1170 -820 1373 -786
rect 1407 -820 1430 -786
rect 1170 -823 1430 -820
rect 1170 -873 1210 -823
rect 1350 -843 1430 -823
rect 1470 -873 1510 -703
rect 2183 -723 2263 -703
rect 1750 -783 1830 -763
rect 1750 -786 2254 -783
rect 1750 -820 1773 -786
rect 1807 -820 2254 -786
rect 1750 -823 2254 -820
rect 1750 -843 1830 -823
rect -1030 -903 -950 -883
rect -1230 -906 -950 -903
rect -1230 -940 -1007 -906
rect -973 -940 -950 -906
rect -1230 -943 -950 -940
rect -1030 -963 -950 -943
rect -880 -906 -800 -883
rect -880 -940 -857 -906
rect -823 -940 -800 -906
rect -880 -986 -800 -940
rect -880 -1020 -857 -986
rect -823 -1020 -800 -986
rect -880 -1066 -800 -1020
rect -1318 -1085 -1238 -1067
rect -1425 -1090 -1238 -1085
rect -1425 -1124 -1295 -1090
rect -1261 -1124 -1238 -1090
rect -1425 -1125 -1238 -1124
rect -4434 -1153 -4354 -1133
rect -3480 -1153 -3400 -1133
rect -3350 -1153 -3270 -1133
rect -4434 -1156 -3270 -1153
rect -4434 -1190 -4411 -1156
rect -4377 -1190 -3457 -1156
rect -3423 -1190 -3327 -1156
rect -3293 -1190 -3270 -1156
rect -4434 -1193 -3270 -1190
rect -4434 -1213 -4354 -1193
rect -3480 -1213 -3400 -1193
rect -3350 -1213 -3270 -1193
rect -2090 -1156 -2010 -1133
rect -1318 -1147 -1238 -1125
rect -880 -1100 -857 -1066
rect -823 -1100 -800 -1066
rect -880 -1133 -800 -1100
rect -730 -906 -650 -873
rect -730 -940 -707 -906
rect -673 -940 -650 -906
rect -730 -986 -650 -940
rect -730 -1020 -707 -986
rect -673 -1020 -650 -986
rect -730 -1066 -650 -1020
rect -730 -1100 -707 -1066
rect -673 -1100 -650 -1066
rect -730 -1133 -650 -1100
rect -580 -906 -500 -883
rect -580 -940 -557 -906
rect -523 -940 -500 -906
rect -580 -986 -500 -940
rect -580 -1020 -557 -986
rect -523 -1020 -500 -986
rect -580 -1066 -500 -1020
rect -580 -1100 -557 -1066
rect -523 -1100 -500 -1066
rect -580 -1133 -500 -1100
rect -430 -906 -350 -873
rect -430 -940 -407 -906
rect -373 -940 -350 -906
rect -430 -986 -350 -940
rect -430 -1020 -407 -986
rect -373 -1020 -350 -986
rect -430 -1066 -350 -1020
rect -430 -1100 -407 -1066
rect -373 -1100 -350 -1066
rect -430 -1133 -350 -1100
rect -280 -906 -200 -883
rect -280 -940 -257 -906
rect -223 -940 -200 -906
rect -280 -986 -200 -940
rect -130 -903 -50 -883
rect 0 -903 80 -883
rect -130 -906 80 -903
rect -130 -940 -107 -906
rect -73 -940 23 -906
rect 57 -940 80 -906
rect -130 -943 80 -940
rect -130 -963 -50 -943
rect 0 -963 80 -943
rect 158 -941 238 -921
rect 272 -941 312 -873
rect 720 -893 800 -873
rect 1000 -906 1080 -883
rect 158 -944 312 -941
rect -280 -1020 -257 -986
rect -223 -1020 -200 -986
rect 158 -978 181 -944
rect 215 -978 312 -944
rect 158 -981 312 -978
rect 420 -933 500 -913
rect 850 -933 930 -913
rect 420 -936 930 -933
rect 420 -970 443 -936
rect 477 -970 873 -936
rect 907 -970 930 -936
rect 420 -973 930 -970
rect 158 -1001 238 -981
rect 420 -993 500 -973
rect 850 -993 930 -973
rect 1000 -940 1023 -906
rect 1057 -940 1080 -906
rect 1000 -986 1080 -940
rect -280 -1066 -200 -1020
rect 1000 -1020 1023 -986
rect 1057 -1020 1080 -986
rect -280 -1100 -257 -1066
rect -223 -1100 -200 -1066
rect -280 -1133 -200 -1100
rect 420 -1053 500 -1034
rect 850 -1053 930 -1033
rect 420 -1056 930 -1053
rect 420 -1057 873 -1056
rect 420 -1091 443 -1057
rect 477 -1090 873 -1057
rect 907 -1090 930 -1056
rect 477 -1091 930 -1090
rect 420 -1093 930 -1091
rect 420 -1114 500 -1093
rect 850 -1113 930 -1093
rect 1000 -1066 1080 -1020
rect 1000 -1100 1023 -1066
rect 1057 -1100 1080 -1066
rect 1000 -1133 1080 -1100
rect 1150 -906 1230 -873
rect 1150 -940 1173 -906
rect 1207 -940 1230 -906
rect 1150 -986 1230 -940
rect 1150 -1020 1173 -986
rect 1207 -1020 1230 -986
rect 1150 -1066 1230 -1020
rect 1150 -1100 1173 -1066
rect 1207 -1100 1230 -1066
rect 1150 -1133 1230 -1100
rect 1300 -906 1380 -883
rect 1300 -940 1323 -906
rect 1357 -940 1380 -906
rect 1300 -986 1380 -940
rect 1300 -1020 1323 -986
rect 1357 -1020 1380 -986
rect 1300 -1066 1380 -1020
rect 1300 -1100 1323 -1066
rect 1357 -1100 1380 -1066
rect 1300 -1133 1380 -1100
rect 1450 -906 1530 -873
rect 1450 -940 1473 -906
rect 1507 -940 1530 -906
rect 1450 -986 1530 -940
rect 1450 -1020 1473 -986
rect 1507 -1020 1530 -986
rect 1450 -1066 1530 -1020
rect 1450 -1100 1473 -1066
rect 1507 -1100 1530 -1066
rect 1450 -1133 1530 -1100
rect 1600 -906 1680 -883
rect 1600 -940 1623 -906
rect 1657 -940 1680 -906
rect 1600 -986 1680 -940
rect 1600 -1020 1623 -986
rect 1657 -1020 1680 -986
rect 1830 -936 1910 -913
rect 1830 -970 1853 -936
rect 1887 -970 1910 -936
rect 1830 -993 1910 -970
rect 1600 -1066 1680 -1020
rect 1600 -1100 1623 -1066
rect 1657 -1100 1680 -1066
rect 1600 -1133 1680 -1100
rect 1980 -1056 2060 -1033
rect 1980 -1090 2003 -1056
rect 2037 -1090 2060 -1056
rect 1980 -1113 2060 -1090
rect -2090 -1190 -2067 -1156
rect -2033 -1190 -2010 -1156
rect -2090 -1213 -2010 -1190
rect -3870 -1286 -1590 -1263
rect -3870 -1320 -3787 -1286
rect -3753 -1320 -3707 -1286
rect -3673 -1320 -3627 -1286
rect -3593 -1320 -3547 -1286
rect -3513 -1320 -3467 -1286
rect -3433 -1320 -3387 -1286
rect -3353 -1320 -3307 -1286
rect -3273 -1320 -3227 -1286
rect -3193 -1320 -3147 -1286
rect -3113 -1320 -3067 -1286
rect -3033 -1320 -2987 -1286
rect -2953 -1320 -2907 -1286
rect -2873 -1320 -2827 -1286
rect -2793 -1320 -2747 -1286
rect -2713 -1320 -2667 -1286
rect -2633 -1320 -2587 -1286
rect -2553 -1320 -2507 -1286
rect -2473 -1320 -2427 -1286
rect -2393 -1320 -2347 -1286
rect -2313 -1320 -2267 -1286
rect -2233 -1320 -2187 -1286
rect -2153 -1320 -2107 -1286
rect -2073 -1320 -2027 -1286
rect -1993 -1320 -1947 -1286
rect -1913 -1320 -1867 -1286
rect -1833 -1320 -1787 -1286
rect -1753 -1320 -1707 -1286
rect -1673 -1320 -1590 -1286
rect -3870 -1343 -1590 -1320
rect -1230 -1286 150 -1263
rect -1230 -1320 -1197 -1286
rect -1163 -1320 -1117 -1286
rect -1083 -1320 -1037 -1286
rect -1003 -1320 -957 -1286
rect -923 -1320 -877 -1286
rect -843 -1320 -797 -1286
rect -763 -1320 -717 -1286
rect -683 -1320 -637 -1286
rect -603 -1320 -557 -1286
rect -523 -1320 -477 -1286
rect -443 -1320 -397 -1286
rect -363 -1320 -317 -1286
rect -283 -1320 -237 -1286
rect -203 -1320 -157 -1286
rect -123 -1320 -77 -1286
rect -43 -1320 3 -1286
rect 37 -1320 83 -1286
rect 117 -1320 150 -1286
rect -1230 -1343 150 -1320
rect 500 -1286 2180 -1263
rect 500 -1320 523 -1286
rect 557 -1320 603 -1286
rect 637 -1320 683 -1286
rect 717 -1320 763 -1286
rect 797 -1320 843 -1286
rect 877 -1320 923 -1286
rect 957 -1320 1003 -1286
rect 1037 -1320 1083 -1286
rect 1117 -1320 1163 -1286
rect 1197 -1320 1243 -1286
rect 1277 -1320 1323 -1286
rect 1357 -1320 1403 -1286
rect 1437 -1320 1483 -1286
rect 1517 -1320 1563 -1286
rect 1597 -1320 1643 -1286
rect 1677 -1320 1723 -1286
rect 1757 -1320 1803 -1286
rect 1837 -1320 1883 -1286
rect 1917 -1320 1963 -1286
rect 1997 -1320 2043 -1286
rect 2077 -1320 2123 -1286
rect 2157 -1320 2180 -1286
rect 500 -1343 2180 -1320
rect 508 -1517 588 -1497
rect 134 -1520 588 -1517
rect 134 -1554 531 -1520
rect 565 -1554 588 -1520
rect 134 -1557 588 -1554
rect -3729 -1746 -1729 -1723
rect -3729 -1780 -3706 -1746
rect -3672 -1780 -3626 -1746
rect -3592 -1780 -3546 -1746
rect -3512 -1780 -3466 -1746
rect -3432 -1780 -3386 -1746
rect -3352 -1780 -3306 -1746
rect -3272 -1780 -3226 -1746
rect -3192 -1780 -3146 -1746
rect -3112 -1780 -3066 -1746
rect -3032 -1780 -2986 -1746
rect -2952 -1780 -2906 -1746
rect -2872 -1780 -2826 -1746
rect -2792 -1780 -2746 -1746
rect -2712 -1780 -2666 -1746
rect -2632 -1780 -2586 -1746
rect -2552 -1780 -2506 -1746
rect -2472 -1780 -2426 -1746
rect -2392 -1780 -2346 -1746
rect -2312 -1780 -2266 -1746
rect -2232 -1780 -2186 -1746
rect -2152 -1780 -2106 -1746
rect -2072 -1780 -2026 -1746
rect -1992 -1780 -1946 -1746
rect -1912 -1780 -1866 -1746
rect -1832 -1780 -1786 -1746
rect -1752 -1780 -1729 -1746
rect -3729 -1803 -1729 -1780
rect -1369 -1746 11 -1723
rect -1369 -1780 -1336 -1746
rect -1302 -1780 -1256 -1746
rect -1222 -1780 -1176 -1746
rect -1142 -1780 -1096 -1746
rect -1062 -1780 -1016 -1746
rect -982 -1780 -936 -1746
rect -902 -1780 -856 -1746
rect -822 -1780 -776 -1746
rect -742 -1780 -696 -1746
rect -662 -1780 -616 -1746
rect -582 -1780 -536 -1746
rect -502 -1780 -456 -1746
rect -422 -1780 -376 -1746
rect -342 -1780 -296 -1746
rect -262 -1780 -216 -1746
rect -182 -1780 -136 -1746
rect -102 -1780 -56 -1746
rect -22 -1780 11 -1746
rect -1369 -1803 11 -1780
rect -4320 -1863 -4240 -1843
rect -3309 -1863 -3229 -1843
rect -4320 -1866 -3229 -1863
rect -4320 -1900 -4297 -1866
rect -4263 -1900 -3286 -1866
rect -3252 -1900 -3229 -1866
rect -4320 -1903 -3229 -1900
rect -4320 -1923 -4240 -1903
rect -3309 -1923 -3229 -1903
rect -1939 -1866 -1859 -1843
rect -1939 -1900 -1916 -1866
rect -1882 -1900 -1859 -1866
rect -1939 -1923 -1859 -1900
rect 134 -1930 174 -1557
rect 508 -1577 588 -1557
rect 2214 -1644 2254 -823
rect 2297 -1551 2337 537
rect 2453 -1551 2533 -1530
rect 2297 -1553 2533 -1551
rect 2297 -1587 2476 -1553
rect 2510 -1587 2533 -1553
rect 2297 -1591 2533 -1587
rect 2453 -1610 2533 -1591
rect 2214 -1684 2539 -1644
rect 361 -1747 2361 -1724
rect 361 -1781 384 -1747
rect 418 -1781 464 -1747
rect 498 -1781 544 -1747
rect 578 -1781 624 -1747
rect 658 -1781 704 -1747
rect 738 -1781 784 -1747
rect 818 -1781 864 -1747
rect 898 -1781 944 -1747
rect 978 -1781 1024 -1747
rect 1058 -1781 1104 -1747
rect 1138 -1781 1184 -1747
rect 1218 -1781 1264 -1747
rect 1298 -1781 1344 -1747
rect 1378 -1781 1424 -1747
rect 1458 -1781 1504 -1747
rect 1538 -1781 1584 -1747
rect 1618 -1781 1664 -1747
rect 1698 -1781 1744 -1747
rect 1778 -1781 1824 -1747
rect 1858 -1781 1904 -1747
rect 1938 -1781 1984 -1747
rect 2018 -1781 2064 -1747
rect 2098 -1781 2144 -1747
rect 2178 -1781 2224 -1747
rect 2258 -1781 2304 -1747
rect 2338 -1781 2361 -1747
rect 361 -1804 2361 -1781
rect 491 -1872 571 -1849
rect 491 -1906 514 -1872
rect 548 -1906 571 -1872
rect 491 -1929 571 -1906
rect 1771 -1874 1851 -1854
rect 2339 -1874 2419 -1854
rect 1771 -1877 2419 -1874
rect 1771 -1911 1794 -1877
rect 1828 -1911 2362 -1877
rect 2396 -1911 2419 -1877
rect 1771 -1914 2419 -1911
rect -4890 -1983 -4810 -1963
rect -3219 -1983 -3139 -1963
rect -4890 -1986 -3139 -1983
rect -4890 -2020 -4867 -1986
rect -4833 -2020 -3196 -1986
rect -3162 -2020 -3139 -1986
rect -4890 -2023 -3139 -2020
rect -4890 -2043 -4810 -2023
rect -3219 -2043 -3139 -2023
rect -3069 -1966 -2989 -1933
rect -3069 -2000 -3046 -1966
rect -3012 -2000 -2989 -1966
rect -3069 -2046 -2989 -2000
rect -4206 -2082 -4126 -2059
rect -4206 -2116 -4183 -2082
rect -4149 -2093 -4126 -2082
rect -3069 -2080 -3046 -2046
rect -3012 -2080 -2989 -2046
rect -3249 -2093 -3169 -2083
rect -4149 -2106 -3169 -2093
rect -4149 -2116 -3226 -2106
rect -4206 -2133 -3226 -2116
rect -4206 -2139 -4126 -2133
rect -4434 -2162 -4354 -2139
rect -4434 -2196 -4411 -2162
rect -4377 -2173 -4354 -2162
rect -3249 -2140 -3226 -2133
rect -3192 -2140 -3169 -2106
rect -3249 -2163 -3169 -2140
rect -3069 -2126 -2989 -2080
rect -3069 -2160 -3046 -2126
rect -3012 -2160 -2989 -2126
rect -4377 -2196 -3289 -2173
rect -3069 -2183 -2989 -2160
rect -2919 -1966 -2839 -1933
rect -2919 -2000 -2896 -1966
rect -2862 -2000 -2839 -1966
rect -2919 -2046 -2839 -2000
rect -2919 -2080 -2896 -2046
rect -2862 -2080 -2839 -2046
rect -2919 -2126 -2839 -2080
rect -2919 -2160 -2896 -2126
rect -2862 -2160 -2839 -2126
rect -2919 -2193 -2839 -2160
rect -2769 -1966 -2689 -1933
rect -2769 -2000 -2746 -1966
rect -2712 -2000 -2689 -1966
rect -2769 -2046 -2689 -2000
rect -2769 -2080 -2746 -2046
rect -2712 -2080 -2689 -2046
rect -2769 -2126 -2689 -2080
rect -2769 -2160 -2746 -2126
rect -2712 -2160 -2689 -2126
rect -2769 -2183 -2689 -2160
rect -2619 -1966 -2539 -1933
rect -2619 -2000 -2596 -1966
rect -2562 -2000 -2539 -1966
rect -2619 -2046 -2539 -2000
rect -2619 -2080 -2596 -2046
rect -2562 -2080 -2539 -2046
rect -2619 -2126 -2539 -2080
rect -2619 -2160 -2596 -2126
rect -2562 -2160 -2539 -2126
rect -2619 -2193 -2539 -2160
rect -2469 -1966 -2389 -1933
rect -2469 -2000 -2446 -1966
rect -2412 -2000 -2389 -1966
rect -2469 -2046 -2389 -2000
rect -2089 -1986 -2009 -1963
rect -2089 -2020 -2066 -1986
rect -2032 -2020 -2009 -1986
rect -2089 -2043 -2009 -2020
rect -1019 -1966 -939 -1933
rect -1019 -2000 -996 -1966
rect -962 -2000 -939 -1966
rect -2469 -2080 -2446 -2046
rect -2412 -2080 -2389 -2046
rect -2469 -2126 -2389 -2080
rect -1019 -2046 -939 -2000
rect -1019 -2080 -996 -2046
rect -962 -2080 -939 -2046
rect -2469 -2160 -2446 -2126
rect -2412 -2160 -2389 -2126
rect -2469 -2183 -2389 -2160
rect -2219 -2106 -2139 -2083
rect -2219 -2140 -2196 -2106
rect -2162 -2140 -2139 -2106
rect -2219 -2163 -2139 -2140
rect -1457 -2123 -1377 -2103
rect -1169 -2123 -1089 -2103
rect -1457 -2126 -1089 -2123
rect -1457 -2160 -1434 -2126
rect -1400 -2160 -1146 -2126
rect -1112 -2160 -1089 -2126
rect -1457 -2163 -1089 -2160
rect -1457 -2183 -1377 -2163
rect -1169 -2183 -1089 -2163
rect -1019 -2126 -939 -2080
rect -1019 -2160 -996 -2126
rect -962 -2160 -939 -2126
rect -1019 -2183 -939 -2160
rect -869 -1966 -789 -1933
rect -869 -2000 -846 -1966
rect -812 -2000 -789 -1966
rect -869 -2046 -789 -2000
rect -869 -2080 -846 -2046
rect -812 -2080 -789 -2046
rect -869 -2126 -789 -2080
rect -869 -2160 -846 -2126
rect -812 -2160 -789 -2126
rect -869 -2193 -789 -2160
rect -719 -1966 -639 -1933
rect -719 -2000 -696 -1966
rect -662 -2000 -639 -1966
rect -719 -2046 -639 -2000
rect -719 -2080 -696 -2046
rect -662 -2080 -639 -2046
rect -719 -2126 -639 -2080
rect -719 -2160 -696 -2126
rect -662 -2160 -639 -2126
rect -719 -2183 -639 -2160
rect -569 -1966 -489 -1933
rect -569 -2000 -546 -1966
rect -512 -2000 -489 -1966
rect -569 -2046 -489 -2000
rect -569 -2080 -546 -2046
rect -512 -2080 -489 -2046
rect -569 -2126 -489 -2080
rect -569 -2160 -546 -2126
rect -512 -2160 -489 -2126
rect -569 -2193 -489 -2160
rect -419 -1966 -339 -1933
rect -419 -2000 -396 -1966
rect -362 -2000 -339 -1966
rect -419 -2046 -339 -2000
rect 114 -1953 194 -1930
rect 1771 -1934 1851 -1914
rect 2339 -1934 2419 -1914
rect 114 -1987 137 -1953
rect 171 -1987 194 -1953
rect 1021 -1967 1101 -1934
rect 114 -2010 194 -1987
rect 591 -1997 671 -1974
rect -419 -2080 -396 -2046
rect -362 -2080 -339 -2046
rect 591 -2031 614 -1997
rect 648 -2031 671 -1997
rect 591 -2054 671 -2031
rect 1021 -2001 1044 -1967
rect 1078 -2001 1101 -1967
rect 1021 -2047 1101 -2001
rect -419 -2126 -339 -2080
rect 791 -2087 871 -2064
rect -419 -2160 -396 -2126
rect -362 -2160 -339 -2126
rect -419 -2183 -339 -2160
rect -269 -2123 -189 -2103
rect -139 -2123 -59 -2103
rect -269 -2126 -59 -2123
rect 791 -2121 814 -2087
rect 848 -2121 871 -2087
rect -269 -2160 -246 -2126
rect -212 -2160 -116 -2126
rect -82 -2160 -59 -2126
rect 290 -2146 370 -2126
rect 791 -2144 871 -2121
rect 1021 -2081 1044 -2047
rect 1078 -2081 1101 -2047
rect 1021 -2127 1101 -2081
rect -269 -2163 -59 -2160
rect -269 -2183 -189 -2163
rect -139 -2183 -59 -2163
rect 176 -2149 370 -2146
rect 176 -2183 313 -2149
rect 347 -2183 370 -2149
rect 176 -2186 370 -2183
rect 1021 -2161 1044 -2127
rect 1078 -2161 1101 -2127
rect 1021 -2184 1101 -2161
rect 1171 -1967 1251 -1934
rect 1171 -2001 1194 -1967
rect 1228 -2001 1251 -1967
rect 1171 -2047 1251 -2001
rect 1171 -2081 1194 -2047
rect 1228 -2081 1251 -2047
rect 1171 -2127 1251 -2081
rect 1171 -2161 1194 -2127
rect 1228 -2161 1251 -2127
rect -4434 -2213 -3289 -2196
rect -4434 -2219 -4354 -2213
rect -3349 -2233 -3289 -2213
rect -4776 -2253 -4696 -2233
rect -4776 -2256 -3439 -2253
rect -4776 -2290 -4753 -2256
rect -4719 -2276 -3439 -2256
rect -4719 -2290 -3496 -2276
rect -4776 -2293 -3496 -2290
rect -4776 -2313 -4696 -2293
rect -3519 -2310 -3496 -2293
rect -3462 -2310 -3439 -2276
rect -3519 -2333 -3439 -2310
rect -3349 -2256 -3269 -2233
rect -3349 -2290 -3326 -2256
rect -3292 -2290 -3269 -2256
rect -3349 -2313 -3269 -2290
rect -2899 -2243 -2859 -2193
rect -2719 -2243 -2639 -2223
rect -2899 -2246 -2639 -2243
rect -2899 -2280 -2696 -2246
rect -2662 -2280 -2639 -2246
rect -2899 -2283 -2639 -2280
rect -4092 -2353 -4012 -2333
rect -3649 -2353 -3569 -2333
rect -4092 -2356 -3569 -2353
rect -4092 -2390 -4069 -2356
rect -4035 -2390 -3626 -2356
rect -3592 -2390 -3569 -2356
rect -4092 -2393 -3569 -2390
rect -4092 -2413 -4012 -2393
rect -3649 -2413 -3569 -2393
rect -2899 -2413 -2859 -2283
rect -2719 -2303 -2639 -2283
rect -3529 -2453 -2859 -2413
rect -2819 -2363 -2739 -2348
rect -2599 -2363 -2559 -2193
rect -2319 -2243 -2239 -2223
rect -849 -2243 -809 -2193
rect -669 -2243 -589 -2223
rect -2319 -2246 -1536 -2243
rect -2319 -2280 -2296 -2246
rect -2262 -2280 -1536 -2246
rect -2319 -2283 -1536 -2280
rect -2319 -2303 -2239 -2283
rect -1739 -2363 -1659 -2342
rect -2819 -2365 -1659 -2363
rect -2819 -2371 -1716 -2365
rect -2819 -2405 -2796 -2371
rect -2762 -2399 -1716 -2371
rect -1682 -2399 -1659 -2365
rect -2762 -2403 -1659 -2399
rect -1576 -2363 -1536 -2283
rect -849 -2246 -589 -2243
rect -849 -2280 -646 -2246
rect -612 -2280 -589 -2246
rect -849 -2283 -589 -2280
rect -1299 -2363 -1219 -2343
rect -1576 -2366 -1219 -2363
rect -1576 -2400 -1276 -2366
rect -1242 -2400 -1219 -2366
rect -1576 -2403 -1219 -2400
rect -2762 -2405 -2739 -2403
rect -2819 -2428 -2739 -2405
rect -3529 -2493 -3489 -2453
rect -3229 -2493 -3189 -2453
rect -2899 -2493 -2859 -2453
rect -2599 -2493 -2559 -2403
rect -2269 -2493 -2229 -2403
rect -1739 -2422 -1659 -2403
rect -1299 -2423 -1219 -2403
rect -849 -2413 -809 -2283
rect -669 -2303 -589 -2283
rect -1179 -2453 -809 -2413
rect -769 -2363 -689 -2348
rect -549 -2363 -509 -2193
rect -269 -2243 -189 -2223
rect 176 -2243 216 -2186
rect 290 -2206 370 -2186
rect 1171 -2194 1251 -2161
rect 1321 -1967 1401 -1934
rect 1321 -2001 1344 -1967
rect 1378 -2001 1401 -1967
rect 1321 -2047 1401 -2001
rect 1321 -2081 1344 -2047
rect 1378 -2081 1401 -2047
rect 1321 -2127 1401 -2081
rect 1321 -2161 1344 -2127
rect 1378 -2161 1401 -2127
rect 1321 -2184 1401 -2161
rect 1471 -1967 1551 -1934
rect 1471 -2001 1494 -1967
rect 1528 -2001 1551 -1967
rect 1471 -2047 1551 -2001
rect 1471 -2081 1494 -2047
rect 1528 -2081 1551 -2047
rect 1471 -2127 1551 -2081
rect 1471 -2161 1494 -2127
rect 1528 -2161 1551 -2127
rect 1471 -2194 1551 -2161
rect 1621 -1967 1701 -1934
rect 1621 -2001 1644 -1967
rect 1678 -2001 1701 -1967
rect 1621 -2047 1701 -2001
rect 1891 -1984 1971 -1964
rect 2143 -1984 2223 -1964
rect 1891 -1987 2351 -1984
rect 1891 -2021 1914 -1987
rect 1948 -2021 2166 -1987
rect 2200 -2021 2351 -1987
rect 1891 -2024 2351 -2021
rect 1891 -2044 1971 -2024
rect 2143 -2044 2223 -2024
rect 1621 -2081 1644 -2047
rect 1678 -2081 1701 -2047
rect 1621 -2127 1701 -2081
rect 1621 -2161 1644 -2127
rect 1678 -2161 1701 -2127
rect 1771 -2084 1851 -2064
rect 1771 -2087 2351 -2084
rect 1771 -2121 1794 -2087
rect 1828 -2121 2351 -2087
rect 1771 -2124 2351 -2121
rect 1771 -2144 1851 -2124
rect 1621 -2184 1701 -2161
rect 2385 -2174 2465 -2152
rect 2191 -2175 2465 -2174
rect -269 -2246 216 -2243
rect -269 -2280 -246 -2246
rect -212 -2280 216 -2246
rect -269 -2283 216 -2280
rect 291 -2244 371 -2240
rect 871 -2244 951 -2224
rect 291 -2247 951 -2244
rect 291 -2263 894 -2247
rect -269 -2303 -189 -2283
rect 291 -2297 314 -2263
rect 348 -2281 894 -2263
rect 928 -2281 951 -2247
rect 348 -2284 951 -2281
rect 348 -2297 371 -2284
rect 291 -2320 371 -2297
rect 871 -2304 951 -2284
rect -769 -2371 -509 -2363
rect -769 -2405 -746 -2371
rect -712 -2403 -509 -2371
rect 291 -2364 371 -2354
rect 1191 -2364 1231 -2194
rect 1271 -2244 1351 -2224
rect 1491 -2244 1531 -2194
rect 1271 -2247 1531 -2244
rect 1271 -2281 1294 -2247
rect 1328 -2281 1531 -2247
rect 2191 -2197 2408 -2175
rect 2191 -2231 2214 -2197
rect 2248 -2209 2408 -2197
rect 2442 -2209 2465 -2175
rect 2248 -2214 2465 -2209
rect 2248 -2231 2271 -2214
rect 2191 -2254 2271 -2231
rect 2385 -2232 2465 -2214
rect 1271 -2284 1531 -2281
rect 1271 -2304 1351 -2284
rect 1371 -2364 1451 -2349
rect 291 -2372 1451 -2364
rect 291 -2377 1394 -2372
rect -712 -2405 -689 -2403
rect -769 -2428 -689 -2405
rect -549 -2413 -509 -2403
rect 25 -2413 105 -2393
rect -549 -2416 105 -2413
rect -549 -2450 48 -2416
rect 82 -2450 105 -2416
rect 291 -2411 314 -2377
rect 348 -2404 1394 -2377
rect 348 -2411 371 -2404
rect 291 -2434 371 -2411
rect -549 -2453 105 -2450
rect -1179 -2493 -1139 -2453
rect -849 -2493 -809 -2453
rect -3699 -2526 -3619 -2493
rect -3699 -2560 -3676 -2526
rect -3642 -2560 -3619 -2526
rect -3699 -2606 -3619 -2560
rect -3699 -2640 -3676 -2606
rect -3642 -2640 -3619 -2606
rect -3699 -2686 -3619 -2640
rect -3699 -2720 -3676 -2686
rect -3642 -2720 -3619 -2686
rect -3699 -2743 -3619 -2720
rect -3549 -2526 -3469 -2493
rect -3549 -2560 -3526 -2526
rect -3492 -2560 -3469 -2526
rect -3549 -2606 -3469 -2560
rect -3549 -2640 -3526 -2606
rect -3492 -2640 -3469 -2606
rect -3549 -2686 -3469 -2640
rect -3549 -2720 -3526 -2686
rect -3492 -2720 -3469 -2686
rect -3549 -2743 -3469 -2720
rect -3399 -2526 -3319 -2493
rect -3399 -2560 -3376 -2526
rect -3342 -2560 -3319 -2526
rect -3399 -2606 -3319 -2560
rect -3399 -2640 -3376 -2606
rect -3342 -2640 -3319 -2606
rect -3399 -2686 -3319 -2640
rect -3399 -2720 -3376 -2686
rect -3342 -2720 -3319 -2686
rect -3399 -2743 -3319 -2720
rect -3249 -2526 -3169 -2493
rect -3249 -2560 -3226 -2526
rect -3192 -2560 -3169 -2526
rect -3249 -2606 -3169 -2560
rect -3249 -2640 -3226 -2606
rect -3192 -2640 -3169 -2606
rect -3249 -2686 -3169 -2640
rect -3249 -2720 -3226 -2686
rect -3192 -2720 -3169 -2686
rect -3249 -2743 -3169 -2720
rect -3069 -2526 -2989 -2493
rect -3069 -2560 -3046 -2526
rect -3012 -2560 -2989 -2526
rect -3069 -2606 -2989 -2560
rect -3069 -2640 -3046 -2606
rect -3012 -2640 -2989 -2606
rect -3069 -2686 -2989 -2640
rect -3069 -2720 -3046 -2686
rect -3012 -2720 -2989 -2686
rect -3069 -2743 -2989 -2720
rect -2919 -2526 -2839 -2493
rect -2919 -2560 -2896 -2526
rect -2862 -2560 -2839 -2526
rect -2919 -2606 -2839 -2560
rect -2919 -2640 -2896 -2606
rect -2862 -2640 -2839 -2606
rect -2919 -2686 -2839 -2640
rect -2919 -2720 -2896 -2686
rect -2862 -2720 -2839 -2686
rect -2919 -2743 -2839 -2720
rect -2769 -2526 -2689 -2493
rect -2769 -2560 -2746 -2526
rect -2712 -2560 -2689 -2526
rect -2769 -2606 -2689 -2560
rect -2769 -2640 -2746 -2606
rect -2712 -2640 -2689 -2606
rect -2769 -2686 -2689 -2640
rect -2769 -2720 -2746 -2686
rect -2712 -2720 -2689 -2686
rect -2769 -2743 -2689 -2720
rect -2619 -2526 -2539 -2493
rect -2619 -2560 -2596 -2526
rect -2562 -2560 -2539 -2526
rect -2619 -2606 -2539 -2560
rect -2619 -2640 -2596 -2606
rect -2562 -2640 -2539 -2606
rect -2619 -2686 -2539 -2640
rect -2619 -2720 -2596 -2686
rect -2562 -2720 -2539 -2686
rect -2619 -2743 -2539 -2720
rect -2469 -2526 -2389 -2493
rect -2469 -2560 -2446 -2526
rect -2412 -2560 -2389 -2526
rect -2469 -2606 -2389 -2560
rect -2469 -2640 -2446 -2606
rect -2412 -2640 -2389 -2606
rect -2469 -2686 -2389 -2640
rect -2469 -2720 -2446 -2686
rect -2412 -2720 -2389 -2686
rect -2469 -2743 -2389 -2720
rect -2289 -2526 -2209 -2493
rect -2289 -2560 -2266 -2526
rect -2232 -2560 -2209 -2526
rect -2289 -2606 -2209 -2560
rect -2289 -2640 -2266 -2606
rect -2232 -2640 -2209 -2606
rect -2289 -2686 -2209 -2640
rect -2289 -2720 -2266 -2686
rect -2232 -2720 -2209 -2686
rect -2289 -2743 -2209 -2720
rect -1839 -2526 -1759 -2493
rect -1839 -2560 -1816 -2526
rect -1782 -2560 -1759 -2526
rect -1839 -2606 -1759 -2560
rect -1839 -2640 -1816 -2606
rect -1782 -2640 -1759 -2606
rect -1839 -2686 -1759 -2640
rect -1839 -2720 -1816 -2686
rect -1782 -2720 -1759 -2686
rect -1839 -2743 -1759 -2720
rect -1349 -2526 -1269 -2493
rect -1349 -2560 -1326 -2526
rect -1292 -2560 -1269 -2526
rect -1349 -2606 -1269 -2560
rect -1349 -2640 -1326 -2606
rect -1292 -2640 -1269 -2606
rect -1349 -2686 -1269 -2640
rect -1349 -2720 -1326 -2686
rect -1292 -2720 -1269 -2686
rect -1349 -2743 -1269 -2720
rect -1199 -2526 -1119 -2493
rect -1199 -2560 -1176 -2526
rect -1142 -2560 -1119 -2526
rect -1199 -2606 -1119 -2560
rect -1199 -2640 -1176 -2606
rect -1142 -2640 -1119 -2606
rect -1199 -2686 -1119 -2640
rect -1199 -2720 -1176 -2686
rect -1142 -2720 -1119 -2686
rect -1199 -2743 -1119 -2720
rect -1019 -2526 -939 -2493
rect -1019 -2560 -996 -2526
rect -962 -2560 -939 -2526
rect -1019 -2606 -939 -2560
rect -1019 -2640 -996 -2606
rect -962 -2640 -939 -2606
rect -1019 -2686 -939 -2640
rect -1019 -2720 -996 -2686
rect -962 -2720 -939 -2686
rect -1019 -2743 -939 -2720
rect -869 -2526 -789 -2493
rect -869 -2560 -846 -2526
rect -812 -2560 -789 -2526
rect -869 -2606 -789 -2560
rect -869 -2640 -846 -2606
rect -812 -2640 -789 -2606
rect -869 -2686 -789 -2640
rect -869 -2720 -846 -2686
rect -812 -2720 -789 -2686
rect -869 -2743 -789 -2720
rect -719 -2526 -639 -2493
rect -719 -2560 -696 -2526
rect -662 -2560 -639 -2526
rect -719 -2606 -639 -2560
rect -719 -2640 -696 -2606
rect -662 -2640 -639 -2606
rect -719 -2686 -639 -2640
rect -719 -2720 -696 -2686
rect -662 -2720 -639 -2686
rect -719 -2743 -639 -2720
rect -569 -2526 -489 -2453
rect -219 -2493 -179 -2453
rect 25 -2473 105 -2453
rect -569 -2560 -546 -2526
rect -512 -2560 -489 -2526
rect -569 -2606 -489 -2560
rect -569 -2640 -546 -2606
rect -512 -2640 -489 -2606
rect -569 -2686 -489 -2640
rect -569 -2720 -546 -2686
rect -512 -2720 -489 -2686
rect -569 -2743 -489 -2720
rect -419 -2526 -339 -2493
rect -419 -2560 -396 -2526
rect -362 -2560 -339 -2526
rect -419 -2606 -339 -2560
rect -419 -2640 -396 -2606
rect -362 -2640 -339 -2606
rect -419 -2686 -339 -2640
rect -419 -2720 -396 -2686
rect -362 -2720 -339 -2686
rect -419 -2743 -339 -2720
rect -239 -2526 -159 -2493
rect -239 -2560 -216 -2526
rect -182 -2560 -159 -2526
rect -239 -2606 -159 -2560
rect -239 -2640 -216 -2606
rect -182 -2640 -159 -2606
rect -239 -2686 -159 -2640
rect -239 -2720 -216 -2686
rect -182 -2720 -159 -2686
rect -239 -2743 -159 -2720
rect -89 -2526 -9 -2493
rect 561 -2494 601 -2404
rect 861 -2494 901 -2404
rect 1191 -2494 1231 -2404
rect 1371 -2406 1394 -2404
rect 1428 -2406 1451 -2372
rect 1371 -2429 1451 -2406
rect 1491 -2414 1531 -2284
rect 2051 -2294 2131 -2274
rect 2499 -2294 2539 -1684
rect 2051 -2297 2539 -2294
rect 2051 -2331 2074 -2297
rect 2108 -2331 2539 -2297
rect 2051 -2334 2539 -2331
rect 2051 -2354 2131 -2334
rect 1901 -2377 1981 -2354
rect 1901 -2411 1924 -2377
rect 1958 -2394 1981 -2377
rect 1958 -2411 2351 -2394
rect 1491 -2454 1841 -2414
rect 1901 -2434 2351 -2411
rect 1491 -2494 1531 -2454
rect 1801 -2494 1841 -2454
rect -89 -2560 -66 -2526
rect -32 -2560 -9 -2526
rect -89 -2606 -9 -2560
rect 108 -2530 188 -2507
rect 108 -2564 131 -2530
rect 165 -2564 188 -2530
rect 108 -2587 188 -2564
rect 391 -2527 471 -2494
rect 391 -2561 414 -2527
rect 448 -2561 471 -2527
rect -89 -2640 -66 -2606
rect -32 -2640 -9 -2606
rect -89 -2686 -9 -2640
rect -89 -2720 -66 -2686
rect -32 -2720 -9 -2686
rect -89 -2743 -9 -2720
rect -3719 -2803 -3639 -2783
rect -2969 -2803 -2889 -2783
rect -2569 -2803 -2489 -2783
rect -919 -2803 -839 -2783
rect -519 -2803 -439 -2783
rect 128 -2803 168 -2587
rect 391 -2607 471 -2561
rect 391 -2641 414 -2607
rect 448 -2641 471 -2607
rect 391 -2687 471 -2641
rect 391 -2721 414 -2687
rect 448 -2721 471 -2687
rect 391 -2744 471 -2721
rect 541 -2527 621 -2494
rect 541 -2561 564 -2527
rect 598 -2561 621 -2527
rect 541 -2607 621 -2561
rect 541 -2641 564 -2607
rect 598 -2641 621 -2607
rect 541 -2687 621 -2641
rect 541 -2721 564 -2687
rect 598 -2721 621 -2687
rect 541 -2744 621 -2721
rect 691 -2527 771 -2494
rect 691 -2561 714 -2527
rect 748 -2561 771 -2527
rect 691 -2607 771 -2561
rect 691 -2641 714 -2607
rect 748 -2641 771 -2607
rect 691 -2687 771 -2641
rect 691 -2721 714 -2687
rect 748 -2721 771 -2687
rect 691 -2744 771 -2721
rect 841 -2527 921 -2494
rect 841 -2561 864 -2527
rect 898 -2561 921 -2527
rect 841 -2607 921 -2561
rect 841 -2641 864 -2607
rect 898 -2641 921 -2607
rect 841 -2687 921 -2641
rect 841 -2721 864 -2687
rect 898 -2721 921 -2687
rect 841 -2744 921 -2721
rect 1021 -2527 1101 -2494
rect 1021 -2561 1044 -2527
rect 1078 -2561 1101 -2527
rect 1021 -2607 1101 -2561
rect 1021 -2641 1044 -2607
rect 1078 -2641 1101 -2607
rect 1021 -2687 1101 -2641
rect 1021 -2721 1044 -2687
rect 1078 -2721 1101 -2687
rect 1021 -2744 1101 -2721
rect 1171 -2527 1251 -2494
rect 1171 -2561 1194 -2527
rect 1228 -2561 1251 -2527
rect 1171 -2607 1251 -2561
rect 1171 -2641 1194 -2607
rect 1228 -2641 1251 -2607
rect 1171 -2687 1251 -2641
rect 1171 -2721 1194 -2687
rect 1228 -2721 1251 -2687
rect 1171 -2744 1251 -2721
rect 1321 -2527 1401 -2494
rect 1321 -2561 1344 -2527
rect 1378 -2561 1401 -2527
rect 1321 -2607 1401 -2561
rect 1321 -2641 1344 -2607
rect 1378 -2641 1401 -2607
rect 1321 -2687 1401 -2641
rect 1321 -2721 1344 -2687
rect 1378 -2721 1401 -2687
rect 1321 -2744 1401 -2721
rect 1471 -2527 1551 -2494
rect 1471 -2561 1494 -2527
rect 1528 -2561 1551 -2527
rect 1471 -2607 1551 -2561
rect 1471 -2641 1494 -2607
rect 1528 -2641 1551 -2607
rect 1471 -2687 1551 -2641
rect 1471 -2721 1494 -2687
rect 1528 -2721 1551 -2687
rect 1471 -2744 1551 -2721
rect 1621 -2527 1701 -2494
rect 1621 -2561 1644 -2527
rect 1678 -2561 1701 -2527
rect 1621 -2607 1701 -2561
rect 1621 -2641 1644 -2607
rect 1678 -2641 1701 -2607
rect 1621 -2687 1701 -2641
rect 1621 -2721 1644 -2687
rect 1678 -2721 1701 -2687
rect 1621 -2744 1701 -2721
rect 1801 -2527 1881 -2494
rect 1801 -2561 1824 -2527
rect 1858 -2561 1881 -2527
rect 1801 -2607 1881 -2561
rect 1801 -2641 1824 -2607
rect 1858 -2641 1881 -2607
rect 1801 -2687 1881 -2641
rect 1801 -2721 1824 -2687
rect 1858 -2721 1881 -2687
rect 1801 -2744 1881 -2721
rect 2251 -2527 2331 -2494
rect 2251 -2561 2274 -2527
rect 2308 -2561 2331 -2527
rect 2251 -2607 2331 -2561
rect 2251 -2641 2274 -2607
rect 2308 -2641 2331 -2607
rect 2251 -2687 2331 -2641
rect 2251 -2721 2274 -2687
rect 2308 -2721 2331 -2687
rect 2251 -2744 2331 -2721
rect -3719 -2806 -2489 -2803
rect -3719 -2840 -3696 -2806
rect -3662 -2840 -2946 -2806
rect -2912 -2840 -2546 -2806
rect -2512 -2840 -2489 -2806
rect -3719 -2843 -2489 -2840
rect -1369 -2806 168 -2803
rect -1369 -2840 -896 -2806
rect -862 -2840 -496 -2806
rect -462 -2840 168 -2806
rect -1369 -2843 168 -2840
rect 202 -2804 282 -2785
rect 1121 -2804 1201 -2784
rect 1521 -2804 1601 -2784
rect 202 -2807 2351 -2804
rect 202 -2808 1144 -2807
rect 202 -2842 225 -2808
rect 259 -2841 1144 -2808
rect 1178 -2841 1544 -2807
rect 1578 -2841 2351 -2807
rect 259 -2842 2351 -2841
rect -3719 -2863 -3639 -2843
rect -2969 -2863 -2889 -2843
rect -2569 -2863 -2489 -2843
rect -919 -2863 -839 -2843
rect -519 -2863 -439 -2843
rect 202 -2844 2351 -2842
rect 202 -2865 282 -2844
rect 1121 -2864 1201 -2844
rect 1521 -2864 1601 -2844
rect -3978 -2926 -1729 -2903
rect -3978 -2960 -3955 -2926
rect -3921 -2960 -3706 -2926
rect -3672 -2960 -3626 -2926
rect -3592 -2960 -3546 -2926
rect -3512 -2960 -3466 -2926
rect -3432 -2960 -3386 -2926
rect -3352 -2960 -3306 -2926
rect -3272 -2960 -3226 -2926
rect -3192 -2960 -3146 -2926
rect -3112 -2960 -3066 -2926
rect -3032 -2960 -2986 -2926
rect -2952 -2960 -2906 -2926
rect -2872 -2960 -2826 -2926
rect -2792 -2960 -2746 -2926
rect -2712 -2960 -2666 -2926
rect -2632 -2960 -2586 -2926
rect -2552 -2960 -2506 -2926
rect -2472 -2960 -2426 -2926
rect -2392 -2960 -2346 -2926
rect -2312 -2960 -2266 -2926
rect -2232 -2960 -2186 -2926
rect -2152 -2960 -2106 -2926
rect -2072 -2960 -2026 -2926
rect -1992 -2960 -1946 -2926
rect -1912 -2960 -1866 -2926
rect -1832 -2960 -1786 -2926
rect -1752 -2960 -1729 -2926
rect -3978 -2983 -1729 -2960
rect -1369 -2926 11 -2903
rect -1369 -2960 -1336 -2926
rect -1302 -2960 -1256 -2926
rect -1222 -2960 -1176 -2926
rect -1142 -2960 -1096 -2926
rect -1062 -2960 -1016 -2926
rect -982 -2960 -936 -2926
rect -902 -2960 -856 -2926
rect -822 -2960 -776 -2926
rect -742 -2960 -696 -2926
rect -662 -2960 -616 -2926
rect -582 -2960 -536 -2926
rect -502 -2960 -456 -2926
rect -422 -2960 -376 -2926
rect -342 -2960 -296 -2926
rect -262 -2960 -216 -2926
rect -182 -2960 -136 -2926
rect -102 -2960 -56 -2926
rect -22 -2960 11 -2926
rect -1369 -2983 11 -2960
rect 361 -2927 2361 -2904
rect 361 -2961 384 -2927
rect 418 -2961 464 -2927
rect 498 -2961 544 -2927
rect 578 -2961 624 -2927
rect 658 -2961 704 -2927
rect 738 -2961 784 -2927
rect 818 -2961 864 -2927
rect 898 -2961 944 -2927
rect 978 -2961 1024 -2927
rect 1058 -2961 1104 -2927
rect 1138 -2961 1184 -2927
rect 1218 -2961 1264 -2927
rect 1298 -2961 1344 -2927
rect 1378 -2961 1424 -2927
rect 1458 -2961 1504 -2927
rect 1538 -2961 1584 -2927
rect 1618 -2961 1664 -2927
rect 1698 -2961 1744 -2927
rect 1778 -2961 1824 -2927
rect 1858 -2961 1904 -2927
rect 1938 -2961 1984 -2927
rect 2018 -2961 2064 -2927
rect 2098 -2961 2144 -2927
rect 2178 -2961 2224 -2927
rect 2258 -2961 2304 -2927
rect 2338 -2961 2361 -2927
rect 361 -2984 2361 -2961
<< viali >>
rect -3787 1040 -3753 1074
rect -3707 1040 -3673 1074
rect -3627 1040 -3593 1074
rect -3547 1040 -3513 1074
rect -3467 1040 -3433 1074
rect -3387 1040 -3353 1074
rect -3307 1040 -3273 1074
rect -3227 1040 -3193 1074
rect -3147 1040 -3113 1074
rect -3067 1040 -3033 1074
rect -2987 1040 -2953 1074
rect -2907 1040 -2873 1074
rect -2827 1040 -2793 1074
rect -2747 1040 -2713 1074
rect -2667 1040 -2633 1074
rect -2587 1040 -2553 1074
rect -2507 1040 -2473 1074
rect -2427 1040 -2393 1074
rect -2347 1040 -2313 1074
rect -2267 1040 -2233 1074
rect -2187 1040 -2153 1074
rect -2107 1040 -2073 1074
rect -2027 1040 -1993 1074
rect -1947 1040 -1913 1074
rect -1867 1040 -1833 1074
rect -1787 1040 -1753 1074
rect -1707 1040 -1673 1074
rect -1197 1040 -1163 1074
rect -1117 1040 -1083 1074
rect -1037 1040 -1003 1074
rect -957 1040 -923 1074
rect -877 1040 -843 1074
rect -797 1040 -763 1074
rect -717 1040 -683 1074
rect -637 1040 -603 1074
rect -557 1040 -523 1074
rect -477 1040 -443 1074
rect -397 1040 -363 1074
rect -317 1040 -283 1074
rect -237 1040 -203 1074
rect -157 1040 -123 1074
rect -77 1040 -43 1074
rect 3 1040 37 1074
rect 83 1040 117 1074
rect 523 1040 557 1074
rect 603 1040 637 1074
rect 683 1040 717 1074
rect 763 1040 797 1074
rect 843 1040 877 1074
rect 923 1040 957 1074
rect 1003 1040 1037 1074
rect 1083 1040 1117 1074
rect 1163 1040 1197 1074
rect 1243 1040 1277 1074
rect 1323 1040 1357 1074
rect 1403 1040 1437 1074
rect 1483 1040 1517 1074
rect 1563 1040 1597 1074
rect 1643 1040 1677 1074
rect 1723 1040 1757 1074
rect 1803 1040 1837 1074
rect 1883 1040 1917 1074
rect 1963 1040 1997 1074
rect 2043 1040 2077 1074
rect 2123 1040 2157 1074
rect -4639 910 -4605 944
rect -3327 910 -3293 944
rect -2067 910 -2033 944
rect -4525 810 -4491 844
rect -3197 810 -3163 844
rect -3047 820 -3013 854
rect -4867 710 -4833 744
rect -3327 710 -3293 744
rect -3047 740 -3013 774
rect -4753 610 -4719 644
rect -3197 610 -3163 644
rect -3047 660 -3013 694
rect -2747 820 -2713 854
rect -2747 740 -2713 774
rect -2747 660 -2713 694
rect -2447 820 -2413 854
rect -1867 810 -1833 844
rect -1295 844 -1261 878
rect -2447 740 -2413 774
rect -2447 660 -2413 694
rect -1717 710 -1683 744
rect -2697 540 -2663 574
rect -2167 610 -2133 644
rect -2327 530 -2293 564
rect -857 820 -823 854
rect -857 740 -823 774
rect -1007 660 -973 694
rect -857 660 -823 694
rect -557 820 -523 854
rect -557 740 -523 774
rect -557 660 -523 694
rect -257 820 -223 854
rect 443 810 477 844
rect 873 810 907 844
rect 1023 820 1057 854
rect -257 740 -223 774
rect -257 660 -223 694
rect -107 660 -73 694
rect -507 540 -473 574
rect -1567 416 -1533 450
rect -3527 260 -3493 294
rect -3527 180 -3493 214
rect -3527 100 -3493 134
rect -3047 260 -3013 294
rect -3047 180 -3013 214
rect -3047 100 -3013 134
rect -2747 260 -2713 294
rect -2747 180 -2713 214
rect -2747 100 -2713 134
rect -2447 260 -2413 294
rect -2447 180 -2413 214
rect -2447 100 -2413 134
rect -1967 260 -1933 294
rect -1967 180 -1933 214
rect -1967 100 -1933 134
rect -107 540 -73 574
rect 181 534 215 568
rect 873 690 907 724
rect 1023 740 1057 774
rect 1023 660 1057 694
rect 1323 820 1357 854
rect 1323 740 1357 774
rect 1323 660 1357 694
rect 1623 820 1657 854
rect 2003 810 2037 844
rect 1623 740 1657 774
rect 1623 660 1657 694
rect 1853 690 1887 724
rect 443 590 477 624
rect 443 470 477 504
rect 1373 540 1407 574
rect 1773 540 1807 574
rect 2206 420 2240 454
rect -1553 212 -1519 246
rect -1187 260 -1153 294
rect -1187 180 -1153 214
rect -1187 100 -1153 134
rect -857 260 -823 294
rect -857 180 -823 214
rect -857 100 -823 134
rect -557 260 -523 294
rect -557 180 -523 214
rect -557 100 -523 134
rect -257 260 -223 294
rect -257 180 -223 214
rect -257 100 -223 134
rect 73 260 107 294
rect 73 180 107 214
rect 73 100 107 134
rect 693 260 727 294
rect 693 180 727 214
rect 693 100 727 134
rect 1023 260 1057 294
rect 1023 180 1057 214
rect 1023 100 1057 134
rect 1323 260 1357 294
rect 1323 180 1357 214
rect 1323 100 1357 134
rect 1623 260 1657 294
rect 1623 180 1657 214
rect 1623 100 1657 134
rect 2103 260 2137 294
rect 2103 180 2137 214
rect 2103 100 2137 134
rect -3696 -20 -3662 14
rect 531 -20 565 14
rect -3955 -140 -3921 -106
rect -3787 -140 -3753 -106
rect -3707 -140 -3673 -106
rect -3627 -140 -3593 -106
rect -3547 -140 -3513 -106
rect -3467 -140 -3433 -106
rect -3387 -140 -3353 -106
rect -3307 -140 -3273 -106
rect -3227 -140 -3193 -106
rect -3147 -140 -3113 -106
rect -3067 -140 -3033 -106
rect -2987 -140 -2953 -106
rect -2907 -140 -2873 -106
rect -2827 -140 -2793 -106
rect -2747 -140 -2713 -106
rect -2667 -140 -2633 -106
rect -2587 -140 -2553 -106
rect -2507 -140 -2473 -106
rect -2427 -140 -2393 -106
rect -2347 -140 -2313 -106
rect -2267 -140 -2233 -106
rect -2187 -140 -2153 -106
rect -2107 -140 -2073 -106
rect -2027 -140 -1993 -106
rect -1947 -140 -1913 -106
rect -1867 -140 -1833 -106
rect -1787 -140 -1753 -106
rect -1707 -140 -1673 -106
rect -1197 -140 -1163 -106
rect -1117 -140 -1083 -106
rect -1037 -140 -1003 -106
rect -957 -140 -923 -106
rect -877 -140 -843 -106
rect -797 -140 -763 -106
rect -717 -140 -683 -106
rect -637 -140 -603 -106
rect -557 -140 -523 -106
rect -477 -140 -443 -106
rect -397 -140 -363 -106
rect -317 -140 -283 -106
rect -237 -140 -203 -106
rect -157 -140 -123 -106
rect -77 -140 -43 -106
rect 3 -140 37 -106
rect 83 -140 117 -106
rect 523 -140 557 -106
rect 603 -140 637 -106
rect 683 -140 717 -106
rect 763 -140 797 -106
rect 843 -140 877 -106
rect 923 -140 957 -106
rect 1003 -140 1037 -106
rect 1083 -140 1117 -106
rect 1163 -140 1197 -106
rect 1243 -140 1277 -106
rect 1323 -140 1357 -106
rect 1403 -140 1437 -106
rect 1483 -140 1517 -106
rect 1563 -140 1597 -106
rect 1643 -140 1677 -106
rect 1723 -140 1757 -106
rect 1803 -140 1837 -106
rect 1883 -140 1917 -106
rect 1963 -140 1997 -106
rect 2043 -140 2077 -106
rect 2123 -140 2157 -106
rect -3696 -260 -3662 -226
rect 531 -259 565 -225
rect -3527 -380 -3493 -346
rect -3527 -460 -3493 -426
rect -3527 -540 -3493 -506
rect -3047 -380 -3013 -346
rect -3047 -460 -3013 -426
rect -3047 -540 -3013 -506
rect -2747 -380 -2713 -346
rect -2747 -460 -2713 -426
rect -2747 -540 -2713 -506
rect -2447 -380 -2413 -346
rect -2447 -460 -2413 -426
rect -2447 -540 -2413 -506
rect -1967 -380 -1933 -346
rect -1967 -460 -1933 -426
rect -1967 -540 -1933 -506
rect -1187 -380 -1153 -346
rect -1553 -483 -1519 -449
rect -1187 -460 -1153 -426
rect -1187 -540 -1153 -506
rect -857 -380 -823 -346
rect -857 -460 -823 -426
rect -857 -540 -823 -506
rect -557 -380 -523 -346
rect -557 -460 -523 -426
rect -557 -540 -523 -506
rect -257 -380 -223 -346
rect -257 -460 -223 -426
rect -257 -540 -223 -506
rect 73 -380 107 -346
rect 73 -460 107 -426
rect 73 -540 107 -506
rect 693 -380 727 -346
rect 693 -460 727 -426
rect 693 -540 727 -506
rect 1023 -380 1057 -346
rect 1023 -460 1057 -426
rect 1023 -540 1057 -506
rect 1323 -380 1357 -346
rect 1323 -460 1357 -426
rect 1323 -540 1357 -506
rect 1623 -380 1657 -346
rect 1623 -460 1657 -426
rect 1623 -540 1657 -506
rect 2103 -380 2137 -346
rect 2103 -460 2137 -426
rect 2103 -540 2137 -506
rect -2697 -820 -2663 -786
rect -4069 -890 -4035 -856
rect -3197 -890 -3163 -856
rect -2327 -810 -2293 -776
rect -1567 -810 -1533 -776
rect -4183 -990 -4149 -956
rect -3327 -990 -3293 -956
rect -3047 -940 -3013 -906
rect -3047 -1020 -3013 -986
rect -4297 -1090 -4263 -1056
rect -3197 -1090 -3163 -1056
rect -3047 -1100 -3013 -1066
rect -2747 -940 -2713 -906
rect -2747 -1020 -2713 -986
rect -2747 -1100 -2713 -1066
rect -2447 -940 -2413 -906
rect -2167 -890 -2133 -856
rect -2447 -1020 -2413 -986
rect -1717 -990 -1683 -956
rect -2447 -1100 -2413 -1066
rect -1867 -1090 -1833 -1056
rect 181 -650 215 -616
rect -507 -820 -473 -786
rect -107 -820 -73 -786
rect 2206 -700 2240 -666
rect 1373 -820 1407 -786
rect 1773 -820 1807 -786
rect -1007 -940 -973 -906
rect -857 -940 -823 -906
rect -857 -1020 -823 -986
rect -1295 -1124 -1261 -1090
rect -4411 -1190 -4377 -1156
rect -3327 -1190 -3293 -1156
rect -857 -1100 -823 -1066
rect -557 -940 -523 -906
rect -557 -1020 -523 -986
rect -557 -1100 -523 -1066
rect -257 -940 -223 -906
rect -107 -940 -73 -906
rect -257 -1020 -223 -986
rect 181 -978 215 -944
rect 443 -970 477 -936
rect 873 -970 907 -936
rect 1023 -940 1057 -906
rect 1023 -1020 1057 -986
rect -257 -1100 -223 -1066
rect 443 -1091 477 -1057
rect 873 -1090 907 -1056
rect 1023 -1100 1057 -1066
rect 1323 -940 1357 -906
rect 1323 -1020 1357 -986
rect 1323 -1100 1357 -1066
rect 1623 -940 1657 -906
rect 1623 -1020 1657 -986
rect 1853 -970 1887 -936
rect 1623 -1100 1657 -1066
rect 2003 -1090 2037 -1056
rect -2067 -1190 -2033 -1156
rect -3787 -1320 -3753 -1286
rect -3707 -1320 -3673 -1286
rect -3627 -1320 -3593 -1286
rect -3547 -1320 -3513 -1286
rect -3467 -1320 -3433 -1286
rect -3387 -1320 -3353 -1286
rect -3307 -1320 -3273 -1286
rect -3227 -1320 -3193 -1286
rect -3147 -1320 -3113 -1286
rect -3067 -1320 -3033 -1286
rect -2987 -1320 -2953 -1286
rect -2907 -1320 -2873 -1286
rect -2827 -1320 -2793 -1286
rect -2747 -1320 -2713 -1286
rect -2667 -1320 -2633 -1286
rect -2587 -1320 -2553 -1286
rect -2507 -1320 -2473 -1286
rect -2427 -1320 -2393 -1286
rect -2347 -1320 -2313 -1286
rect -2267 -1320 -2233 -1286
rect -2187 -1320 -2153 -1286
rect -2107 -1320 -2073 -1286
rect -2027 -1320 -1993 -1286
rect -1947 -1320 -1913 -1286
rect -1867 -1320 -1833 -1286
rect -1787 -1320 -1753 -1286
rect -1707 -1320 -1673 -1286
rect -1197 -1320 -1163 -1286
rect -1117 -1320 -1083 -1286
rect -1037 -1320 -1003 -1286
rect -957 -1320 -923 -1286
rect -877 -1320 -843 -1286
rect -797 -1320 -763 -1286
rect -717 -1320 -683 -1286
rect -637 -1320 -603 -1286
rect -557 -1320 -523 -1286
rect -477 -1320 -443 -1286
rect -397 -1320 -363 -1286
rect -317 -1320 -283 -1286
rect -237 -1320 -203 -1286
rect -157 -1320 -123 -1286
rect -77 -1320 -43 -1286
rect 3 -1320 37 -1286
rect 83 -1320 117 -1286
rect 523 -1320 557 -1286
rect 603 -1320 637 -1286
rect 683 -1320 717 -1286
rect 763 -1320 797 -1286
rect 843 -1320 877 -1286
rect 923 -1320 957 -1286
rect 1003 -1320 1037 -1286
rect 1083 -1320 1117 -1286
rect 1163 -1320 1197 -1286
rect 1243 -1320 1277 -1286
rect 1323 -1320 1357 -1286
rect 1403 -1320 1437 -1286
rect 1483 -1320 1517 -1286
rect 1563 -1320 1597 -1286
rect 1643 -1320 1677 -1286
rect 1723 -1320 1757 -1286
rect 1803 -1320 1837 -1286
rect 1883 -1320 1917 -1286
rect 1963 -1320 1997 -1286
rect 2043 -1320 2077 -1286
rect 2123 -1320 2157 -1286
rect 531 -1554 565 -1520
rect -3706 -1780 -3672 -1746
rect -3626 -1780 -3592 -1746
rect -3546 -1780 -3512 -1746
rect -3466 -1780 -3432 -1746
rect -3386 -1780 -3352 -1746
rect -3306 -1780 -3272 -1746
rect -3226 -1780 -3192 -1746
rect -3146 -1780 -3112 -1746
rect -3066 -1780 -3032 -1746
rect -2986 -1780 -2952 -1746
rect -2906 -1780 -2872 -1746
rect -2826 -1780 -2792 -1746
rect -2746 -1780 -2712 -1746
rect -2666 -1780 -2632 -1746
rect -2586 -1780 -2552 -1746
rect -2506 -1780 -2472 -1746
rect -2426 -1780 -2392 -1746
rect -2346 -1780 -2312 -1746
rect -2266 -1780 -2232 -1746
rect -2186 -1780 -2152 -1746
rect -2106 -1780 -2072 -1746
rect -2026 -1780 -1992 -1746
rect -1946 -1780 -1912 -1746
rect -1866 -1780 -1832 -1746
rect -1786 -1780 -1752 -1746
rect -1336 -1780 -1302 -1746
rect -1256 -1780 -1222 -1746
rect -1176 -1780 -1142 -1746
rect -1096 -1780 -1062 -1746
rect -1016 -1780 -982 -1746
rect -936 -1780 -902 -1746
rect -856 -1780 -822 -1746
rect -776 -1780 -742 -1746
rect -696 -1780 -662 -1746
rect -616 -1780 -582 -1746
rect -536 -1780 -502 -1746
rect -456 -1780 -422 -1746
rect -376 -1780 -342 -1746
rect -296 -1780 -262 -1746
rect -216 -1780 -182 -1746
rect -136 -1780 -102 -1746
rect -56 -1780 -22 -1746
rect -4297 -1900 -4263 -1866
rect -3286 -1900 -3252 -1866
rect -1916 -1900 -1882 -1866
rect 2476 -1587 2510 -1553
rect 384 -1781 418 -1747
rect 464 -1781 498 -1747
rect 544 -1781 578 -1747
rect 624 -1781 658 -1747
rect 704 -1781 738 -1747
rect 784 -1781 818 -1747
rect 864 -1781 898 -1747
rect 944 -1781 978 -1747
rect 1024 -1781 1058 -1747
rect 1104 -1781 1138 -1747
rect 1184 -1781 1218 -1747
rect 1264 -1781 1298 -1747
rect 1344 -1781 1378 -1747
rect 1424 -1781 1458 -1747
rect 1504 -1781 1538 -1747
rect 1584 -1781 1618 -1747
rect 1664 -1781 1698 -1747
rect 1744 -1781 1778 -1747
rect 1824 -1781 1858 -1747
rect 1904 -1781 1938 -1747
rect 1984 -1781 2018 -1747
rect 2064 -1781 2098 -1747
rect 2144 -1781 2178 -1747
rect 2224 -1781 2258 -1747
rect 2304 -1781 2338 -1747
rect 514 -1906 548 -1872
rect 1794 -1911 1828 -1877
rect 2362 -1911 2396 -1877
rect -4867 -2020 -4833 -1986
rect -3196 -2020 -3162 -1986
rect -3046 -2000 -3012 -1966
rect -4183 -2116 -4149 -2082
rect -3046 -2080 -3012 -2046
rect -4411 -2196 -4377 -2162
rect -3226 -2140 -3192 -2106
rect -3046 -2160 -3012 -2126
rect -2746 -2000 -2712 -1966
rect -2746 -2080 -2712 -2046
rect -2746 -2160 -2712 -2126
rect -2446 -2000 -2412 -1966
rect -2066 -2020 -2032 -1986
rect -996 -2000 -962 -1966
rect -2446 -2080 -2412 -2046
rect -996 -2080 -962 -2046
rect -2446 -2160 -2412 -2126
rect -2196 -2140 -2162 -2106
rect -1434 -2160 -1400 -2126
rect -1146 -2160 -1112 -2126
rect -996 -2160 -962 -2126
rect -696 -2000 -662 -1966
rect -696 -2080 -662 -2046
rect -696 -2160 -662 -2126
rect -396 -2000 -362 -1966
rect 137 -1987 171 -1953
rect -396 -2080 -362 -2046
rect 614 -2031 648 -1997
rect 1044 -2001 1078 -1967
rect -396 -2160 -362 -2126
rect 814 -2121 848 -2087
rect -246 -2160 -212 -2126
rect 1044 -2081 1078 -2047
rect 313 -2183 347 -2149
rect 1044 -2161 1078 -2127
rect -4753 -2290 -4719 -2256
rect -2696 -2280 -2662 -2246
rect -4069 -2390 -4035 -2356
rect -2296 -2280 -2262 -2246
rect -1716 -2399 -1682 -2365
rect -646 -2280 -612 -2246
rect 1344 -2001 1378 -1967
rect 1344 -2081 1378 -2047
rect 1344 -2161 1378 -2127
rect 1644 -2001 1678 -1967
rect 1914 -2021 1948 -1987
rect 2166 -2021 2200 -1987
rect 1644 -2081 1678 -2047
rect 1644 -2161 1678 -2127
rect 1794 -2121 1828 -2087
rect -246 -2280 -212 -2246
rect 314 -2297 348 -2263
rect 894 -2281 928 -2247
rect 1294 -2281 1328 -2247
rect 2408 -2209 2442 -2175
rect 48 -2450 82 -2416
rect 314 -2411 348 -2377
rect -3676 -2560 -3642 -2526
rect -3676 -2640 -3642 -2606
rect -3676 -2720 -3642 -2686
rect -3376 -2560 -3342 -2526
rect -3376 -2640 -3342 -2606
rect -3376 -2720 -3342 -2686
rect -3046 -2560 -3012 -2526
rect -3046 -2640 -3012 -2606
rect -3046 -2720 -3012 -2686
rect -2746 -2560 -2712 -2526
rect -2746 -2640 -2712 -2606
rect -2746 -2720 -2712 -2686
rect -2446 -2560 -2412 -2526
rect -2446 -2640 -2412 -2606
rect -2446 -2720 -2412 -2686
rect -1816 -2560 -1782 -2526
rect -1816 -2640 -1782 -2606
rect -1816 -2720 -1782 -2686
rect -1326 -2560 -1292 -2526
rect -1326 -2640 -1292 -2606
rect -1326 -2720 -1292 -2686
rect -996 -2560 -962 -2526
rect -996 -2640 -962 -2606
rect -996 -2720 -962 -2686
rect -696 -2560 -662 -2526
rect -696 -2640 -662 -2606
rect -696 -2720 -662 -2686
rect -396 -2560 -362 -2526
rect -396 -2640 -362 -2606
rect -396 -2720 -362 -2686
rect 1924 -2411 1958 -2377
rect -66 -2560 -32 -2526
rect 131 -2564 165 -2530
rect 414 -2561 448 -2527
rect -66 -2640 -32 -2606
rect -66 -2720 -32 -2686
rect 414 -2641 448 -2607
rect 414 -2721 448 -2687
rect 714 -2561 748 -2527
rect 714 -2641 748 -2607
rect 714 -2721 748 -2687
rect 1044 -2561 1078 -2527
rect 1044 -2641 1078 -2607
rect 1044 -2721 1078 -2687
rect 1344 -2561 1378 -2527
rect 1344 -2641 1378 -2607
rect 1344 -2721 1378 -2687
rect 1644 -2561 1678 -2527
rect 1644 -2641 1678 -2607
rect 1644 -2721 1678 -2687
rect 2274 -2561 2308 -2527
rect 2274 -2641 2308 -2607
rect 2274 -2721 2308 -2687
rect -3696 -2840 -3662 -2806
rect 225 -2842 259 -2808
rect -3955 -2960 -3921 -2926
rect -3706 -2960 -3672 -2926
rect -3626 -2960 -3592 -2926
rect -3546 -2960 -3512 -2926
rect -3466 -2960 -3432 -2926
rect -3386 -2960 -3352 -2926
rect -3306 -2960 -3272 -2926
rect -3226 -2960 -3192 -2926
rect -3146 -2960 -3112 -2926
rect -3066 -2960 -3032 -2926
rect -2986 -2960 -2952 -2926
rect -2906 -2960 -2872 -2926
rect -2826 -2960 -2792 -2926
rect -2746 -2960 -2712 -2926
rect -2666 -2960 -2632 -2926
rect -2586 -2960 -2552 -2926
rect -2506 -2960 -2472 -2926
rect -2426 -2960 -2392 -2926
rect -2346 -2960 -2312 -2926
rect -2266 -2960 -2232 -2926
rect -2186 -2960 -2152 -2926
rect -2106 -2960 -2072 -2926
rect -2026 -2960 -1992 -2926
rect -1946 -2960 -1912 -2926
rect -1866 -2960 -1832 -2926
rect -1786 -2960 -1752 -2926
rect -1336 -2960 -1302 -2926
rect -1256 -2960 -1222 -2926
rect -1176 -2960 -1142 -2926
rect -1096 -2960 -1062 -2926
rect -1016 -2960 -982 -2926
rect -936 -2960 -902 -2926
rect -856 -2960 -822 -2926
rect -776 -2960 -742 -2926
rect -696 -2960 -662 -2926
rect -616 -2960 -582 -2926
rect -536 -2960 -502 -2926
rect -456 -2960 -422 -2926
rect -376 -2960 -342 -2926
rect -296 -2960 -262 -2926
rect -216 -2960 -182 -2926
rect -136 -2960 -102 -2926
rect -56 -2960 -22 -2926
rect 384 -2961 418 -2927
rect 464 -2961 498 -2927
rect 544 -2961 578 -2927
rect 624 -2961 658 -2927
rect 704 -2961 738 -2927
rect 784 -2961 818 -2927
rect 864 -2961 898 -2927
rect 944 -2961 978 -2927
rect 1024 -2961 1058 -2927
rect 1104 -2961 1138 -2927
rect 1184 -2961 1218 -2927
rect 1264 -2961 1298 -2927
rect 1344 -2961 1378 -2927
rect 1424 -2961 1458 -2927
rect 1504 -2961 1538 -2927
rect 1584 -2961 1618 -2927
rect 1664 -2961 1698 -2927
rect 1744 -2961 1778 -2927
rect 1824 -2961 1858 -2927
rect 1904 -2961 1938 -2927
rect 1984 -2961 2018 -2927
rect 2064 -2961 2098 -2927
rect 2144 -2961 2178 -2927
rect 2224 -2961 2258 -2927
rect 2304 -2961 2338 -2927
<< metal1 >>
rect -3870 1083 150 1107
rect -3870 1031 -3820 1083
rect -3768 1074 150 1083
rect -3753 1040 -3707 1074
rect -3673 1040 -3627 1074
rect -3593 1040 -3547 1074
rect -3513 1040 -3467 1074
rect -3433 1040 -3387 1074
rect -3353 1040 -3307 1074
rect -3273 1040 -3227 1074
rect -3193 1040 -3147 1074
rect -3113 1040 -3067 1074
rect -3033 1040 -2987 1074
rect -2953 1040 -2907 1074
rect -2873 1040 -2827 1074
rect -2793 1040 -2747 1074
rect -2713 1040 -2667 1074
rect -2633 1040 -2587 1074
rect -2553 1040 -2507 1074
rect -2473 1040 -2427 1074
rect -2393 1040 -2347 1074
rect -2313 1040 -2267 1074
rect -2233 1040 -2187 1074
rect -2153 1040 -2107 1074
rect -2073 1040 -2027 1074
rect -1993 1040 -1947 1074
rect -1913 1040 -1867 1074
rect -1833 1040 -1787 1074
rect -1753 1040 -1707 1074
rect -1673 1040 -1197 1074
rect -1163 1040 -1117 1074
rect -1083 1040 -1037 1074
rect -1003 1040 -957 1074
rect -923 1040 -877 1074
rect -843 1040 -797 1074
rect -763 1040 -717 1074
rect -683 1040 -637 1074
rect -603 1040 -557 1074
rect -523 1040 -477 1074
rect -443 1040 -397 1074
rect -363 1040 -317 1074
rect -283 1040 -237 1074
rect -203 1040 -157 1074
rect -123 1040 -77 1074
rect -43 1040 3 1074
rect 37 1040 83 1074
rect 117 1040 150 1074
rect -3768 1031 150 1040
rect -3870 1007 150 1031
rect 500 1083 2180 1107
rect 500 1074 2114 1083
rect 500 1040 523 1074
rect 557 1040 603 1074
rect 637 1040 683 1074
rect 717 1040 763 1074
rect 797 1040 843 1074
rect 877 1040 923 1074
rect 957 1040 1003 1074
rect 1037 1040 1083 1074
rect 1117 1040 1163 1074
rect 1197 1040 1243 1074
rect 1277 1040 1323 1074
rect 1357 1040 1403 1074
rect 1437 1040 1483 1074
rect 1517 1040 1563 1074
rect 1597 1040 1643 1074
rect 1677 1040 1723 1074
rect 1757 1040 1803 1074
rect 1837 1040 1883 1074
rect 1917 1040 1963 1074
rect 1997 1040 2043 1074
rect 2077 1040 2114 1074
rect 500 1031 2114 1040
rect 2166 1031 2180 1083
rect 500 1007 2180 1031
rect -4890 744 -4810 947
rect -4890 710 -4867 744
rect -4833 710 -4810 744
rect -4890 -1986 -4810 710
rect -4890 -2020 -4867 -1986
rect -4833 -2020 -4810 -1986
rect -4890 -3000 -4810 -2020
rect -4776 644 -4696 947
rect -4776 610 -4753 644
rect -4719 610 -4696 644
rect -4776 -2256 -4696 610
rect -4776 -2290 -4753 -2256
rect -4719 -2290 -4696 -2256
rect -4776 -3000 -4696 -2290
rect -4662 944 -4582 967
rect -4092 955 -4012 968
rect -4662 910 -4639 944
rect -4605 910 -4582 944
rect -4662 -1148 -4582 910
rect -4662 -1200 -4648 -1148
rect -4596 -1200 -4582 -1148
rect -4662 -3000 -4582 -1200
rect -4548 844 -4468 947
rect -4548 810 -4525 844
rect -4491 810 -4468 844
rect -4548 -441 -4468 810
rect -4548 -493 -4534 -441
rect -4482 -493 -4468 -441
rect -4548 -3000 -4468 -493
rect -4434 -1156 -4354 947
rect -4434 -1190 -4411 -1156
rect -4377 -1190 -4354 -1156
rect -4434 -2162 -4354 -1190
rect -4434 -2196 -4411 -2162
rect -4377 -2196 -4354 -2162
rect -4434 -3000 -4354 -2196
rect -4320 -1056 -4240 947
rect -4320 -1090 -4297 -1056
rect -4263 -1090 -4240 -1056
rect -4320 -1866 -4240 -1090
rect -4320 -1900 -4297 -1866
rect -4263 -1900 -4240 -1866
rect -4320 -3000 -4240 -1900
rect -4206 255 -4126 947
rect -4206 203 -4192 255
rect -4140 203 -4126 255
rect -4206 -956 -4126 203
rect -4206 -990 -4183 -956
rect -4149 -990 -4126 -956
rect -4206 -2082 -4126 -990
rect -4206 -2116 -4183 -2082
rect -4149 -2116 -4126 -2082
rect -4206 -3000 -4126 -2116
rect -4092 903 -4078 955
rect -4026 903 -4012 955
rect -4092 -856 -4012 903
rect -3530 327 -3490 1007
rect -3350 953 -3270 967
rect -3350 901 -3336 953
rect -3284 901 -3270 953
rect -3350 887 -3270 901
rect -3220 853 -3140 867
rect -3220 801 -3206 853
rect -3154 801 -3140 853
rect -3220 787 -3140 801
rect -3070 854 -2990 1007
rect -3070 820 -3047 854
rect -3013 820 -2990 854
rect -3070 774 -2990 820
rect -3350 753 -3270 767
rect -3350 701 -3336 753
rect -3284 701 -3270 753
rect -3350 687 -3270 701
rect -3070 740 -3047 774
rect -3013 740 -2990 774
rect -3070 694 -2990 740
rect -3220 653 -3140 667
rect -3220 601 -3206 653
rect -3154 601 -3140 653
rect -3070 660 -3047 694
rect -3013 660 -2990 694
rect -3070 637 -2990 660
rect -2770 854 -2690 1007
rect -2770 820 -2747 854
rect -2713 820 -2690 854
rect -2770 774 -2690 820
rect -2770 740 -2747 774
rect -2713 740 -2690 774
rect -2770 694 -2690 740
rect -2770 660 -2747 694
rect -2713 660 -2690 694
rect -2770 637 -2690 660
rect -2470 854 -2390 1007
rect -2090 953 -2010 967
rect -2090 901 -2076 953
rect -2024 901 -2010 953
rect -2090 887 -2010 901
rect -2470 820 -2447 854
rect -2413 820 -2390 854
rect -2470 774 -2390 820
rect -2470 740 -2447 774
rect -2413 740 -2390 774
rect -2470 694 -2390 740
rect -2470 660 -2447 694
rect -2413 660 -2390 694
rect -2470 637 -2390 660
rect -2190 653 -2110 667
rect -3220 587 -3140 601
rect -2190 601 -2176 653
rect -2124 601 -2110 653
rect -2720 574 -2640 597
rect -2190 587 -2110 601
rect -2720 540 -2697 574
rect -2663 557 -2640 574
rect -2350 564 -2270 587
rect -2350 557 -2327 564
rect -2663 540 -2327 557
rect -2720 530 -2327 540
rect -2293 530 -2270 564
rect -2720 517 -2270 530
rect -2350 507 -2270 517
rect -1970 327 -1930 1007
rect -1318 887 -1238 901
rect -1890 853 -1810 867
rect -1890 801 -1876 853
rect -1824 801 -1810 853
rect -1318 835 -1304 887
rect -1252 835 -1238 887
rect -1318 821 -1238 835
rect -1890 787 -1810 801
rect -1318 776 -1238 790
rect -1740 753 -1660 767
rect -1740 701 -1726 753
rect -1674 701 -1660 753
rect -1318 724 -1304 776
rect -1252 724 -1238 776
rect -1318 710 -1238 724
rect -1740 687 -1660 701
rect -1590 452 -1510 473
rect -1299 452 -1259 710
rect -1590 450 -1259 452
rect -1590 416 -1567 450
rect -1533 416 -1259 450
rect -1590 412 -1259 416
rect -1590 393 -1510 412
rect -3550 294 -3470 327
rect -3550 260 -3527 294
rect -3493 260 -3470 294
rect -3550 214 -3470 260
rect -3550 180 -3527 214
rect -3493 180 -3470 214
rect -3550 134 -3470 180
rect -3550 100 -3527 134
rect -3493 100 -3470 134
rect -3550 77 -3470 100
rect -3070 294 -2990 327
rect -3070 260 -3047 294
rect -3013 260 -2990 294
rect -3070 214 -2990 260
rect -3070 180 -3047 214
rect -3013 180 -2990 214
rect -3070 134 -2990 180
rect -3070 100 -3047 134
rect -3013 100 -2990 134
rect -3070 77 -2990 100
rect -2770 294 -2690 327
rect -2770 260 -2747 294
rect -2713 260 -2690 294
rect -2770 214 -2690 260
rect -2770 180 -2747 214
rect -2713 180 -2690 214
rect -2770 134 -2690 180
rect -2770 100 -2747 134
rect -2713 100 -2690 134
rect -2770 77 -2690 100
rect -2470 294 -2390 327
rect -2470 260 -2447 294
rect -2413 260 -2390 294
rect -2470 214 -2390 260
rect -2470 180 -2447 214
rect -2413 180 -2390 214
rect -2470 134 -2390 180
rect -2470 100 -2447 134
rect -2413 100 -2390 134
rect -2470 77 -2390 100
rect -1990 294 -1910 327
rect -1990 260 -1967 294
rect -1933 260 -1910 294
rect -1210 294 -1130 1007
rect -1030 956 -950 969
rect -1030 904 -1016 956
rect -964 904 -950 956
rect -1030 889 -950 904
rect -1010 717 -970 889
rect -880 854 -800 1007
rect -880 820 -857 854
rect -823 820 -800 854
rect -880 774 -800 820
rect -880 740 -857 774
rect -823 740 -800 774
rect -1030 703 -950 717
rect -1030 651 -1016 703
rect -964 651 -950 703
rect -1030 637 -950 651
rect -880 694 -800 740
rect -880 660 -857 694
rect -823 660 -800 694
rect -880 637 -800 660
rect -580 854 -500 1007
rect -580 820 -557 854
rect -523 820 -500 854
rect -580 774 -500 820
rect -580 740 -557 774
rect -523 740 -500 774
rect -580 694 -500 740
rect -580 660 -557 694
rect -523 660 -500 694
rect -580 637 -500 660
rect -280 854 -200 1007
rect -280 820 -257 854
rect -223 820 -200 854
rect -280 774 -200 820
rect -280 740 -257 774
rect -223 740 -200 774
rect -280 694 -200 740
rect -280 660 -257 694
rect -223 660 -200 694
rect -280 637 -200 660
rect -130 703 -50 717
rect -130 651 -116 703
rect -64 651 -50 703
rect -130 637 -50 651
rect -530 577 -450 597
rect -130 577 -50 597
rect -530 574 -50 577
rect -530 540 -507 574
rect -473 540 -107 574
rect -73 540 -50 574
rect -530 537 -50 540
rect -530 517 -450 537
rect -130 517 -50 537
rect -1990 214 -1910 260
rect -1990 180 -1967 214
rect -1933 180 -1910 214
rect -1576 255 -1496 268
rect -1576 203 -1562 255
rect -1510 203 -1496 255
rect -1576 188 -1496 203
rect -1210 260 -1187 294
rect -1153 260 -1130 294
rect -1210 214 -1130 260
rect -1990 134 -1910 180
rect -1990 100 -1967 134
rect -1933 100 -1910 134
rect -1990 77 -1910 100
rect -1210 180 -1187 214
rect -1153 180 -1130 214
rect -1210 134 -1130 180
rect -1210 100 -1187 134
rect -1153 100 -1130 134
rect -1210 77 -1130 100
rect -880 294 -800 327
rect -880 260 -857 294
rect -823 260 -800 294
rect -880 214 -800 260
rect -880 180 -857 214
rect -823 180 -800 214
rect -880 134 -800 180
rect -880 100 -857 134
rect -823 100 -800 134
rect -880 77 -800 100
rect -580 294 -500 327
rect -580 260 -557 294
rect -523 260 -500 294
rect -580 214 -500 260
rect -580 180 -557 214
rect -523 180 -500 214
rect -580 134 -500 180
rect -580 100 -557 134
rect -523 100 -500 134
rect -580 77 -500 100
rect -280 294 -200 327
rect -280 260 -257 294
rect -223 260 -200 294
rect -280 214 -200 260
rect -280 180 -257 214
rect -223 180 -200 214
rect -280 134 -200 180
rect -280 100 -257 134
rect -223 100 -200 134
rect -280 77 -200 100
rect 50 294 130 1007
rect 158 866 238 880
rect 158 814 172 866
rect 224 852 238 866
rect 420 852 500 867
rect 224 844 500 852
rect 224 814 443 844
rect 158 812 443 814
rect 158 800 238 812
rect 420 810 443 812
rect 477 810 500 844
rect 420 787 500 810
rect 158 757 238 771
rect 158 705 172 757
rect 224 751 238 757
rect 224 711 480 751
rect 224 705 238 711
rect 158 691 238 705
rect 440 647 480 711
rect 420 624 500 647
rect 158 568 238 591
rect 158 534 181 568
rect 215 534 238 568
rect 420 590 443 624
rect 477 590 500 624
rect 420 567 500 590
rect 158 511 238 534
rect 420 511 500 527
rect 158 504 500 511
rect 158 471 443 504
rect 420 470 443 471
rect 477 470 500 504
rect 420 447 500 470
rect 690 327 730 1007
rect 850 853 930 867
rect 850 801 864 853
rect 916 801 930 853
rect 850 787 930 801
rect 1000 854 1080 1007
rect 1000 820 1023 854
rect 1057 820 1080 854
rect 1000 774 1080 820
rect 850 733 930 747
rect 850 681 864 733
rect 916 681 930 733
rect 850 667 930 681
rect 1000 740 1023 774
rect 1057 740 1080 774
rect 1000 694 1080 740
rect 1000 660 1023 694
rect 1057 660 1080 694
rect 1000 637 1080 660
rect 1300 854 1380 1007
rect 1300 820 1323 854
rect 1357 820 1380 854
rect 1300 774 1380 820
rect 1300 740 1323 774
rect 1357 740 1380 774
rect 1300 694 1380 740
rect 1300 660 1323 694
rect 1357 660 1380 694
rect 1300 637 1380 660
rect 1600 854 1680 1007
rect 1600 820 1623 854
rect 1657 820 1680 854
rect 1600 774 1680 820
rect 1980 853 2060 867
rect 1980 801 1994 853
rect 2046 801 2060 853
rect 1980 787 2060 801
rect 1600 740 1623 774
rect 1657 740 1680 774
rect 1600 694 1680 740
rect 1600 660 1623 694
rect 1657 660 1680 694
rect 1830 733 1910 747
rect 1830 681 1844 733
rect 1896 681 1910 733
rect 1830 667 1910 681
rect 1600 637 1680 660
rect 1350 577 1430 597
rect 1750 577 1830 597
rect 1350 574 1830 577
rect 1350 540 1373 574
rect 1407 540 1773 574
rect 1807 540 1830 574
rect 1350 537 1830 540
rect 1350 517 1430 537
rect 1750 517 1830 537
rect 2100 327 2140 1007
rect 2183 463 2263 477
rect 2183 411 2197 463
rect 2249 411 2263 463
rect 2183 397 2263 411
rect 50 260 73 294
rect 107 260 130 294
rect 50 214 130 260
rect 50 180 73 214
rect 107 180 130 214
rect 50 134 130 180
rect 50 100 73 134
rect 107 100 130 134
rect 50 77 130 100
rect 670 294 750 327
rect 670 260 693 294
rect 727 260 750 294
rect 670 214 750 260
rect 670 180 693 214
rect 727 180 750 214
rect 670 134 750 180
rect 670 100 693 134
rect 727 100 750 134
rect 670 77 750 100
rect 1000 294 1080 327
rect 1000 260 1023 294
rect 1057 260 1080 294
rect 1000 214 1080 260
rect 1000 180 1023 214
rect 1057 180 1080 214
rect 1000 134 1080 180
rect 1000 100 1023 134
rect 1057 100 1080 134
rect 1000 77 1080 100
rect 1300 294 1380 327
rect 1300 260 1323 294
rect 1357 260 1380 294
rect 1300 214 1380 260
rect 1300 180 1323 214
rect 1357 180 1380 214
rect 1300 134 1380 180
rect 1300 100 1323 134
rect 1357 100 1380 134
rect 1300 77 1380 100
rect 1600 294 1680 327
rect 1600 260 1623 294
rect 1657 260 1680 294
rect 1600 214 1680 260
rect 1600 180 1623 214
rect 1657 180 1680 214
rect 1600 134 1680 180
rect 1600 100 1623 134
rect 1657 100 1680 134
rect 1600 77 1680 100
rect 2080 294 2160 327
rect 2080 260 2103 294
rect 2137 260 2160 294
rect 2080 214 2160 260
rect 2080 180 2103 214
rect 2137 180 2160 214
rect 2080 143 2160 180
rect 2080 91 2094 143
rect 2146 91 2160 143
rect 2080 77 2160 91
rect -3719 23 -3639 37
rect -3719 -29 -3705 23
rect -3653 -29 -3639 23
rect -3719 -43 -3639 -29
rect -3050 -73 -3010 77
rect -2750 -73 -2710 77
rect -2450 -73 -2410 77
rect -860 -73 -820 77
rect -560 -73 -520 77
rect -260 -73 -220 77
rect 508 23 588 37
rect 508 -29 522 23
rect 574 -29 588 23
rect 508 -43 588 -29
rect 1020 -73 1060 77
rect 1320 -73 1360 77
rect 1620 -73 1660 77
rect -4092 -890 -4069 -856
rect -4035 -890 -4012 -856
rect -4092 -2356 -4012 -890
rect -4092 -2390 -4069 -2356
rect -4035 -2390 -4012 -2356
rect -4092 -2999 -4012 -2390
rect -3978 -106 -3898 -83
rect -3978 -140 -3955 -106
rect -3921 -140 -3898 -106
rect -3978 -2926 -3898 -140
rect -3870 -106 2180 -73
rect -3870 -140 -3787 -106
rect -3753 -140 -3707 -106
rect -3673 -140 -3627 -106
rect -3593 -140 -3547 -106
rect -3513 -140 -3467 -106
rect -3433 -140 -3387 -106
rect -3353 -140 -3307 -106
rect -3273 -140 -3227 -106
rect -3193 -140 -3147 -106
rect -3113 -140 -3067 -106
rect -3033 -140 -2987 -106
rect -2953 -140 -2907 -106
rect -2873 -140 -2827 -106
rect -2793 -140 -2747 -106
rect -2713 -140 -2667 -106
rect -2633 -140 -2587 -106
rect -2553 -140 -2507 -106
rect -2473 -140 -2427 -106
rect -2393 -140 -2347 -106
rect -2313 -140 -2267 -106
rect -2233 -140 -2187 -106
rect -2153 -140 -2107 -106
rect -2073 -140 -2027 -106
rect -1993 -140 -1947 -106
rect -1913 -140 -1867 -106
rect -1833 -140 -1787 -106
rect -1753 -140 -1707 -106
rect -1673 -140 -1197 -106
rect -1163 -140 -1117 -106
rect -1083 -140 -1037 -106
rect -1003 -140 -957 -106
rect -923 -140 -877 -106
rect -843 -140 -797 -106
rect -763 -140 -717 -106
rect -683 -140 -637 -106
rect -603 -140 -557 -106
rect -523 -140 -477 -106
rect -443 -140 -397 -106
rect -363 -140 -317 -106
rect -283 -140 -237 -106
rect -203 -140 -157 -106
rect -123 -140 -77 -106
rect -43 -140 3 -106
rect 37 -140 83 -106
rect 117 -140 523 -106
rect 557 -140 603 -106
rect 637 -140 683 -106
rect 717 -140 763 -106
rect 797 -140 843 -106
rect 877 -140 923 -106
rect 957 -140 1003 -106
rect 1037 -140 1083 -106
rect 1117 -140 1163 -106
rect 1197 -140 1243 -106
rect 1277 -140 1323 -106
rect 1357 -140 1403 -106
rect 1437 -140 1483 -106
rect 1517 -140 1563 -106
rect 1597 -140 1643 -106
rect 1677 -140 1723 -106
rect 1757 -140 1803 -106
rect 1837 -140 1883 -106
rect 1917 -140 1963 -106
rect 1997 -140 2043 -106
rect 2077 -140 2123 -106
rect 2157 -140 2180 -106
rect -3870 -173 2180 -140
rect -3719 -217 -3639 -203
rect -3719 -269 -3705 -217
rect -3653 -269 -3639 -217
rect -3719 -283 -3639 -269
rect -3050 -323 -3010 -173
rect -2750 -323 -2710 -173
rect -2450 -323 -2410 -173
rect -860 -323 -820 -173
rect -560 -323 -520 -173
rect -260 -323 -220 -173
rect 508 -216 588 -202
rect 508 -268 522 -216
rect 574 -268 588 -216
rect 508 -282 588 -268
rect 1020 -323 1060 -173
rect 1320 -323 1360 -173
rect 1620 -323 1660 -173
rect -3550 -346 -3470 -323
rect -3550 -380 -3527 -346
rect -3493 -380 -3470 -346
rect -3550 -426 -3470 -380
rect -3550 -460 -3527 -426
rect -3493 -460 -3470 -426
rect -3550 -506 -3470 -460
rect -3550 -540 -3527 -506
rect -3493 -540 -3470 -506
rect -3550 -573 -3470 -540
rect -3070 -346 -2990 -323
rect -3070 -380 -3047 -346
rect -3013 -380 -2990 -346
rect -3070 -426 -2990 -380
rect -3070 -460 -3047 -426
rect -3013 -460 -2990 -426
rect -3070 -506 -2990 -460
rect -3070 -540 -3047 -506
rect -3013 -540 -2990 -506
rect -3070 -573 -2990 -540
rect -2770 -346 -2690 -323
rect -2770 -380 -2747 -346
rect -2713 -380 -2690 -346
rect -2770 -426 -2690 -380
rect -2770 -460 -2747 -426
rect -2713 -460 -2690 -426
rect -2770 -506 -2690 -460
rect -2770 -540 -2747 -506
rect -2713 -540 -2690 -506
rect -2770 -573 -2690 -540
rect -2470 -346 -2390 -323
rect -2470 -380 -2447 -346
rect -2413 -380 -2390 -346
rect -2470 -426 -2390 -380
rect -2470 -460 -2447 -426
rect -2413 -460 -2390 -426
rect -2470 -506 -2390 -460
rect -2470 -540 -2447 -506
rect -2413 -540 -2390 -506
rect -2470 -573 -2390 -540
rect -1990 -346 -1910 -323
rect -1990 -380 -1967 -346
rect -1933 -380 -1910 -346
rect -1990 -426 -1910 -380
rect -1990 -460 -1967 -426
rect -1933 -460 -1910 -426
rect -1210 -346 -1130 -323
rect -1210 -380 -1187 -346
rect -1153 -380 -1130 -346
rect -1210 -426 -1130 -380
rect -1990 -506 -1910 -460
rect -1990 -540 -1967 -506
rect -1933 -540 -1910 -506
rect -1576 -440 -1496 -427
rect -1576 -492 -1562 -440
rect -1510 -492 -1496 -440
rect -1576 -507 -1496 -492
rect -1210 -460 -1187 -426
rect -1153 -460 -1130 -426
rect -1210 -506 -1130 -460
rect -1990 -573 -1910 -540
rect -1210 -540 -1187 -506
rect -1153 -540 -1130 -506
rect -3530 -1253 -3490 -573
rect -2350 -763 -2270 -753
rect -2720 -776 -2270 -763
rect -2720 -786 -2327 -776
rect -2720 -820 -2697 -786
rect -2663 -803 -2327 -786
rect -2663 -820 -2640 -803
rect -3220 -847 -3140 -833
rect -2720 -843 -2640 -820
rect -2350 -810 -2327 -803
rect -2293 -810 -2270 -776
rect -2350 -833 -2270 -810
rect -3220 -899 -3206 -847
rect -3154 -899 -3140 -847
rect -2190 -847 -2110 -833
rect -3220 -913 -3140 -899
rect -3070 -906 -2990 -883
rect -3350 -947 -3270 -933
rect -3350 -999 -3336 -947
rect -3284 -999 -3270 -947
rect -3350 -1013 -3270 -999
rect -3070 -940 -3047 -906
rect -3013 -940 -2990 -906
rect -3070 -986 -2990 -940
rect -3070 -1020 -3047 -986
rect -3013 -1020 -2990 -986
rect -3220 -1047 -3140 -1033
rect -3220 -1099 -3206 -1047
rect -3154 -1099 -3140 -1047
rect -3220 -1113 -3140 -1099
rect -3070 -1066 -2990 -1020
rect -3070 -1100 -3047 -1066
rect -3013 -1100 -2990 -1066
rect -3350 -1147 -3270 -1133
rect -3350 -1199 -3336 -1147
rect -3284 -1199 -3270 -1147
rect -3350 -1213 -3270 -1199
rect -3070 -1253 -2990 -1100
rect -2770 -906 -2690 -883
rect -2770 -940 -2747 -906
rect -2713 -940 -2690 -906
rect -2770 -986 -2690 -940
rect -2770 -1020 -2747 -986
rect -2713 -1020 -2690 -986
rect -2770 -1066 -2690 -1020
rect -2770 -1100 -2747 -1066
rect -2713 -1100 -2690 -1066
rect -2770 -1253 -2690 -1100
rect -2470 -906 -2390 -883
rect -2470 -940 -2447 -906
rect -2413 -940 -2390 -906
rect -2190 -899 -2176 -847
rect -2124 -899 -2110 -847
rect -2190 -913 -2110 -899
rect -2470 -986 -2390 -940
rect -2470 -1020 -2447 -986
rect -2413 -1020 -2390 -986
rect -2470 -1066 -2390 -1020
rect -2470 -1100 -2447 -1066
rect -2413 -1100 -2390 -1066
rect -2470 -1253 -2390 -1100
rect -2090 -1147 -2010 -1133
rect -2090 -1199 -2076 -1147
rect -2024 -1199 -2010 -1147
rect -2090 -1213 -2010 -1199
rect -1970 -1253 -1930 -573
rect -1590 -776 -1259 -753
rect -1590 -810 -1567 -776
rect -1533 -793 -1259 -776
rect -1533 -810 -1510 -793
rect -1590 -833 -1510 -810
rect -1740 -947 -1660 -933
rect -1740 -999 -1726 -947
rect -1674 -999 -1660 -947
rect -1299 -954 -1259 -793
rect -1740 -1013 -1660 -999
rect -1318 -968 -1238 -954
rect -1318 -1020 -1304 -968
rect -1252 -1020 -1238 -968
rect -1890 -1047 -1810 -1033
rect -1318 -1034 -1238 -1020
rect -1890 -1099 -1876 -1047
rect -1824 -1099 -1810 -1047
rect -1890 -1113 -1810 -1099
rect -1318 -1081 -1238 -1067
rect -1318 -1133 -1304 -1081
rect -1252 -1133 -1238 -1081
rect -1318 -1147 -1238 -1133
rect -1210 -1253 -1130 -540
rect -880 -346 -800 -323
rect -880 -380 -857 -346
rect -823 -380 -800 -346
rect -880 -426 -800 -380
rect -880 -460 -857 -426
rect -823 -460 -800 -426
rect -880 -506 -800 -460
rect -880 -540 -857 -506
rect -823 -540 -800 -506
rect -880 -573 -800 -540
rect -580 -346 -500 -323
rect -580 -380 -557 -346
rect -523 -380 -500 -346
rect -580 -426 -500 -380
rect -580 -460 -557 -426
rect -523 -460 -500 -426
rect -580 -506 -500 -460
rect -580 -540 -557 -506
rect -523 -540 -500 -506
rect -580 -573 -500 -540
rect -280 -346 -200 -323
rect -280 -380 -257 -346
rect -223 -380 -200 -346
rect -280 -426 -200 -380
rect -280 -460 -257 -426
rect -223 -460 -200 -426
rect -280 -506 -200 -460
rect -280 -540 -257 -506
rect -223 -540 -200 -506
rect -280 -573 -200 -540
rect 50 -346 130 -323
rect 50 -380 73 -346
rect 107 -380 130 -346
rect 50 -426 130 -380
rect 50 -460 73 -426
rect 107 -460 130 -426
rect 50 -506 130 -460
rect 50 -540 73 -506
rect 107 -540 130 -506
rect -530 -783 -450 -763
rect -130 -783 -50 -763
rect -530 -786 -50 -783
rect -530 -820 -507 -786
rect -473 -820 -107 -786
rect -73 -820 -50 -786
rect -530 -823 -50 -820
rect -530 -843 -450 -823
rect -130 -843 -50 -823
rect -1030 -897 -950 -883
rect -1030 -949 -1016 -897
rect -964 -949 -950 -897
rect -1030 -963 -950 -949
rect -880 -906 -800 -883
rect -880 -940 -857 -906
rect -823 -940 -800 -906
rect -1010 -1135 -970 -963
rect -880 -986 -800 -940
rect -880 -1020 -857 -986
rect -823 -1020 -800 -986
rect -880 -1066 -800 -1020
rect -880 -1100 -857 -1066
rect -823 -1100 -800 -1066
rect -1030 -1148 -950 -1135
rect -1030 -1200 -1016 -1148
rect -964 -1200 -950 -1148
rect -1030 -1215 -950 -1200
rect -880 -1253 -800 -1100
rect -580 -906 -500 -883
rect -580 -940 -557 -906
rect -523 -940 -500 -906
rect -580 -986 -500 -940
rect -580 -1020 -557 -986
rect -523 -1020 -500 -986
rect -580 -1066 -500 -1020
rect -580 -1100 -557 -1066
rect -523 -1100 -500 -1066
rect -580 -1253 -500 -1100
rect -280 -906 -200 -883
rect -280 -940 -257 -906
rect -223 -940 -200 -906
rect -280 -986 -200 -940
rect -130 -897 -50 -883
rect -130 -949 -116 -897
rect -64 -949 -50 -897
rect -130 -963 -50 -949
rect -280 -1020 -257 -986
rect -223 -1020 -200 -986
rect -280 -1066 -200 -1020
rect -280 -1100 -257 -1066
rect -223 -1100 -200 -1066
rect -280 -1253 -200 -1100
rect 50 -1253 130 -540
rect 670 -346 750 -323
rect 670 -380 693 -346
rect 727 -380 750 -346
rect 670 -426 750 -380
rect 670 -460 693 -426
rect 727 -460 750 -426
rect 670 -506 750 -460
rect 670 -540 693 -506
rect 727 -540 750 -506
rect 670 -573 750 -540
rect 1000 -346 1080 -323
rect 1000 -380 1023 -346
rect 1057 -380 1080 -346
rect 1000 -426 1080 -380
rect 1000 -460 1023 -426
rect 1057 -460 1080 -426
rect 1000 -506 1080 -460
rect 1000 -540 1023 -506
rect 1057 -540 1080 -506
rect 1000 -573 1080 -540
rect 1300 -346 1380 -323
rect 1300 -380 1323 -346
rect 1357 -380 1380 -346
rect 1300 -426 1380 -380
rect 1300 -460 1323 -426
rect 1357 -460 1380 -426
rect 1300 -506 1380 -460
rect 1300 -540 1323 -506
rect 1357 -540 1380 -506
rect 1300 -573 1380 -540
rect 1600 -346 1680 -323
rect 1600 -380 1623 -346
rect 1657 -380 1680 -346
rect 1600 -426 1680 -380
rect 1600 -460 1623 -426
rect 1657 -460 1680 -426
rect 1600 -506 1680 -460
rect 1600 -540 1623 -506
rect 1657 -540 1680 -506
rect 1600 -573 1680 -540
rect 2080 -337 2160 -323
rect 2080 -389 2094 -337
rect 2146 -389 2160 -337
rect 2080 -426 2160 -389
rect 2080 -460 2103 -426
rect 2137 -460 2160 -426
rect 2080 -506 2160 -460
rect 2080 -540 2103 -506
rect 2137 -540 2160 -506
rect 2080 -573 2160 -540
rect 158 -613 238 -593
rect 158 -616 480 -613
rect 158 -650 181 -616
rect 215 -650 480 -616
rect 158 -653 480 -650
rect 158 -673 238 -653
rect 440 -913 480 -653
rect 158 -935 238 -921
rect 158 -987 172 -935
rect 224 -987 238 -935
rect 158 -1001 238 -987
rect 420 -936 500 -913
rect 420 -970 443 -936
rect 477 -970 500 -936
rect 420 -993 500 -970
rect 158 -1043 238 -1029
rect 158 -1095 172 -1043
rect 224 -1048 238 -1043
rect 420 -1048 500 -1034
rect 224 -1057 500 -1048
rect 224 -1088 443 -1057
rect 224 -1095 238 -1088
rect 158 -1109 238 -1095
rect 420 -1091 443 -1088
rect 477 -1091 500 -1057
rect 420 -1114 500 -1091
rect 690 -1253 730 -573
rect 1350 -783 1430 -763
rect 1750 -783 1830 -763
rect 1350 -786 1830 -783
rect 1350 -820 1373 -786
rect 1407 -820 1773 -786
rect 1807 -820 1830 -786
rect 1350 -823 1830 -820
rect 1350 -843 1430 -823
rect 1750 -843 1830 -823
rect 1000 -906 1080 -883
rect 850 -927 930 -913
rect 850 -979 864 -927
rect 916 -979 930 -927
rect 850 -993 930 -979
rect 1000 -940 1023 -906
rect 1057 -940 1080 -906
rect 1000 -986 1080 -940
rect 1000 -1020 1023 -986
rect 1057 -1020 1080 -986
rect 850 -1047 930 -1033
rect 850 -1099 864 -1047
rect 916 -1099 930 -1047
rect 850 -1113 930 -1099
rect 1000 -1066 1080 -1020
rect 1000 -1100 1023 -1066
rect 1057 -1100 1080 -1066
rect 1000 -1253 1080 -1100
rect 1300 -906 1380 -883
rect 1300 -940 1323 -906
rect 1357 -940 1380 -906
rect 1300 -986 1380 -940
rect 1300 -1020 1323 -986
rect 1357 -1020 1380 -986
rect 1300 -1066 1380 -1020
rect 1300 -1100 1323 -1066
rect 1357 -1100 1380 -1066
rect 1300 -1253 1380 -1100
rect 1600 -906 1680 -883
rect 1600 -940 1623 -906
rect 1657 -940 1680 -906
rect 1600 -986 1680 -940
rect 1600 -1020 1623 -986
rect 1657 -1020 1680 -986
rect 1830 -927 1910 -913
rect 1830 -979 1844 -927
rect 1896 -979 1910 -927
rect 1830 -993 1910 -979
rect 1600 -1066 1680 -1020
rect 1600 -1100 1623 -1066
rect 1657 -1100 1680 -1066
rect 1600 -1253 1680 -1100
rect 1980 -1047 2060 -1033
rect 1980 -1099 1994 -1047
rect 2046 -1099 2060 -1047
rect 1980 -1113 2060 -1099
rect 2100 -1253 2140 -573
rect 2183 -657 2263 -643
rect 2183 -709 2197 -657
rect 2249 -709 2263 -657
rect 2183 -723 2263 -709
rect -3870 -1277 150 -1253
rect -3870 -1329 -3821 -1277
rect -3769 -1286 150 -1277
rect -3753 -1320 -3707 -1286
rect -3673 -1320 -3627 -1286
rect -3593 -1320 -3547 -1286
rect -3513 -1320 -3467 -1286
rect -3433 -1320 -3387 -1286
rect -3353 -1320 -3307 -1286
rect -3273 -1320 -3227 -1286
rect -3193 -1320 -3147 -1286
rect -3113 -1320 -3067 -1286
rect -3033 -1320 -2987 -1286
rect -2953 -1320 -2907 -1286
rect -2873 -1320 -2827 -1286
rect -2793 -1320 -2747 -1286
rect -2713 -1320 -2667 -1286
rect -2633 -1320 -2587 -1286
rect -2553 -1320 -2507 -1286
rect -2473 -1320 -2427 -1286
rect -2393 -1320 -2347 -1286
rect -2313 -1320 -2267 -1286
rect -2233 -1320 -2187 -1286
rect -2153 -1320 -2107 -1286
rect -2073 -1320 -2027 -1286
rect -1993 -1320 -1947 -1286
rect -1913 -1320 -1867 -1286
rect -1833 -1320 -1787 -1286
rect -1753 -1320 -1707 -1286
rect -1673 -1320 -1197 -1286
rect -1163 -1320 -1117 -1286
rect -1083 -1320 -1037 -1286
rect -1003 -1320 -957 -1286
rect -923 -1320 -877 -1286
rect -843 -1320 -797 -1286
rect -763 -1320 -717 -1286
rect -683 -1320 -637 -1286
rect -603 -1320 -557 -1286
rect -523 -1320 -477 -1286
rect -443 -1320 -397 -1286
rect -363 -1320 -317 -1286
rect -283 -1320 -237 -1286
rect -203 -1320 -157 -1286
rect -123 -1320 -77 -1286
rect -43 -1320 3 -1286
rect 37 -1320 83 -1286
rect 117 -1320 150 -1286
rect -3769 -1329 150 -1320
rect -3870 -1353 150 -1329
rect 280 -1286 2180 -1253
rect 280 -1320 523 -1286
rect 557 -1320 603 -1286
rect 637 -1320 683 -1286
rect 717 -1320 763 -1286
rect 797 -1320 843 -1286
rect 877 -1320 923 -1286
rect 957 -1320 1003 -1286
rect 1037 -1320 1083 -1286
rect 1117 -1320 1163 -1286
rect 1197 -1320 1243 -1286
rect 1277 -1320 1323 -1286
rect 1357 -1320 1403 -1286
rect 1437 -1320 1483 -1286
rect 1517 -1320 1563 -1286
rect 1597 -1320 1643 -1286
rect 1677 -1320 1723 -1286
rect 1757 -1320 1803 -1286
rect 1837 -1320 1883 -1286
rect 1917 -1320 1963 -1286
rect 1997 -1320 2043 -1286
rect 2077 -1320 2123 -1286
rect 2157 -1320 2180 -1286
rect 280 -1353 2180 -1320
rect 280 -1483 380 -1353
rect -89 -1583 380 -1483
rect 508 -1511 588 -1497
rect 508 -1563 522 -1511
rect 574 -1563 588 -1511
rect 508 -1577 588 -1563
rect 2453 -1544 2533 -1530
rect -89 -1713 11 -1583
rect 2453 -1596 2467 -1544
rect 2519 -1596 2533 -1544
rect 2453 -1610 2533 -1596
rect -3835 -1738 -1729 -1713
rect -3835 -1790 -3821 -1738
rect -3769 -1746 -1729 -1738
rect -3769 -1780 -3706 -1746
rect -3672 -1780 -3626 -1746
rect -3592 -1780 -3546 -1746
rect -3512 -1780 -3466 -1746
rect -3432 -1780 -3386 -1746
rect -3352 -1780 -3306 -1746
rect -3272 -1780 -3226 -1746
rect -3192 -1780 -3146 -1746
rect -3112 -1780 -3066 -1746
rect -3032 -1780 -2986 -1746
rect -2952 -1780 -2906 -1746
rect -2872 -1780 -2826 -1746
rect -2792 -1780 -2746 -1746
rect -2712 -1780 -2666 -1746
rect -2632 -1780 -2586 -1746
rect -2552 -1780 -2506 -1746
rect -2472 -1780 -2426 -1746
rect -2392 -1780 -2346 -1746
rect -2312 -1780 -2266 -1746
rect -2232 -1780 -2186 -1746
rect -2152 -1780 -2106 -1746
rect -2072 -1780 -2026 -1746
rect -1992 -1780 -1946 -1746
rect -1912 -1780 -1866 -1746
rect -1832 -1780 -1786 -1746
rect -1752 -1780 -1729 -1746
rect -3769 -1790 -1729 -1780
rect -3835 -1813 -1729 -1790
rect -1369 -1746 11 -1713
rect -1369 -1780 -1336 -1746
rect -1302 -1780 -1256 -1746
rect -1222 -1780 -1176 -1746
rect -1142 -1780 -1096 -1746
rect -1062 -1780 -1016 -1746
rect -982 -1780 -936 -1746
rect -902 -1780 -856 -1746
rect -822 -1780 -776 -1746
rect -742 -1780 -696 -1746
rect -662 -1780 -616 -1746
rect -582 -1780 -536 -1746
rect -502 -1780 -456 -1746
rect -422 -1780 -376 -1746
rect -342 -1780 -296 -1746
rect -262 -1780 -216 -1746
rect -182 -1780 -136 -1746
rect -102 -1780 -56 -1746
rect -22 -1780 11 -1746
rect -1369 -1813 11 -1780
rect 361 -1738 2361 -1714
rect 361 -1790 375 -1738
rect 427 -1747 2361 -1738
rect 427 -1781 464 -1747
rect 498 -1781 544 -1747
rect 578 -1781 624 -1747
rect 658 -1781 704 -1747
rect 738 -1781 784 -1747
rect 818 -1781 864 -1747
rect 898 -1781 944 -1747
rect 978 -1781 1024 -1747
rect 1058 -1781 1104 -1747
rect 1138 -1781 1184 -1747
rect 1218 -1781 1264 -1747
rect 1298 -1781 1344 -1747
rect 1378 -1781 1424 -1747
rect 1458 -1781 1504 -1747
rect 1538 -1781 1584 -1747
rect 1618 -1781 1664 -1747
rect 1698 -1781 1744 -1747
rect 1778 -1781 1824 -1747
rect 1858 -1781 1904 -1747
rect 1938 -1781 1984 -1747
rect 2018 -1781 2064 -1747
rect 2098 -1781 2144 -1747
rect 2178 -1781 2224 -1747
rect 2258 -1781 2304 -1747
rect 2338 -1781 2361 -1747
rect 427 -1790 2361 -1781
rect -3679 -2493 -3639 -1813
rect -3379 -2493 -3339 -1813
rect -3309 -1857 -3229 -1843
rect -3309 -1909 -3295 -1857
rect -3243 -1909 -3229 -1857
rect -3309 -1923 -3229 -1909
rect -3219 -1977 -3139 -1963
rect -3219 -2029 -3205 -1977
rect -3153 -2029 -3139 -1977
rect -3219 -2043 -3139 -2029
rect -3069 -1966 -2989 -1813
rect -3069 -2000 -3046 -1966
rect -3012 -2000 -2989 -1966
rect -3069 -2046 -2989 -2000
rect -3069 -2080 -3046 -2046
rect -3012 -2080 -2989 -2046
rect -3249 -2097 -3169 -2083
rect -3249 -2149 -3235 -2097
rect -3183 -2149 -3169 -2097
rect -3249 -2163 -3169 -2149
rect -3069 -2126 -2989 -2080
rect -3069 -2160 -3046 -2126
rect -3012 -2160 -2989 -2126
rect -3069 -2183 -2989 -2160
rect -2769 -1966 -2689 -1813
rect -2769 -2000 -2746 -1966
rect -2712 -2000 -2689 -1966
rect -2769 -2046 -2689 -2000
rect -2769 -2080 -2746 -2046
rect -2712 -2080 -2689 -2046
rect -2769 -2126 -2689 -2080
rect -2769 -2160 -2746 -2126
rect -2712 -2160 -2689 -2126
rect -2769 -2183 -2689 -2160
rect -2469 -1966 -2389 -1813
rect -1939 -1857 -1859 -1843
rect -1939 -1909 -1925 -1857
rect -1873 -1909 -1859 -1857
rect -1939 -1923 -1859 -1909
rect -2469 -2000 -2446 -1966
rect -2412 -2000 -2389 -1966
rect -2469 -2046 -2389 -2000
rect -2089 -1977 -2009 -1963
rect -2089 -2029 -2075 -1977
rect -2023 -2029 -2009 -1977
rect -2089 -2043 -2009 -2029
rect -2469 -2080 -2446 -2046
rect -2412 -2080 -2389 -2046
rect -2469 -2126 -2389 -2080
rect -2469 -2160 -2446 -2126
rect -2412 -2160 -2389 -2126
rect -2469 -2183 -2389 -2160
rect -2219 -2097 -2139 -2083
rect -2219 -2149 -2205 -2097
rect -2153 -2149 -2139 -2097
rect -2219 -2163 -2139 -2149
rect -2719 -2243 -2639 -2223
rect -2319 -2243 -2239 -2223
rect -2719 -2246 -2239 -2243
rect -2719 -2280 -2696 -2246
rect -2662 -2280 -2296 -2246
rect -2262 -2280 -2239 -2246
rect -2719 -2283 -2239 -2280
rect -2719 -2303 -2639 -2283
rect -2319 -2303 -2239 -2283
rect -1819 -2493 -1779 -1813
rect -1457 -2123 -1377 -2103
rect -1718 -2126 -1377 -2123
rect -1718 -2160 -1434 -2126
rect -1400 -2160 -1377 -2126
rect -1718 -2163 -1377 -2160
rect -1718 -2342 -1678 -2163
rect -1457 -2183 -1377 -2163
rect -1739 -2365 -1659 -2342
rect -1739 -2399 -1716 -2365
rect -1682 -2399 -1659 -2365
rect -1739 -2422 -1659 -2399
rect -3699 -2526 -3619 -2493
rect -3699 -2560 -3676 -2526
rect -3642 -2560 -3619 -2526
rect -3699 -2606 -3619 -2560
rect -3699 -2640 -3676 -2606
rect -3642 -2640 -3619 -2606
rect -3699 -2686 -3619 -2640
rect -3699 -2720 -3676 -2686
rect -3642 -2720 -3619 -2686
rect -3699 -2743 -3619 -2720
rect -3399 -2526 -3319 -2493
rect -3399 -2560 -3376 -2526
rect -3342 -2560 -3319 -2526
rect -3399 -2606 -3319 -2560
rect -3399 -2640 -3376 -2606
rect -3342 -2640 -3319 -2606
rect -3399 -2686 -3319 -2640
rect -3399 -2720 -3376 -2686
rect -3342 -2720 -3319 -2686
rect -3399 -2743 -3319 -2720
rect -3069 -2526 -2989 -2493
rect -3069 -2560 -3046 -2526
rect -3012 -2560 -2989 -2526
rect -3069 -2606 -2989 -2560
rect -3069 -2640 -3046 -2606
rect -3012 -2640 -2989 -2606
rect -3069 -2686 -2989 -2640
rect -3069 -2720 -3046 -2686
rect -3012 -2720 -2989 -2686
rect -3069 -2743 -2989 -2720
rect -2769 -2526 -2689 -2493
rect -2769 -2560 -2746 -2526
rect -2712 -2560 -2689 -2526
rect -2769 -2606 -2689 -2560
rect -2769 -2640 -2746 -2606
rect -2712 -2640 -2689 -2606
rect -2769 -2686 -2689 -2640
rect -2769 -2720 -2746 -2686
rect -2712 -2720 -2689 -2686
rect -2769 -2743 -2689 -2720
rect -2469 -2526 -2389 -2493
rect -2469 -2560 -2446 -2526
rect -2412 -2560 -2389 -2526
rect -2469 -2606 -2389 -2560
rect -2469 -2640 -2446 -2606
rect -2412 -2640 -2389 -2606
rect -2469 -2686 -2389 -2640
rect -2469 -2720 -2446 -2686
rect -2412 -2720 -2389 -2686
rect -2469 -2743 -2389 -2720
rect -1839 -2526 -1759 -2493
rect -1839 -2560 -1816 -2526
rect -1782 -2560 -1759 -2526
rect -1839 -2606 -1759 -2560
rect -1839 -2640 -1816 -2606
rect -1782 -2640 -1759 -2606
rect -1839 -2686 -1759 -2640
rect -1839 -2720 -1816 -2686
rect -1782 -2720 -1759 -2686
rect -1839 -2743 -1759 -2720
rect -1349 -2526 -1269 -1813
rect -1019 -1966 -939 -1813
rect -1019 -2000 -996 -1966
rect -962 -2000 -939 -1966
rect -1019 -2046 -939 -2000
rect -1019 -2080 -996 -2046
rect -962 -2080 -939 -2046
rect -1169 -2117 -1089 -2103
rect -1169 -2169 -1155 -2117
rect -1103 -2169 -1089 -2117
rect -1169 -2183 -1089 -2169
rect -1019 -2126 -939 -2080
rect -1019 -2160 -996 -2126
rect -962 -2160 -939 -2126
rect -1019 -2183 -939 -2160
rect -719 -1966 -639 -1813
rect -719 -2000 -696 -1966
rect -662 -2000 -639 -1966
rect -719 -2046 -639 -2000
rect -719 -2080 -696 -2046
rect -662 -2080 -639 -2046
rect -719 -2126 -639 -2080
rect -719 -2160 -696 -2126
rect -662 -2160 -639 -2126
rect -719 -2183 -639 -2160
rect -419 -1966 -339 -1813
rect -419 -2000 -396 -1966
rect -362 -2000 -339 -1966
rect -419 -2046 -339 -2000
rect -419 -2080 -396 -2046
rect -362 -2080 -339 -2046
rect -419 -2126 -339 -2080
rect -419 -2160 -396 -2126
rect -362 -2160 -339 -2126
rect -419 -2183 -339 -2160
rect -269 -2117 -189 -2103
rect -269 -2169 -255 -2117
rect -203 -2169 -189 -2117
rect -269 -2183 -189 -2169
rect -669 -2243 -589 -2223
rect -269 -2243 -189 -2223
rect -669 -2246 -189 -2243
rect -669 -2280 -646 -2246
rect -612 -2280 -246 -2246
rect -212 -2280 -189 -2246
rect -669 -2283 -189 -2280
rect -669 -2303 -589 -2283
rect -269 -2303 -189 -2283
rect -1349 -2560 -1326 -2526
rect -1292 -2560 -1269 -2526
rect -1349 -2606 -1269 -2560
rect -1349 -2640 -1326 -2606
rect -1292 -2640 -1269 -2606
rect -1349 -2686 -1269 -2640
rect -1349 -2720 -1326 -2686
rect -1292 -2720 -1269 -2686
rect -1349 -2743 -1269 -2720
rect -1019 -2526 -939 -2493
rect -1019 -2560 -996 -2526
rect -962 -2560 -939 -2526
rect -1019 -2606 -939 -2560
rect -1019 -2640 -996 -2606
rect -962 -2640 -939 -2606
rect -1019 -2686 -939 -2640
rect -1019 -2720 -996 -2686
rect -962 -2720 -939 -2686
rect -1019 -2743 -939 -2720
rect -719 -2526 -639 -2493
rect -719 -2560 -696 -2526
rect -662 -2560 -639 -2526
rect -719 -2606 -639 -2560
rect -719 -2640 -696 -2606
rect -662 -2640 -639 -2606
rect -719 -2686 -639 -2640
rect -719 -2720 -696 -2686
rect -662 -2720 -639 -2686
rect -719 -2743 -639 -2720
rect -419 -2526 -339 -2493
rect -419 -2560 -396 -2526
rect -362 -2560 -339 -2526
rect -419 -2606 -339 -2560
rect -419 -2640 -396 -2606
rect -362 -2640 -339 -2606
rect -419 -2686 -339 -2640
rect -419 -2720 -396 -2686
rect -362 -2720 -339 -2686
rect -419 -2743 -339 -2720
rect -89 -2526 -9 -1813
rect 361 -1814 2361 -1790
rect 114 -1944 194 -1930
rect 114 -1996 128 -1944
rect 180 -1996 194 -1944
rect 114 -2010 194 -1996
rect 290 -2030 370 -2016
rect 290 -2038 304 -2030
rect 45 -2078 304 -2038
rect 45 -2393 85 -2078
rect 290 -2082 304 -2078
rect 356 -2082 370 -2030
rect 290 -2096 370 -2082
rect 290 -2140 370 -2126
rect 290 -2192 304 -2140
rect 356 -2192 370 -2140
rect 290 -2206 370 -2192
rect 291 -2254 371 -2240
rect 291 -2306 305 -2254
rect 357 -2306 371 -2254
rect 291 -2320 371 -2306
rect 291 -2368 371 -2354
rect 25 -2416 105 -2393
rect 25 -2450 48 -2416
rect 82 -2450 105 -2416
rect 291 -2420 305 -2368
rect 357 -2420 371 -2368
rect 291 -2434 371 -2420
rect 25 -2473 105 -2450
rect 411 -2494 451 -1814
rect 491 -1863 571 -1849
rect 491 -1915 505 -1863
rect 557 -1915 571 -1863
rect 491 -1929 571 -1915
rect 591 -1988 671 -1974
rect 591 -2040 605 -1988
rect 657 -2040 671 -1988
rect 591 -2054 671 -2040
rect 711 -2494 751 -1814
rect 1021 -1967 1101 -1814
rect 1021 -2001 1044 -1967
rect 1078 -2001 1101 -1967
rect 1021 -2047 1101 -2001
rect 791 -2078 871 -2064
rect 791 -2130 805 -2078
rect 857 -2130 871 -2078
rect 791 -2144 871 -2130
rect 1021 -2081 1044 -2047
rect 1078 -2081 1101 -2047
rect 1021 -2127 1101 -2081
rect 1021 -2161 1044 -2127
rect 1078 -2161 1101 -2127
rect 1021 -2184 1101 -2161
rect 1321 -1967 1401 -1814
rect 1321 -2001 1344 -1967
rect 1378 -2001 1401 -1967
rect 1321 -2047 1401 -2001
rect 1321 -2081 1344 -2047
rect 1378 -2081 1401 -2047
rect 1321 -2127 1401 -2081
rect 1321 -2161 1344 -2127
rect 1378 -2161 1401 -2127
rect 1321 -2184 1401 -2161
rect 1621 -1967 1701 -1814
rect 1771 -1868 1851 -1854
rect 1771 -1920 1785 -1868
rect 1837 -1920 1851 -1868
rect 1771 -1934 1851 -1920
rect 1621 -2001 1644 -1967
rect 1678 -2001 1701 -1967
rect 1621 -2047 1701 -2001
rect 1891 -1978 1971 -1964
rect 1891 -2030 1905 -1978
rect 1957 -2030 1971 -1978
rect 1891 -2044 1971 -2030
rect 2143 -1978 2223 -1964
rect 2143 -2030 2157 -1978
rect 2209 -2030 2223 -1978
rect 2143 -2044 2223 -2030
rect 1621 -2081 1644 -2047
rect 1678 -2081 1701 -2047
rect 1621 -2127 1701 -2081
rect 1621 -2161 1644 -2127
rect 1678 -2161 1701 -2127
rect 1771 -2078 1851 -2064
rect 1771 -2130 1785 -2078
rect 1837 -2130 1851 -2078
rect 1771 -2144 1851 -2130
rect 1621 -2184 1701 -2161
rect 1901 -2166 1981 -2152
rect 1901 -2218 1915 -2166
rect 1967 -2218 1981 -2166
rect 871 -2244 951 -2224
rect 1271 -2244 1351 -2224
rect 1901 -2232 1981 -2218
rect 871 -2247 1351 -2244
rect 871 -2281 894 -2247
rect 928 -2281 1294 -2247
rect 1328 -2281 1351 -2247
rect 871 -2284 1351 -2281
rect 871 -2304 951 -2284
rect 1271 -2304 1351 -2284
rect 1921 -2354 1961 -2232
rect 1901 -2377 1981 -2354
rect 1901 -2411 1924 -2377
rect 1958 -2411 1981 -2377
rect 1901 -2434 1981 -2411
rect 2271 -2494 2311 -1814
rect 2339 -1868 2419 -1854
rect 2339 -1920 2353 -1868
rect 2405 -1920 2419 -1868
rect 2339 -1934 2419 -1920
rect 2385 -2166 2465 -2152
rect 2385 -2218 2399 -2166
rect 2451 -2218 2465 -2166
rect 2385 -2232 2465 -2218
rect -89 -2560 -66 -2526
rect -32 -2560 -9 -2526
rect -89 -2606 -9 -2560
rect 108 -2521 188 -2507
rect 108 -2573 122 -2521
rect 174 -2573 188 -2521
rect 108 -2587 188 -2573
rect 391 -2527 471 -2494
rect 391 -2561 414 -2527
rect 448 -2561 471 -2527
rect -89 -2640 -66 -2606
rect -32 -2640 -9 -2606
rect -89 -2686 -9 -2640
rect -89 -2720 -66 -2686
rect -32 -2720 -9 -2686
rect -89 -2743 -9 -2720
rect 391 -2607 471 -2561
rect 391 -2641 414 -2607
rect 448 -2641 471 -2607
rect 391 -2687 471 -2641
rect 391 -2721 414 -2687
rect 448 -2721 471 -2687
rect -3719 -2797 -3639 -2783
rect -3719 -2849 -3705 -2797
rect -3653 -2849 -3639 -2797
rect -3719 -2863 -3639 -2849
rect -3049 -2893 -3009 -2743
rect -2749 -2893 -2709 -2743
rect -2449 -2893 -2409 -2743
rect -999 -2893 -959 -2743
rect -699 -2893 -659 -2743
rect -399 -2893 -359 -2743
rect 391 -2744 471 -2721
rect 691 -2527 771 -2494
rect 691 -2561 714 -2527
rect 748 -2561 771 -2527
rect 691 -2607 771 -2561
rect 691 -2641 714 -2607
rect 748 -2641 771 -2607
rect 691 -2687 771 -2641
rect 691 -2721 714 -2687
rect 748 -2721 771 -2687
rect 691 -2744 771 -2721
rect 1021 -2527 1101 -2494
rect 1021 -2561 1044 -2527
rect 1078 -2561 1101 -2527
rect 1021 -2607 1101 -2561
rect 1021 -2641 1044 -2607
rect 1078 -2641 1101 -2607
rect 1021 -2687 1101 -2641
rect 1021 -2721 1044 -2687
rect 1078 -2721 1101 -2687
rect 1021 -2744 1101 -2721
rect 1321 -2527 1401 -2494
rect 1321 -2561 1344 -2527
rect 1378 -2561 1401 -2527
rect 1321 -2607 1401 -2561
rect 1321 -2641 1344 -2607
rect 1378 -2641 1401 -2607
rect 1321 -2687 1401 -2641
rect 1321 -2721 1344 -2687
rect 1378 -2721 1401 -2687
rect 1321 -2744 1401 -2721
rect 1621 -2527 1701 -2494
rect 1621 -2561 1644 -2527
rect 1678 -2561 1701 -2527
rect 1621 -2607 1701 -2561
rect 1621 -2641 1644 -2607
rect 1678 -2641 1701 -2607
rect 1621 -2687 1701 -2641
rect 1621 -2721 1644 -2687
rect 1678 -2721 1701 -2687
rect 1621 -2744 1701 -2721
rect 2251 -2527 2331 -2494
rect 2251 -2561 2274 -2527
rect 2308 -2561 2331 -2527
rect 2251 -2607 2331 -2561
rect 2251 -2641 2274 -2607
rect 2308 -2641 2331 -2607
rect 2251 -2687 2331 -2641
rect 2251 -2721 2274 -2687
rect 2308 -2721 2331 -2687
rect 2251 -2744 2331 -2721
rect 202 -2799 282 -2785
rect 202 -2851 216 -2799
rect 268 -2851 282 -2799
rect 202 -2865 282 -2851
rect -3978 -2960 -3955 -2926
rect -3921 -2960 -3898 -2926
rect -3978 -2983 -3898 -2960
rect -3729 -2894 361 -2893
rect 1041 -2894 1081 -2744
rect 1341 -2894 1381 -2744
rect 1641 -2894 1681 -2744
rect -3729 -2926 2361 -2894
rect -3729 -2960 -3706 -2926
rect -3672 -2960 -3626 -2926
rect -3592 -2960 -3546 -2926
rect -3512 -2960 -3466 -2926
rect -3432 -2960 -3386 -2926
rect -3352 -2960 -3306 -2926
rect -3272 -2960 -3226 -2926
rect -3192 -2960 -3146 -2926
rect -3112 -2960 -3066 -2926
rect -3032 -2960 -2986 -2926
rect -2952 -2960 -2906 -2926
rect -2872 -2960 -2826 -2926
rect -2792 -2960 -2746 -2926
rect -2712 -2960 -2666 -2926
rect -2632 -2960 -2586 -2926
rect -2552 -2960 -2506 -2926
rect -2472 -2960 -2426 -2926
rect -2392 -2960 -2346 -2926
rect -2312 -2960 -2266 -2926
rect -2232 -2960 -2186 -2926
rect -2152 -2960 -2106 -2926
rect -2072 -2960 -2026 -2926
rect -1992 -2960 -1946 -2926
rect -1912 -2960 -1866 -2926
rect -1832 -2960 -1786 -2926
rect -1752 -2960 -1336 -2926
rect -1302 -2960 -1256 -2926
rect -1222 -2960 -1176 -2926
rect -1142 -2960 -1096 -2926
rect -1062 -2960 -1016 -2926
rect -982 -2960 -936 -2926
rect -902 -2960 -856 -2926
rect -822 -2960 -776 -2926
rect -742 -2960 -696 -2926
rect -662 -2960 -616 -2926
rect -582 -2960 -536 -2926
rect -502 -2960 -456 -2926
rect -422 -2960 -376 -2926
rect -342 -2960 -296 -2926
rect -262 -2960 -216 -2926
rect -182 -2960 -136 -2926
rect -102 -2960 -56 -2926
rect -22 -2927 2361 -2926
rect -22 -2960 384 -2927
rect -3729 -2961 384 -2960
rect 418 -2961 464 -2927
rect 498 -2961 544 -2927
rect 578 -2961 624 -2927
rect 658 -2961 704 -2927
rect 738 -2961 784 -2927
rect 818 -2961 864 -2927
rect 898 -2961 944 -2927
rect 978 -2961 1024 -2927
rect 1058 -2961 1104 -2927
rect 1138 -2961 1184 -2927
rect 1218 -2961 1264 -2927
rect 1298 -2961 1344 -2927
rect 1378 -2961 1424 -2927
rect 1458 -2961 1504 -2927
rect 1538 -2961 1584 -2927
rect 1618 -2961 1664 -2927
rect 1698 -2961 1744 -2927
rect 1778 -2961 1824 -2927
rect 1858 -2961 1904 -2927
rect 1938 -2961 1984 -2927
rect 2018 -2961 2064 -2927
rect 2098 -2961 2144 -2927
rect 2178 -2961 2224 -2927
rect 2258 -2961 2304 -2927
rect 2338 -2961 2361 -2927
rect -3729 -2993 2361 -2961
rect 361 -2994 2361 -2993
<< via1 >>
rect -3820 1074 -3768 1083
rect -3820 1040 -3787 1074
rect -3787 1040 -3768 1074
rect -3820 1031 -3768 1040
rect 2114 1074 2166 1083
rect 2114 1040 2123 1074
rect 2123 1040 2157 1074
rect 2157 1040 2166 1074
rect 2114 1031 2166 1040
rect -4648 -1200 -4596 -1148
rect -4534 -493 -4482 -441
rect -4192 203 -4140 255
rect -4078 903 -4026 955
rect -3336 944 -3284 953
rect -3336 910 -3327 944
rect -3327 910 -3293 944
rect -3293 910 -3284 944
rect -3336 901 -3284 910
rect -3206 844 -3154 853
rect -3206 810 -3197 844
rect -3197 810 -3163 844
rect -3163 810 -3154 844
rect -3206 801 -3154 810
rect -3336 744 -3284 753
rect -3336 710 -3327 744
rect -3327 710 -3293 744
rect -3293 710 -3284 744
rect -3336 701 -3284 710
rect -3206 644 -3154 653
rect -3206 610 -3197 644
rect -3197 610 -3163 644
rect -3163 610 -3154 644
rect -3206 601 -3154 610
rect -2076 944 -2024 953
rect -2076 910 -2067 944
rect -2067 910 -2033 944
rect -2033 910 -2024 944
rect -2076 901 -2024 910
rect -2176 644 -2124 653
rect -2176 610 -2167 644
rect -2167 610 -2133 644
rect -2133 610 -2124 644
rect -2176 601 -2124 610
rect -1876 844 -1824 853
rect -1876 810 -1867 844
rect -1867 810 -1833 844
rect -1833 810 -1824 844
rect -1876 801 -1824 810
rect -1304 878 -1252 887
rect -1304 844 -1295 878
rect -1295 844 -1261 878
rect -1261 844 -1252 878
rect -1304 835 -1252 844
rect -1726 744 -1674 753
rect -1726 710 -1717 744
rect -1717 710 -1683 744
rect -1683 710 -1674 744
rect -1726 701 -1674 710
rect -1304 724 -1252 776
rect -1016 904 -964 956
rect -1016 694 -964 703
rect -1016 660 -1007 694
rect -1007 660 -973 694
rect -973 660 -964 694
rect -1016 651 -964 660
rect -116 694 -64 703
rect -116 660 -107 694
rect -107 660 -73 694
rect -73 660 -64 694
rect -116 651 -64 660
rect -1562 246 -1510 255
rect -1562 212 -1553 246
rect -1553 212 -1519 246
rect -1519 212 -1510 246
rect -1562 203 -1510 212
rect 172 814 224 866
rect 172 705 224 757
rect 864 844 916 853
rect 864 810 873 844
rect 873 810 907 844
rect 907 810 916 844
rect 864 801 916 810
rect 864 724 916 733
rect 864 690 873 724
rect 873 690 907 724
rect 907 690 916 724
rect 864 681 916 690
rect 1994 844 2046 853
rect 1994 810 2003 844
rect 2003 810 2037 844
rect 2037 810 2046 844
rect 1994 801 2046 810
rect 1844 724 1896 733
rect 1844 690 1853 724
rect 1853 690 1887 724
rect 1887 690 1896 724
rect 1844 681 1896 690
rect 2197 454 2249 463
rect 2197 420 2206 454
rect 2206 420 2240 454
rect 2240 420 2249 454
rect 2197 411 2249 420
rect 2094 134 2146 143
rect 2094 100 2103 134
rect 2103 100 2137 134
rect 2137 100 2146 134
rect 2094 91 2146 100
rect -3705 14 -3653 23
rect -3705 -20 -3696 14
rect -3696 -20 -3662 14
rect -3662 -20 -3653 14
rect -3705 -29 -3653 -20
rect 522 14 574 23
rect 522 -20 531 14
rect 531 -20 565 14
rect 565 -20 574 14
rect 522 -29 574 -20
rect -3705 -226 -3653 -217
rect -3705 -260 -3696 -226
rect -3696 -260 -3662 -226
rect -3662 -260 -3653 -226
rect -3705 -269 -3653 -260
rect 522 -225 574 -216
rect 522 -259 531 -225
rect 531 -259 565 -225
rect 565 -259 574 -225
rect 522 -268 574 -259
rect -1562 -449 -1510 -440
rect -1562 -483 -1553 -449
rect -1553 -483 -1519 -449
rect -1519 -483 -1510 -449
rect -1562 -492 -1510 -483
rect -3206 -856 -3154 -847
rect -3206 -890 -3197 -856
rect -3197 -890 -3163 -856
rect -3163 -890 -3154 -856
rect -3206 -899 -3154 -890
rect -3336 -956 -3284 -947
rect -3336 -990 -3327 -956
rect -3327 -990 -3293 -956
rect -3293 -990 -3284 -956
rect -3336 -999 -3284 -990
rect -3206 -1056 -3154 -1047
rect -3206 -1090 -3197 -1056
rect -3197 -1090 -3163 -1056
rect -3163 -1090 -3154 -1056
rect -3206 -1099 -3154 -1090
rect -3336 -1156 -3284 -1147
rect -3336 -1190 -3327 -1156
rect -3327 -1190 -3293 -1156
rect -3293 -1190 -3284 -1156
rect -3336 -1199 -3284 -1190
rect -2176 -856 -2124 -847
rect -2176 -890 -2167 -856
rect -2167 -890 -2133 -856
rect -2133 -890 -2124 -856
rect -2176 -899 -2124 -890
rect -2076 -1156 -2024 -1147
rect -2076 -1190 -2067 -1156
rect -2067 -1190 -2033 -1156
rect -2033 -1190 -2024 -1156
rect -2076 -1199 -2024 -1190
rect -1726 -956 -1674 -947
rect -1726 -990 -1717 -956
rect -1717 -990 -1683 -956
rect -1683 -990 -1674 -956
rect -1726 -999 -1674 -990
rect -1304 -1020 -1252 -968
rect -1876 -1056 -1824 -1047
rect -1876 -1090 -1867 -1056
rect -1867 -1090 -1833 -1056
rect -1833 -1090 -1824 -1056
rect -1876 -1099 -1824 -1090
rect -1304 -1090 -1252 -1081
rect -1304 -1124 -1295 -1090
rect -1295 -1124 -1261 -1090
rect -1261 -1124 -1252 -1090
rect -1304 -1133 -1252 -1124
rect -1016 -906 -964 -897
rect -1016 -940 -1007 -906
rect -1007 -940 -973 -906
rect -973 -940 -964 -906
rect -1016 -949 -964 -940
rect -1016 -1200 -964 -1148
rect -116 -906 -64 -897
rect -116 -940 -107 -906
rect -107 -940 -73 -906
rect -73 -940 -64 -906
rect -116 -949 -64 -940
rect 2094 -346 2146 -337
rect 2094 -380 2103 -346
rect 2103 -380 2137 -346
rect 2137 -380 2146 -346
rect 2094 -389 2146 -380
rect 172 -944 224 -935
rect 172 -978 181 -944
rect 181 -978 215 -944
rect 215 -978 224 -944
rect 172 -987 224 -978
rect 172 -1095 224 -1043
rect 864 -936 916 -927
rect 864 -970 873 -936
rect 873 -970 907 -936
rect 907 -970 916 -936
rect 864 -979 916 -970
rect 864 -1056 916 -1047
rect 864 -1090 873 -1056
rect 873 -1090 907 -1056
rect 907 -1090 916 -1056
rect 864 -1099 916 -1090
rect 1844 -936 1896 -927
rect 1844 -970 1853 -936
rect 1853 -970 1887 -936
rect 1887 -970 1896 -936
rect 1844 -979 1896 -970
rect 1994 -1056 2046 -1047
rect 1994 -1090 2003 -1056
rect 2003 -1090 2037 -1056
rect 2037 -1090 2046 -1056
rect 1994 -1099 2046 -1090
rect 2197 -666 2249 -657
rect 2197 -700 2206 -666
rect 2206 -700 2240 -666
rect 2240 -700 2249 -666
rect 2197 -709 2249 -700
rect -3821 -1286 -3769 -1277
rect -3821 -1320 -3787 -1286
rect -3787 -1320 -3769 -1286
rect -3821 -1329 -3769 -1320
rect 522 -1520 574 -1511
rect 522 -1554 531 -1520
rect 531 -1554 565 -1520
rect 565 -1554 574 -1520
rect 522 -1563 574 -1554
rect 2467 -1553 2519 -1544
rect 2467 -1587 2476 -1553
rect 2476 -1587 2510 -1553
rect 2510 -1587 2519 -1553
rect 2467 -1596 2519 -1587
rect -3821 -1790 -3769 -1738
rect 375 -1747 427 -1738
rect 375 -1781 384 -1747
rect 384 -1781 418 -1747
rect 418 -1781 427 -1747
rect 375 -1790 427 -1781
rect -3295 -1866 -3243 -1857
rect -3295 -1900 -3286 -1866
rect -3286 -1900 -3252 -1866
rect -3252 -1900 -3243 -1866
rect -3295 -1909 -3243 -1900
rect -3205 -1986 -3153 -1977
rect -3205 -2020 -3196 -1986
rect -3196 -2020 -3162 -1986
rect -3162 -2020 -3153 -1986
rect -3205 -2029 -3153 -2020
rect -3235 -2106 -3183 -2097
rect -3235 -2140 -3226 -2106
rect -3226 -2140 -3192 -2106
rect -3192 -2140 -3183 -2106
rect -3235 -2149 -3183 -2140
rect -1925 -1866 -1873 -1857
rect -1925 -1900 -1916 -1866
rect -1916 -1900 -1882 -1866
rect -1882 -1900 -1873 -1866
rect -1925 -1909 -1873 -1900
rect -2075 -1986 -2023 -1977
rect -2075 -2020 -2066 -1986
rect -2066 -2020 -2032 -1986
rect -2032 -2020 -2023 -1986
rect -2075 -2029 -2023 -2020
rect -2205 -2106 -2153 -2097
rect -2205 -2140 -2196 -2106
rect -2196 -2140 -2162 -2106
rect -2162 -2140 -2153 -2106
rect -2205 -2149 -2153 -2140
rect -1155 -2126 -1103 -2117
rect -1155 -2160 -1146 -2126
rect -1146 -2160 -1112 -2126
rect -1112 -2160 -1103 -2126
rect -1155 -2169 -1103 -2160
rect -255 -2126 -203 -2117
rect -255 -2160 -246 -2126
rect -246 -2160 -212 -2126
rect -212 -2160 -203 -2126
rect -255 -2169 -203 -2160
rect 128 -1953 180 -1944
rect 128 -1987 137 -1953
rect 137 -1987 171 -1953
rect 171 -1987 180 -1953
rect 128 -1996 180 -1987
rect 304 -2082 356 -2030
rect 304 -2149 356 -2140
rect 304 -2183 313 -2149
rect 313 -2183 347 -2149
rect 347 -2183 356 -2149
rect 304 -2192 356 -2183
rect 305 -2263 357 -2254
rect 305 -2297 314 -2263
rect 314 -2297 348 -2263
rect 348 -2297 357 -2263
rect 305 -2306 357 -2297
rect 305 -2377 357 -2368
rect 305 -2411 314 -2377
rect 314 -2411 348 -2377
rect 348 -2411 357 -2377
rect 305 -2420 357 -2411
rect 505 -1872 557 -1863
rect 505 -1906 514 -1872
rect 514 -1906 548 -1872
rect 548 -1906 557 -1872
rect 505 -1915 557 -1906
rect 605 -1997 657 -1988
rect 605 -2031 614 -1997
rect 614 -2031 648 -1997
rect 648 -2031 657 -1997
rect 605 -2040 657 -2031
rect 805 -2087 857 -2078
rect 805 -2121 814 -2087
rect 814 -2121 848 -2087
rect 848 -2121 857 -2087
rect 805 -2130 857 -2121
rect 1785 -1877 1837 -1868
rect 1785 -1911 1794 -1877
rect 1794 -1911 1828 -1877
rect 1828 -1911 1837 -1877
rect 1785 -1920 1837 -1911
rect 1905 -1987 1957 -1978
rect 1905 -2021 1914 -1987
rect 1914 -2021 1948 -1987
rect 1948 -2021 1957 -1987
rect 1905 -2030 1957 -2021
rect 2157 -1987 2209 -1978
rect 2157 -2021 2166 -1987
rect 2166 -2021 2200 -1987
rect 2200 -2021 2209 -1987
rect 2157 -2030 2209 -2021
rect 1785 -2087 1837 -2078
rect 1785 -2121 1794 -2087
rect 1794 -2121 1828 -2087
rect 1828 -2121 1837 -2087
rect 1785 -2130 1837 -2121
rect 1915 -2218 1967 -2166
rect 2353 -1877 2405 -1868
rect 2353 -1911 2362 -1877
rect 2362 -1911 2396 -1877
rect 2396 -1911 2405 -1877
rect 2353 -1920 2405 -1911
rect 2399 -2175 2451 -2166
rect 2399 -2209 2408 -2175
rect 2408 -2209 2442 -2175
rect 2442 -2209 2451 -2175
rect 2399 -2218 2451 -2209
rect 122 -2530 174 -2521
rect 122 -2564 131 -2530
rect 131 -2564 165 -2530
rect 165 -2564 174 -2530
rect 122 -2573 174 -2564
rect -3705 -2806 -3653 -2797
rect -3705 -2840 -3696 -2806
rect -3696 -2840 -3662 -2806
rect -3662 -2840 -3653 -2806
rect -3705 -2849 -3653 -2840
rect 216 -2808 268 -2799
rect 216 -2842 225 -2808
rect 225 -2842 259 -2808
rect 259 -2842 268 -2808
rect 216 -2851 268 -2842
<< metal2 >>
rect -3835 1097 -3755 1200
rect -3835 1083 -3754 1097
rect -3835 1031 -3820 1083
rect -3768 1031 -3754 1083
rect -3835 1017 -3754 1031
rect -4092 957 -4012 968
rect -4092 901 -4080 957
rect -4024 901 -4012 957
rect -4092 888 -4012 901
rect -4206 257 -4126 268
rect -4206 201 -4194 257
rect -4138 201 -4126 257
rect -4206 188 -4126 201
rect -4548 -439 -4468 -428
rect -4548 -495 -4536 -439
rect -4480 -495 -4468 -439
rect -4548 -508 -4468 -495
rect -4662 -1146 -4582 -1135
rect -4662 -1202 -4650 -1146
rect -4594 -1202 -4582 -1146
rect -4662 -1215 -4582 -1202
rect -3835 -1277 -3755 1017
rect -3699 37 -3659 1200
rect -3350 953 -3270 967
rect -3350 901 -3336 953
rect -3284 947 -3270 953
rect -2090 953 -2010 967
rect -2090 947 -2076 953
rect -3284 907 -2076 947
rect -3284 901 -3270 907
rect -3350 887 -3270 901
rect -2090 901 -2076 907
rect -2024 901 -2010 953
rect -1030 958 -950 969
rect -1030 902 -1018 958
rect -962 902 -950 958
rect -2090 887 -2010 901
rect -1318 887 -1238 901
rect -1030 889 -950 902
rect -3220 853 -3140 867
rect -3220 801 -3206 853
rect -3154 847 -3140 853
rect -1890 853 -1810 867
rect -1890 847 -1876 853
rect -3154 807 -1876 847
rect -3154 801 -3140 807
rect -3220 787 -3140 801
rect -1890 801 -1876 807
rect -1824 801 -1810 853
rect -1318 835 -1304 887
rect -1252 861 -1238 887
rect 158 866 238 880
rect 158 861 172 866
rect -1252 835 172 861
rect -1318 821 172 835
rect -1890 787 -1810 801
rect 158 814 172 821
rect 224 814 238 866
rect 158 800 238 814
rect -1318 776 106 790
rect -3350 753 -3270 767
rect -3350 701 -3336 753
rect -3284 747 -3270 753
rect -1740 753 -1660 767
rect -1740 747 -1726 753
rect -3284 707 -1726 747
rect -3284 701 -3270 707
rect -3350 687 -3270 701
rect -1740 701 -1726 707
rect -1674 701 -1660 753
rect -1318 724 -1304 776
rect -1252 750 106 776
rect -1252 724 -1238 750
rect -1318 710 -1238 724
rect 66 749 106 750
rect 158 757 238 771
rect 158 749 172 757
rect -1740 687 -1660 701
rect -1030 703 -950 717
rect -3220 653 -3140 667
rect -3220 601 -3206 653
rect -3154 647 -3140 653
rect -2190 653 -2110 667
rect -2190 647 -2176 653
rect -3154 607 -2176 647
rect -3154 601 -3140 607
rect -3220 587 -3140 601
rect -2190 601 -2176 607
rect -2124 601 -2110 653
rect -1030 651 -1016 703
rect -964 697 -950 703
rect -130 703 -50 717
rect 66 709 172 749
rect -130 697 -116 703
rect -964 657 -116 697
rect -964 651 -950 657
rect -1030 637 -950 651
rect -130 651 -116 657
rect -64 651 -50 703
rect 158 705 172 709
rect 224 705 238 757
rect 158 691 238 705
rect -130 637 -50 651
rect -2190 587 -2110 601
rect -1576 257 -1496 268
rect -1576 201 -1564 257
rect -1508 201 -1496 257
rect -1576 188 -1496 201
rect -3719 23 -3639 37
rect -3719 -29 -3705 23
rect -3653 -29 -3639 23
rect -3719 -43 -3639 -29
rect -3699 -203 -3659 -43
rect -3719 -217 -3639 -203
rect -3719 -269 -3705 -217
rect -3653 -269 -3639 -217
rect -3719 -283 -3639 -269
rect -3835 -1329 -3821 -1277
rect -3769 -1329 -3755 -1277
rect -3835 -1738 -3755 -1329
rect -3835 -1790 -3821 -1738
rect -3769 -1790 -3755 -1738
rect -3835 -1804 -3755 -1790
rect -3699 -2783 -3659 -283
rect -1576 -438 -1496 -427
rect -1576 -494 -1564 -438
rect -1508 -494 -1496 -438
rect -1576 -507 -1496 -494
rect -3220 -847 -3140 -833
rect -3220 -899 -3206 -847
rect -3154 -853 -3140 -847
rect -2190 -847 -2110 -833
rect -2190 -853 -2176 -847
rect -3154 -893 -2176 -853
rect -3154 -899 -3140 -893
rect -3220 -913 -3140 -899
rect -2190 -899 -2176 -893
rect -2124 -899 -2110 -847
rect -2190 -913 -2110 -899
rect -1030 -897 -950 -883
rect -3350 -947 -3270 -933
rect -3350 -999 -3336 -947
rect -3284 -953 -3270 -947
rect -1740 -947 -1660 -933
rect -1740 -953 -1726 -947
rect -3284 -993 -1726 -953
rect -3284 -999 -3270 -993
rect -3350 -1013 -3270 -999
rect -1740 -999 -1726 -993
rect -1674 -999 -1660 -947
rect -1030 -949 -1016 -897
rect -964 -903 -950 -897
rect -130 -897 -50 -883
rect -130 -903 -116 -897
rect -964 -943 -116 -903
rect -964 -949 -950 -943
rect -1740 -1013 -1660 -999
rect -1318 -968 -1238 -954
rect -1030 -963 -950 -949
rect -130 -949 -116 -943
rect -64 -949 -50 -897
rect 158 -935 238 -921
rect 158 -941 172 -935
rect -130 -963 -50 -949
rect -1318 -1020 -1304 -968
rect -1252 -994 -1238 -968
rect 10 -981 172 -941
rect 10 -994 50 -981
rect -1252 -1020 50 -994
rect 158 -987 172 -981
rect 224 -987 238 -935
rect 158 -1001 238 -987
rect -3220 -1047 -3140 -1033
rect -3220 -1099 -3206 -1047
rect -3154 -1053 -3140 -1047
rect -1890 -1047 -1810 -1033
rect -1318 -1034 50 -1020
rect -1890 -1053 -1876 -1047
rect -3154 -1093 -1876 -1053
rect -3154 -1099 -3140 -1093
rect -3220 -1113 -3140 -1099
rect -1890 -1099 -1876 -1093
rect -1824 -1099 -1810 -1047
rect 158 -1043 238 -1029
rect 158 -1067 172 -1043
rect -1890 -1113 -1810 -1099
rect -1318 -1081 172 -1067
rect -1318 -1133 -1304 -1081
rect -1252 -1095 172 -1081
rect 224 -1095 238 -1043
rect -1252 -1107 238 -1095
rect -1252 -1133 -1238 -1107
rect 158 -1109 238 -1107
rect -3350 -1147 -3270 -1133
rect -3350 -1199 -3336 -1147
rect -3284 -1153 -3270 -1147
rect -2090 -1147 -2010 -1133
rect -1318 -1147 -1238 -1133
rect -1030 -1146 -950 -1135
rect -2090 -1153 -2076 -1147
rect -3284 -1193 -2076 -1153
rect -3284 -1199 -3270 -1193
rect -3350 -1213 -3270 -1199
rect -2090 -1199 -2076 -1193
rect -2024 -1199 -2010 -1147
rect -2090 -1213 -2010 -1199
rect -1030 -1202 -1018 -1146
rect -962 -1202 -950 -1146
rect 266 -1160 306 1200
rect -1030 -1215 -950 -1202
rect 222 -1200 306 -1160
rect -3309 -1857 -3229 -1843
rect -3309 -1909 -3295 -1857
rect -3243 -1863 -3229 -1857
rect -1939 -1857 -1859 -1843
rect -1939 -1863 -1925 -1857
rect -3243 -1903 -1925 -1863
rect -3243 -1909 -3229 -1903
rect -3309 -1923 -3229 -1909
rect -1939 -1909 -1925 -1903
rect -1873 -1909 -1859 -1857
rect -1939 -1923 -1859 -1909
rect 114 -1944 194 -1930
rect -3219 -1977 -3139 -1963
rect -3219 -2029 -3205 -1977
rect -3153 -1983 -3139 -1977
rect -2089 -1977 -2009 -1963
rect -2089 -1983 -2075 -1977
rect -3153 -2023 -2075 -1983
rect -3153 -2029 -3139 -2023
rect -3219 -2043 -3139 -2029
rect -2089 -2029 -2075 -2023
rect -2023 -2029 -2009 -1977
rect 114 -1996 128 -1944
rect 180 -1996 194 -1944
rect 114 -2010 194 -1996
rect -2089 -2043 -2009 -2029
rect -3249 -2097 -3169 -2083
rect -3249 -2149 -3235 -2097
rect -3183 -2103 -3169 -2097
rect -2219 -2097 -2139 -2083
rect -2219 -2103 -2205 -2097
rect -3183 -2143 -2205 -2103
rect -3183 -2149 -3169 -2143
rect -3249 -2163 -3169 -2149
rect -2219 -2149 -2205 -2143
rect -2153 -2149 -2139 -2097
rect -2219 -2163 -2139 -2149
rect -1169 -2117 -1089 -2103
rect -1169 -2169 -1155 -2117
rect -1103 -2123 -1089 -2117
rect -269 -2117 -189 -2103
rect -269 -2123 -255 -2117
rect -1103 -2163 -255 -2123
rect -1103 -2169 -1089 -2163
rect -1169 -2183 -1089 -2169
rect -269 -2169 -255 -2163
rect -203 -2169 -189 -2117
rect -269 -2183 -189 -2169
rect 133 -2507 173 -2010
rect 108 -2521 188 -2507
rect 108 -2573 122 -2521
rect 174 -2573 188 -2521
rect 108 -2587 188 -2573
rect -3719 -2797 -3639 -2783
rect 222 -2785 262 -1200
rect 381 -1724 421 1200
rect 528 37 568 1200
rect 2100 1083 2180 1200
rect 2100 1031 2114 1083
rect 2166 1031 2180 1083
rect 2100 1017 2180 1031
rect 850 853 930 867
rect 850 801 864 853
rect 916 847 930 853
rect 1980 853 2060 867
rect 1980 847 1994 853
rect 916 807 1994 847
rect 916 801 930 807
rect 850 787 930 801
rect 1980 801 1994 807
rect 2046 801 2060 853
rect 1980 787 2060 801
rect 850 733 930 747
rect 850 681 864 733
rect 916 727 930 733
rect 1830 733 1910 747
rect 1830 727 1844 733
rect 916 687 1844 727
rect 916 681 930 687
rect 850 667 930 681
rect 1830 681 1844 687
rect 1896 681 1910 733
rect 1830 667 1910 681
rect 2183 463 2263 477
rect 2183 411 2197 463
rect 2249 457 2263 463
rect 2249 417 2379 457
rect 2249 411 2263 417
rect 2183 397 2263 411
rect 2080 143 2160 157
rect 2080 91 2094 143
rect 2146 91 2160 143
rect 508 23 588 37
rect 508 -29 522 23
rect 574 -29 588 23
rect 508 -43 588 -29
rect 528 -202 568 -43
rect 508 -216 588 -202
rect 508 -268 522 -216
rect 574 -268 588 -216
rect 508 -282 588 -268
rect 528 -1497 568 -282
rect 2080 -337 2160 91
rect 2080 -389 2094 -337
rect 2146 -389 2160 -337
rect 2080 -403 2160 -389
rect 2183 -657 2263 -643
rect 2183 -709 2197 -657
rect 2249 -709 2263 -657
rect 2183 -723 2263 -709
rect 850 -927 930 -913
rect 850 -979 864 -927
rect 916 -933 930 -927
rect 1830 -927 1910 -913
rect 1830 -933 1844 -927
rect 916 -973 1844 -933
rect 916 -979 930 -973
rect 850 -993 930 -979
rect 1830 -979 1844 -973
rect 1896 -979 1910 -927
rect 1830 -993 1910 -979
rect 850 -1047 930 -1033
rect 850 -1099 864 -1047
rect 916 -1053 930 -1047
rect 1980 -1047 2060 -1033
rect 1980 -1053 1994 -1047
rect 916 -1093 1994 -1053
rect 916 -1099 930 -1093
rect 850 -1113 930 -1099
rect 1980 -1099 1994 -1093
rect 2046 -1099 2060 -1047
rect 1980 -1113 2060 -1099
rect 508 -1511 588 -1497
rect 508 -1563 522 -1511
rect 574 -1563 588 -1511
rect 508 -1577 588 -1563
rect 361 -1738 441 -1724
rect 361 -1790 375 -1738
rect 427 -1790 441 -1738
rect 361 -1804 441 -1790
rect 491 -1863 571 -1849
rect 491 -1915 505 -1863
rect 557 -1874 571 -1863
rect 1771 -1868 1851 -1854
rect 1771 -1874 1785 -1868
rect 557 -1914 1785 -1874
rect 557 -1915 571 -1914
rect 491 -1929 571 -1915
rect 1771 -1920 1785 -1914
rect 1837 -1920 1851 -1868
rect 1771 -1934 1851 -1920
rect 2183 -1964 2223 -723
rect 2339 -1854 2379 417
rect 2453 -1544 2533 -1530
rect 2453 -1596 2467 -1544
rect 2519 -1596 2533 -1544
rect 2453 -1610 2533 -1596
rect 2339 -1868 2419 -1854
rect 2339 -1920 2353 -1868
rect 2405 -1920 2419 -1868
rect 2339 -1934 2419 -1920
rect 591 -1984 671 -1974
rect 1891 -1978 1971 -1964
rect 1891 -1984 1905 -1978
rect 591 -1988 1905 -1984
rect 290 -2030 370 -2016
rect 290 -2082 304 -2030
rect 356 -2036 370 -2030
rect 356 -2076 463 -2036
rect 591 -2040 605 -1988
rect 657 -2024 1905 -1988
rect 657 -2040 671 -2024
rect 591 -2054 671 -2040
rect 1891 -2030 1905 -2024
rect 1957 -2030 1971 -1978
rect 1891 -2044 1971 -2030
rect 2143 -1978 2223 -1964
rect 2143 -2030 2157 -1978
rect 2209 -2030 2223 -1978
rect 2143 -2044 2223 -2030
rect 356 -2082 370 -2076
rect 290 -2096 370 -2082
rect 423 -2084 463 -2076
rect 791 -2078 871 -2064
rect 791 -2084 805 -2078
rect 423 -2124 805 -2084
rect 290 -2140 370 -2126
rect 290 -2192 304 -2140
rect 356 -2172 370 -2140
rect 791 -2130 805 -2124
rect 857 -2084 871 -2078
rect 1771 -2078 1851 -2064
rect 1771 -2084 1785 -2078
rect 857 -2124 1785 -2084
rect 857 -2130 871 -2124
rect 791 -2144 871 -2130
rect 1771 -2130 1785 -2124
rect 1837 -2130 1851 -2078
rect 1771 -2144 1851 -2130
rect 1901 -2166 1981 -2152
rect 1901 -2172 1915 -2166
rect 356 -2192 1915 -2172
rect 290 -2212 1915 -2192
rect 1901 -2218 1915 -2212
rect 1967 -2218 1981 -2166
rect 1901 -2232 1981 -2218
rect 2385 -2166 2465 -2152
rect 2385 -2218 2399 -2166
rect 2451 -2174 2465 -2166
rect 2493 -2174 2533 -1610
rect 2451 -2214 2533 -2174
rect 2451 -2218 2465 -2214
rect 2385 -2232 2465 -2218
rect 291 -2254 371 -2240
rect 291 -2306 305 -2254
rect 357 -2260 371 -2254
rect 357 -2300 2401 -2260
rect 357 -2306 371 -2300
rect 291 -2320 371 -2306
rect 291 -2364 371 -2354
rect 291 -2368 2401 -2364
rect 291 -2420 305 -2368
rect 357 -2404 2401 -2368
rect 357 -2420 371 -2404
rect 291 -2434 371 -2420
rect -3719 -2849 -3705 -2797
rect -3653 -2849 -3639 -2797
rect -3719 -2863 -3639 -2849
rect 202 -2799 282 -2785
rect 202 -2851 216 -2799
rect 268 -2851 282 -2799
rect 202 -2865 282 -2851
<< via2 >>
rect -4080 955 -4024 957
rect -4080 903 -4078 955
rect -4078 903 -4026 955
rect -4026 903 -4024 955
rect -4080 901 -4024 903
rect -4194 255 -4138 257
rect -4194 203 -4192 255
rect -4192 203 -4140 255
rect -4140 203 -4138 255
rect -4194 201 -4138 203
rect -4536 -441 -4480 -439
rect -4536 -493 -4534 -441
rect -4534 -493 -4482 -441
rect -4482 -493 -4480 -441
rect -4536 -495 -4480 -493
rect -4650 -1148 -4594 -1146
rect -4650 -1200 -4648 -1148
rect -4648 -1200 -4596 -1148
rect -4596 -1200 -4594 -1148
rect -4650 -1202 -4594 -1200
rect -1018 956 -962 958
rect -1018 904 -1016 956
rect -1016 904 -964 956
rect -964 904 -962 956
rect -1018 902 -962 904
rect -1564 255 -1508 257
rect -1564 203 -1562 255
rect -1562 203 -1510 255
rect -1510 203 -1508 255
rect -1564 201 -1508 203
rect -1564 -440 -1508 -438
rect -1564 -492 -1562 -440
rect -1562 -492 -1510 -440
rect -1510 -492 -1508 -440
rect -1564 -494 -1508 -492
rect -1018 -1148 -962 -1146
rect -1018 -1200 -1016 -1148
rect -1016 -1200 -964 -1148
rect -964 -1200 -962 -1148
rect -1018 -1202 -962 -1200
<< metal3 >>
rect -4102 959 -4002 978
rect -1040 959 -940 979
rect -4102 958 -940 959
rect -4102 957 -1018 958
rect -4102 901 -4080 957
rect -4024 902 -1018 957
rect -962 902 -940 958
rect -4024 901 -940 902
rect -4102 899 -940 901
rect -4102 878 -4002 899
rect -1040 879 -940 899
rect -4216 258 -4116 278
rect -1586 258 -1486 278
rect -4216 257 -1486 258
rect -4216 201 -4194 257
rect -4138 201 -1564 257
rect -1508 201 -1486 257
rect -4216 198 -1486 201
rect -4216 178 -4116 198
rect -1586 178 -1486 198
rect -4558 -436 -4458 -418
rect -1586 -436 -1486 -417
rect -4558 -438 -1486 -436
rect -4558 -439 -1564 -438
rect -4558 -495 -4536 -439
rect -4480 -494 -1564 -439
rect -1508 -494 -1486 -438
rect -4480 -495 -1486 -494
rect -4558 -496 -1486 -495
rect -4558 -518 -4458 -496
rect -1586 -517 -1486 -496
rect -4672 -1145 -4572 -1125
rect -1040 -1145 -940 -1125
rect -4672 -1146 -940 -1145
rect -4672 -1202 -4650 -1146
rect -4594 -1202 -1018 -1146
rect -962 -1202 -940 -1146
rect -4672 -1205 -940 -1202
rect -4672 -1225 -4572 -1205
rect -1040 -1225 -940 -1205
<< labels >>
flabel metal1 s -3960 -146 -3916 -100 2 FreeSans 2000 0 0 0 GND
port 1 nsew
flabel metal1 s -4880 873 -4819 933 2 FreeSans 2500 0 0 0 x0
port 2 nsew
flabel metal1 s -4767 812 -4706 872 2 FreeSans 2500 0 0 0 x0_bar
port 3 nsew
flabel metal1 s -4652 873 -4591 933 2 FreeSans 2500 0 0 0 x1
port 4 nsew
flabel metal1 s -4538 812 -4477 872 2 FreeSans 2500 0 0 0 x1_bar
port 5 nsew
flabel metal1 s -4423 877 -4362 937 2 FreeSans 2500 0 0 0 x2
port 6 nsew
flabel metal1 s -4311 813 -4250 873 2 FreeSans 2500 0 0 0 x2_bar
port 7 nsew
flabel metal1 s -4196 874 -4135 934 2 FreeSans 2500 0 0 0 x3
port 8 nsew
flabel metal1 s -4082 813 -4021 873 2 FreeSans 2500 0 0 0 x3_bar
port 9 nsew
flabel metal2 s 2370 -2290 2390 -2270 2 FreeSans 2000 0 0 0 s3_bar
port 10 nsew
flabel metal2 s -3810 1159 -3779 1190 2 FreeSans 2000 0 0 0 CLK1
port 11 nsew
flabel metal2 s 2370 -2396 2390 -2375 2 FreeSans 2000 0 0 0 s3
port 12 nsew
flabel metal2 s -3690 1165 -3667 1189 2 FreeSans 2000 0 0 0 Dis1
port 13 nsew
flabel metal2 s 277 1172 296 1193 2 FreeSans 2000 0 0 0 Dis3
port 14 nsew
flabel metal2 s 388 1169 413 1194 2 FreeSans 2000 0 0 0 CLK3
port 15 nsew
flabel metal2 s 536 1171 561 1195 2 FreeSans 2000 0 0 0 Dis2
port 16 nsew
flabel metal2 s 2124 1161 2158 1195 2 FreeSans 2000 0 0 0 CLK2
port 17 nsew
rlabel metal1 -2699 -2283 -2659 -2243 4 EESPFAL_3in_NAND_v2_0/OUT_bar
rlabel metal1 -2749 -2963 -2709 -2923 4 EESPFAL_3in_NAND_v2_0/GND!
rlabel metal1 -2749 -1783 -2709 -1743 4 EESPFAL_3in_NAND_v2_0/CLK
rlabel locali -2799 -2408 -2759 -2368 4 EESPFAL_3in_NAND_v2_0/OUT
rlabel locali -3709 -1893 -3689 -1873 4 EESPFAL_3in_NAND_v2_0/A
rlabel locali -3709 -2203 -3689 -2183 4 EESPFAL_3in_NAND_v2_0/A_bar
rlabel locali -3709 -2013 -3689 -1993 4 EESPFAL_3in_NAND_v2_0/B
rlabel locali -3709 -2283 -3689 -2263 4 EESPFAL_3in_NAND_v2_0/B_bar
rlabel locali -3709 -2123 -3689 -2103 4 EESPFAL_3in_NAND_v2_0/C
rlabel locali -3709 -2383 -3689 -2363 4 EESPFAL_3in_NAND_v2_0/C_bar
rlabel locali -2949 -2843 -2909 -2803 4 EESPFAL_3in_NAND_v2_0/Dis
rlabel metal1 -649 -2283 -609 -2243 4 EESPFAL_INV4_0/OUT
rlabel metal1 -699 -2963 -659 -2923 4 EESPFAL_INV4_0/GND!
rlabel metal1 -699 -1783 -659 -1743 4 EESPFAL_INV4_0/CLK
rlabel locali -749 -2408 -709 -2368 4 EESPFAL_INV4_0/OUT_bar
rlabel locali -119 -2163 -79 -2123 4 EESPFAL_INV4_0/A
rlabel locali -1279 -2403 -1239 -2363 4 EESPFAL_INV4_0/A_bar
rlabel locali -899 -2843 -859 -2803 4 EESPFAL_INV4_0/Dis
rlabel metal1 1291 -2284 1331 -2244 6 EESPFAL_3in_NOR_v2_0/OUT_bar
rlabel metal1 1341 -2964 1381 -2924 6 EESPFAL_3in_NOR_v2_0/GND!
rlabel metal1 1341 -1784 1381 -1744 6 EESPFAL_3in_NOR_v2_0/CLK
rlabel locali 1391 -2409 1431 -2369 6 EESPFAL_3in_NOR_v2_0/OUT
rlabel locali 2321 -1904 2341 -1884 6 EESPFAL_3in_NOR_v2_0/A
rlabel locali 2321 -2204 2341 -2184 6 EESPFAL_3in_NOR_v2_0/A_bar
rlabel locali 2321 -2014 2341 -1994 6 EESPFAL_3in_NOR_v2_0/B
rlabel locali 2321 -2324 2341 -2304 6 EESPFAL_3in_NOR_v2_0/B_bar
rlabel locali 2321 -2114 2341 -2094 6 EESPFAL_3in_NOR_v2_0/C
rlabel locali 2321 -2424 2341 -2404 6 EESPFAL_3in_NOR_v2_0/C_bar
rlabel locali 1541 -2844 1581 -2804 6 EESPFAL_3in_NOR_v2_0/Dis
rlabel metal1 -2700 -823 -2660 -783 2 EESPFAL_XOR_v3_1/OUT_bar
rlabel metal1 -2750 -143 -2710 -103 2 EESPFAL_XOR_v3_1/GND!
rlabel metal1 -2750 -1323 -2710 -1283 2 EESPFAL_XOR_v3_1/CLK
rlabel locali -2800 -698 -2760 -658 2 EESPFAL_XOR_v3_1/OUT
rlabel locali -3860 -1183 -3840 -1163 2 EESPFAL_XOR_v3_1/A
rlabel locali -3860 -1083 -3840 -1063 2 EESPFAL_XOR_v3_1/A_bar
rlabel locali -3860 -983 -3840 -963 2 EESPFAL_XOR_v3_1/B
rlabel locali -3860 -883 -3840 -863 2 EESPFAL_XOR_v3_1/B_bar
rlabel locali -2950 -263 -2910 -223 2 EESPFAL_XOR_v3_1/Dis
rlabel metal1 -510 -823 -470 -783 2 EESPFAL_INV4_1/OUT
rlabel metal1 -560 -143 -520 -103 2 EESPFAL_INV4_1/GND!
rlabel metal1 -560 -1323 -520 -1283 2 EESPFAL_INV4_1/CLK
rlabel locali -610 -698 -570 -658 2 EESPFAL_INV4_1/OUT_bar
rlabel locali 20 -943 60 -903 2 EESPFAL_INV4_1/A
rlabel locali -1140 -703 -1100 -663 2 EESPFAL_INV4_1/A_bar
rlabel locali -760 -263 -720 -223 2 EESPFAL_INV4_1/Dis
rlabel metal1 1370 -823 1410 -783 2 EESPFAL_NAND_v3_1/OUT_bar
rlabel metal1 1320 -143 1360 -103 2 EESPFAL_NAND_v3_1/GND!
rlabel metal1 1320 -1323 1360 -1283 2 EESPFAL_NAND_v3_1/CLK
rlabel locali 1270 -698 1310 -658 2 EESPFAL_NAND_v3_1/OUT
rlabel locali 510 -1083 530 -1063 2 EESPFAL_NAND_v3_1/A
rlabel locali 510 -863 530 -843 2 EESPFAL_NAND_v3_1/A_bar
rlabel locali 510 -963 530 -943 2 EESPFAL_NAND_v3_1/B
rlabel locali 510 -763 530 -743 2 EESPFAL_NAND_v3_1/B_bar
rlabel locali 1120 -263 1160 -223 2 EESPFAL_NAND_v3_1/Dis
rlabel metal1 -2700 537 -2660 577 4 EESPFAL_XOR_v3_0/OUT_bar
rlabel metal1 -2750 -143 -2710 -103 4 EESPFAL_XOR_v3_0/GND!
rlabel metal1 -2750 1037 -2710 1077 4 EESPFAL_XOR_v3_0/CLK
rlabel locali -2800 412 -2760 452 4 EESPFAL_XOR_v3_0/OUT
rlabel locali -3860 917 -3840 937 4 EESPFAL_XOR_v3_0/A
rlabel locali -3860 817 -3840 837 4 EESPFAL_XOR_v3_0/A_bar
rlabel locali -3860 717 -3840 737 4 EESPFAL_XOR_v3_0/B
rlabel locali -3860 617 -3840 637 4 EESPFAL_XOR_v3_0/B_bar
rlabel locali -2950 -23 -2910 17 4 EESPFAL_XOR_v3_0/Dis
rlabel metal1 -510 537 -470 577 4 EESPFAL_INV4_2/OUT
rlabel metal1 -560 -143 -520 -103 4 EESPFAL_INV4_2/GND!
rlabel metal1 -560 1037 -520 1077 4 EESPFAL_INV4_2/CLK
rlabel locali -610 412 -570 452 4 EESPFAL_INV4_2/OUT_bar
rlabel locali 20 657 60 697 4 EESPFAL_INV4_2/A
rlabel locali -1140 417 -1100 457 4 EESPFAL_INV4_2/A_bar
rlabel locali -760 -23 -720 17 4 EESPFAL_INV4_2/Dis
rlabel metal1 1370 537 1410 577 4 EESPFAL_NAND_v3_0/OUT_bar
rlabel metal1 1320 -143 1360 -103 4 EESPFAL_NAND_v3_0/GND!
rlabel metal1 1320 1037 1360 1077 4 EESPFAL_NAND_v3_0/CLK
rlabel locali 1270 412 1310 452 4 EESPFAL_NAND_v3_0/OUT
rlabel locali 510 817 530 837 4 EESPFAL_NAND_v3_0/A
rlabel locali 510 597 530 617 4 EESPFAL_NAND_v3_0/A_bar
rlabel locali 510 697 530 717 4 EESPFAL_NAND_v3_0/B
rlabel locali 510 497 530 517 4 EESPFAL_NAND_v3_0/B_bar
rlabel locali 1120 -23 1160 17 4 EESPFAL_NAND_v3_0/Dis
<< end >>
