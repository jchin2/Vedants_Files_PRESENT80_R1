magic
tech sky130A
magscale 1 2
timestamp 1677167062
<< locali >>
rect -1487 1258 -1407 1281
rect -1487 1224 -1464 1258
rect -1430 1224 -1407 1258
rect -1487 1189 -1407 1224
rect 1660 1189 1740 1205
rect -1487 1186 247 1189
rect -1487 1152 -1464 1186
rect -1430 1152 247 1186
rect -1487 1149 247 1152
rect 1660 1182 1805 1189
rect -1487 1114 -1407 1149
rect 1660 1148 1683 1182
rect 1717 1149 1805 1182
rect 1717 1148 1740 1149
rect 1660 1125 1740 1148
rect -1487 1080 -1464 1114
rect -1430 1080 -1407 1114
rect -1487 1057 -1407 1080
rect -1373 524 -1293 547
rect -1373 490 -1350 524
rect -1316 490 -1293 524
rect -1373 455 -1293 490
rect -1373 452 -233 455
rect -1373 418 -1350 452
rect -1316 418 -233 452
rect -1373 415 -233 418
rect -1373 380 -1293 415
rect 3212 408 3319 431
rect -1373 346 -1350 380
rect -1316 346 -1293 380
rect 2056 360 2136 383
rect -1373 323 -1293 346
rect -1259 333 -1179 356
rect -1259 299 -1236 333
rect -1202 299 -1179 333
rect 2056 326 2079 360
rect 2113 326 2136 360
rect 2056 303 2136 326
rect 3212 374 3262 408
rect 3296 374 3319 408
rect 3212 336 3319 374
rect -1259 264 -1179 299
rect -1259 261 -203 264
rect -1259 227 -1236 261
rect -1202 227 -203 261
rect -1259 224 -203 227
rect -1259 189 -1179 224
rect -1259 155 -1236 189
rect -1202 155 -1179 189
rect -1259 132 -1179 155
rect -1145 -92 -1065 -69
rect 828 -91 958 -51
rect -1145 -126 -1122 -92
rect -1088 -126 -1065 -92
rect -1145 -161 -1065 -126
rect -649 -149 -421 -109
rect -649 -161 -609 -149
rect -1145 -164 -609 -161
rect -1145 -198 -1122 -164
rect -1088 -198 -609 -164
rect -461 -161 -421 -149
rect -1145 -201 -609 -198
rect -1145 -236 -1065 -201
rect -1145 -270 -1122 -236
rect -1088 -270 -1065 -236
rect -1145 -293 -1065 -270
rect -575 -206 -495 -183
rect -461 -201 247 -161
rect -575 -240 -552 -206
rect -518 -240 -495 -206
rect -575 -255 -495 -240
rect -575 -278 -353 -255
rect -575 -312 -552 -278
rect -518 -312 -353 -278
rect -575 -335 -353 -312
rect -1487 -372 -1407 -349
rect -1487 -406 -1464 -372
rect -1430 -406 -1407 -372
rect -1487 -441 -1407 -406
rect -575 -350 -495 -335
rect -575 -384 -552 -350
rect -518 -384 -495 -350
rect -575 -407 -495 -384
rect 918 -389 958 -91
rect 1660 -160 1740 -137
rect 1660 -194 1683 -160
rect 1717 -161 1740 -160
rect 2077 -161 2117 303
rect 3212 302 3262 336
rect 3296 302 3319 336
rect 3212 279 3319 302
rect 1717 -194 1805 -161
rect 1660 -201 1805 -194
rect 2077 -201 2662 -161
rect 1660 -217 1740 -201
rect -461 -431 -108 -391
rect 918 -429 1450 -389
rect 3239 -393 3319 -373
rect 2742 -396 3319 -393
rect 2742 -430 3262 -396
rect 3296 -430 3319 -396
rect -461 -441 -421 -431
rect 2742 -433 3319 -430
rect -1487 -444 -421 -441
rect -1487 -478 -1464 -444
rect -1430 -478 -421 -444
rect 3239 -453 3319 -433
rect -1487 -481 -421 -478
rect -1487 -516 -1407 -481
rect -1487 -550 -1464 -516
rect -1430 -550 -1407 -516
rect -1487 -573 -1407 -550
rect 3303 -883 3383 -860
rect -803 -920 -723 -897
rect -803 -954 -780 -920
rect -746 -954 -723 -920
rect -803 -989 -723 -954
rect 3303 -917 3326 -883
rect 3360 -917 3383 -883
rect 3303 -955 3383 -917
rect 3303 -989 3326 -955
rect 3360 -989 3383 -955
rect -803 -992 -258 -989
rect -803 -1026 -780 -992
rect -746 -1026 -258 -992
rect -803 -1029 -258 -1026
rect -803 -1064 -723 -1029
rect 2000 -1029 2512 -989
rect 3303 -1012 3383 -989
rect -803 -1098 -780 -1064
rect -746 -1098 -723 -1064
rect -803 -1121 -723 -1098
rect 230 -1738 310 -1715
rect 230 -1739 253 -1738
rect 172 -1772 253 -1739
rect 287 -1772 310 -1738
rect 172 -1779 310 -1772
rect 552 -1739 592 -1669
rect 552 -1779 2832 -1739
rect 230 -1795 310 -1779
<< viali >>
rect -1464 1224 -1430 1258
rect -1464 1152 -1430 1186
rect 1683 1148 1717 1182
rect -1464 1080 -1430 1114
rect -1350 490 -1316 524
rect -1350 418 -1316 452
rect 1348 418 1382 452
rect 2505 412 2539 446
rect -1350 346 -1316 380
rect -1236 299 -1202 333
rect 2079 326 2113 360
rect 3262 374 3296 408
rect -1236 227 -1202 261
rect 1378 227 1412 261
rect -1236 155 -1202 189
rect -1122 -126 -1088 -92
rect -1122 -198 -1088 -164
rect -1122 -270 -1088 -236
rect -552 -240 -518 -206
rect -552 -312 -518 -278
rect -1464 -406 -1430 -372
rect -552 -384 -518 -350
rect 1683 -194 1717 -160
rect 3262 302 3296 336
rect 3262 -430 3296 -396
rect -1464 -478 -1430 -444
rect -1464 -550 -1430 -516
rect -780 -954 -746 -920
rect 3326 -917 3360 -883
rect 3326 -989 3360 -955
rect -780 -1026 -746 -992
rect 1293 -1036 1327 -1002
rect -780 -1098 -746 -1064
rect 253 -1772 287 -1738
<< metal1 >>
rect -1487 1258 -1407 1333
rect -1487 1224 -1464 1258
rect -1430 1224 -1407 1258
rect -1487 1186 -1407 1224
rect -1487 1152 -1464 1186
rect -1430 1152 -1407 1186
rect -1487 1114 -1407 1152
rect -1487 1080 -1464 1114
rect -1430 1080 -1407 1114
rect -1487 -372 -1407 1080
rect -1487 -406 -1464 -372
rect -1430 -406 -1407 -372
rect -1487 -444 -1407 -406
rect -1487 -478 -1464 -444
rect -1430 -478 -1407 -444
rect -1487 -516 -1407 -478
rect -1487 -550 -1464 -516
rect -1430 -550 -1407 -516
rect -1487 -1924 -1407 -550
rect -1373 524 -1293 1333
rect -1373 490 -1350 524
rect -1316 490 -1293 524
rect -1373 452 -1293 490
rect -1373 418 -1350 452
rect -1316 418 -1293 452
rect -1373 380 -1293 418
rect -1373 346 -1350 380
rect -1316 346 -1293 380
rect -1373 -1924 -1293 346
rect -1259 333 -1179 1333
rect -1259 299 -1236 333
rect -1202 299 -1179 333
rect -1259 261 -1179 299
rect -1259 227 -1236 261
rect -1202 227 -1179 261
rect -1259 189 -1179 227
rect -1259 155 -1236 189
rect -1202 155 -1179 189
rect -1259 -628 -1179 155
rect -1259 -680 -1245 -628
rect -1193 -680 -1179 -628
rect -1259 -696 -1179 -680
rect -1259 -748 -1245 -696
rect -1193 -748 -1179 -696
rect -1259 -764 -1179 -748
rect -1259 -816 -1245 -764
rect -1193 -816 -1179 -764
rect -1259 -1924 -1179 -816
rect -1145 -92 -1065 1333
rect -1145 -126 -1122 -92
rect -1088 -126 -1065 -92
rect -1145 -164 -1065 -126
rect -1145 -198 -1122 -164
rect -1088 -198 -1065 -164
rect -1145 -236 -1065 -198
rect -1145 -270 -1122 -236
rect -1088 -270 -1065 -236
rect -1145 -1924 -1065 -270
rect -1031 -316 -951 1333
rect -1031 -368 -1017 -316
rect -965 -368 -951 -316
rect -1031 -384 -951 -368
rect -1031 -436 -1017 -384
rect -965 -436 -951 -384
rect -1031 -452 -951 -436
rect -1031 -504 -1017 -452
rect -965 -504 -951 -452
rect -1031 -1923 -951 -504
rect -917 -472 -837 1333
rect -917 -524 -903 -472
rect -851 -524 -837 -472
rect -917 -540 -837 -524
rect -917 -592 -903 -540
rect -851 -592 -837 -540
rect -917 -608 -837 -592
rect -917 -660 -903 -608
rect -851 -660 -837 -608
rect -917 -1665 -837 -660
rect -917 -1717 -903 -1665
rect -851 -1717 -837 -1665
rect -917 -1733 -837 -1717
rect -917 -1785 -903 -1733
rect -851 -1785 -837 -1733
rect -917 -1801 -837 -1785
rect -917 -1853 -903 -1801
rect -851 -1853 -837 -1801
rect -917 -1924 -837 -1853
rect -803 1259 -723 1333
rect -803 1207 -789 1259
rect -737 1207 -723 1259
rect -803 1191 -723 1207
rect -803 1139 -789 1191
rect -737 1139 -723 1191
rect -803 1123 -723 1139
rect -803 1071 -789 1123
rect -737 1071 -723 1123
rect -803 -920 -723 1071
rect -803 -954 -780 -920
rect -746 -954 -723 -920
rect -803 -992 -723 -954
rect -803 -1026 -780 -992
rect -746 -1026 -723 -992
rect -803 -1064 -723 -1026
rect -803 -1098 -780 -1064
rect -746 -1098 -723 -1064
rect -803 -1923 -723 -1098
rect -689 -87 -609 1333
rect -689 -139 -675 -87
rect -623 -139 -609 -87
rect -689 -155 -609 -139
rect -689 -207 -675 -155
rect -623 -207 -609 -155
rect -689 -223 -609 -207
rect -689 -275 -675 -223
rect -623 -275 -609 -223
rect -689 -926 -609 -275
rect -689 -978 -675 -926
rect -623 -978 -609 -926
rect -689 -994 -609 -978
rect -689 -1046 -675 -994
rect -623 -1046 -609 -994
rect -689 -1062 -609 -1046
rect -689 -1114 -675 -1062
rect -623 -1114 -609 -1062
rect -689 -1923 -609 -1114
rect -575 -206 -495 1333
rect -575 -240 -552 -206
rect -518 -240 -495 -206
rect -575 -278 -495 -240
rect -575 -312 -552 -278
rect -518 -312 -495 -278
rect -575 -350 -495 -312
rect -575 -384 -552 -350
rect -518 -384 -495 -350
rect -575 -1923 -495 -384
rect -461 1233 -353 1333
rect 873 1233 1205 1333
rect 2121 1233 2417 1333
rect -461 -1823 -381 1233
rect 1660 1191 1740 1205
rect 1660 1139 1674 1191
rect 1726 1139 1740 1191
rect 1660 1125 1740 1139
rect 1325 461 1405 475
rect 1325 409 1339 461
rect 1391 409 1405 461
rect 1325 395 1405 409
rect 2482 455 2562 469
rect 2482 403 2496 455
rect 2548 403 2562 455
rect 2482 389 2562 403
rect 3239 417 3319 431
rect 2056 369 2136 383
rect 2056 317 2070 369
rect 2122 317 2136 369
rect 2056 303 2136 317
rect 3239 365 3253 417
rect 3305 365 3319 417
rect 3239 345 3319 365
rect 3239 293 3253 345
rect 3305 293 3319 345
rect 1355 270 1435 284
rect 3239 279 3319 293
rect 1355 218 1369 270
rect 1421 218 1435 270
rect 1355 204 1435 218
rect 1660 -151 1740 -137
rect 1660 -203 1674 -151
rect 1726 -203 1740 -151
rect 1660 -217 1740 -203
rect 884 -345 1205 -245
rect 2085 -345 2417 -245
rect 556 -387 636 -373
rect 556 -439 570 -387
rect 622 -439 636 -387
rect 556 -453 636 -439
rect 3239 -387 3319 -373
rect 3239 -439 3253 -387
rect 3305 -439 3319 -387
rect 3239 -453 3319 -439
rect 3303 -874 3383 -860
rect 3303 -926 3317 -874
rect 3369 -926 3383 -874
rect 3303 -946 3383 -926
rect 1270 -993 1350 -979
rect 1270 -1045 1284 -993
rect 1336 -1045 1350 -993
rect 3303 -998 3317 -946
rect 3369 -998 3383 -946
rect 3303 -1012 3383 -998
rect 1270 -1059 1350 -1045
rect 230 -1729 310 -1715
rect 230 -1781 244 -1729
rect 296 -1781 310 -1729
rect 230 -1795 310 -1781
rect -461 -1923 -353 -1823
rect 657 -1923 1169 -1823
rect 2085 -1923 2417 -1823
<< via1 >>
rect -1245 -680 -1193 -628
rect -1245 -748 -1193 -696
rect -1245 -816 -1193 -764
rect -1017 -368 -965 -316
rect -1017 -436 -965 -384
rect -1017 -504 -965 -452
rect -903 -524 -851 -472
rect -903 -592 -851 -540
rect -903 -660 -851 -608
rect -903 -1717 -851 -1665
rect -903 -1785 -851 -1733
rect -903 -1853 -851 -1801
rect -789 1207 -737 1259
rect -789 1139 -737 1191
rect -789 1071 -737 1123
rect -675 -139 -623 -87
rect -675 -207 -623 -155
rect -675 -275 -623 -223
rect -675 -978 -623 -926
rect -675 -1046 -623 -994
rect -675 -1114 -623 -1062
rect 1674 1182 1726 1191
rect 1674 1148 1683 1182
rect 1683 1148 1717 1182
rect 1717 1148 1726 1182
rect 1674 1139 1726 1148
rect 1339 452 1391 461
rect 1339 418 1348 452
rect 1348 418 1382 452
rect 1382 418 1391 452
rect 1339 409 1391 418
rect 2496 446 2548 455
rect 2496 412 2505 446
rect 2505 412 2539 446
rect 2539 412 2548 446
rect 2496 403 2548 412
rect 2070 360 2122 369
rect 2070 326 2079 360
rect 2079 326 2113 360
rect 2113 326 2122 360
rect 2070 317 2122 326
rect 3253 408 3305 417
rect 3253 374 3262 408
rect 3262 374 3296 408
rect 3296 374 3305 408
rect 3253 365 3305 374
rect 3253 336 3305 345
rect 3253 302 3262 336
rect 3262 302 3296 336
rect 3296 302 3305 336
rect 3253 293 3305 302
rect 1369 261 1421 270
rect 1369 227 1378 261
rect 1378 227 1412 261
rect 1412 227 1421 261
rect 1369 218 1421 227
rect 1674 -160 1726 -151
rect 1674 -194 1683 -160
rect 1683 -194 1717 -160
rect 1717 -194 1726 -160
rect 1674 -203 1726 -194
rect 570 -439 622 -387
rect 3253 -396 3305 -387
rect 3253 -430 3262 -396
rect 3262 -430 3296 -396
rect 3296 -430 3305 -396
rect 3253 -439 3305 -430
rect 3317 -883 3369 -874
rect 3317 -917 3326 -883
rect 3326 -917 3360 -883
rect 3360 -917 3369 -883
rect 3317 -926 3369 -917
rect 1284 -1002 1336 -993
rect 1284 -1036 1293 -1002
rect 1293 -1036 1327 -1002
rect 1327 -1036 1336 -1002
rect 1284 -1045 1336 -1036
rect 3317 -955 3369 -946
rect 3317 -989 3326 -955
rect 3326 -989 3360 -955
rect 3360 -989 3369 -955
rect 3317 -998 3369 -989
rect 244 -1738 296 -1729
rect 244 -1772 253 -1738
rect 253 -1772 287 -1738
rect 287 -1772 296 -1738
rect 244 -1781 296 -1772
<< metal2 >>
rect -803 1259 -723 1273
rect -803 1207 -789 1259
rect -737 1207 -723 1259
rect -803 1191 -723 1207
rect -803 1139 -789 1191
rect -737 1185 -723 1191
rect 1660 1191 1740 1205
rect 1660 1185 1674 1191
rect -737 1145 1674 1185
rect -737 1139 -723 1145
rect -803 1123 -723 1139
rect 1660 1139 1674 1145
rect 1726 1139 1740 1191
rect 1660 1125 1740 1139
rect -803 1071 -789 1123
rect -737 1071 -723 1123
rect -803 1057 -723 1071
rect 1325 461 1405 475
rect 1325 455 1339 461
rect 980 415 1339 455
rect -689 -87 -609 -73
rect -689 -139 -675 -87
rect -623 -139 -609 -87
rect -689 -155 -609 -139
rect -689 -207 -675 -155
rect -623 -161 -609 -155
rect 980 -161 1020 415
rect 1325 409 1339 415
rect 1391 409 1405 461
rect 2482 455 2562 469
rect 2482 449 2496 455
rect 1325 395 1405 409
rect 2164 409 2496 449
rect 2056 369 2136 383
rect 2056 317 2070 369
rect 2122 317 2136 369
rect 2056 303 2136 317
rect 1355 270 1435 284
rect 1355 218 1369 270
rect 1421 218 1435 270
rect 1355 204 1435 218
rect -623 -201 1020 -161
rect -623 -207 -609 -201
rect -689 -223 -609 -207
rect -689 -275 -675 -223
rect -623 -275 -609 -223
rect -689 -289 -609 -275
rect -1031 -316 -951 -302
rect -1031 -368 -1017 -316
rect -965 -368 -951 -316
rect -1031 -384 -951 -368
rect -1031 -436 -1017 -384
rect -965 -390 -951 -384
rect 556 -387 636 -373
rect 556 -390 570 -387
rect -965 -430 570 -390
rect -965 -436 -951 -430
rect -1031 -452 -951 -436
rect -1031 -504 -1017 -452
rect -965 -504 -951 -452
rect 556 -439 570 -430
rect 622 -393 636 -387
rect 1375 -393 1415 204
rect 1660 -151 1740 -137
rect 1660 -203 1674 -151
rect 1726 -203 1740 -151
rect 1660 -217 1740 -203
rect 622 -433 1415 -393
rect 622 -439 636 -433
rect 556 -453 636 -439
rect -1031 -518 -951 -504
rect -917 -472 -837 -458
rect -917 -524 -903 -472
rect -851 -481 -837 -472
rect 1680 -481 1720 -217
rect -851 -521 1720 -481
rect -851 -524 -837 -521
rect -917 -540 -837 -524
rect -917 -592 -903 -540
rect -851 -592 -837 -540
rect -917 -608 -837 -592
rect -1259 -628 -1179 -614
rect -1259 -680 -1245 -628
rect -1193 -680 -1179 -628
rect -917 -660 -903 -608
rect -851 -660 -837 -608
rect -917 -674 -837 -660
rect -1259 -696 -1179 -680
rect -1259 -748 -1245 -696
rect -1193 -702 -1179 -696
rect 2164 -702 2204 409
rect 2482 403 2496 409
rect 2548 403 2562 455
rect 2482 389 2562 403
rect 3239 417 3319 431
rect 3239 365 3253 417
rect 3305 365 3319 417
rect 3239 345 3319 365
rect 3239 293 3253 345
rect 3305 293 3319 345
rect 3239 279 3319 293
rect 3259 -373 3299 279
rect 3239 -387 3319 -373
rect 3239 -439 3253 -387
rect 3305 -439 3319 -387
rect 3239 -453 3319 -439
rect -1193 -742 2204 -702
rect -1193 -748 -1179 -742
rect -1259 -764 -1179 -748
rect -1259 -816 -1245 -764
rect -1193 -816 -1179 -764
rect -1259 -830 -1179 -816
rect 3303 -874 3383 -860
rect -689 -926 -609 -912
rect -689 -978 -675 -926
rect -623 -978 -609 -926
rect -689 -994 -609 -978
rect 3303 -926 3317 -874
rect 3369 -916 3383 -874
rect 3369 -926 3428 -916
rect 3303 -946 3428 -926
rect -689 -1046 -675 -994
rect -623 -1000 -609 -994
rect 1270 -993 1350 -979
rect 1270 -1000 1284 -993
rect -623 -1040 1284 -1000
rect -623 -1046 -609 -1040
rect -689 -1062 -609 -1046
rect 1270 -1045 1284 -1040
rect 1336 -1045 1350 -993
rect 3303 -998 3317 -946
rect 3369 -956 3428 -946
rect 3369 -998 3383 -956
rect 3303 -1012 3383 -998
rect 1270 -1059 1350 -1045
rect -689 -1114 -675 -1062
rect -623 -1114 -609 -1062
rect -689 -1128 -609 -1114
rect -917 -1665 -837 -1651
rect -917 -1717 -903 -1665
rect -851 -1717 -837 -1665
rect -917 -1733 -837 -1717
rect -917 -1785 -903 -1733
rect -851 -1739 -837 -1733
rect 230 -1729 310 -1715
rect 230 -1739 244 -1729
rect -851 -1779 244 -1739
rect -851 -1785 -837 -1779
rect -917 -1801 -837 -1785
rect 230 -1781 244 -1779
rect 296 -1781 310 -1729
rect 230 -1795 310 -1781
rect -917 -1853 -903 -1801
rect -851 -1853 -837 -1801
rect -917 -1867 -837 -1853
use CMOS_3in_AND  CMOS_3in_AND_0
timestamp 1505768449
transform 1 0 152 0 -1 -1089
box -541 -870 542 870
use CMOS_3in_OR  CMOS_3in_OR_0
timestamp 1505768449
transform 1 0 2922 0 -1 -1089
box -541 -870 542 870
use CMOS_AND  CMOS_AND_0
timestamp 1505768449
transform 1 0 2857 0 1 499
box -476 -870 476 870
use CMOS_AND  CMOS_AND_1
timestamp 1505768449
transform 1 0 1645 0 -1 -1089
box -476 -870 476 870
use CMOS_XNOR  CMOS_XNOR_0
timestamp 1505768449
transform 1 0 260 0 1 499
box -649 -870 650 870
use CMOS_XOR  CMOS_XOR_0
timestamp 1505768449
transform 1 0 1645 0 1 499
box -476 -870 476 870
<< labels >>
flabel metal1 s -552 -312 -518 -278 2 FreeSans 2500 0 0 0 GND
port 1 nsew
flabel metal1 s -1477 1267 -1416 1327 2 FreeSans 3126 0 0 0 x0
port 2 nsew
flabel metal1 s -1364 1206 -1303 1266 2 FreeSans 3126 0 0 0 x0_bar
port 3 nsew
flabel metal1 s -1249 1267 -1188 1327 2 FreeSans 3126 0 0 0 x1
port 4 nsew
flabel metal1 s -1135 1206 -1074 1266 2 FreeSans 3126 0 0 0 x1_bar
port 5 nsew
flabel metal1 s -1021 1268 -960 1328 2 FreeSans 3126 0 0 0 x2
port 6 nsew
flabel metal1 s -908 1207 -847 1267 2 FreeSans 3126 0 0 0 x2_bar
port 7 nsew
flabel metal1 s -793 1268 -732 1328 2 FreeSans 3126 0 0 0 x3
port 8 nsew
flabel metal1 s -443 1267 -409 1301 2 FreeSans 2500 0 0 0 VDD
port 9 nsew
flabel metal1 s -678 1208 -617 1268 2 FreeSans 3126 0 0 0 x3_bar
port 10 nsew
flabel metal2 s 3326 -917 3360 -883 2 FreeSans 2500 0 0 0 s3
port 11 nsew
<< properties >>
string path -29.475 -18.050 55.100 -18.050 
<< end >>
