magic
tech sky130A
magscale 1 2
timestamp 1671306811
<< locali >>
rect -450 37 -370 60
rect -450 3 -427 37
rect -393 3 -370 37
rect -450 -20 -370 3
rect -330 37 -250 60
rect -330 3 -307 37
rect -273 3 -250 37
rect -330 -20 -250 3
rect -450 -83 -370 -60
rect -450 -117 -427 -83
rect -393 -117 -370 -83
rect -450 -140 -370 -117
rect -330 -83 -250 -60
rect -330 -117 -307 -83
rect -273 -117 -250 -83
rect -330 -140 -250 -117
<< viali >>
rect -427 3 -393 37
rect -307 3 -273 37
rect -427 -117 -393 -83
rect -307 -117 -273 -83
<< metal1 >>
rect -480 46 -220 90
rect -480 -6 -436 46
rect -384 -6 -316 46
rect -264 -6 -220 46
rect -480 -74 -220 -6
rect -480 -126 -436 -74
rect -384 -126 -316 -74
rect -264 -126 -220 -74
rect -480 -170 -220 -126
<< via1 >>
rect -436 37 -384 46
rect -436 3 -427 37
rect -427 3 -393 37
rect -393 3 -384 37
rect -436 -6 -384 3
rect -316 37 -264 46
rect -316 3 -307 37
rect -307 3 -273 37
rect -273 3 -264 37
rect -316 -6 -264 3
rect -436 -83 -384 -74
rect -436 -117 -427 -83
rect -427 -117 -393 -83
rect -393 -117 -384 -83
rect -436 -126 -384 -117
rect -316 -83 -264 -74
rect -316 -117 -307 -83
rect -307 -117 -273 -83
rect -273 -117 -264 -83
rect -316 -126 -264 -117
<< metal2 >>
rect -480 48 -220 90
rect -480 -8 -438 48
rect -382 -8 -318 48
rect -262 -8 -220 48
rect -480 -72 -220 -8
rect -480 -128 -438 -72
rect -382 -128 -318 -72
rect -262 -128 -220 -72
rect -480 -170 -220 -128
<< via2 >>
rect -438 46 -382 48
rect -438 -6 -436 46
rect -436 -6 -384 46
rect -384 -6 -382 46
rect -438 -8 -382 -6
rect -318 46 -262 48
rect -318 -6 -316 46
rect -316 -6 -264 46
rect -264 -6 -262 46
rect -318 -8 -262 -6
rect -438 -74 -382 -72
rect -438 -126 -436 -74
rect -436 -126 -384 -74
rect -384 -126 -382 -74
rect -438 -128 -382 -126
rect -318 -74 -262 -72
rect -318 -126 -316 -74
rect -316 -126 -264 -74
rect -264 -126 -262 -74
rect -318 -128 -262 -126
<< metal3 >>
rect -480 52 -220 90
rect -480 -12 -442 52
rect -378 -12 -322 52
rect -258 -12 -220 52
rect -480 -68 -220 -12
rect -480 -132 -442 -68
rect -378 -132 -322 -68
rect -258 -132 -220 -68
rect -480 -170 -220 -132
<< via3 >>
rect -442 48 -378 52
rect -442 -8 -438 48
rect -438 -8 -382 48
rect -382 -8 -378 48
rect -442 -12 -378 -8
rect -322 48 -258 52
rect -322 -8 -318 48
rect -318 -8 -262 48
rect -262 -8 -258 48
rect -322 -12 -258 -8
rect -442 -72 -378 -68
rect -442 -128 -438 -72
rect -438 -128 -382 -72
rect -382 -128 -378 -72
rect -442 -132 -378 -128
rect -322 -72 -258 -68
rect -322 -128 -318 -72
rect -318 -128 -262 -72
rect -262 -128 -258 -72
rect -322 -132 -258 -128
<< metal4 >>
rect -480 52 -220 90
rect -480 -12 -442 52
rect -378 -12 -322 52
rect -258 -12 -220 52
rect -480 -68 -220 -12
rect -480 -132 -442 -68
rect -378 -132 -322 -68
rect -258 -132 -220 -68
rect -480 -170 -220 -132
<< end >>
