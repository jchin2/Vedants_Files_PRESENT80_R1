magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -33 -15 863 505
<< l67d20 >>
rect 135 475 755 495
rect 735 455 755 475
rect 585 455 605 475
rect 435 455 455 475
rect 285 455 305 475
rect 135 455 155 475
rect 800 25 840 455
rect 725 25 765 455
rect 650 25 690 455
rect 575 25 615 455
rect 500 25 540 455
rect 425 25 465 455
rect 350 25 390 455
rect 275 25 315 455
rect 200 25 240 455
rect 125 25 165 455
rect 50 25 90 455
rect 810 5 830 25
rect 660 5 680 25
rect 510 5 530 25
rect 360 5 380 25
rect 210 5 230 25
rect 60 5 80 25
rect 60 -15 830 5
rect -10 25 30 455
<< l66d20 >>
rect 100 490 790 505
rect 775 0 790 490
rect 700 0 715 490
rect 625 0 640 490
rect 550 0 565 490
rect 475 0 490 490
rect 400 0 415 490
rect 325 0 340 490
rect 250 0 265 490
rect 175 0 190 490
rect 100 0 115 490
<< l66d44 >>
rect 437 419 454 436
rect 437 385 454 402
rect 437 351 454 368
rect 437 317 454 334
rect 437 283 454 300
rect 437 249 454 266
rect 812 351 829 368
rect 737 346 754 363
rect 812 283 829 300
rect 737 278 754 295
rect 662 283 679 300
rect 587 283 604 300
rect 512 283 529 300
rect 662 351 679 368
rect 587 351 604 368
rect 512 351 529 368
rect 737 380 754 397
rect 662 385 679 402
rect 587 385 604 402
rect 812 249 829 266
rect 737 244 754 261
rect 662 249 679 266
rect 587 249 604 266
rect 512 249 529 266
rect 512 385 529 402
rect 737 414 754 431
rect 662 419 679 436
rect 812 317 829 334
rect 737 312 754 329
rect 662 317 679 334
rect 587 317 604 334
rect 512 317 529 334
rect 587 419 604 436
rect 512 419 529 436
rect 812 419 829 436
rect 812 385 829 402
rect 287 419 304 436
rect 362 351 379 368
rect 287 351 304 368
rect 212 351 229 368
rect 137 351 154 368
rect 62 351 79 368
rect 212 419 229 436
rect 362 317 379 334
rect 287 317 304 334
rect 212 317 229 334
rect 137 317 154 334
rect 62 317 79 334
rect 137 419 154 436
rect 362 283 379 300
rect 287 283 304 300
rect 212 283 229 300
rect 137 283 154 300
rect 62 283 79 300
rect 62 419 79 436
rect 362 249 379 266
rect 287 249 304 266
rect 212 249 229 266
rect 137 249 154 266
rect 62 249 79 266
rect 362 419 379 436
rect 362 385 379 402
rect 287 385 304 402
rect 212 385 229 402
rect 137 385 154 402
rect 62 385 79 402
rect 2 351 19 368
rect 2 317 19 334
rect 2 283 19 300
rect 2 419 19 436
rect 2 249 19 266
rect 2 385 19 402
rect 212 181 229 198
rect 362 113 379 130
rect 287 113 304 130
rect 212 113 229 130
rect 137 113 154 130
rect 62 113 79 130
rect 137 181 154 198
rect 62 181 79 198
rect 212 215 229 232
rect 137 215 154 232
rect 62 215 79 232
rect 287 45 304 62
rect 362 79 379 96
rect 287 79 304 96
rect 212 79 229 96
rect 137 79 154 96
rect 62 79 79 96
rect 212 45 229 62
rect 137 45 154 62
rect 362 147 379 164
rect 287 147 304 164
rect 212 147 229 164
rect 137 147 154 164
rect 362 45 379 62
rect 62 147 79 164
rect 62 45 79 62
rect 362 215 379 232
rect 287 215 304 232
rect 362 181 379 198
rect 287 181 304 198
rect 2 147 19 164
rect 2 45 19 62
rect 2 113 19 130
rect 2 181 19 198
rect 2 215 19 232
rect 2 79 19 96
rect 812 147 829 164
rect 737 142 754 159
rect 662 147 679 164
rect 587 147 604 164
rect 512 147 529 164
rect 662 215 679 232
rect 812 113 829 130
rect 737 108 754 125
rect 662 113 679 130
rect 587 113 604 130
rect 512 113 529 130
rect 587 215 604 232
rect 812 79 829 96
rect 737 74 754 91
rect 662 79 679 96
rect 587 79 604 96
rect 512 79 529 96
rect 512 215 529 232
rect 812 45 829 62
rect 737 40 754 57
rect 662 45 679 62
rect 587 45 604 62
rect 512 45 529 62
rect 812 215 829 232
rect 437 215 454 232
rect 437 181 454 198
rect 437 147 454 164
rect 437 113 454 130
rect 437 79 454 96
rect 437 45 454 62
rect 812 181 829 198
rect 737 176 754 193
rect 662 181 679 198
rect 587 181 604 198
rect 512 181 529 198
rect 737 210 754 227
<< l65d20 >>
rect 40 15 850 465
<< l93d44 >>
rect 40 3 863 478
<< l125d44 >>
rect 82 -3 808 483
<< l94d20 >>
rect -33 3 40 478
<< l65d44 >>
rect -20 15 40 465
<< end >>
