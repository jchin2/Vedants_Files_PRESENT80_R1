magic
tech sky130A
timestamp 1667076306
<< nwell >>
rect -1440 720 -560 815
rect -1205 525 -795 720
<< nmos >>
rect -1360 165 -1345 315
rect -1285 165 -1270 315
rect -1120 165 -1105 315
rect -1045 165 -1030 315
rect -970 165 -955 315
rect -895 165 -880 315
rect -730 165 -715 315
rect -655 165 -640 315
<< pmos >>
rect -1120 550 -1105 700
rect -1045 550 -1030 700
rect -970 550 -955 700
rect -895 550 -880 700
<< ndiff >>
rect -1420 280 -1360 315
rect -1420 260 -1400 280
rect -1380 260 -1360 280
rect -1420 240 -1360 260
rect -1420 220 -1400 240
rect -1380 220 -1360 240
rect -1420 200 -1360 220
rect -1420 180 -1400 200
rect -1380 180 -1360 200
rect -1420 165 -1360 180
rect -1345 165 -1285 315
rect -1270 280 -1210 315
rect -1270 260 -1250 280
rect -1230 260 -1210 280
rect -1270 240 -1210 260
rect -1270 220 -1250 240
rect -1230 220 -1210 240
rect -1270 200 -1210 220
rect -1270 180 -1250 200
rect -1230 180 -1210 200
rect -1270 165 -1210 180
rect -1180 280 -1120 315
rect -1180 260 -1160 280
rect -1140 260 -1120 280
rect -1180 240 -1120 260
rect -1180 220 -1160 240
rect -1140 220 -1120 240
rect -1180 200 -1120 220
rect -1180 180 -1160 200
rect -1140 180 -1120 200
rect -1180 165 -1120 180
rect -1105 280 -1045 315
rect -1105 260 -1085 280
rect -1065 260 -1045 280
rect -1105 240 -1045 260
rect -1105 220 -1085 240
rect -1065 220 -1045 240
rect -1105 200 -1045 220
rect -1105 180 -1085 200
rect -1065 180 -1045 200
rect -1105 165 -1045 180
rect -1030 280 -970 315
rect -1030 260 -1010 280
rect -990 260 -970 280
rect -1030 240 -970 260
rect -1030 220 -1010 240
rect -990 220 -970 240
rect -1030 200 -970 220
rect -1030 180 -1010 200
rect -990 180 -970 200
rect -1030 165 -970 180
rect -955 280 -895 315
rect -955 260 -935 280
rect -915 260 -895 280
rect -955 240 -895 260
rect -955 220 -935 240
rect -915 220 -895 240
rect -955 200 -895 220
rect -955 180 -935 200
rect -915 180 -895 200
rect -955 165 -895 180
rect -880 280 -820 315
rect -880 260 -860 280
rect -840 260 -820 280
rect -880 240 -820 260
rect -880 220 -860 240
rect -840 220 -820 240
rect -880 200 -820 220
rect -880 180 -860 200
rect -840 180 -820 200
rect -880 165 -820 180
rect -790 280 -730 315
rect -790 260 -770 280
rect -750 260 -730 280
rect -790 240 -730 260
rect -790 220 -770 240
rect -750 220 -730 240
rect -790 200 -730 220
rect -790 180 -770 200
rect -750 180 -730 200
rect -790 165 -730 180
rect -715 280 -655 315
rect -715 260 -695 280
rect -675 260 -655 280
rect -715 240 -655 260
rect -715 220 -695 240
rect -675 220 -655 240
rect -715 200 -655 220
rect -715 180 -695 200
rect -675 180 -655 200
rect -715 165 -655 180
rect -640 280 -580 315
rect -640 260 -620 280
rect -600 260 -580 280
rect -640 240 -580 260
rect -640 220 -620 240
rect -600 220 -580 240
rect -640 200 -580 220
rect -640 180 -620 200
rect -600 180 -580 200
rect -640 165 -580 180
<< pdiff >>
rect -1180 665 -1120 700
rect -1180 645 -1160 665
rect -1140 645 -1120 665
rect -1180 625 -1120 645
rect -1180 605 -1160 625
rect -1140 605 -1120 625
rect -1180 585 -1120 605
rect -1180 565 -1160 585
rect -1140 565 -1120 585
rect -1180 550 -1120 565
rect -1105 665 -1045 700
rect -1105 645 -1085 665
rect -1065 645 -1045 665
rect -1105 625 -1045 645
rect -1105 605 -1085 625
rect -1065 605 -1045 625
rect -1105 585 -1045 605
rect -1105 565 -1085 585
rect -1065 565 -1045 585
rect -1105 550 -1045 565
rect -1030 665 -970 700
rect -1030 645 -1010 665
rect -990 645 -970 665
rect -1030 625 -970 645
rect -1030 605 -1010 625
rect -990 605 -970 625
rect -1030 585 -970 605
rect -1030 565 -1010 585
rect -990 565 -970 585
rect -1030 550 -970 565
rect -955 665 -895 700
rect -955 645 -935 665
rect -915 645 -895 665
rect -955 625 -895 645
rect -955 605 -935 625
rect -915 605 -895 625
rect -955 585 -895 605
rect -955 565 -935 585
rect -915 565 -895 585
rect -955 550 -895 565
rect -880 665 -820 700
rect -880 645 -860 665
rect -840 645 -820 665
rect -880 625 -820 645
rect -880 605 -860 625
rect -840 605 -820 625
rect -880 585 -820 605
rect -880 565 -860 585
rect -840 565 -820 585
rect -880 550 -820 565
<< ndiffc >>
rect -1400 260 -1380 280
rect -1400 220 -1380 240
rect -1400 180 -1380 200
rect -1250 260 -1230 280
rect -1250 220 -1230 240
rect -1250 180 -1230 200
rect -1160 260 -1140 280
rect -1160 220 -1140 240
rect -1160 180 -1140 200
rect -1085 260 -1065 280
rect -1085 220 -1065 240
rect -1085 180 -1065 200
rect -1010 260 -990 280
rect -1010 220 -990 240
rect -1010 180 -990 200
rect -935 260 -915 280
rect -935 220 -915 240
rect -935 180 -915 200
rect -860 260 -840 280
rect -860 220 -840 240
rect -860 180 -840 200
rect -770 260 -750 280
rect -770 220 -750 240
rect -770 180 -750 200
rect -695 260 -675 280
rect -695 220 -675 240
rect -695 180 -675 200
rect -620 260 -600 280
rect -620 220 -600 240
rect -620 180 -600 200
<< pdiffc >>
rect -1160 645 -1140 665
rect -1160 605 -1140 625
rect -1160 565 -1140 585
rect -1085 645 -1065 665
rect -1085 605 -1065 625
rect -1085 565 -1065 585
rect -1010 645 -990 665
rect -1010 605 -990 625
rect -1010 565 -990 585
rect -935 645 -915 665
rect -935 605 -915 625
rect -935 565 -915 585
rect -860 645 -840 665
rect -860 605 -840 625
rect -860 565 -840 585
<< psubdiff >>
rect -1420 80 -580 95
rect -1420 60 -1410 80
rect -1390 60 -1370 80
rect -1350 60 -1330 80
rect -1310 60 -1290 80
rect -1270 60 -1250 80
rect -1230 60 -1210 80
rect -1190 60 -1170 80
rect -1150 60 -1130 80
rect -1110 60 -1090 80
rect -1070 60 -1050 80
rect -1030 60 -1010 80
rect -990 60 -970 80
rect -950 60 -930 80
rect -910 60 -890 80
rect -870 60 -850 80
rect -830 60 -810 80
rect -790 60 -770 80
rect -750 60 -730 80
rect -710 60 -690 80
rect -670 60 -650 80
rect -630 60 -610 80
rect -590 60 -580 80
rect -1420 45 -580 60
<< nsubdiff >>
rect -1420 775 -580 790
rect -1420 755 -1410 775
rect -1390 755 -1370 775
rect -1350 755 -1330 775
rect -1310 755 -1290 775
rect -1270 755 -1250 775
rect -1230 755 -1210 775
rect -1190 755 -1170 775
rect -1150 755 -1130 775
rect -1110 755 -1090 775
rect -1070 755 -1050 775
rect -1030 755 -1010 775
rect -990 755 -970 775
rect -950 755 -930 775
rect -910 755 -890 775
rect -870 755 -850 775
rect -830 755 -810 775
rect -790 755 -770 775
rect -750 755 -730 775
rect -710 755 -690 775
rect -670 755 -650 775
rect -630 755 -610 775
rect -590 755 -580 775
rect -1420 740 -580 755
<< psubdiffcont >>
rect -1410 60 -1390 80
rect -1370 60 -1350 80
rect -1330 60 -1310 80
rect -1290 60 -1270 80
rect -1250 60 -1230 80
rect -1210 60 -1190 80
rect -1170 60 -1150 80
rect -1130 60 -1110 80
rect -1090 60 -1070 80
rect -1050 60 -1030 80
rect -1010 60 -990 80
rect -970 60 -950 80
rect -930 60 -910 80
rect -890 60 -870 80
rect -850 60 -830 80
rect -810 60 -790 80
rect -770 60 -750 80
rect -730 60 -710 80
rect -690 60 -670 80
rect -650 60 -630 80
rect -610 60 -590 80
<< nsubdiffcont >>
rect -1410 755 -1390 775
rect -1370 755 -1350 775
rect -1330 755 -1310 775
rect -1290 755 -1270 775
rect -1250 755 -1230 775
rect -1210 755 -1190 775
rect -1170 755 -1150 775
rect -1130 755 -1110 775
rect -1090 755 -1070 775
rect -1050 755 -1030 775
rect -1010 755 -990 775
rect -970 755 -950 775
rect -930 755 -910 775
rect -890 755 -870 775
rect -850 755 -830 775
rect -810 755 -790 775
rect -770 755 -750 775
rect -730 755 -710 775
rect -690 755 -670 775
rect -650 755 -630 775
rect -610 755 -590 775
<< poly >>
rect -1120 715 -1030 730
rect -1120 700 -1105 715
rect -1045 700 -1030 715
rect -970 715 -880 730
rect -970 700 -955 715
rect -895 700 -880 715
rect -1120 535 -1105 550
rect -1045 475 -1030 550
rect -970 535 -955 550
rect -895 535 -880 550
rect -995 525 -955 535
rect -995 505 -985 525
rect -965 505 -955 525
rect -995 495 -955 505
rect -1045 465 -1005 475
rect -1045 445 -1035 465
rect -1015 445 -1005 465
rect -1045 435 -1005 445
rect -1385 385 -1345 395
rect -1385 365 -1375 385
rect -1355 365 -1345 385
rect -1385 355 -1345 365
rect -1310 385 -1270 395
rect -1310 365 -1300 385
rect -1280 365 -1270 385
rect -1310 355 -1270 365
rect -1360 315 -1345 355
rect -1285 315 -1270 355
rect -1120 315 -1105 330
rect -1045 315 -1030 435
rect -970 315 -955 495
rect -655 415 -615 425
rect -655 395 -645 415
rect -625 395 -615 415
rect -655 385 -615 395
rect -895 315 -880 330
rect -730 315 -715 335
rect -655 315 -640 385
rect -1360 150 -1345 165
rect -1285 150 -1270 165
rect -1120 150 -1105 165
rect -1045 150 -1030 165
rect -970 150 -955 165
rect -895 150 -880 165
rect -730 150 -715 165
rect -655 150 -640 165
rect -1120 140 -1080 150
rect -1120 120 -1110 140
rect -1090 120 -1080 140
rect -1120 110 -1080 120
rect -920 140 -880 150
rect -920 120 -910 140
rect -890 120 -880 140
rect -920 110 -880 120
rect -755 140 -715 150
rect -755 120 -745 140
rect -725 120 -715 140
rect -755 110 -715 120
<< polycont >>
rect -985 505 -965 525
rect -1035 445 -1015 465
rect -1375 365 -1355 385
rect -1300 365 -1280 385
rect -645 395 -625 415
rect -1110 120 -1090 140
rect -910 120 -890 140
rect -745 120 -725 140
<< locali >>
rect -1420 775 -580 785
rect -1420 755 -1410 775
rect -1390 755 -1370 775
rect -1350 755 -1330 775
rect -1310 755 -1290 775
rect -1270 755 -1250 775
rect -1230 755 -1210 775
rect -1190 755 -1170 775
rect -1150 755 -1130 775
rect -1110 755 -1090 775
rect -1070 755 -1050 775
rect -1030 755 -1010 775
rect -990 755 -970 775
rect -950 755 -930 775
rect -910 755 -890 775
rect -870 755 -850 775
rect -830 755 -810 775
rect -790 755 -770 775
rect -750 755 -730 775
rect -710 755 -690 775
rect -670 755 -650 775
rect -630 755 -610 775
rect -590 755 -580 775
rect -1420 745 -580 755
rect -1170 665 -1130 680
rect -1170 645 -1160 665
rect -1140 645 -1130 665
rect -1170 625 -1130 645
rect -1170 605 -1160 625
rect -1140 605 -1130 625
rect -1170 585 -1130 605
rect -1170 565 -1160 585
rect -1140 565 -1130 585
rect -1170 555 -1130 565
rect -1095 665 -1055 680
rect -1095 645 -1085 665
rect -1065 645 -1055 665
rect -1095 625 -1055 645
rect -1095 605 -1085 625
rect -1065 605 -1055 625
rect -1095 585 -1055 605
rect -1095 565 -1085 585
rect -1065 565 -1055 585
rect -1095 550 -1055 565
rect -1020 665 -980 680
rect -1020 645 -1010 665
rect -990 645 -980 665
rect -1020 625 -980 645
rect -1020 605 -1010 625
rect -990 605 -980 625
rect -1020 585 -980 605
rect -1020 565 -1010 585
rect -990 565 -980 585
rect -1020 555 -980 565
rect -945 665 -905 680
rect -945 645 -935 665
rect -915 645 -905 665
rect -945 625 -905 645
rect -945 605 -935 625
rect -915 605 -905 625
rect -945 585 -905 605
rect -945 565 -935 585
rect -915 565 -905 585
rect -945 550 -905 565
rect -870 665 -830 680
rect -870 645 -860 665
rect -840 645 -830 665
rect -870 625 -830 645
rect -870 605 -860 625
rect -840 605 -830 625
rect -870 585 -830 605
rect -870 565 -860 585
rect -840 565 -830 585
rect -870 555 -830 565
rect -1085 525 -1065 550
rect -995 525 -955 535
rect -1420 505 -1160 525
rect -1200 495 -1160 505
rect -1260 475 -1220 485
rect -1420 455 -1250 475
rect -1230 455 -1220 475
rect -1200 475 -1190 495
rect -1170 475 -1160 495
rect -1200 465 -1160 475
rect -1085 505 -985 525
rect -965 505 -955 525
rect -1260 445 -1220 455
rect -1420 415 -1280 435
rect -1300 395 -1280 415
rect -1385 385 -1345 395
rect -1420 365 -1375 385
rect -1355 365 -1345 385
rect -1385 355 -1345 365
rect -1310 385 -1270 395
rect -1310 365 -1300 385
rect -1280 365 -1270 385
rect -1310 355 -1270 365
rect -1085 335 -1065 505
rect -995 495 -955 505
rect -1045 465 -1005 475
rect -935 465 -915 550
rect -795 525 -755 535
rect -795 505 -785 525
rect -765 505 -580 525
rect -795 495 -755 505
rect -1045 445 -1035 465
rect -1015 445 -580 465
rect -1045 435 -1005 445
rect -935 335 -915 445
rect -795 415 -755 425
rect -655 415 -615 425
rect -795 395 -785 415
rect -765 395 -645 415
rect -625 395 -615 415
rect -795 385 -755 395
rect -655 385 -615 395
rect -1250 315 -1055 335
rect -1250 295 -1230 315
rect -1410 280 -1370 295
rect -1410 260 -1400 280
rect -1380 260 -1370 280
rect -1410 240 -1370 260
rect -1410 220 -1400 240
rect -1380 220 -1370 240
rect -1410 200 -1370 220
rect -1410 180 -1400 200
rect -1380 180 -1370 200
rect -1410 170 -1370 180
rect -1260 280 -1220 295
rect -1260 260 -1250 280
rect -1230 260 -1220 280
rect -1260 240 -1220 260
rect -1260 220 -1250 240
rect -1230 220 -1220 240
rect -1260 200 -1220 220
rect -1260 180 -1250 200
rect -1230 180 -1220 200
rect -1260 170 -1220 180
rect -1170 280 -1130 295
rect -1170 260 -1160 280
rect -1140 260 -1130 280
rect -1170 240 -1130 260
rect -1170 220 -1160 240
rect -1140 220 -1130 240
rect -1170 200 -1130 220
rect -1170 180 -1160 200
rect -1140 180 -1130 200
rect -1170 170 -1130 180
rect -1095 280 -1055 315
rect -945 315 -600 335
rect -1095 260 -1085 280
rect -1065 260 -1055 280
rect -1095 240 -1055 260
rect -1095 220 -1085 240
rect -1065 220 -1055 240
rect -1095 200 -1055 220
rect -1095 180 -1085 200
rect -1065 180 -1055 200
rect -1095 170 -1055 180
rect -1020 280 -980 295
rect -1020 260 -1010 280
rect -990 260 -980 280
rect -1020 240 -980 260
rect -1020 220 -1010 240
rect -990 220 -980 240
rect -1020 200 -980 220
rect -1020 180 -1010 200
rect -990 180 -980 200
rect -1020 170 -980 180
rect -945 280 -905 315
rect -780 295 -760 315
rect -620 295 -600 315
rect -945 260 -935 280
rect -915 260 -905 280
rect -945 240 -905 260
rect -945 220 -935 240
rect -915 220 -905 240
rect -945 200 -905 220
rect -945 180 -935 200
rect -915 180 -905 200
rect -945 170 -905 180
rect -870 280 -830 295
rect -870 260 -860 280
rect -840 260 -830 280
rect -870 240 -830 260
rect -870 220 -860 240
rect -840 220 -830 240
rect -870 200 -830 220
rect -870 180 -860 200
rect -840 180 -830 200
rect -870 170 -830 180
rect -780 280 -740 295
rect -780 260 -770 280
rect -750 260 -740 280
rect -780 240 -740 260
rect -780 220 -770 240
rect -750 220 -740 240
rect -780 200 -740 220
rect -780 180 -770 200
rect -750 180 -740 200
rect -780 170 -740 180
rect -705 280 -665 295
rect -705 260 -695 280
rect -675 260 -665 280
rect -705 240 -665 260
rect -705 220 -695 240
rect -675 220 -665 240
rect -705 200 -665 220
rect -705 180 -695 200
rect -675 180 -665 200
rect -705 170 -665 180
rect -630 280 -590 295
rect -630 260 -620 280
rect -600 260 -590 280
rect -630 240 -590 260
rect -630 220 -620 240
rect -600 220 -590 240
rect -630 200 -590 220
rect -630 180 -620 200
rect -600 180 -590 200
rect -630 170 -590 180
rect -1120 140 -1080 150
rect -920 140 -880 150
rect -1420 120 -1110 140
rect -1090 120 -910 140
rect -890 120 -880 140
rect -1120 110 -1080 120
rect -920 110 -880 120
rect -755 140 -715 150
rect -755 120 -745 140
rect -725 120 -715 140
rect -755 110 -715 120
rect -1420 80 -580 90
rect -1420 60 -1410 80
rect -1390 60 -1370 80
rect -1350 60 -1330 80
rect -1310 60 -1290 80
rect -1270 60 -1250 80
rect -1230 60 -1210 80
rect -1190 60 -1170 80
rect -1150 60 -1130 80
rect -1110 60 -1090 80
rect -1070 60 -1050 80
rect -1030 60 -1010 80
rect -990 60 -970 80
rect -950 60 -930 80
rect -910 60 -890 80
rect -870 60 -850 80
rect -830 60 -810 80
rect -790 60 -770 80
rect -750 60 -730 80
rect -710 60 -690 80
rect -670 60 -650 80
rect -630 60 -610 80
rect -590 60 -580 80
rect -1420 50 -580 60
<< viali >>
rect -1410 755 -1390 775
rect -1370 755 -1350 775
rect -1330 755 -1310 775
rect -1290 755 -1270 775
rect -1250 755 -1230 775
rect -1210 755 -1190 775
rect -1170 755 -1150 775
rect -1130 755 -1110 775
rect -1090 755 -1070 775
rect -1050 755 -1030 775
rect -1010 755 -990 775
rect -970 755 -950 775
rect -930 755 -910 775
rect -890 755 -870 775
rect -850 755 -830 775
rect -810 755 -790 775
rect -770 755 -750 775
rect -730 755 -710 775
rect -690 755 -670 775
rect -650 755 -630 775
rect -610 755 -590 775
rect -1160 645 -1140 665
rect -1160 605 -1140 625
rect -1160 565 -1140 585
rect -1010 645 -990 665
rect -1010 605 -990 625
rect -1010 565 -990 585
rect -860 645 -840 665
rect -860 605 -840 625
rect -860 565 -840 585
rect -1250 455 -1230 475
rect -1190 475 -1170 495
rect -985 505 -965 525
rect -785 505 -765 525
rect -785 395 -765 415
rect -1400 260 -1380 280
rect -1400 220 -1380 240
rect -1400 180 -1380 200
rect -1160 260 -1140 280
rect -1160 220 -1140 240
rect -1160 180 -1140 200
rect -1010 260 -990 280
rect -1010 220 -990 240
rect -1010 180 -990 200
rect -860 260 -840 280
rect -860 220 -840 240
rect -860 180 -840 200
rect -695 260 -675 280
rect -695 220 -675 240
rect -695 180 -675 200
rect -745 120 -725 140
rect -1410 60 -1390 80
rect -1370 60 -1350 80
rect -1330 60 -1310 80
rect -1290 60 -1270 80
rect -1250 60 -1230 80
rect -1210 60 -1190 80
rect -1170 60 -1150 80
rect -1130 60 -1110 80
rect -1090 60 -1070 80
rect -1050 60 -1030 80
rect -1010 60 -990 80
rect -970 60 -950 80
rect -930 60 -910 80
rect -890 60 -870 80
rect -850 60 -830 80
rect -810 60 -790 80
rect -770 60 -750 80
rect -730 60 -710 80
rect -690 60 -670 80
rect -650 60 -630 80
rect -610 60 -590 80
<< metal1 >>
rect -1420 775 -580 790
rect -1420 755 -1410 775
rect -1390 755 -1370 775
rect -1350 755 -1330 775
rect -1310 755 -1290 775
rect -1270 755 -1250 775
rect -1230 755 -1210 775
rect -1190 755 -1170 775
rect -1150 755 -1130 775
rect -1110 755 -1090 775
rect -1070 755 -1050 775
rect -1030 755 -1010 775
rect -990 755 -970 775
rect -950 755 -930 775
rect -910 755 -890 775
rect -870 755 -850 775
rect -830 755 -810 775
rect -790 755 -770 775
rect -750 755 -730 775
rect -710 755 -690 775
rect -670 755 -650 775
rect -630 755 -610 775
rect -590 755 -580 775
rect -1420 740 -580 755
rect -1400 295 -1380 740
rect -1170 665 -1130 740
rect -1170 645 -1160 665
rect -1140 645 -1130 665
rect -1170 625 -1130 645
rect -1170 605 -1160 625
rect -1140 605 -1130 625
rect -1170 585 -1130 605
rect -1170 565 -1160 585
rect -1140 565 -1130 585
rect -1170 555 -1130 565
rect -1020 665 -980 740
rect -1020 645 -1010 665
rect -990 645 -980 665
rect -1020 625 -980 645
rect -1020 605 -1010 625
rect -990 605 -980 625
rect -1020 585 -980 605
rect -1020 565 -1010 585
rect -990 565 -980 585
rect -1020 555 -980 565
rect -870 665 -830 740
rect -870 645 -860 665
rect -840 645 -830 665
rect -870 625 -830 645
rect -870 605 -860 625
rect -840 605 -830 625
rect -870 585 -830 605
rect -870 565 -860 585
rect -840 565 -830 585
rect -870 555 -830 565
rect -995 525 -955 535
rect -795 525 -755 535
rect -995 505 -985 525
rect -965 505 -785 525
rect -765 505 -755 525
rect -1200 495 -1160 505
rect -995 495 -955 505
rect -795 495 -755 505
rect -1260 475 -1220 485
rect -1260 455 -1250 475
rect -1230 455 -1220 475
rect -1200 475 -1190 495
rect -1170 475 -1160 495
rect -1200 465 -1160 475
rect -1260 445 -1220 455
rect -1250 365 -1230 445
rect -1190 415 -1170 465
rect -795 415 -755 425
rect -1190 395 -785 415
rect -765 395 -755 415
rect -795 385 -755 395
rect -1250 345 -785 365
rect -1410 280 -1370 295
rect -1410 260 -1400 280
rect -1380 260 -1370 280
rect -1410 240 -1370 260
rect -1410 220 -1400 240
rect -1380 220 -1370 240
rect -1410 200 -1370 220
rect -1410 180 -1400 200
rect -1380 180 -1370 200
rect -1410 170 -1370 180
rect -1170 280 -1130 295
rect -1170 260 -1160 280
rect -1140 260 -1130 280
rect -1170 240 -1130 260
rect -1170 220 -1160 240
rect -1140 220 -1130 240
rect -1170 200 -1130 220
rect -1170 180 -1160 200
rect -1140 180 -1130 200
rect -1170 170 -1130 180
rect -1020 280 -980 295
rect -1020 260 -1010 280
rect -990 260 -980 280
rect -1020 240 -980 260
rect -1020 220 -1010 240
rect -990 220 -980 240
rect -1020 200 -980 220
rect -1020 180 -1010 200
rect -990 180 -980 200
rect -1020 170 -980 180
rect -870 280 -830 295
rect -870 260 -860 280
rect -840 260 -830 280
rect -870 240 -830 260
rect -870 220 -860 240
rect -840 220 -830 240
rect -870 200 -830 220
rect -870 180 -860 200
rect -840 180 -830 200
rect -870 170 -830 180
rect -1160 95 -1140 170
rect -1010 95 -990 170
rect -860 95 -840 170
rect -805 140 -785 345
rect -695 295 -675 740
rect -705 280 -665 295
rect -705 260 -695 280
rect -675 260 -665 280
rect -705 240 -665 260
rect -705 220 -695 240
rect -675 220 -665 240
rect -705 200 -665 220
rect -705 180 -695 200
rect -675 180 -665 200
rect -705 170 -665 180
rect -755 140 -715 150
rect -805 120 -745 140
rect -725 120 -715 140
rect -755 110 -715 120
rect -1420 80 -580 95
rect -1420 60 -1410 80
rect -1390 60 -1370 80
rect -1350 60 -1330 80
rect -1310 60 -1290 80
rect -1270 60 -1250 80
rect -1230 60 -1210 80
rect -1190 60 -1170 80
rect -1150 60 -1130 80
rect -1110 60 -1090 80
rect -1070 60 -1050 80
rect -1030 60 -1010 80
rect -990 60 -970 80
rect -950 60 -930 80
rect -910 60 -890 80
rect -870 60 -850 80
rect -830 60 -810 80
rect -790 60 -770 80
rect -750 60 -730 80
rect -710 60 -690 80
rect -670 60 -650 80
rect -630 60 -610 80
rect -590 60 -580 80
rect -1420 45 -580 60
<< labels >>
rlabel locali -1415 510 -1405 520 7 A
port 1 w
rlabel locali -1415 460 -1405 470 7 B
port 3 w
rlabel viali -985 505 -965 525 7 OUT_bar
port 6 w
rlabel locali -1035 445 -1015 465 7 OUT
port 5 w
rlabel locali -1110 120 -1090 140 7 Dis
port 7 w
rlabel metal1 -1010 755 -990 775 7 CLK
port 9 w
rlabel locali -1415 420 -1405 430 7 B_bar
port 4 w
rlabel locali -1415 370 -1405 380 7 A_bar
port 2 w
rlabel metal1 -1010 60 -990 80 7 GND!
port 8 w
<< end >>
