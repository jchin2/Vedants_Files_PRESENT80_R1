magic
tech sky130A
magscale 1 2
timestamp 1677185616
<< nwell >>
rect -2556 1280 -1604 1510
rect -998 1280 -46 1510
rect 214 1280 1166 1510
rect 1426 1280 2378 1510
rect -2500 590 -1650 1280
rect -977 590 -87 1280
rect 235 590 1125 1280
rect 1447 590 2337 1280
rect -2500 -1588 -1279 -898
rect -977 -1588 -87 -898
rect 235 -1588 1125 -898
rect -2556 -1818 -1258 -1588
rect -998 -1818 -46 -1588
rect 214 -1818 1166 -1588
<< pwell >>
rect -2466 -78 -1694 356
rect -963 -78 -101 356
rect 249 -78 1111 356
rect 1461 -78 2323 356
rect -2546 -230 -1257 -78
rect -988 -230 -56 -78
rect 224 -230 1156 -78
rect 1436 -230 2368 -78
rect -2466 -664 -1293 -230
rect -963 -664 -101 -230
rect 249 -664 1111 -230
<< nmos >>
rect -2320 30 -2290 330
rect -2170 30 -2140 330
rect -2020 30 -1990 330
rect -1870 30 -1840 330
rect -817 30 -787 330
rect -667 30 -637 330
rect -277 30 -247 330
rect 395 30 425 330
rect 545 30 575 330
rect 935 30 965 330
rect 1607 30 1637 330
rect 1757 30 1787 330
rect 2147 30 2177 330
rect -2320 -638 -2290 -338
rect -2170 -638 -2140 -338
rect -2020 -638 -1990 -338
rect -1870 -638 -1840 -338
rect -1469 -638 -1439 -338
rect -817 -638 -787 -338
rect -667 -638 -637 -338
rect -277 -638 -247 -338
rect 395 -638 425 -338
rect 545 -638 575 -338
rect 935 -638 965 -338
<< pmos >>
rect -2320 640 -2290 1240
rect -2170 640 -2140 1240
rect -2020 640 -1990 1240
rect -1870 640 -1840 1240
rect -817 640 -787 1240
rect -667 640 -637 1240
rect -277 640 -247 1240
rect 395 640 425 1240
rect 545 640 575 1240
rect 935 640 965 1240
rect 1607 640 1637 1240
rect 1757 640 1787 1240
rect 2147 640 2177 1240
rect -2320 -1548 -2290 -948
rect -2170 -1548 -2140 -948
rect -2020 -1548 -1990 -948
rect -1870 -1548 -1840 -948
rect -1469 -1548 -1439 -948
rect -817 -1548 -787 -948
rect -667 -1548 -637 -948
rect -277 -1548 -247 -948
rect 395 -1548 425 -948
rect 545 -1548 575 -948
rect 935 -1548 965 -948
<< ndiff >>
rect -2440 299 -2320 330
rect -2440 265 -2397 299
rect -2363 265 -2320 299
rect -2440 231 -2320 265
rect -2440 197 -2397 231
rect -2363 197 -2320 231
rect -2440 163 -2320 197
rect -2440 129 -2397 163
rect -2363 129 -2320 163
rect -2440 95 -2320 129
rect -2440 61 -2397 95
rect -2363 61 -2320 95
rect -2440 30 -2320 61
rect -2290 30 -2170 330
rect -2140 299 -2020 330
rect -2140 265 -2097 299
rect -2063 265 -2020 299
rect -2140 231 -2020 265
rect -2140 197 -2097 231
rect -2063 197 -2020 231
rect -2140 163 -2020 197
rect -2140 129 -2097 163
rect -2063 129 -2020 163
rect -2140 95 -2020 129
rect -2140 61 -2097 95
rect -2063 61 -2020 95
rect -2140 30 -2020 61
rect -1990 30 -1870 330
rect -1840 299 -1720 330
rect -1840 265 -1797 299
rect -1763 265 -1720 299
rect -1840 231 -1720 265
rect -1840 197 -1797 231
rect -1763 197 -1720 231
rect -1840 163 -1720 197
rect -1840 129 -1797 163
rect -1763 129 -1720 163
rect -1840 95 -1720 129
rect -1840 61 -1797 95
rect -1763 61 -1720 95
rect -1840 30 -1720 61
rect -937 299 -817 330
rect -937 265 -894 299
rect -860 265 -817 299
rect -937 231 -817 265
rect -937 197 -894 231
rect -860 197 -817 231
rect -937 163 -817 197
rect -937 129 -894 163
rect -860 129 -817 163
rect -937 95 -817 129
rect -937 61 -894 95
rect -860 61 -817 95
rect -937 30 -817 61
rect -787 299 -667 330
rect -787 265 -744 299
rect -710 265 -667 299
rect -787 231 -667 265
rect -787 197 -744 231
rect -710 197 -667 231
rect -787 163 -667 197
rect -787 129 -744 163
rect -710 129 -667 163
rect -787 95 -667 129
rect -787 61 -744 95
rect -710 61 -667 95
rect -787 30 -667 61
rect -637 299 -517 330
rect -637 265 -594 299
rect -560 265 -517 299
rect -637 231 -517 265
rect -637 197 -594 231
rect -560 197 -517 231
rect -637 163 -517 197
rect -637 129 -594 163
rect -560 129 -517 163
rect -637 95 -517 129
rect -637 61 -594 95
rect -560 61 -517 95
rect -637 30 -517 61
rect -397 299 -277 330
rect -397 265 -354 299
rect -320 265 -277 299
rect -397 231 -277 265
rect -397 197 -354 231
rect -320 197 -277 231
rect -397 163 -277 197
rect -397 129 -354 163
rect -320 129 -277 163
rect -397 95 -277 129
rect -397 61 -354 95
rect -320 61 -277 95
rect -397 30 -277 61
rect -247 299 -127 330
rect -247 265 -204 299
rect -170 265 -127 299
rect -247 231 -127 265
rect -247 197 -204 231
rect -170 197 -127 231
rect -247 163 -127 197
rect -247 129 -204 163
rect -170 129 -127 163
rect -247 95 -127 129
rect -247 61 -204 95
rect -170 61 -127 95
rect -247 30 -127 61
rect 275 299 395 330
rect 275 265 318 299
rect 352 265 395 299
rect 275 231 395 265
rect 275 197 318 231
rect 352 197 395 231
rect 275 163 395 197
rect 275 129 318 163
rect 352 129 395 163
rect 275 95 395 129
rect 275 61 318 95
rect 352 61 395 95
rect 275 30 395 61
rect 425 30 545 330
rect 575 299 695 330
rect 575 265 618 299
rect 652 265 695 299
rect 575 231 695 265
rect 575 197 618 231
rect 652 197 695 231
rect 575 163 695 197
rect 575 129 618 163
rect 652 129 695 163
rect 575 95 695 129
rect 575 61 618 95
rect 652 61 695 95
rect 575 30 695 61
rect 815 299 935 330
rect 815 265 858 299
rect 892 265 935 299
rect 815 231 935 265
rect 815 197 858 231
rect 892 197 935 231
rect 815 163 935 197
rect 815 129 858 163
rect 892 129 935 163
rect 815 95 935 129
rect 815 61 858 95
rect 892 61 935 95
rect 815 30 935 61
rect 965 299 1085 330
rect 965 265 1008 299
rect 1042 265 1085 299
rect 965 231 1085 265
rect 965 197 1008 231
rect 1042 197 1085 231
rect 965 163 1085 197
rect 965 129 1008 163
rect 1042 129 1085 163
rect 965 95 1085 129
rect 965 61 1008 95
rect 1042 61 1085 95
rect 965 30 1085 61
rect 1487 299 1607 330
rect 1487 265 1530 299
rect 1564 265 1607 299
rect 1487 231 1607 265
rect 1487 197 1530 231
rect 1564 197 1607 231
rect 1487 163 1607 197
rect 1487 129 1530 163
rect 1564 129 1607 163
rect 1487 95 1607 129
rect 1487 61 1530 95
rect 1564 61 1607 95
rect 1487 30 1607 61
rect 1637 299 1757 330
rect 1637 265 1680 299
rect 1714 265 1757 299
rect 1637 231 1757 265
rect 1637 197 1680 231
rect 1714 197 1757 231
rect 1637 163 1757 197
rect 1637 129 1680 163
rect 1714 129 1757 163
rect 1637 95 1757 129
rect 1637 61 1680 95
rect 1714 61 1757 95
rect 1637 30 1757 61
rect 1787 299 1907 330
rect 1787 265 1830 299
rect 1864 265 1907 299
rect 1787 231 1907 265
rect 1787 197 1830 231
rect 1864 197 1907 231
rect 1787 163 1907 197
rect 1787 129 1830 163
rect 1864 129 1907 163
rect 1787 95 1907 129
rect 1787 61 1830 95
rect 1864 61 1907 95
rect 1787 30 1907 61
rect 2027 299 2147 330
rect 2027 265 2070 299
rect 2104 265 2147 299
rect 2027 231 2147 265
rect 2027 197 2070 231
rect 2104 197 2147 231
rect 2027 163 2147 197
rect 2027 129 2070 163
rect 2104 129 2147 163
rect 2027 95 2147 129
rect 2027 61 2070 95
rect 2104 61 2147 95
rect 2027 30 2147 61
rect 2177 299 2297 330
rect 2177 265 2220 299
rect 2254 265 2297 299
rect 2177 231 2297 265
rect 2177 197 2220 231
rect 2254 197 2297 231
rect 2177 163 2297 197
rect 2177 129 2220 163
rect 2254 129 2297 163
rect 2177 95 2297 129
rect 2177 61 2220 95
rect 2254 61 2297 95
rect 2177 30 2297 61
rect -2440 -369 -2320 -338
rect -2440 -403 -2397 -369
rect -2363 -403 -2320 -369
rect -2440 -437 -2320 -403
rect -2440 -471 -2397 -437
rect -2363 -471 -2320 -437
rect -2440 -505 -2320 -471
rect -2440 -539 -2397 -505
rect -2363 -539 -2320 -505
rect -2440 -573 -2320 -539
rect -2440 -607 -2397 -573
rect -2363 -607 -2320 -573
rect -2440 -638 -2320 -607
rect -2290 -638 -2170 -338
rect -2140 -369 -2020 -338
rect -2140 -403 -2097 -369
rect -2063 -403 -2020 -369
rect -2140 -437 -2020 -403
rect -2140 -471 -2097 -437
rect -2063 -471 -2020 -437
rect -2140 -505 -2020 -471
rect -2140 -539 -2097 -505
rect -2063 -539 -2020 -505
rect -2140 -573 -2020 -539
rect -2140 -607 -2097 -573
rect -2063 -607 -2020 -573
rect -2140 -638 -2020 -607
rect -1990 -638 -1870 -338
rect -1840 -369 -1720 -338
rect -1840 -403 -1797 -369
rect -1763 -403 -1720 -369
rect -1840 -437 -1720 -403
rect -1840 -471 -1797 -437
rect -1763 -471 -1720 -437
rect -1840 -505 -1720 -471
rect -1840 -539 -1797 -505
rect -1763 -539 -1720 -505
rect -1840 -573 -1720 -539
rect -1840 -607 -1797 -573
rect -1763 -607 -1720 -573
rect -1840 -638 -1720 -607
rect -1589 -369 -1469 -338
rect -1589 -403 -1546 -369
rect -1512 -403 -1469 -369
rect -1589 -437 -1469 -403
rect -1589 -471 -1546 -437
rect -1512 -471 -1469 -437
rect -1589 -505 -1469 -471
rect -1589 -539 -1546 -505
rect -1512 -539 -1469 -505
rect -1589 -573 -1469 -539
rect -1589 -607 -1546 -573
rect -1512 -607 -1469 -573
rect -1589 -638 -1469 -607
rect -1439 -369 -1319 -338
rect -1439 -403 -1396 -369
rect -1362 -403 -1319 -369
rect -1439 -437 -1319 -403
rect -1439 -471 -1396 -437
rect -1362 -471 -1319 -437
rect -1439 -505 -1319 -471
rect -1439 -539 -1396 -505
rect -1362 -539 -1319 -505
rect -1439 -573 -1319 -539
rect -1439 -607 -1396 -573
rect -1362 -607 -1319 -573
rect -1439 -638 -1319 -607
rect -937 -369 -817 -338
rect -937 -403 -894 -369
rect -860 -403 -817 -369
rect -937 -437 -817 -403
rect -937 -471 -894 -437
rect -860 -471 -817 -437
rect -937 -505 -817 -471
rect -937 -539 -894 -505
rect -860 -539 -817 -505
rect -937 -573 -817 -539
rect -937 -607 -894 -573
rect -860 -607 -817 -573
rect -937 -638 -817 -607
rect -787 -638 -667 -338
rect -637 -369 -517 -338
rect -637 -403 -594 -369
rect -560 -403 -517 -369
rect -637 -437 -517 -403
rect -637 -471 -594 -437
rect -560 -471 -517 -437
rect -637 -505 -517 -471
rect -637 -539 -594 -505
rect -560 -539 -517 -505
rect -637 -573 -517 -539
rect -637 -607 -594 -573
rect -560 -607 -517 -573
rect -637 -638 -517 -607
rect -397 -369 -277 -338
rect -397 -403 -354 -369
rect -320 -403 -277 -369
rect -397 -437 -277 -403
rect -397 -471 -354 -437
rect -320 -471 -277 -437
rect -397 -505 -277 -471
rect -397 -539 -354 -505
rect -320 -539 -277 -505
rect -397 -573 -277 -539
rect -397 -607 -354 -573
rect -320 -607 -277 -573
rect -397 -638 -277 -607
rect -247 -369 -127 -338
rect -247 -403 -204 -369
rect -170 -403 -127 -369
rect -247 -437 -127 -403
rect -247 -471 -204 -437
rect -170 -471 -127 -437
rect -247 -505 -127 -471
rect -247 -539 -204 -505
rect -170 -539 -127 -505
rect -247 -573 -127 -539
rect -247 -607 -204 -573
rect -170 -607 -127 -573
rect -247 -638 -127 -607
rect 275 -369 395 -338
rect 275 -403 318 -369
rect 352 -403 395 -369
rect 275 -437 395 -403
rect 275 -471 318 -437
rect 352 -471 395 -437
rect 275 -505 395 -471
rect 275 -539 318 -505
rect 352 -539 395 -505
rect 275 -573 395 -539
rect 275 -607 318 -573
rect 352 -607 395 -573
rect 275 -638 395 -607
rect 425 -638 545 -338
rect 575 -369 695 -338
rect 575 -403 618 -369
rect 652 -403 695 -369
rect 575 -437 695 -403
rect 575 -471 618 -437
rect 652 -471 695 -437
rect 575 -505 695 -471
rect 575 -539 618 -505
rect 652 -539 695 -505
rect 575 -573 695 -539
rect 575 -607 618 -573
rect 652 -607 695 -573
rect 575 -638 695 -607
rect 815 -369 935 -338
rect 815 -403 858 -369
rect 892 -403 935 -369
rect 815 -437 935 -403
rect 815 -471 858 -437
rect 892 -471 935 -437
rect 815 -505 935 -471
rect 815 -539 858 -505
rect 892 -539 935 -505
rect 815 -573 935 -539
rect 815 -607 858 -573
rect 892 -607 935 -573
rect 815 -638 935 -607
rect 965 -369 1085 -338
rect 965 -403 1008 -369
rect 1042 -403 1085 -369
rect 965 -437 1085 -403
rect 965 -471 1008 -437
rect 1042 -471 1085 -437
rect 965 -505 1085 -471
rect 965 -539 1008 -505
rect 1042 -539 1085 -505
rect 965 -573 1085 -539
rect 965 -607 1008 -573
rect 1042 -607 1085 -573
rect 965 -638 1085 -607
<< pdiff >>
rect -2440 1195 -2320 1240
rect -2440 1161 -2397 1195
rect -2363 1161 -2320 1195
rect -2440 1127 -2320 1161
rect -2440 1093 -2397 1127
rect -2363 1093 -2320 1127
rect -2440 1059 -2320 1093
rect -2440 1025 -2397 1059
rect -2363 1025 -2320 1059
rect -2440 991 -2320 1025
rect -2440 957 -2397 991
rect -2363 957 -2320 991
rect -2440 923 -2320 957
rect -2440 889 -2397 923
rect -2363 889 -2320 923
rect -2440 855 -2320 889
rect -2440 821 -2397 855
rect -2363 821 -2320 855
rect -2440 787 -2320 821
rect -2440 753 -2397 787
rect -2363 753 -2320 787
rect -2440 719 -2320 753
rect -2440 685 -2397 719
rect -2363 685 -2320 719
rect -2440 640 -2320 685
rect -2290 640 -2170 1240
rect -2140 1195 -2020 1240
rect -2140 1161 -2097 1195
rect -2063 1161 -2020 1195
rect -2140 1127 -2020 1161
rect -2140 1093 -2097 1127
rect -2063 1093 -2020 1127
rect -2140 1059 -2020 1093
rect -2140 1025 -2097 1059
rect -2063 1025 -2020 1059
rect -2140 991 -2020 1025
rect -2140 957 -2097 991
rect -2063 957 -2020 991
rect -2140 923 -2020 957
rect -2140 889 -2097 923
rect -2063 889 -2020 923
rect -2140 855 -2020 889
rect -2140 821 -2097 855
rect -2063 821 -2020 855
rect -2140 787 -2020 821
rect -2140 753 -2097 787
rect -2063 753 -2020 787
rect -2140 719 -2020 753
rect -2140 685 -2097 719
rect -2063 685 -2020 719
rect -2140 640 -2020 685
rect -1990 640 -1870 1240
rect -1840 1195 -1720 1240
rect -1840 1161 -1797 1195
rect -1763 1161 -1720 1195
rect -1840 1127 -1720 1161
rect -1840 1093 -1797 1127
rect -1763 1093 -1720 1127
rect -1840 1059 -1720 1093
rect -1840 1025 -1797 1059
rect -1763 1025 -1720 1059
rect -1840 991 -1720 1025
rect -1840 957 -1797 991
rect -1763 957 -1720 991
rect -1840 923 -1720 957
rect -1840 889 -1797 923
rect -1763 889 -1720 923
rect -1840 855 -1720 889
rect -1840 821 -1797 855
rect -1763 821 -1720 855
rect -1840 787 -1720 821
rect -1840 753 -1797 787
rect -1763 753 -1720 787
rect -1840 719 -1720 753
rect -1840 685 -1797 719
rect -1763 685 -1720 719
rect -1840 640 -1720 685
rect -937 1195 -817 1240
rect -937 1161 -894 1195
rect -860 1161 -817 1195
rect -937 1127 -817 1161
rect -937 1093 -894 1127
rect -860 1093 -817 1127
rect -937 1059 -817 1093
rect -937 1025 -894 1059
rect -860 1025 -817 1059
rect -937 991 -817 1025
rect -937 957 -894 991
rect -860 957 -817 991
rect -937 923 -817 957
rect -937 889 -894 923
rect -860 889 -817 923
rect -937 855 -817 889
rect -937 821 -894 855
rect -860 821 -817 855
rect -937 787 -817 821
rect -937 753 -894 787
rect -860 753 -817 787
rect -937 719 -817 753
rect -937 685 -894 719
rect -860 685 -817 719
rect -937 640 -817 685
rect -787 640 -667 1240
rect -637 1195 -517 1240
rect -637 1161 -594 1195
rect -560 1161 -517 1195
rect -637 1127 -517 1161
rect -637 1093 -594 1127
rect -560 1093 -517 1127
rect -637 1059 -517 1093
rect -637 1025 -594 1059
rect -560 1025 -517 1059
rect -637 991 -517 1025
rect -637 957 -594 991
rect -560 957 -517 991
rect -637 923 -517 957
rect -637 889 -594 923
rect -560 889 -517 923
rect -637 855 -517 889
rect -637 821 -594 855
rect -560 821 -517 855
rect -637 787 -517 821
rect -637 753 -594 787
rect -560 753 -517 787
rect -637 719 -517 753
rect -637 685 -594 719
rect -560 685 -517 719
rect -637 640 -517 685
rect -397 1195 -277 1240
rect -397 1161 -354 1195
rect -320 1161 -277 1195
rect -397 1127 -277 1161
rect -397 1093 -354 1127
rect -320 1093 -277 1127
rect -397 1059 -277 1093
rect -397 1025 -354 1059
rect -320 1025 -277 1059
rect -397 991 -277 1025
rect -397 957 -354 991
rect -320 957 -277 991
rect -397 923 -277 957
rect -397 889 -354 923
rect -320 889 -277 923
rect -397 855 -277 889
rect -397 821 -354 855
rect -320 821 -277 855
rect -397 787 -277 821
rect -397 753 -354 787
rect -320 753 -277 787
rect -397 719 -277 753
rect -397 685 -354 719
rect -320 685 -277 719
rect -397 640 -277 685
rect -247 1195 -127 1240
rect -247 1161 -204 1195
rect -170 1161 -127 1195
rect -247 1127 -127 1161
rect -247 1093 -204 1127
rect -170 1093 -127 1127
rect -247 1059 -127 1093
rect -247 1025 -204 1059
rect -170 1025 -127 1059
rect -247 991 -127 1025
rect -247 957 -204 991
rect -170 957 -127 991
rect -247 923 -127 957
rect -247 889 -204 923
rect -170 889 -127 923
rect -247 855 -127 889
rect -247 821 -204 855
rect -170 821 -127 855
rect -247 787 -127 821
rect -247 753 -204 787
rect -170 753 -127 787
rect -247 719 -127 753
rect -247 685 -204 719
rect -170 685 -127 719
rect -247 640 -127 685
rect 275 1195 395 1240
rect 275 1161 318 1195
rect 352 1161 395 1195
rect 275 1127 395 1161
rect 275 1093 318 1127
rect 352 1093 395 1127
rect 275 1059 395 1093
rect 275 1025 318 1059
rect 352 1025 395 1059
rect 275 991 395 1025
rect 275 957 318 991
rect 352 957 395 991
rect 275 923 395 957
rect 275 889 318 923
rect 352 889 395 923
rect 275 855 395 889
rect 275 821 318 855
rect 352 821 395 855
rect 275 787 395 821
rect 275 753 318 787
rect 352 753 395 787
rect 275 719 395 753
rect 275 685 318 719
rect 352 685 395 719
rect 275 640 395 685
rect 425 1195 545 1240
rect 425 1161 468 1195
rect 502 1161 545 1195
rect 425 1127 545 1161
rect 425 1093 468 1127
rect 502 1093 545 1127
rect 425 1059 545 1093
rect 425 1025 468 1059
rect 502 1025 545 1059
rect 425 991 545 1025
rect 425 957 468 991
rect 502 957 545 991
rect 425 923 545 957
rect 425 889 468 923
rect 502 889 545 923
rect 425 855 545 889
rect 425 821 468 855
rect 502 821 545 855
rect 425 787 545 821
rect 425 753 468 787
rect 502 753 545 787
rect 425 719 545 753
rect 425 685 468 719
rect 502 685 545 719
rect 425 640 545 685
rect 575 1195 695 1240
rect 575 1161 618 1195
rect 652 1161 695 1195
rect 575 1127 695 1161
rect 575 1093 618 1127
rect 652 1093 695 1127
rect 575 1059 695 1093
rect 575 1025 618 1059
rect 652 1025 695 1059
rect 575 991 695 1025
rect 575 957 618 991
rect 652 957 695 991
rect 575 923 695 957
rect 575 889 618 923
rect 652 889 695 923
rect 575 855 695 889
rect 575 821 618 855
rect 652 821 695 855
rect 575 787 695 821
rect 575 753 618 787
rect 652 753 695 787
rect 575 719 695 753
rect 575 685 618 719
rect 652 685 695 719
rect 575 640 695 685
rect 815 1195 935 1240
rect 815 1161 858 1195
rect 892 1161 935 1195
rect 815 1127 935 1161
rect 815 1093 858 1127
rect 892 1093 935 1127
rect 815 1059 935 1093
rect 815 1025 858 1059
rect 892 1025 935 1059
rect 815 991 935 1025
rect 815 957 858 991
rect 892 957 935 991
rect 815 923 935 957
rect 815 889 858 923
rect 892 889 935 923
rect 815 855 935 889
rect 815 821 858 855
rect 892 821 935 855
rect 815 787 935 821
rect 815 753 858 787
rect 892 753 935 787
rect 815 719 935 753
rect 815 685 858 719
rect 892 685 935 719
rect 815 640 935 685
rect 965 1195 1085 1240
rect 965 1161 1008 1195
rect 1042 1161 1085 1195
rect 965 1127 1085 1161
rect 965 1093 1008 1127
rect 1042 1093 1085 1127
rect 965 1059 1085 1093
rect 965 1025 1008 1059
rect 1042 1025 1085 1059
rect 965 991 1085 1025
rect 965 957 1008 991
rect 1042 957 1085 991
rect 965 923 1085 957
rect 965 889 1008 923
rect 1042 889 1085 923
rect 965 855 1085 889
rect 965 821 1008 855
rect 1042 821 1085 855
rect 965 787 1085 821
rect 965 753 1008 787
rect 1042 753 1085 787
rect 965 719 1085 753
rect 965 685 1008 719
rect 1042 685 1085 719
rect 965 640 1085 685
rect 1487 1195 1607 1240
rect 1487 1161 1530 1195
rect 1564 1161 1607 1195
rect 1487 1127 1607 1161
rect 1487 1093 1530 1127
rect 1564 1093 1607 1127
rect 1487 1059 1607 1093
rect 1487 1025 1530 1059
rect 1564 1025 1607 1059
rect 1487 991 1607 1025
rect 1487 957 1530 991
rect 1564 957 1607 991
rect 1487 923 1607 957
rect 1487 889 1530 923
rect 1564 889 1607 923
rect 1487 855 1607 889
rect 1487 821 1530 855
rect 1564 821 1607 855
rect 1487 787 1607 821
rect 1487 753 1530 787
rect 1564 753 1607 787
rect 1487 719 1607 753
rect 1487 685 1530 719
rect 1564 685 1607 719
rect 1487 640 1607 685
rect 1637 640 1757 1240
rect 1787 1195 1907 1240
rect 1787 1161 1830 1195
rect 1864 1161 1907 1195
rect 1787 1127 1907 1161
rect 1787 1093 1830 1127
rect 1864 1093 1907 1127
rect 1787 1059 1907 1093
rect 1787 1025 1830 1059
rect 1864 1025 1907 1059
rect 1787 991 1907 1025
rect 1787 957 1830 991
rect 1864 957 1907 991
rect 1787 923 1907 957
rect 1787 889 1830 923
rect 1864 889 1907 923
rect 1787 855 1907 889
rect 1787 821 1830 855
rect 1864 821 1907 855
rect 1787 787 1907 821
rect 1787 753 1830 787
rect 1864 753 1907 787
rect 1787 719 1907 753
rect 1787 685 1830 719
rect 1864 685 1907 719
rect 1787 640 1907 685
rect 2027 1195 2147 1240
rect 2027 1161 2070 1195
rect 2104 1161 2147 1195
rect 2027 1127 2147 1161
rect 2027 1093 2070 1127
rect 2104 1093 2147 1127
rect 2027 1059 2147 1093
rect 2027 1025 2070 1059
rect 2104 1025 2147 1059
rect 2027 991 2147 1025
rect 2027 957 2070 991
rect 2104 957 2147 991
rect 2027 923 2147 957
rect 2027 889 2070 923
rect 2104 889 2147 923
rect 2027 855 2147 889
rect 2027 821 2070 855
rect 2104 821 2147 855
rect 2027 787 2147 821
rect 2027 753 2070 787
rect 2104 753 2147 787
rect 2027 719 2147 753
rect 2027 685 2070 719
rect 2104 685 2147 719
rect 2027 640 2147 685
rect 2177 1195 2297 1240
rect 2177 1161 2220 1195
rect 2254 1161 2297 1195
rect 2177 1127 2297 1161
rect 2177 1093 2220 1127
rect 2254 1093 2297 1127
rect 2177 1059 2297 1093
rect 2177 1025 2220 1059
rect 2254 1025 2297 1059
rect 2177 991 2297 1025
rect 2177 957 2220 991
rect 2254 957 2297 991
rect 2177 923 2297 957
rect 2177 889 2220 923
rect 2254 889 2297 923
rect 2177 855 2297 889
rect 2177 821 2220 855
rect 2254 821 2297 855
rect 2177 787 2297 821
rect 2177 753 2220 787
rect 2254 753 2297 787
rect 2177 719 2297 753
rect 2177 685 2220 719
rect 2254 685 2297 719
rect 2177 640 2297 685
rect -2440 -993 -2320 -948
rect -2440 -1027 -2397 -993
rect -2363 -1027 -2320 -993
rect -2440 -1061 -2320 -1027
rect -2440 -1095 -2397 -1061
rect -2363 -1095 -2320 -1061
rect -2440 -1129 -2320 -1095
rect -2440 -1163 -2397 -1129
rect -2363 -1163 -2320 -1129
rect -2440 -1197 -2320 -1163
rect -2440 -1231 -2397 -1197
rect -2363 -1231 -2320 -1197
rect -2440 -1265 -2320 -1231
rect -2440 -1299 -2397 -1265
rect -2363 -1299 -2320 -1265
rect -2440 -1333 -2320 -1299
rect -2440 -1367 -2397 -1333
rect -2363 -1367 -2320 -1333
rect -2440 -1401 -2320 -1367
rect -2440 -1435 -2397 -1401
rect -2363 -1435 -2320 -1401
rect -2440 -1469 -2320 -1435
rect -2440 -1503 -2397 -1469
rect -2363 -1503 -2320 -1469
rect -2440 -1548 -2320 -1503
rect -2290 -1548 -2170 -948
rect -2140 -993 -2020 -948
rect -2140 -1027 -2097 -993
rect -2063 -1027 -2020 -993
rect -2140 -1061 -2020 -1027
rect -2140 -1095 -2097 -1061
rect -2063 -1095 -2020 -1061
rect -2140 -1129 -2020 -1095
rect -2140 -1163 -2097 -1129
rect -2063 -1163 -2020 -1129
rect -2140 -1197 -2020 -1163
rect -2140 -1231 -2097 -1197
rect -2063 -1231 -2020 -1197
rect -2140 -1265 -2020 -1231
rect -2140 -1299 -2097 -1265
rect -2063 -1299 -2020 -1265
rect -2140 -1333 -2020 -1299
rect -2140 -1367 -2097 -1333
rect -2063 -1367 -2020 -1333
rect -2140 -1401 -2020 -1367
rect -2140 -1435 -2097 -1401
rect -2063 -1435 -2020 -1401
rect -2140 -1469 -2020 -1435
rect -2140 -1503 -2097 -1469
rect -2063 -1503 -2020 -1469
rect -2140 -1548 -2020 -1503
rect -1990 -1548 -1870 -948
rect -1840 -993 -1720 -948
rect -1840 -1027 -1797 -993
rect -1763 -1027 -1720 -993
rect -1840 -1061 -1720 -1027
rect -1840 -1095 -1797 -1061
rect -1763 -1095 -1720 -1061
rect -1840 -1129 -1720 -1095
rect -1840 -1163 -1797 -1129
rect -1763 -1163 -1720 -1129
rect -1840 -1197 -1720 -1163
rect -1840 -1231 -1797 -1197
rect -1763 -1231 -1720 -1197
rect -1840 -1265 -1720 -1231
rect -1840 -1299 -1797 -1265
rect -1763 -1299 -1720 -1265
rect -1840 -1333 -1720 -1299
rect -1840 -1367 -1797 -1333
rect -1763 -1367 -1720 -1333
rect -1840 -1401 -1720 -1367
rect -1840 -1435 -1797 -1401
rect -1763 -1435 -1720 -1401
rect -1840 -1469 -1720 -1435
rect -1840 -1503 -1797 -1469
rect -1763 -1503 -1720 -1469
rect -1840 -1548 -1720 -1503
rect -1589 -993 -1469 -948
rect -1589 -1027 -1546 -993
rect -1512 -1027 -1469 -993
rect -1589 -1061 -1469 -1027
rect -1589 -1095 -1546 -1061
rect -1512 -1095 -1469 -1061
rect -1589 -1129 -1469 -1095
rect -1589 -1163 -1546 -1129
rect -1512 -1163 -1469 -1129
rect -1589 -1197 -1469 -1163
rect -1589 -1231 -1546 -1197
rect -1512 -1231 -1469 -1197
rect -1589 -1265 -1469 -1231
rect -1589 -1299 -1546 -1265
rect -1512 -1299 -1469 -1265
rect -1589 -1333 -1469 -1299
rect -1589 -1367 -1546 -1333
rect -1512 -1367 -1469 -1333
rect -1589 -1401 -1469 -1367
rect -1589 -1435 -1546 -1401
rect -1512 -1435 -1469 -1401
rect -1589 -1469 -1469 -1435
rect -1589 -1503 -1546 -1469
rect -1512 -1503 -1469 -1469
rect -1589 -1548 -1469 -1503
rect -1439 -993 -1319 -948
rect -1439 -1027 -1396 -993
rect -1362 -1027 -1319 -993
rect -1439 -1061 -1319 -1027
rect -1439 -1095 -1396 -1061
rect -1362 -1095 -1319 -1061
rect -1439 -1129 -1319 -1095
rect -1439 -1163 -1396 -1129
rect -1362 -1163 -1319 -1129
rect -1439 -1197 -1319 -1163
rect -1439 -1231 -1396 -1197
rect -1362 -1231 -1319 -1197
rect -1439 -1265 -1319 -1231
rect -1439 -1299 -1396 -1265
rect -1362 -1299 -1319 -1265
rect -1439 -1333 -1319 -1299
rect -1439 -1367 -1396 -1333
rect -1362 -1367 -1319 -1333
rect -1439 -1401 -1319 -1367
rect -1439 -1435 -1396 -1401
rect -1362 -1435 -1319 -1401
rect -1439 -1469 -1319 -1435
rect -1439 -1503 -1396 -1469
rect -1362 -1503 -1319 -1469
rect -1439 -1548 -1319 -1503
rect -937 -993 -817 -948
rect -937 -1027 -894 -993
rect -860 -1027 -817 -993
rect -937 -1061 -817 -1027
rect -937 -1095 -894 -1061
rect -860 -1095 -817 -1061
rect -937 -1129 -817 -1095
rect -937 -1163 -894 -1129
rect -860 -1163 -817 -1129
rect -937 -1197 -817 -1163
rect -937 -1231 -894 -1197
rect -860 -1231 -817 -1197
rect -937 -1265 -817 -1231
rect -937 -1299 -894 -1265
rect -860 -1299 -817 -1265
rect -937 -1333 -817 -1299
rect -937 -1367 -894 -1333
rect -860 -1367 -817 -1333
rect -937 -1401 -817 -1367
rect -937 -1435 -894 -1401
rect -860 -1435 -817 -1401
rect -937 -1469 -817 -1435
rect -937 -1503 -894 -1469
rect -860 -1503 -817 -1469
rect -937 -1548 -817 -1503
rect -787 -993 -667 -948
rect -787 -1027 -744 -993
rect -710 -1027 -667 -993
rect -787 -1061 -667 -1027
rect -787 -1095 -744 -1061
rect -710 -1095 -667 -1061
rect -787 -1129 -667 -1095
rect -787 -1163 -744 -1129
rect -710 -1163 -667 -1129
rect -787 -1197 -667 -1163
rect -787 -1231 -744 -1197
rect -710 -1231 -667 -1197
rect -787 -1265 -667 -1231
rect -787 -1299 -744 -1265
rect -710 -1299 -667 -1265
rect -787 -1333 -667 -1299
rect -787 -1367 -744 -1333
rect -710 -1367 -667 -1333
rect -787 -1401 -667 -1367
rect -787 -1435 -744 -1401
rect -710 -1435 -667 -1401
rect -787 -1469 -667 -1435
rect -787 -1503 -744 -1469
rect -710 -1503 -667 -1469
rect -787 -1548 -667 -1503
rect -637 -993 -517 -948
rect -637 -1027 -594 -993
rect -560 -1027 -517 -993
rect -637 -1061 -517 -1027
rect -637 -1095 -594 -1061
rect -560 -1095 -517 -1061
rect -637 -1129 -517 -1095
rect -637 -1163 -594 -1129
rect -560 -1163 -517 -1129
rect -637 -1197 -517 -1163
rect -637 -1231 -594 -1197
rect -560 -1231 -517 -1197
rect -637 -1265 -517 -1231
rect -637 -1299 -594 -1265
rect -560 -1299 -517 -1265
rect -637 -1333 -517 -1299
rect -637 -1367 -594 -1333
rect -560 -1367 -517 -1333
rect -637 -1401 -517 -1367
rect -637 -1435 -594 -1401
rect -560 -1435 -517 -1401
rect -637 -1469 -517 -1435
rect -637 -1503 -594 -1469
rect -560 -1503 -517 -1469
rect -637 -1548 -517 -1503
rect -397 -993 -277 -948
rect -397 -1027 -354 -993
rect -320 -1027 -277 -993
rect -397 -1061 -277 -1027
rect -397 -1095 -354 -1061
rect -320 -1095 -277 -1061
rect -397 -1129 -277 -1095
rect -397 -1163 -354 -1129
rect -320 -1163 -277 -1129
rect -397 -1197 -277 -1163
rect -397 -1231 -354 -1197
rect -320 -1231 -277 -1197
rect -397 -1265 -277 -1231
rect -397 -1299 -354 -1265
rect -320 -1299 -277 -1265
rect -397 -1333 -277 -1299
rect -397 -1367 -354 -1333
rect -320 -1367 -277 -1333
rect -397 -1401 -277 -1367
rect -397 -1435 -354 -1401
rect -320 -1435 -277 -1401
rect -397 -1469 -277 -1435
rect -397 -1503 -354 -1469
rect -320 -1503 -277 -1469
rect -397 -1548 -277 -1503
rect -247 -993 -127 -948
rect -247 -1027 -204 -993
rect -170 -1027 -127 -993
rect -247 -1061 -127 -1027
rect -247 -1095 -204 -1061
rect -170 -1095 -127 -1061
rect -247 -1129 -127 -1095
rect -247 -1163 -204 -1129
rect -170 -1163 -127 -1129
rect -247 -1197 -127 -1163
rect -247 -1231 -204 -1197
rect -170 -1231 -127 -1197
rect -247 -1265 -127 -1231
rect -247 -1299 -204 -1265
rect -170 -1299 -127 -1265
rect -247 -1333 -127 -1299
rect -247 -1367 -204 -1333
rect -170 -1367 -127 -1333
rect -247 -1401 -127 -1367
rect -247 -1435 -204 -1401
rect -170 -1435 -127 -1401
rect -247 -1469 -127 -1435
rect -247 -1503 -204 -1469
rect -170 -1503 -127 -1469
rect -247 -1548 -127 -1503
rect 275 -993 395 -948
rect 275 -1027 318 -993
rect 352 -1027 395 -993
rect 275 -1061 395 -1027
rect 275 -1095 318 -1061
rect 352 -1095 395 -1061
rect 275 -1129 395 -1095
rect 275 -1163 318 -1129
rect 352 -1163 395 -1129
rect 275 -1197 395 -1163
rect 275 -1231 318 -1197
rect 352 -1231 395 -1197
rect 275 -1265 395 -1231
rect 275 -1299 318 -1265
rect 352 -1299 395 -1265
rect 275 -1333 395 -1299
rect 275 -1367 318 -1333
rect 352 -1367 395 -1333
rect 275 -1401 395 -1367
rect 275 -1435 318 -1401
rect 352 -1435 395 -1401
rect 275 -1469 395 -1435
rect 275 -1503 318 -1469
rect 352 -1503 395 -1469
rect 275 -1548 395 -1503
rect 425 -993 545 -948
rect 425 -1027 468 -993
rect 502 -1027 545 -993
rect 425 -1061 545 -1027
rect 425 -1095 468 -1061
rect 502 -1095 545 -1061
rect 425 -1129 545 -1095
rect 425 -1163 468 -1129
rect 502 -1163 545 -1129
rect 425 -1197 545 -1163
rect 425 -1231 468 -1197
rect 502 -1231 545 -1197
rect 425 -1265 545 -1231
rect 425 -1299 468 -1265
rect 502 -1299 545 -1265
rect 425 -1333 545 -1299
rect 425 -1367 468 -1333
rect 502 -1367 545 -1333
rect 425 -1401 545 -1367
rect 425 -1435 468 -1401
rect 502 -1435 545 -1401
rect 425 -1469 545 -1435
rect 425 -1503 468 -1469
rect 502 -1503 545 -1469
rect 425 -1548 545 -1503
rect 575 -993 695 -948
rect 575 -1027 618 -993
rect 652 -1027 695 -993
rect 575 -1061 695 -1027
rect 575 -1095 618 -1061
rect 652 -1095 695 -1061
rect 575 -1129 695 -1095
rect 575 -1163 618 -1129
rect 652 -1163 695 -1129
rect 575 -1197 695 -1163
rect 575 -1231 618 -1197
rect 652 -1231 695 -1197
rect 575 -1265 695 -1231
rect 575 -1299 618 -1265
rect 652 -1299 695 -1265
rect 575 -1333 695 -1299
rect 575 -1367 618 -1333
rect 652 -1367 695 -1333
rect 575 -1401 695 -1367
rect 575 -1435 618 -1401
rect 652 -1435 695 -1401
rect 575 -1469 695 -1435
rect 575 -1503 618 -1469
rect 652 -1503 695 -1469
rect 575 -1548 695 -1503
rect 815 -993 935 -948
rect 815 -1027 858 -993
rect 892 -1027 935 -993
rect 815 -1061 935 -1027
rect 815 -1095 858 -1061
rect 892 -1095 935 -1061
rect 815 -1129 935 -1095
rect 815 -1163 858 -1129
rect 892 -1163 935 -1129
rect 815 -1197 935 -1163
rect 815 -1231 858 -1197
rect 892 -1231 935 -1197
rect 815 -1265 935 -1231
rect 815 -1299 858 -1265
rect 892 -1299 935 -1265
rect 815 -1333 935 -1299
rect 815 -1367 858 -1333
rect 892 -1367 935 -1333
rect 815 -1401 935 -1367
rect 815 -1435 858 -1401
rect 892 -1435 935 -1401
rect 815 -1469 935 -1435
rect 815 -1503 858 -1469
rect 892 -1503 935 -1469
rect 815 -1548 935 -1503
rect 965 -993 1085 -948
rect 965 -1027 1008 -993
rect 1042 -1027 1085 -993
rect 965 -1061 1085 -1027
rect 965 -1095 1008 -1061
rect 1042 -1095 1085 -1061
rect 965 -1129 1085 -1095
rect 965 -1163 1008 -1129
rect 1042 -1163 1085 -1129
rect 965 -1197 1085 -1163
rect 965 -1231 1008 -1197
rect 1042 -1231 1085 -1197
rect 965 -1265 1085 -1231
rect 965 -1299 1008 -1265
rect 1042 -1299 1085 -1265
rect 965 -1333 1085 -1299
rect 965 -1367 1008 -1333
rect 1042 -1367 1085 -1333
rect 965 -1401 1085 -1367
rect 965 -1435 1008 -1401
rect 1042 -1435 1085 -1401
rect 965 -1469 1085 -1435
rect 965 -1503 1008 -1469
rect 1042 -1503 1085 -1469
rect 965 -1548 1085 -1503
<< ndiffc >>
rect -2397 265 -2363 299
rect -2397 197 -2363 231
rect -2397 129 -2363 163
rect -2397 61 -2363 95
rect -2097 265 -2063 299
rect -2097 197 -2063 231
rect -2097 129 -2063 163
rect -2097 61 -2063 95
rect -1797 265 -1763 299
rect -1797 197 -1763 231
rect -1797 129 -1763 163
rect -1797 61 -1763 95
rect -894 265 -860 299
rect -894 197 -860 231
rect -894 129 -860 163
rect -894 61 -860 95
rect -744 265 -710 299
rect -744 197 -710 231
rect -744 129 -710 163
rect -744 61 -710 95
rect -594 265 -560 299
rect -594 197 -560 231
rect -594 129 -560 163
rect -594 61 -560 95
rect -354 265 -320 299
rect -354 197 -320 231
rect -354 129 -320 163
rect -354 61 -320 95
rect -204 265 -170 299
rect -204 197 -170 231
rect -204 129 -170 163
rect -204 61 -170 95
rect 318 265 352 299
rect 318 197 352 231
rect 318 129 352 163
rect 318 61 352 95
rect 618 265 652 299
rect 618 197 652 231
rect 618 129 652 163
rect 618 61 652 95
rect 858 265 892 299
rect 858 197 892 231
rect 858 129 892 163
rect 858 61 892 95
rect 1008 265 1042 299
rect 1008 197 1042 231
rect 1008 129 1042 163
rect 1008 61 1042 95
rect 1530 265 1564 299
rect 1530 197 1564 231
rect 1530 129 1564 163
rect 1530 61 1564 95
rect 1680 265 1714 299
rect 1680 197 1714 231
rect 1680 129 1714 163
rect 1680 61 1714 95
rect 1830 265 1864 299
rect 1830 197 1864 231
rect 1830 129 1864 163
rect 1830 61 1864 95
rect 2070 265 2104 299
rect 2070 197 2104 231
rect 2070 129 2104 163
rect 2070 61 2104 95
rect 2220 265 2254 299
rect 2220 197 2254 231
rect 2220 129 2254 163
rect 2220 61 2254 95
rect -2397 -403 -2363 -369
rect -2397 -471 -2363 -437
rect -2397 -539 -2363 -505
rect -2397 -607 -2363 -573
rect -2097 -403 -2063 -369
rect -2097 -471 -2063 -437
rect -2097 -539 -2063 -505
rect -2097 -607 -2063 -573
rect -1797 -403 -1763 -369
rect -1797 -471 -1763 -437
rect -1797 -539 -1763 -505
rect -1797 -607 -1763 -573
rect -1546 -403 -1512 -369
rect -1546 -471 -1512 -437
rect -1546 -539 -1512 -505
rect -1546 -607 -1512 -573
rect -1396 -403 -1362 -369
rect -1396 -471 -1362 -437
rect -1396 -539 -1362 -505
rect -1396 -607 -1362 -573
rect -894 -403 -860 -369
rect -894 -471 -860 -437
rect -894 -539 -860 -505
rect -894 -607 -860 -573
rect -594 -403 -560 -369
rect -594 -471 -560 -437
rect -594 -539 -560 -505
rect -594 -607 -560 -573
rect -354 -403 -320 -369
rect -354 -471 -320 -437
rect -354 -539 -320 -505
rect -354 -607 -320 -573
rect -204 -403 -170 -369
rect -204 -471 -170 -437
rect -204 -539 -170 -505
rect -204 -607 -170 -573
rect 318 -403 352 -369
rect 318 -471 352 -437
rect 318 -539 352 -505
rect 318 -607 352 -573
rect 618 -403 652 -369
rect 618 -471 652 -437
rect 618 -539 652 -505
rect 618 -607 652 -573
rect 858 -403 892 -369
rect 858 -471 892 -437
rect 858 -539 892 -505
rect 858 -607 892 -573
rect 1008 -403 1042 -369
rect 1008 -471 1042 -437
rect 1008 -539 1042 -505
rect 1008 -607 1042 -573
<< pdiffc >>
rect -2397 1161 -2363 1195
rect -2397 1093 -2363 1127
rect -2397 1025 -2363 1059
rect -2397 957 -2363 991
rect -2397 889 -2363 923
rect -2397 821 -2363 855
rect -2397 753 -2363 787
rect -2397 685 -2363 719
rect -2097 1161 -2063 1195
rect -2097 1093 -2063 1127
rect -2097 1025 -2063 1059
rect -2097 957 -2063 991
rect -2097 889 -2063 923
rect -2097 821 -2063 855
rect -2097 753 -2063 787
rect -2097 685 -2063 719
rect -1797 1161 -1763 1195
rect -1797 1093 -1763 1127
rect -1797 1025 -1763 1059
rect -1797 957 -1763 991
rect -1797 889 -1763 923
rect -1797 821 -1763 855
rect -1797 753 -1763 787
rect -1797 685 -1763 719
rect -894 1161 -860 1195
rect -894 1093 -860 1127
rect -894 1025 -860 1059
rect -894 957 -860 991
rect -894 889 -860 923
rect -894 821 -860 855
rect -894 753 -860 787
rect -894 685 -860 719
rect -594 1161 -560 1195
rect -594 1093 -560 1127
rect -594 1025 -560 1059
rect -594 957 -560 991
rect -594 889 -560 923
rect -594 821 -560 855
rect -594 753 -560 787
rect -594 685 -560 719
rect -354 1161 -320 1195
rect -354 1093 -320 1127
rect -354 1025 -320 1059
rect -354 957 -320 991
rect -354 889 -320 923
rect -354 821 -320 855
rect -354 753 -320 787
rect -354 685 -320 719
rect -204 1161 -170 1195
rect -204 1093 -170 1127
rect -204 1025 -170 1059
rect -204 957 -170 991
rect -204 889 -170 923
rect -204 821 -170 855
rect -204 753 -170 787
rect -204 685 -170 719
rect 318 1161 352 1195
rect 318 1093 352 1127
rect 318 1025 352 1059
rect 318 957 352 991
rect 318 889 352 923
rect 318 821 352 855
rect 318 753 352 787
rect 318 685 352 719
rect 468 1161 502 1195
rect 468 1093 502 1127
rect 468 1025 502 1059
rect 468 957 502 991
rect 468 889 502 923
rect 468 821 502 855
rect 468 753 502 787
rect 468 685 502 719
rect 618 1161 652 1195
rect 618 1093 652 1127
rect 618 1025 652 1059
rect 618 957 652 991
rect 618 889 652 923
rect 618 821 652 855
rect 618 753 652 787
rect 618 685 652 719
rect 858 1161 892 1195
rect 858 1093 892 1127
rect 858 1025 892 1059
rect 858 957 892 991
rect 858 889 892 923
rect 858 821 892 855
rect 858 753 892 787
rect 858 685 892 719
rect 1008 1161 1042 1195
rect 1008 1093 1042 1127
rect 1008 1025 1042 1059
rect 1008 957 1042 991
rect 1008 889 1042 923
rect 1008 821 1042 855
rect 1008 753 1042 787
rect 1008 685 1042 719
rect 1530 1161 1564 1195
rect 1530 1093 1564 1127
rect 1530 1025 1564 1059
rect 1530 957 1564 991
rect 1530 889 1564 923
rect 1530 821 1564 855
rect 1530 753 1564 787
rect 1530 685 1564 719
rect 1830 1161 1864 1195
rect 1830 1093 1864 1127
rect 1830 1025 1864 1059
rect 1830 957 1864 991
rect 1830 889 1864 923
rect 1830 821 1864 855
rect 1830 753 1864 787
rect 1830 685 1864 719
rect 2070 1161 2104 1195
rect 2070 1093 2104 1127
rect 2070 1025 2104 1059
rect 2070 957 2104 991
rect 2070 889 2104 923
rect 2070 821 2104 855
rect 2070 753 2104 787
rect 2070 685 2104 719
rect 2220 1161 2254 1195
rect 2220 1093 2254 1127
rect 2220 1025 2254 1059
rect 2220 957 2254 991
rect 2220 889 2254 923
rect 2220 821 2254 855
rect 2220 753 2254 787
rect 2220 685 2254 719
rect -2397 -1027 -2363 -993
rect -2397 -1095 -2363 -1061
rect -2397 -1163 -2363 -1129
rect -2397 -1231 -2363 -1197
rect -2397 -1299 -2363 -1265
rect -2397 -1367 -2363 -1333
rect -2397 -1435 -2363 -1401
rect -2397 -1503 -2363 -1469
rect -2097 -1027 -2063 -993
rect -2097 -1095 -2063 -1061
rect -2097 -1163 -2063 -1129
rect -2097 -1231 -2063 -1197
rect -2097 -1299 -2063 -1265
rect -2097 -1367 -2063 -1333
rect -2097 -1435 -2063 -1401
rect -2097 -1503 -2063 -1469
rect -1797 -1027 -1763 -993
rect -1797 -1095 -1763 -1061
rect -1797 -1163 -1763 -1129
rect -1797 -1231 -1763 -1197
rect -1797 -1299 -1763 -1265
rect -1797 -1367 -1763 -1333
rect -1797 -1435 -1763 -1401
rect -1797 -1503 -1763 -1469
rect -1546 -1027 -1512 -993
rect -1546 -1095 -1512 -1061
rect -1546 -1163 -1512 -1129
rect -1546 -1231 -1512 -1197
rect -1546 -1299 -1512 -1265
rect -1546 -1367 -1512 -1333
rect -1546 -1435 -1512 -1401
rect -1546 -1503 -1512 -1469
rect -1396 -1027 -1362 -993
rect -1396 -1095 -1362 -1061
rect -1396 -1163 -1362 -1129
rect -1396 -1231 -1362 -1197
rect -1396 -1299 -1362 -1265
rect -1396 -1367 -1362 -1333
rect -1396 -1435 -1362 -1401
rect -1396 -1503 -1362 -1469
rect -894 -1027 -860 -993
rect -894 -1095 -860 -1061
rect -894 -1163 -860 -1129
rect -894 -1231 -860 -1197
rect -894 -1299 -860 -1265
rect -894 -1367 -860 -1333
rect -894 -1435 -860 -1401
rect -894 -1503 -860 -1469
rect -744 -1027 -710 -993
rect -744 -1095 -710 -1061
rect -744 -1163 -710 -1129
rect -744 -1231 -710 -1197
rect -744 -1299 -710 -1265
rect -744 -1367 -710 -1333
rect -744 -1435 -710 -1401
rect -744 -1503 -710 -1469
rect -594 -1027 -560 -993
rect -594 -1095 -560 -1061
rect -594 -1163 -560 -1129
rect -594 -1231 -560 -1197
rect -594 -1299 -560 -1265
rect -594 -1367 -560 -1333
rect -594 -1435 -560 -1401
rect -594 -1503 -560 -1469
rect -354 -1027 -320 -993
rect -354 -1095 -320 -1061
rect -354 -1163 -320 -1129
rect -354 -1231 -320 -1197
rect -354 -1299 -320 -1265
rect -354 -1367 -320 -1333
rect -354 -1435 -320 -1401
rect -354 -1503 -320 -1469
rect -204 -1027 -170 -993
rect -204 -1095 -170 -1061
rect -204 -1163 -170 -1129
rect -204 -1231 -170 -1197
rect -204 -1299 -170 -1265
rect -204 -1367 -170 -1333
rect -204 -1435 -170 -1401
rect -204 -1503 -170 -1469
rect 318 -1027 352 -993
rect 318 -1095 352 -1061
rect 318 -1163 352 -1129
rect 318 -1231 352 -1197
rect 318 -1299 352 -1265
rect 318 -1367 352 -1333
rect 318 -1435 352 -1401
rect 318 -1503 352 -1469
rect 468 -1027 502 -993
rect 468 -1095 502 -1061
rect 468 -1163 502 -1129
rect 468 -1231 502 -1197
rect 468 -1299 502 -1265
rect 468 -1367 502 -1333
rect 468 -1435 502 -1401
rect 468 -1503 502 -1469
rect 618 -1027 652 -993
rect 618 -1095 652 -1061
rect 618 -1163 652 -1129
rect 618 -1231 652 -1197
rect 618 -1299 652 -1265
rect 618 -1367 652 -1333
rect 618 -1435 652 -1401
rect 618 -1503 652 -1469
rect 858 -1027 892 -993
rect 858 -1095 892 -1061
rect 858 -1163 892 -1129
rect 858 -1231 892 -1197
rect 858 -1299 892 -1265
rect 858 -1367 892 -1333
rect 858 -1435 892 -1401
rect 858 -1503 892 -1469
rect 1008 -1027 1042 -993
rect 1008 -1095 1042 -1061
rect 1008 -1163 1042 -1129
rect 1008 -1231 1042 -1197
rect 1008 -1299 1042 -1265
rect 1008 -1367 1042 -1333
rect 1008 -1435 1042 -1401
rect 1008 -1503 1042 -1469
<< psubdiff >>
rect -2520 -137 -1283 -104
rect -2520 -171 -2497 -137
rect -2463 -171 -2425 -137
rect -2391 -171 -2353 -137
rect -2319 -171 -2281 -137
rect -2247 -171 -2209 -137
rect -2175 -171 -2137 -137
rect -2103 -171 -2065 -137
rect -2031 -171 -1993 -137
rect -1959 -171 -1921 -137
rect -1887 -171 -1849 -137
rect -1815 -171 -1777 -137
rect -1743 -171 -1705 -137
rect -1671 -171 -1633 -137
rect -1599 -171 -1561 -137
rect -1527 -171 -1489 -137
rect -1455 -171 -1417 -137
rect -1383 -171 -1345 -137
rect -1311 -171 -1283 -137
rect -2520 -204 -1283 -171
rect -962 -137 -82 -104
rect -962 -171 -939 -137
rect -905 -171 -867 -137
rect -833 -171 -795 -137
rect -761 -171 -723 -137
rect -689 -171 -651 -137
rect -617 -171 -579 -137
rect -545 -171 -507 -137
rect -473 -171 -435 -137
rect -401 -171 -363 -137
rect -329 -171 -291 -137
rect -257 -171 -219 -137
rect -185 -171 -147 -137
rect -113 -171 -82 -137
rect -962 -204 -82 -171
rect 250 -137 1130 -104
rect 250 -171 273 -137
rect 307 -171 345 -137
rect 379 -171 417 -137
rect 451 -171 489 -137
rect 523 -171 561 -137
rect 595 -171 633 -137
rect 667 -171 705 -137
rect 739 -171 777 -137
rect 811 -171 849 -137
rect 883 -171 921 -137
rect 955 -171 993 -137
rect 1027 -171 1065 -137
rect 1099 -171 1130 -137
rect 250 -204 1130 -171
rect 1462 -137 2342 -104
rect 1462 -171 1485 -137
rect 1519 -171 1557 -137
rect 1591 -171 1629 -137
rect 1663 -171 1701 -137
rect 1735 -171 1773 -137
rect 1807 -171 1845 -137
rect 1879 -171 1917 -137
rect 1951 -171 1989 -137
rect 2023 -171 2061 -137
rect 2095 -171 2133 -137
rect 2167 -171 2205 -137
rect 2239 -171 2277 -137
rect 2311 -171 2342 -137
rect 1462 -204 2342 -171
<< nsubdiff >>
rect -2520 1441 -1640 1474
rect -2520 1407 -2497 1441
rect -2463 1407 -2425 1441
rect -2391 1407 -2353 1441
rect -2319 1407 -2281 1441
rect -2247 1407 -2209 1441
rect -2175 1407 -2137 1441
rect -2103 1407 -2065 1441
rect -2031 1407 -1993 1441
rect -1959 1407 -1921 1441
rect -1887 1407 -1849 1441
rect -1815 1407 -1777 1441
rect -1743 1407 -1705 1441
rect -1671 1407 -1640 1441
rect -2520 1374 -1640 1407
rect -962 1441 -82 1474
rect -962 1407 -939 1441
rect -905 1407 -867 1441
rect -833 1407 -795 1441
rect -761 1407 -723 1441
rect -689 1407 -651 1441
rect -617 1407 -579 1441
rect -545 1407 -507 1441
rect -473 1407 -435 1441
rect -401 1407 -363 1441
rect -329 1407 -291 1441
rect -257 1407 -219 1441
rect -185 1407 -147 1441
rect -113 1407 -82 1441
rect -962 1374 -82 1407
rect 250 1441 1130 1474
rect 250 1407 273 1441
rect 307 1407 345 1441
rect 379 1407 417 1441
rect 451 1407 489 1441
rect 523 1407 561 1441
rect 595 1407 633 1441
rect 667 1407 705 1441
rect 739 1407 777 1441
rect 811 1407 849 1441
rect 883 1407 921 1441
rect 955 1407 993 1441
rect 1027 1407 1065 1441
rect 1099 1407 1130 1441
rect 250 1374 1130 1407
rect 1462 1441 2342 1474
rect 1462 1407 1485 1441
rect 1519 1407 1557 1441
rect 1591 1407 1629 1441
rect 1663 1407 1701 1441
rect 1735 1407 1773 1441
rect 1807 1407 1845 1441
rect 1879 1407 1917 1441
rect 1951 1407 1989 1441
rect 2023 1407 2061 1441
rect 2095 1407 2133 1441
rect 2167 1407 2205 1441
rect 2239 1407 2277 1441
rect 2311 1407 2342 1441
rect 1462 1374 2342 1407
rect -2520 -1715 -1294 -1682
rect -2520 -1749 -2497 -1715
rect -2463 -1749 -2425 -1715
rect -2391 -1749 -2353 -1715
rect -2319 -1749 -2281 -1715
rect -2247 -1749 -2209 -1715
rect -2175 -1749 -2137 -1715
rect -2103 -1749 -2065 -1715
rect -2031 -1749 -1993 -1715
rect -1959 -1749 -1921 -1715
rect -1887 -1749 -1849 -1715
rect -1815 -1749 -1777 -1715
rect -1743 -1749 -1705 -1715
rect -1671 -1749 -1633 -1715
rect -1599 -1749 -1561 -1715
rect -1527 -1749 -1489 -1715
rect -1455 -1749 -1417 -1715
rect -1383 -1749 -1345 -1715
rect -1311 -1749 -1294 -1715
rect -2520 -1782 -1294 -1749
rect -962 -1715 -82 -1682
rect -962 -1749 -939 -1715
rect -905 -1749 -867 -1715
rect -833 -1749 -795 -1715
rect -761 -1749 -723 -1715
rect -689 -1749 -651 -1715
rect -617 -1749 -579 -1715
rect -545 -1749 -507 -1715
rect -473 -1749 -435 -1715
rect -401 -1749 -363 -1715
rect -329 -1749 -291 -1715
rect -257 -1749 -219 -1715
rect -185 -1749 -147 -1715
rect -113 -1749 -82 -1715
rect -962 -1782 -82 -1749
rect 250 -1715 1130 -1682
rect 250 -1749 273 -1715
rect 307 -1749 345 -1715
rect 379 -1749 417 -1715
rect 451 -1749 489 -1715
rect 523 -1749 561 -1715
rect 595 -1749 633 -1715
rect 667 -1749 705 -1715
rect 739 -1749 777 -1715
rect 811 -1749 849 -1715
rect 883 -1749 921 -1715
rect 955 -1749 993 -1715
rect 1027 -1749 1065 -1715
rect 1099 -1749 1130 -1715
rect 250 -1782 1130 -1749
<< psubdiffcont >>
rect -2497 -171 -2463 -137
rect -2425 -171 -2391 -137
rect -2353 -171 -2319 -137
rect -2281 -171 -2247 -137
rect -2209 -171 -2175 -137
rect -2137 -171 -2103 -137
rect -2065 -171 -2031 -137
rect -1993 -171 -1959 -137
rect -1921 -171 -1887 -137
rect -1849 -171 -1815 -137
rect -1777 -171 -1743 -137
rect -1705 -171 -1671 -137
rect -1633 -171 -1599 -137
rect -1561 -171 -1527 -137
rect -1489 -171 -1455 -137
rect -1417 -171 -1383 -137
rect -1345 -171 -1311 -137
rect -939 -171 -905 -137
rect -867 -171 -833 -137
rect -795 -171 -761 -137
rect -723 -171 -689 -137
rect -651 -171 -617 -137
rect -579 -171 -545 -137
rect -507 -171 -473 -137
rect -435 -171 -401 -137
rect -363 -171 -329 -137
rect -291 -171 -257 -137
rect -219 -171 -185 -137
rect -147 -171 -113 -137
rect 273 -171 307 -137
rect 345 -171 379 -137
rect 417 -171 451 -137
rect 489 -171 523 -137
rect 561 -171 595 -137
rect 633 -171 667 -137
rect 705 -171 739 -137
rect 777 -171 811 -137
rect 849 -171 883 -137
rect 921 -171 955 -137
rect 993 -171 1027 -137
rect 1065 -171 1099 -137
rect 1485 -171 1519 -137
rect 1557 -171 1591 -137
rect 1629 -171 1663 -137
rect 1701 -171 1735 -137
rect 1773 -171 1807 -137
rect 1845 -171 1879 -137
rect 1917 -171 1951 -137
rect 1989 -171 2023 -137
rect 2061 -171 2095 -137
rect 2133 -171 2167 -137
rect 2205 -171 2239 -137
rect 2277 -171 2311 -137
<< nsubdiffcont >>
rect -2497 1407 -2463 1441
rect -2425 1407 -2391 1441
rect -2353 1407 -2319 1441
rect -2281 1407 -2247 1441
rect -2209 1407 -2175 1441
rect -2137 1407 -2103 1441
rect -2065 1407 -2031 1441
rect -1993 1407 -1959 1441
rect -1921 1407 -1887 1441
rect -1849 1407 -1815 1441
rect -1777 1407 -1743 1441
rect -1705 1407 -1671 1441
rect -939 1407 -905 1441
rect -867 1407 -833 1441
rect -795 1407 -761 1441
rect -723 1407 -689 1441
rect -651 1407 -617 1441
rect -579 1407 -545 1441
rect -507 1407 -473 1441
rect -435 1407 -401 1441
rect -363 1407 -329 1441
rect -291 1407 -257 1441
rect -219 1407 -185 1441
rect -147 1407 -113 1441
rect 273 1407 307 1441
rect 345 1407 379 1441
rect 417 1407 451 1441
rect 489 1407 523 1441
rect 561 1407 595 1441
rect 633 1407 667 1441
rect 705 1407 739 1441
rect 777 1407 811 1441
rect 849 1407 883 1441
rect 921 1407 955 1441
rect 993 1407 1027 1441
rect 1065 1407 1099 1441
rect 1485 1407 1519 1441
rect 1557 1407 1591 1441
rect 1629 1407 1663 1441
rect 1701 1407 1735 1441
rect 1773 1407 1807 1441
rect 1845 1407 1879 1441
rect 1917 1407 1951 1441
rect 1989 1407 2023 1441
rect 2061 1407 2095 1441
rect 2133 1407 2167 1441
rect 2205 1407 2239 1441
rect 2277 1407 2311 1441
rect -2497 -1749 -2463 -1715
rect -2425 -1749 -2391 -1715
rect -2353 -1749 -2319 -1715
rect -2281 -1749 -2247 -1715
rect -2209 -1749 -2175 -1715
rect -2137 -1749 -2103 -1715
rect -2065 -1749 -2031 -1715
rect -1993 -1749 -1959 -1715
rect -1921 -1749 -1887 -1715
rect -1849 -1749 -1815 -1715
rect -1777 -1749 -1743 -1715
rect -1705 -1749 -1671 -1715
rect -1633 -1749 -1599 -1715
rect -1561 -1749 -1527 -1715
rect -1489 -1749 -1455 -1715
rect -1417 -1749 -1383 -1715
rect -1345 -1749 -1311 -1715
rect -939 -1749 -905 -1715
rect -867 -1749 -833 -1715
rect -795 -1749 -761 -1715
rect -723 -1749 -689 -1715
rect -651 -1749 -617 -1715
rect -579 -1749 -545 -1715
rect -507 -1749 -473 -1715
rect -435 -1749 -401 -1715
rect -363 -1749 -329 -1715
rect -291 -1749 -257 -1715
rect -219 -1749 -185 -1715
rect -147 -1749 -113 -1715
rect 273 -1749 307 -1715
rect 345 -1749 379 -1715
rect 417 -1749 451 -1715
rect 489 -1749 523 -1715
rect 561 -1749 595 -1715
rect 633 -1749 667 -1715
rect 705 -1749 739 -1715
rect 777 -1749 811 -1715
rect 849 -1749 883 -1715
rect 921 -1749 955 -1715
rect 993 -1749 1027 -1715
rect 1065 -1749 1099 -1715
<< poly >>
rect -1920 1327 -1840 1350
rect -1920 1293 -1897 1327
rect -1863 1293 -1840 1327
rect -1920 1270 -1840 1293
rect -2320 1240 -2290 1270
rect -2170 1240 -2140 1270
rect -2020 1240 -1990 1270
rect -1870 1240 -1840 1270
rect -817 1240 -787 1270
rect -667 1240 -637 1270
rect -277 1240 -247 1270
rect 395 1240 425 1270
rect 545 1240 575 1270
rect 935 1240 965 1270
rect 1607 1240 1637 1270
rect 1757 1240 1787 1270
rect 2147 1240 2177 1270
rect -2320 616 -2290 640
rect -2400 593 -2290 616
rect -2400 559 -2377 593
rect -2343 559 -2290 593
rect -2400 539 -2290 559
rect -2400 536 -2320 539
rect -2170 497 -2140 640
rect -2292 467 -2140 497
rect -2020 497 -1990 640
rect -1870 616 -1840 640
rect -1870 593 -1760 616
rect -817 610 -787 640
rect -1870 559 -1817 593
rect -1783 559 -1760 593
rect -1870 539 -1760 559
rect -1840 536 -1760 539
rect -897 587 -787 610
rect -897 553 -874 587
rect -840 553 -787 587
rect -897 530 -787 553
rect -2020 467 -1868 497
rect -2292 425 -2262 467
rect -2370 402 -2262 425
rect -2370 368 -2347 402
rect -2313 368 -2262 402
rect -2370 360 -2262 368
rect -2220 402 -2140 425
rect -2220 368 -2197 402
rect -2163 368 -2140 402
rect -2370 345 -2290 360
rect -2220 345 -2140 368
rect -2320 330 -2290 345
rect -2170 330 -2140 345
rect -2020 402 -1940 425
rect -2020 368 -1997 402
rect -1963 368 -1940 402
rect -2020 345 -1940 368
rect -1898 382 -1868 467
rect -1898 352 -1840 382
rect -2020 330 -1990 345
rect -1870 330 -1840 352
rect -817 330 -787 530
rect -667 330 -637 640
rect -277 610 -247 640
rect 395 610 425 640
rect -357 587 -247 610
rect -357 553 -334 587
rect -300 553 -247 587
rect -357 530 -247 553
rect 315 587 425 610
rect 315 553 338 587
rect 372 553 425 587
rect 315 530 425 553
rect -277 330 -247 530
rect 395 330 425 530
rect 545 330 575 640
rect 935 610 965 640
rect 1607 610 1637 640
rect 855 587 965 610
rect 855 553 878 587
rect 912 553 965 587
rect 855 530 965 553
rect 1527 587 1637 610
rect 1527 553 1550 587
rect 1584 553 1637 587
rect 1527 530 1637 553
rect 935 330 965 530
rect 1607 330 1637 530
rect 1757 330 1787 640
rect 2147 610 2177 640
rect 2067 587 2177 610
rect 2067 553 2090 587
rect 2124 553 2177 587
rect 2067 530 2177 553
rect 2147 330 2177 530
rect -2320 0 -2290 30
rect -2170 0 -2140 30
rect -2020 0 -1990 30
rect -1870 0 -1840 30
rect -817 0 -787 30
rect -667 0 -637 30
rect -277 0 -247 30
rect 395 0 425 30
rect 545 0 575 30
rect 935 0 965 30
rect 1607 0 1637 30
rect 1757 0 1787 30
rect 2147 0 2177 30
rect -1920 -23 -1840 0
rect -1920 -57 -1897 -23
rect -1863 -57 -1840 -23
rect -1920 -80 -1840 -57
rect -717 -23 -637 0
rect -717 -57 -694 -23
rect -660 -57 -637 -23
rect -717 -80 -637 -57
rect 495 -23 575 0
rect 495 -57 518 -23
rect 552 -57 575 -23
rect 495 -80 575 -57
rect 1707 -23 1787 0
rect 1707 -57 1730 -23
rect 1764 -57 1787 -23
rect 1707 -80 1787 -57
rect -1920 -251 -1840 -228
rect -1920 -285 -1897 -251
rect -1863 -285 -1840 -251
rect -1920 -308 -1840 -285
rect -717 -251 -637 -228
rect -717 -285 -694 -251
rect -660 -285 -637 -251
rect -717 -308 -637 -285
rect 495 -251 575 -228
rect 495 -285 518 -251
rect 552 -285 575 -251
rect 495 -308 575 -285
rect -2320 -338 -2290 -308
rect -2170 -338 -2140 -308
rect -2020 -338 -1990 -308
rect -1870 -338 -1840 -308
rect -1469 -338 -1439 -308
rect -817 -338 -787 -308
rect -667 -338 -637 -308
rect -277 -338 -247 -308
rect 395 -338 425 -308
rect 545 -338 575 -308
rect 935 -338 965 -308
rect -2320 -653 -2290 -638
rect -2170 -653 -2140 -638
rect -2370 -668 -2290 -653
rect -2370 -676 -2262 -668
rect -2370 -710 -2347 -676
rect -2313 -710 -2262 -676
rect -2370 -733 -2262 -710
rect -2220 -676 -2140 -653
rect -2220 -710 -2197 -676
rect -2163 -710 -2140 -676
rect -2220 -733 -2140 -710
rect -2020 -653 -1990 -638
rect -2020 -676 -1940 -653
rect -1870 -660 -1840 -638
rect -2020 -710 -1997 -676
rect -1963 -710 -1940 -676
rect -2020 -733 -1940 -710
rect -1898 -690 -1840 -660
rect -2292 -775 -2262 -733
rect -1898 -775 -1868 -690
rect -2292 -805 -2140 -775
rect -2400 -847 -2320 -844
rect -2400 -867 -2290 -847
rect -2400 -901 -2377 -867
rect -2343 -901 -2290 -867
rect -2400 -924 -2290 -901
rect -2320 -948 -2290 -924
rect -2170 -948 -2140 -805
rect -2020 -805 -1868 -775
rect -2020 -948 -1990 -805
rect -1469 -838 -1439 -638
rect -817 -838 -787 -638
rect -1840 -847 -1760 -844
rect -1870 -867 -1760 -847
rect -1870 -901 -1817 -867
rect -1783 -901 -1760 -867
rect -1870 -924 -1760 -901
rect -1549 -861 -1439 -838
rect -1549 -895 -1526 -861
rect -1492 -895 -1439 -861
rect -1549 -918 -1439 -895
rect -897 -861 -787 -838
rect -897 -895 -874 -861
rect -840 -895 -787 -861
rect -897 -918 -787 -895
rect -1870 -948 -1840 -924
rect -1469 -948 -1439 -918
rect -817 -948 -787 -918
rect -667 -948 -637 -638
rect -277 -838 -247 -638
rect 395 -838 425 -638
rect -357 -861 -247 -838
rect -357 -895 -334 -861
rect -300 -895 -247 -861
rect -357 -918 -247 -895
rect 315 -861 425 -838
rect 315 -895 338 -861
rect 372 -895 425 -861
rect 315 -918 425 -895
rect -277 -948 -247 -918
rect 395 -948 425 -918
rect 545 -948 575 -638
rect 935 -838 965 -638
rect 855 -861 965 -838
rect 855 -895 878 -861
rect 912 -895 965 -861
rect 855 -918 965 -895
rect 935 -948 965 -918
rect -2320 -1578 -2290 -1548
rect -2170 -1578 -2140 -1548
rect -2020 -1578 -1990 -1548
rect -1870 -1578 -1840 -1548
rect -1469 -1578 -1439 -1548
rect -817 -1578 -787 -1548
rect -667 -1578 -637 -1548
rect -277 -1578 -247 -1548
rect 395 -1578 425 -1548
rect 545 -1578 575 -1548
rect 935 -1578 965 -1548
rect -1920 -1601 -1840 -1578
rect -1920 -1635 -1897 -1601
rect -1863 -1635 -1840 -1601
rect -1920 -1658 -1840 -1635
<< polycont >>
rect -1897 1293 -1863 1327
rect -2377 559 -2343 593
rect -1817 559 -1783 593
rect -874 553 -840 587
rect -2347 368 -2313 402
rect -2197 368 -2163 402
rect -1997 368 -1963 402
rect -334 553 -300 587
rect 338 553 372 587
rect 878 553 912 587
rect 1550 553 1584 587
rect 2090 553 2124 587
rect -1897 -57 -1863 -23
rect -694 -57 -660 -23
rect 518 -57 552 -23
rect 1730 -57 1764 -23
rect -1897 -285 -1863 -251
rect -694 -285 -660 -251
rect 518 -285 552 -251
rect -2347 -710 -2313 -676
rect -2197 -710 -2163 -676
rect -1997 -710 -1963 -676
rect -2377 -901 -2343 -867
rect -1817 -901 -1783 -867
rect -1526 -895 -1492 -861
rect -874 -895 -840 -861
rect -334 -895 -300 -861
rect 338 -895 372 -861
rect 878 -895 912 -861
rect -1897 -1635 -1863 -1601
<< locali >>
rect -2520 1441 -1640 1464
rect -2970 1399 -2890 1422
rect -2970 1365 -2947 1399
rect -2913 1365 -2890 1399
rect -2520 1407 -2497 1441
rect -2463 1407 -2425 1441
rect -2391 1407 -2353 1441
rect -2319 1407 -2281 1441
rect -2247 1407 -2209 1441
rect -2175 1407 -2137 1441
rect -2103 1407 -2065 1441
rect -2031 1407 -1993 1441
rect -1959 1407 -1921 1441
rect -1887 1407 -1849 1441
rect -1815 1407 -1777 1441
rect -1743 1407 -1705 1441
rect -1671 1407 -1640 1441
rect -2520 1384 -1640 1407
rect -962 1441 -82 1464
rect -962 1407 -939 1441
rect -905 1407 -867 1441
rect -833 1407 -795 1441
rect -761 1407 -723 1441
rect -689 1407 -651 1441
rect -617 1407 -579 1441
rect -545 1407 -507 1441
rect -473 1407 -435 1441
rect -401 1407 -363 1441
rect -329 1407 -291 1441
rect -257 1407 -219 1441
rect -185 1407 -147 1441
rect -113 1407 -82 1441
rect -962 1384 -82 1407
rect 250 1441 1130 1464
rect 250 1407 273 1441
rect 307 1407 345 1441
rect 379 1407 417 1441
rect 451 1407 489 1441
rect 523 1407 561 1441
rect 595 1407 633 1441
rect 667 1407 705 1441
rect 739 1407 777 1441
rect 811 1407 849 1441
rect 883 1407 921 1441
rect 955 1407 993 1441
rect 1027 1407 1065 1441
rect 1099 1407 1130 1441
rect 250 1384 1130 1407
rect 1462 1441 2342 1464
rect 1462 1407 1485 1441
rect 1519 1407 1557 1441
rect 1591 1407 1629 1441
rect 1663 1407 1701 1441
rect 1735 1407 1773 1441
rect 1807 1407 1845 1441
rect 1879 1407 1917 1441
rect 1951 1407 1989 1441
rect 2023 1407 2061 1441
rect 2095 1407 2133 1441
rect 2167 1407 2205 1441
rect 2239 1407 2277 1441
rect 2311 1407 2342 1441
rect 1462 1384 2342 1407
rect -2970 1330 -2890 1365
rect -1920 1330 -1840 1350
rect -2970 1327 -1840 1330
rect -2970 1293 -2947 1327
rect -2913 1293 -1897 1327
rect -1863 1293 -1840 1327
rect -2970 1290 -1840 1293
rect -2970 1255 -2890 1290
rect -1920 1270 -1840 1290
rect -1706 1326 -1554 1346
rect -1706 1323 -1480 1326
rect -1706 1289 -1683 1323
rect -1649 1289 -1611 1323
rect -1577 1289 -1480 1323
rect -1706 1286 -1480 1289
rect -1706 1266 -1554 1286
rect -2970 1221 -2947 1255
rect -2913 1221 -2890 1255
rect -2970 1198 -2890 1221
rect -2420 1209 -2340 1220
rect -2420 1161 -2397 1209
rect -2363 1161 -2340 1209
rect -2420 1137 -2340 1161
rect -2420 1093 -2397 1137
rect -2363 1093 -2340 1137
rect -2420 1065 -2340 1093
rect -2420 1025 -2397 1065
rect -2363 1025 -2340 1065
rect -2420 993 -2340 1025
rect -2420 957 -2397 993
rect -2363 957 -2340 993
rect -2420 923 -2340 957
rect -2420 887 -2397 923
rect -2363 887 -2340 923
rect -2420 855 -2340 887
rect -2420 815 -2397 855
rect -2363 815 -2340 855
rect -2420 787 -2340 815
rect -2420 743 -2397 787
rect -2363 743 -2340 787
rect -2420 719 -2340 743
rect -2856 665 -2776 688
rect -2856 631 -2833 665
rect -2799 631 -2776 665
rect -2420 671 -2397 719
rect -2363 671 -2340 719
rect -2420 660 -2340 671
rect -2120 1209 -2040 1220
rect -2120 1161 -2097 1209
rect -2063 1161 -2040 1209
rect -2120 1137 -2040 1161
rect -2120 1093 -2097 1137
rect -2063 1093 -2040 1137
rect -2120 1065 -2040 1093
rect -2120 1025 -2097 1065
rect -2063 1025 -2040 1065
rect -2120 993 -2040 1025
rect -2120 957 -2097 993
rect -2063 957 -2040 993
rect -2120 923 -2040 957
rect -2120 887 -2097 923
rect -2063 887 -2040 923
rect -2120 855 -2040 887
rect -2120 815 -2097 855
rect -2063 815 -2040 855
rect -2120 787 -2040 815
rect -2120 743 -2097 787
rect -2063 743 -2040 787
rect -2120 719 -2040 743
rect -2120 671 -2097 719
rect -2063 671 -2040 719
rect -2120 660 -2040 671
rect -1820 1209 -1740 1220
rect -1820 1161 -1797 1209
rect -1763 1161 -1740 1209
rect -1820 1137 -1740 1161
rect -1820 1093 -1797 1137
rect -1763 1093 -1740 1137
rect -1820 1065 -1740 1093
rect -1820 1025 -1797 1065
rect -1763 1025 -1740 1065
rect -1820 993 -1740 1025
rect -1820 957 -1797 993
rect -1763 957 -1740 993
rect -1820 923 -1740 957
rect -1820 887 -1797 923
rect -1763 887 -1740 923
rect -1820 855 -1740 887
rect -1820 815 -1797 855
rect -1763 815 -1740 855
rect -1820 787 -1740 815
rect -1820 743 -1797 787
rect -1763 743 -1740 787
rect -1820 719 -1740 743
rect -1820 671 -1797 719
rect -1763 671 -1740 719
rect -1820 660 -1740 671
rect -2856 596 -2776 631
rect -2400 596 -2320 616
rect -2856 593 -1960 596
rect -2856 559 -2833 593
rect -2799 559 -2377 593
rect -2343 559 -1960 593
rect -2856 556 -1960 559
rect -2856 521 -2776 556
rect -2400 536 -2320 556
rect -3654 474 -3574 497
rect -3654 440 -3631 474
rect -3597 440 -3574 474
rect -2856 487 -2833 521
rect -2799 487 -2776 521
rect -2856 464 -2776 487
rect -3654 405 -3574 440
rect -2000 425 -1960 556
rect -1840 593 -1760 616
rect -1840 559 -1817 593
rect -1783 559 -1760 593
rect -1840 536 -1760 559
rect -1520 590 -1480 1286
rect -917 1209 -837 1220
rect -917 1161 -894 1209
rect -860 1161 -837 1209
rect -917 1137 -837 1161
rect -917 1093 -894 1137
rect -860 1093 -837 1137
rect -917 1065 -837 1093
rect -917 1025 -894 1065
rect -860 1025 -837 1065
rect -917 993 -837 1025
rect -917 957 -894 993
rect -860 957 -837 993
rect -917 923 -837 957
rect -917 887 -894 923
rect -860 887 -837 923
rect -917 855 -837 887
rect -917 815 -894 855
rect -860 815 -837 855
rect -917 787 -837 815
rect -917 743 -894 787
rect -860 743 -837 787
rect -917 719 -837 743
rect -917 671 -894 719
rect -860 671 -837 719
rect -917 660 -837 671
rect -617 1195 -537 1220
rect -617 1161 -594 1195
rect -560 1161 -537 1195
rect -617 1127 -537 1161
rect -617 1093 -594 1127
rect -560 1093 -537 1127
rect -617 1059 -537 1093
rect -617 1025 -594 1059
rect -560 1025 -537 1059
rect -617 991 -537 1025
rect -617 957 -594 991
rect -560 957 -537 991
rect -617 923 -537 957
rect -617 889 -594 923
rect -560 889 -537 923
rect -617 855 -537 889
rect -617 821 -594 855
rect -560 821 -537 855
rect -617 787 -537 821
rect -617 753 -594 787
rect -560 753 -537 787
rect -617 719 -537 753
rect -617 685 -594 719
rect -560 685 -537 719
rect -617 660 -537 685
rect -377 1209 -297 1220
rect -377 1161 -354 1209
rect -320 1161 -297 1209
rect -377 1137 -297 1161
rect -377 1093 -354 1137
rect -320 1093 -297 1137
rect -377 1065 -297 1093
rect -377 1025 -354 1065
rect -320 1025 -297 1065
rect -377 993 -297 1025
rect -377 957 -354 993
rect -320 957 -297 993
rect -377 923 -297 957
rect -377 887 -354 923
rect -320 887 -297 923
rect -377 855 -297 887
rect -377 815 -354 855
rect -320 815 -297 855
rect -377 787 -297 815
rect -377 743 -354 787
rect -320 743 -297 787
rect -377 719 -297 743
rect -377 671 -354 719
rect -320 671 -297 719
rect -377 660 -297 671
rect -227 1195 -147 1220
rect -227 1161 -204 1195
rect -170 1161 -147 1195
rect -227 1127 -147 1161
rect -227 1093 -204 1127
rect -170 1093 -147 1127
rect -227 1059 -147 1093
rect -227 1025 -204 1059
rect -170 1025 -147 1059
rect -227 991 -147 1025
rect -227 957 -204 991
rect -170 957 -147 991
rect -227 923 -147 957
rect -227 889 -204 923
rect -170 889 -147 923
rect -227 855 -147 889
rect -227 821 -204 855
rect -170 821 -147 855
rect -227 787 -147 821
rect -227 753 -204 787
rect -170 753 -147 787
rect -227 719 -147 753
rect -227 685 -204 719
rect -170 685 -147 719
rect -227 660 -147 685
rect 295 1209 375 1220
rect 295 1161 318 1209
rect 352 1161 375 1209
rect 295 1137 375 1161
rect 295 1093 318 1137
rect 352 1093 375 1137
rect 295 1065 375 1093
rect 295 1025 318 1065
rect 352 1025 375 1065
rect 295 993 375 1025
rect 295 957 318 993
rect 352 957 375 993
rect 295 923 375 957
rect 295 887 318 923
rect 352 887 375 923
rect 295 855 375 887
rect 295 815 318 855
rect 352 815 375 855
rect 295 787 375 815
rect 295 743 318 787
rect 352 743 375 787
rect 295 719 375 743
rect 295 671 318 719
rect 352 671 375 719
rect 295 660 375 671
rect 445 1195 525 1220
rect 445 1161 468 1195
rect 502 1161 525 1195
rect 445 1127 525 1161
rect 445 1093 468 1127
rect 502 1093 525 1127
rect 445 1059 525 1093
rect 445 1025 468 1059
rect 502 1025 525 1059
rect 445 991 525 1025
rect 445 957 468 991
rect 502 957 525 991
rect 445 923 525 957
rect 445 889 468 923
rect 502 889 525 923
rect 445 855 525 889
rect 445 821 468 855
rect 502 821 525 855
rect 445 787 525 821
rect 445 753 468 787
rect 502 753 525 787
rect 445 719 525 753
rect 445 685 468 719
rect 502 685 525 719
rect 445 660 525 685
rect 595 1209 675 1220
rect 595 1161 618 1209
rect 652 1161 675 1209
rect 595 1137 675 1161
rect 595 1093 618 1137
rect 652 1093 675 1137
rect 595 1065 675 1093
rect 595 1025 618 1065
rect 652 1025 675 1065
rect 595 993 675 1025
rect 595 957 618 993
rect 652 957 675 993
rect 595 923 675 957
rect 595 887 618 923
rect 652 887 675 923
rect 595 855 675 887
rect 595 815 618 855
rect 652 815 675 855
rect 595 787 675 815
rect 595 743 618 787
rect 652 743 675 787
rect 595 719 675 743
rect 595 671 618 719
rect 652 671 675 719
rect 595 660 675 671
rect 835 1209 915 1220
rect 835 1161 858 1209
rect 892 1161 915 1209
rect 835 1137 915 1161
rect 835 1093 858 1137
rect 892 1093 915 1137
rect 835 1065 915 1093
rect 835 1025 858 1065
rect 892 1025 915 1065
rect 835 993 915 1025
rect 835 957 858 993
rect 892 957 915 993
rect 835 923 915 957
rect 835 887 858 923
rect 892 887 915 923
rect 835 855 915 887
rect 835 815 858 855
rect 892 815 915 855
rect 835 787 915 815
rect 835 743 858 787
rect 892 743 915 787
rect 835 719 915 743
rect 835 671 858 719
rect 892 671 915 719
rect 835 660 915 671
rect 985 1195 1065 1220
rect 985 1161 1008 1195
rect 1042 1161 1065 1195
rect 985 1127 1065 1161
rect 985 1093 1008 1127
rect 1042 1093 1065 1127
rect 985 1059 1065 1093
rect 985 1025 1008 1059
rect 1042 1025 1065 1059
rect 985 991 1065 1025
rect 985 957 1008 991
rect 1042 957 1065 991
rect 985 923 1065 957
rect 985 889 1008 923
rect 1042 889 1065 923
rect 985 855 1065 889
rect 985 821 1008 855
rect 1042 821 1065 855
rect 985 787 1065 821
rect 985 753 1008 787
rect 1042 753 1065 787
rect 985 719 1065 753
rect 985 685 1008 719
rect 1042 685 1065 719
rect 985 660 1065 685
rect 1507 1209 1587 1220
rect 1507 1161 1530 1209
rect 1564 1161 1587 1209
rect 1507 1137 1587 1161
rect 1507 1093 1530 1137
rect 1564 1093 1587 1137
rect 1507 1065 1587 1093
rect 1507 1025 1530 1065
rect 1564 1025 1587 1065
rect 1507 993 1587 1025
rect 1507 957 1530 993
rect 1564 957 1587 993
rect 1507 923 1587 957
rect 1507 887 1530 923
rect 1564 887 1587 923
rect 1507 855 1587 887
rect 1507 815 1530 855
rect 1564 815 1587 855
rect 1507 787 1587 815
rect 1507 743 1530 787
rect 1564 743 1587 787
rect 1507 719 1587 743
rect 1507 671 1530 719
rect 1564 671 1587 719
rect 1507 660 1587 671
rect 1807 1195 1887 1220
rect 1807 1161 1830 1195
rect 1864 1161 1887 1195
rect 1807 1127 1887 1161
rect 1807 1093 1830 1127
rect 1864 1093 1887 1127
rect 1807 1059 1887 1093
rect 1807 1025 1830 1059
rect 1864 1025 1887 1059
rect 1807 991 1887 1025
rect 1807 957 1830 991
rect 1864 957 1887 991
rect 1807 923 1887 957
rect 1807 889 1830 923
rect 1864 889 1887 923
rect 1807 855 1887 889
rect 1807 821 1830 855
rect 1864 821 1887 855
rect 1807 787 1887 821
rect 1807 753 1830 787
rect 1864 753 1887 787
rect 1807 719 1887 753
rect 1807 685 1830 719
rect 1864 685 1887 719
rect 1807 660 1887 685
rect 2047 1209 2127 1220
rect 2047 1161 2070 1209
rect 2104 1161 2127 1209
rect 2047 1137 2127 1161
rect 2047 1093 2070 1137
rect 2104 1093 2127 1137
rect 2047 1065 2127 1093
rect 2047 1025 2070 1065
rect 2104 1025 2127 1065
rect 2047 993 2127 1025
rect 2047 957 2070 993
rect 2104 957 2127 993
rect 2047 923 2127 957
rect 2047 887 2070 923
rect 2104 887 2127 923
rect 2047 855 2127 887
rect 2047 815 2070 855
rect 2104 815 2127 855
rect 2047 787 2127 815
rect 2047 743 2070 787
rect 2104 743 2127 787
rect 2047 719 2127 743
rect 2047 671 2070 719
rect 2104 671 2127 719
rect 2047 660 2127 671
rect 2197 1195 2277 1220
rect 2197 1161 2220 1195
rect 2254 1161 2277 1195
rect 2197 1127 2277 1161
rect 2197 1093 2220 1127
rect 2254 1093 2277 1127
rect 2197 1059 2277 1093
rect 2197 1025 2220 1059
rect 2254 1025 2277 1059
rect 2197 991 2277 1025
rect 2197 957 2220 991
rect 2254 957 2277 991
rect 2197 923 2277 957
rect 2197 889 2220 923
rect 2254 889 2277 923
rect 2197 855 2277 889
rect 2197 821 2220 855
rect 2254 821 2277 855
rect 2197 787 2277 821
rect 2197 753 2220 787
rect 2254 753 2277 787
rect 2197 719 2277 753
rect 2197 685 2220 719
rect 2254 685 2277 719
rect 2197 660 2277 685
rect -897 590 -817 610
rect -597 590 -557 660
rect -357 590 -277 610
rect -1520 587 -817 590
rect -1520 553 -874 587
rect -840 553 -817 587
rect -1520 550 -817 553
rect -897 530 -817 550
rect -747 587 -277 590
rect -747 553 -334 587
rect -300 553 -277 587
rect -747 550 -277 553
rect -2370 405 -2290 425
rect -3654 402 -2290 405
rect -3654 368 -3631 402
rect -3597 368 -2347 402
rect -2313 368 -2290 402
rect -3654 365 -2290 368
rect -3654 330 -3574 365
rect -2370 345 -2290 365
rect -2220 402 -2140 425
rect -2220 368 -2197 402
rect -2163 368 -2140 402
rect -2220 345 -2140 368
rect -2020 402 -1940 425
rect -2020 368 -1997 402
rect -1963 368 -1940 402
rect -2020 345 -1940 368
rect -3654 296 -3631 330
rect -3597 296 -3574 330
rect -747 310 -707 550
rect -357 530 -277 550
rect -207 596 -167 660
rect 315 596 395 610
rect -207 587 395 596
rect -207 556 338 587
rect -207 310 -167 556
rect 315 553 338 556
rect 372 553 395 587
rect 315 530 395 553
rect 465 590 505 660
rect 855 590 935 610
rect 465 587 935 590
rect 465 553 878 587
rect 912 553 935 587
rect 465 550 935 553
rect -81 499 -1 522
rect -81 465 -58 499
rect -24 465 -1 499
rect -81 442 -1 465
rect -3654 273 -3574 296
rect -2420 299 -2340 310
rect -2420 235 -2397 299
rect -2363 235 -2340 299
rect -2420 231 -2340 235
rect -2420 129 -2397 231
rect -2363 129 -2340 231
rect -2420 125 -2340 129
rect -3540 49 -3460 72
rect -2420 61 -2397 125
rect -2363 61 -2340 125
rect -2420 50 -2340 61
rect -2120 299 -2040 310
rect -2120 235 -2097 299
rect -2063 235 -2040 299
rect -2120 231 -2040 235
rect -2120 129 -2097 231
rect -2063 129 -2040 231
rect -2120 125 -2040 129
rect -2120 61 -2097 125
rect -2063 61 -2040 125
rect -2120 50 -2040 61
rect -1820 299 -1740 310
rect -1820 235 -1797 299
rect -1763 235 -1740 299
rect -1820 231 -1740 235
rect -1820 129 -1797 231
rect -1763 129 -1740 231
rect -1820 125 -1740 129
rect -1820 61 -1797 125
rect -1763 61 -1740 125
rect -1820 50 -1740 61
rect -917 299 -837 310
rect -917 235 -894 299
rect -860 235 -837 299
rect -917 231 -837 235
rect -917 129 -894 231
rect -860 129 -837 231
rect -917 125 -837 129
rect -917 61 -894 125
rect -860 61 -837 125
rect -917 50 -837 61
rect -767 299 -687 310
rect -767 265 -744 299
rect -710 265 -687 299
rect -767 231 -687 265
rect -767 197 -744 231
rect -710 197 -687 231
rect -767 163 -687 197
rect -767 129 -744 163
rect -710 129 -687 163
rect -767 95 -687 129
rect -767 61 -744 95
rect -710 61 -687 95
rect -767 50 -687 61
rect -617 299 -537 310
rect -617 235 -594 299
rect -560 235 -537 299
rect -617 231 -537 235
rect -617 129 -594 231
rect -560 129 -537 231
rect -617 125 -537 129
rect -617 61 -594 125
rect -560 61 -537 125
rect -617 50 -537 61
rect -377 299 -297 310
rect -377 235 -354 299
rect -320 235 -297 299
rect -377 231 -297 235
rect -377 129 -354 231
rect -320 129 -297 231
rect -377 125 -297 129
rect -377 61 -354 125
rect -320 61 -297 125
rect -377 50 -297 61
rect -227 299 -147 310
rect -227 265 -204 299
rect -170 265 -147 299
rect -227 231 -147 265
rect -227 197 -204 231
rect -170 197 -147 231
rect -227 163 -147 197
rect -227 129 -204 163
rect -170 129 -147 163
rect -227 95 -147 129
rect -227 61 -204 95
rect -170 61 -147 95
rect -227 50 -147 61
rect -3540 15 -3517 49
rect -3483 15 -3460 49
rect -3540 -20 -3460 15
rect -2816 -8 -2588 32
rect -2816 -20 -2776 -8
rect -3540 -23 -2776 -20
rect -3540 -57 -3517 -23
rect -3483 -57 -2776 -23
rect -2628 -20 -2588 -8
rect -1920 -20 -1840 0
rect -2628 -23 -1840 -20
rect -3540 -60 -2776 -57
rect -3540 -95 -3460 -60
rect -3540 -129 -3517 -95
rect -3483 -129 -3460 -95
rect -3540 -152 -3460 -129
rect -2742 -65 -2662 -42
rect -2628 -57 -1897 -23
rect -1863 -57 -1840 -23
rect -2628 -60 -1840 -57
rect -2742 -99 -2719 -65
rect -2685 -99 -2662 -65
rect -1920 -80 -1840 -60
rect -1706 -19 -1554 4
rect -1706 -53 -1683 -19
rect -1649 -53 -1611 -19
rect -1577 -20 -1554 -19
rect -717 -20 -637 0
rect -1577 -23 -637 -20
rect -1577 -53 -694 -23
rect -1706 -57 -694 -53
rect -660 -57 -637 -23
rect -1706 -60 -637 -57
rect -61 -20 -21 442
rect 615 310 655 550
rect 855 530 935 550
rect 1005 590 1045 660
rect 1527 590 1607 610
rect 1827 590 1867 660
rect 2067 590 2147 610
rect 1005 587 1607 590
rect 1005 553 1550 587
rect 1584 553 1607 587
rect 1005 550 1607 553
rect 1005 310 1045 550
rect 1527 530 1607 550
rect 1677 587 2147 590
rect 1677 553 2090 587
rect 2124 553 2147 587
rect 1677 550 2147 553
rect 1677 310 1717 550
rect 2067 530 2147 550
rect 2217 548 2257 660
rect 2197 525 2277 548
rect 2197 491 2220 525
rect 2254 491 2277 525
rect 2197 453 2277 491
rect 2197 419 2220 453
rect 2254 419 2277 453
rect 2197 396 2277 419
rect 2217 310 2257 396
rect 295 299 375 310
rect 295 235 318 299
rect 352 235 375 299
rect 295 231 375 235
rect 295 129 318 231
rect 352 129 375 231
rect 295 125 375 129
rect 295 61 318 125
rect 352 61 375 125
rect 295 50 375 61
rect 595 299 675 310
rect 595 265 618 299
rect 652 265 675 299
rect 595 231 675 265
rect 595 197 618 231
rect 652 197 675 231
rect 595 163 675 197
rect 595 129 618 163
rect 652 129 675 163
rect 595 95 675 129
rect 595 61 618 95
rect 652 61 675 95
rect 595 50 675 61
rect 835 299 915 310
rect 835 235 858 299
rect 892 235 915 299
rect 835 231 915 235
rect 835 129 858 231
rect 892 129 915 231
rect 835 125 915 129
rect 835 61 858 125
rect 892 61 915 125
rect 835 50 915 61
rect 985 299 1065 310
rect 985 265 1008 299
rect 1042 265 1065 299
rect 985 231 1065 265
rect 985 197 1008 231
rect 1042 197 1065 231
rect 985 163 1065 197
rect 985 129 1008 163
rect 1042 129 1065 163
rect 985 95 1065 129
rect 985 61 1008 95
rect 1042 61 1065 95
rect 985 50 1065 61
rect 1507 299 1587 310
rect 1507 235 1530 299
rect 1564 235 1587 299
rect 1507 231 1587 235
rect 1507 129 1530 231
rect 1564 129 1587 231
rect 1507 125 1587 129
rect 1507 61 1530 125
rect 1564 61 1587 125
rect 1507 50 1587 61
rect 1657 299 1737 310
rect 1657 265 1680 299
rect 1714 265 1737 299
rect 1657 231 1737 265
rect 1657 197 1680 231
rect 1714 197 1737 231
rect 1657 163 1737 197
rect 1657 129 1680 163
rect 1714 129 1737 163
rect 1657 95 1737 129
rect 1657 61 1680 95
rect 1714 61 1737 95
rect 1657 50 1737 61
rect 1807 299 1887 310
rect 1807 235 1830 299
rect 1864 235 1887 299
rect 1807 231 1887 235
rect 1807 129 1830 231
rect 1864 129 1887 231
rect 1807 125 1887 129
rect 1807 61 1830 125
rect 1864 61 1887 125
rect 1807 50 1887 61
rect 2047 299 2127 310
rect 2047 235 2070 299
rect 2104 235 2127 299
rect 2047 231 2127 235
rect 2047 129 2070 231
rect 2104 129 2127 231
rect 2047 125 2127 129
rect 2047 61 2070 125
rect 2104 61 2127 125
rect 2047 50 2127 61
rect 2197 299 2277 310
rect 2197 265 2220 299
rect 2254 265 2277 299
rect 2197 231 2277 265
rect 2197 197 2220 231
rect 2254 197 2277 231
rect 2197 163 2277 197
rect 2197 129 2220 163
rect 2254 129 2277 163
rect 2197 95 2277 129
rect 2197 61 2220 95
rect 2254 61 2277 95
rect 2197 50 2277 61
rect 495 -20 575 0
rect 1707 -20 1787 0
rect -61 -23 575 -20
rect -61 -57 518 -23
rect 552 -57 575 -23
rect -61 -60 575 -57
rect -1706 -76 -1554 -60
rect -717 -80 -637 -60
rect 495 -80 575 -60
rect 1164 -23 1787 -20
rect 1164 -57 1730 -23
rect 1764 -57 1787 -23
rect 1164 -60 1787 -57
rect -2742 -114 -2662 -99
rect -2742 -137 -1283 -114
rect -2856 -179 -2776 -156
rect -2856 -213 -2833 -179
rect -2799 -213 -2776 -179
rect -2856 -251 -2776 -213
rect -2856 -285 -2833 -251
rect -2799 -285 -2776 -251
rect -2742 -171 -2719 -137
rect -2685 -171 -2497 -137
rect -2463 -171 -2425 -137
rect -2391 -171 -2353 -137
rect -2319 -171 -2281 -137
rect -2247 -171 -2209 -137
rect -2175 -171 -2137 -137
rect -2103 -171 -2065 -137
rect -2031 -171 -1993 -137
rect -1959 -171 -1921 -137
rect -1887 -171 -1849 -137
rect -1815 -171 -1777 -137
rect -1743 -171 -1705 -137
rect -1671 -171 -1633 -137
rect -1599 -171 -1561 -137
rect -1527 -171 -1489 -137
rect -1455 -171 -1417 -137
rect -1383 -171 -1345 -137
rect -1311 -171 -1283 -137
rect -2742 -194 -1283 -171
rect -962 -137 -82 -114
rect -962 -171 -939 -137
rect -905 -171 -867 -137
rect -833 -171 -795 -137
rect -761 -171 -723 -137
rect -689 -171 -651 -137
rect -617 -171 -579 -137
rect -545 -171 -507 -137
rect -473 -171 -435 -137
rect -401 -171 -363 -137
rect -329 -171 -291 -137
rect -257 -171 -219 -137
rect -185 -171 -147 -137
rect -113 -171 -82 -137
rect -962 -194 -82 -171
rect 250 -137 1130 -114
rect 250 -171 273 -137
rect 307 -171 345 -137
rect 379 -171 417 -137
rect 451 -171 489 -137
rect 523 -171 561 -137
rect 595 -171 633 -137
rect 667 -171 705 -137
rect 739 -171 777 -137
rect 811 -171 849 -137
rect 883 -171 921 -137
rect 955 -171 993 -137
rect 1027 -171 1065 -137
rect 1099 -171 1130 -137
rect 250 -194 1130 -171
rect -2742 -209 -2662 -194
rect -2742 -243 -2719 -209
rect -2685 -243 -2662 -209
rect -2742 -266 -2662 -243
rect -1920 -248 -1840 -228
rect -2628 -251 -1840 -248
rect -2856 -300 -2776 -285
rect -2628 -285 -1897 -251
rect -1863 -285 -1840 -251
rect -2628 -288 -1840 -285
rect -2628 -300 -2588 -288
rect -2856 -323 -2588 -300
rect -1920 -308 -1840 -288
rect -1481 -248 -1329 -232
rect -717 -248 -637 -228
rect 495 -248 575 -228
rect -1481 -251 -637 -248
rect -1481 -255 -694 -251
rect -1481 -289 -1458 -255
rect -1424 -289 -1386 -255
rect -1352 -285 -694 -255
rect -660 -285 -637 -251
rect -1352 -288 -637 -285
rect -1352 -289 -1329 -288
rect -1481 -312 -1329 -289
rect -717 -308 -637 -288
rect -60 -251 575 -248
rect -60 -285 518 -251
rect 552 -285 575 -251
rect -60 -288 575 -285
rect -2856 -357 -2833 -323
rect -2799 -340 -2588 -323
rect -2799 -357 -2776 -340
rect -2856 -380 -2776 -357
rect -60 -358 -20 -288
rect 495 -308 575 -288
rect 1164 -358 1204 -60
rect 1707 -80 1787 -60
rect 1462 -137 2342 -114
rect 1462 -171 1485 -137
rect 1519 -171 1557 -137
rect 1591 -171 1629 -137
rect 1663 -171 1701 -137
rect 1735 -171 1773 -137
rect 1807 -171 1845 -137
rect 1879 -171 1917 -137
rect 1951 -171 1989 -137
rect 2023 -171 2061 -137
rect 2095 -171 2133 -137
rect 2167 -171 2205 -137
rect 2239 -171 2277 -137
rect 2311 -171 2342 -137
rect 1462 -194 2342 -171
rect -2420 -369 -2340 -358
rect -2420 -433 -2397 -369
rect -2363 -433 -2340 -369
rect -2420 -437 -2340 -433
rect -2420 -539 -2397 -437
rect -2363 -539 -2340 -437
rect -2420 -543 -2340 -539
rect -2970 -604 -2890 -581
rect -2970 -638 -2947 -604
rect -2913 -638 -2890 -604
rect -2420 -607 -2397 -543
rect -2363 -607 -2340 -543
rect -2420 -618 -2340 -607
rect -2120 -369 -2040 -358
rect -2120 -433 -2097 -369
rect -2063 -433 -2040 -369
rect -2120 -437 -2040 -433
rect -2120 -539 -2097 -437
rect -2063 -539 -2040 -437
rect -2120 -543 -2040 -539
rect -2120 -607 -2097 -543
rect -2063 -607 -2040 -543
rect -2120 -618 -2040 -607
rect -1820 -369 -1740 -358
rect -1820 -433 -1797 -369
rect -1763 -433 -1740 -369
rect -1820 -437 -1740 -433
rect -1820 -539 -1797 -437
rect -1763 -539 -1740 -437
rect -1820 -543 -1740 -539
rect -1820 -607 -1797 -543
rect -1763 -607 -1740 -543
rect -1820 -618 -1740 -607
rect -1569 -369 -1489 -358
rect -1569 -433 -1546 -369
rect -1512 -433 -1489 -369
rect -1569 -437 -1489 -433
rect -1569 -539 -1546 -437
rect -1512 -539 -1489 -437
rect -1569 -543 -1489 -539
rect -1569 -607 -1546 -543
rect -1512 -607 -1489 -543
rect -1569 -618 -1489 -607
rect -1419 -369 -1339 -358
rect -1419 -403 -1396 -369
rect -1362 -403 -1339 -369
rect -1419 -437 -1339 -403
rect -1419 -471 -1396 -437
rect -1362 -471 -1339 -437
rect -1419 -505 -1339 -471
rect -1419 -539 -1396 -505
rect -1362 -539 -1339 -505
rect -1419 -573 -1339 -539
rect -1419 -607 -1396 -573
rect -1362 -607 -1339 -573
rect -1419 -618 -1339 -607
rect -917 -369 -837 -358
rect -917 -433 -894 -369
rect -860 -433 -837 -369
rect -917 -437 -837 -433
rect -917 -539 -894 -437
rect -860 -539 -837 -437
rect -917 -543 -837 -539
rect -917 -607 -894 -543
rect -860 -607 -837 -543
rect -917 -618 -837 -607
rect -617 -369 -537 -358
rect -617 -403 -594 -369
rect -560 -403 -537 -369
rect -617 -437 -537 -403
rect -617 -471 -594 -437
rect -560 -471 -537 -437
rect -617 -505 -537 -471
rect -617 -539 -594 -505
rect -560 -539 -537 -505
rect -617 -573 -537 -539
rect -617 -607 -594 -573
rect -560 -607 -537 -573
rect -617 -618 -537 -607
rect -377 -369 -297 -358
rect -377 -433 -354 -369
rect -320 -433 -297 -369
rect -377 -437 -297 -433
rect -377 -539 -354 -437
rect -320 -539 -297 -437
rect -377 -543 -297 -539
rect -377 -607 -354 -543
rect -320 -607 -297 -543
rect -377 -618 -297 -607
rect -227 -369 -20 -358
rect -227 -403 -204 -369
rect -170 -398 -20 -369
rect 295 -369 375 -358
rect -170 -403 -147 -398
rect -227 -437 -147 -403
rect -227 -471 -204 -437
rect -170 -471 -147 -437
rect -227 -505 -147 -471
rect -227 -539 -204 -505
rect -170 -539 -147 -505
rect -227 -573 -147 -539
rect -227 -607 -204 -573
rect -170 -607 -147 -573
rect -227 -618 -147 -607
rect 295 -433 318 -369
rect 352 -433 375 -369
rect 295 -437 375 -433
rect 295 -539 318 -437
rect 352 -539 375 -437
rect 295 -543 375 -539
rect 295 -607 318 -543
rect 352 -607 375 -543
rect 295 -618 375 -607
rect 595 -369 675 -358
rect 595 -403 618 -369
rect 652 -403 675 -369
rect 595 -437 675 -403
rect 595 -471 618 -437
rect 652 -471 675 -437
rect 595 -505 675 -471
rect 595 -539 618 -505
rect 652 -539 675 -505
rect 595 -573 675 -539
rect 595 -607 618 -573
rect 652 -607 675 -573
rect 595 -618 675 -607
rect 835 -369 915 -358
rect 835 -433 858 -369
rect 892 -433 915 -369
rect 835 -437 915 -433
rect 835 -539 858 -437
rect 892 -539 915 -437
rect 835 -543 915 -539
rect 835 -607 858 -543
rect 892 -607 915 -543
rect 835 -618 915 -607
rect 985 -369 1204 -358
rect 985 -403 1008 -369
rect 1042 -398 1204 -369
rect 1042 -403 1065 -398
rect 985 -437 1065 -403
rect 985 -471 1008 -437
rect 1042 -471 1065 -437
rect 985 -505 1065 -471
rect 985 -539 1008 -505
rect 1042 -539 1065 -505
rect 985 -573 1065 -539
rect 985 -607 1008 -573
rect 1042 -607 1065 -573
rect 985 -618 1065 -607
rect -2970 -673 -2890 -638
rect -2370 -673 -2290 -653
rect -2970 -676 -2290 -673
rect -2970 -710 -2947 -676
rect -2913 -710 -2347 -676
rect -2313 -710 -2290 -676
rect -2970 -713 -2290 -710
rect -2970 -748 -2890 -713
rect -2370 -733 -2290 -713
rect -2220 -676 -2140 -653
rect -2220 -710 -2197 -676
rect -2163 -710 -2140 -676
rect -2220 -733 -2140 -710
rect -2020 -676 -1940 -653
rect -2020 -710 -1997 -676
rect -1963 -710 -1940 -676
rect -1399 -678 -1359 -618
rect -2020 -733 -1940 -710
rect -1419 -701 -1339 -678
rect -3540 -795 -3460 -772
rect -3540 -829 -3517 -795
rect -3483 -829 -3460 -795
rect -2970 -782 -2947 -748
rect -2913 -782 -2890 -748
rect -2970 -805 -2890 -782
rect -3540 -864 -3460 -829
rect -2400 -864 -2320 -844
rect -2000 -864 -1960 -733
rect -1691 -755 -1611 -732
rect -1691 -789 -1668 -755
rect -1634 -789 -1611 -755
rect -1691 -827 -1611 -789
rect -3540 -867 -1960 -864
rect -3540 -901 -3517 -867
rect -3483 -901 -2377 -867
rect -2343 -901 -1960 -867
rect -3540 -904 -1960 -901
rect -1840 -867 -1760 -844
rect -1840 -901 -1817 -867
rect -1783 -901 -1760 -867
rect -1691 -861 -1668 -827
rect -1634 -858 -1611 -827
rect -1419 -735 -1396 -701
rect -1362 -735 -1339 -701
rect -1419 -773 -1339 -735
rect -1419 -807 -1396 -773
rect -1362 -807 -1339 -773
rect -1419 -830 -1339 -807
rect -1549 -858 -1469 -838
rect -1634 -861 -1469 -858
rect -1691 -895 -1526 -861
rect -1492 -895 -1469 -861
rect -1691 -898 -1469 -895
rect -3540 -939 -3460 -904
rect -2400 -924 -2320 -904
rect -1840 -924 -1760 -901
rect -1549 -918 -1469 -898
rect -3540 -973 -3517 -939
rect -3483 -973 -3460 -939
rect -1399 -968 -1359 -830
rect -897 -858 -817 -838
rect -597 -858 -557 -618
rect -357 -858 -277 -838
rect -1295 -861 -817 -858
rect -1295 -895 -874 -861
rect -840 -895 -817 -861
rect -1295 -898 -817 -895
rect -3540 -996 -3460 -973
rect -2420 -979 -2340 -968
rect -2420 -1027 -2397 -979
rect -2363 -1027 -2340 -979
rect -2420 -1051 -2340 -1027
rect -2420 -1095 -2397 -1051
rect -2363 -1095 -2340 -1051
rect -2420 -1123 -2340 -1095
rect -2420 -1163 -2397 -1123
rect -2363 -1163 -2340 -1123
rect -2420 -1195 -2340 -1163
rect -2420 -1231 -2397 -1195
rect -2363 -1231 -2340 -1195
rect -2420 -1265 -2340 -1231
rect -2420 -1301 -2397 -1265
rect -2363 -1301 -2340 -1265
rect -2420 -1333 -2340 -1301
rect -2420 -1373 -2397 -1333
rect -2363 -1373 -2340 -1333
rect -2420 -1401 -2340 -1373
rect -2420 -1445 -2397 -1401
rect -2363 -1445 -2340 -1401
rect -2420 -1469 -2340 -1445
rect -3654 -1529 -3574 -1506
rect -2420 -1517 -2397 -1469
rect -2363 -1517 -2340 -1469
rect -2420 -1528 -2340 -1517
rect -2120 -979 -2040 -968
rect -2120 -1027 -2097 -979
rect -2063 -1027 -2040 -979
rect -2120 -1051 -2040 -1027
rect -2120 -1095 -2097 -1051
rect -2063 -1095 -2040 -1051
rect -2120 -1123 -2040 -1095
rect -2120 -1163 -2097 -1123
rect -2063 -1163 -2040 -1123
rect -2120 -1195 -2040 -1163
rect -2120 -1231 -2097 -1195
rect -2063 -1231 -2040 -1195
rect -2120 -1265 -2040 -1231
rect -2120 -1301 -2097 -1265
rect -2063 -1301 -2040 -1265
rect -2120 -1333 -2040 -1301
rect -2120 -1373 -2097 -1333
rect -2063 -1373 -2040 -1333
rect -2120 -1401 -2040 -1373
rect -2120 -1445 -2097 -1401
rect -2063 -1445 -2040 -1401
rect -2120 -1469 -2040 -1445
rect -2120 -1517 -2097 -1469
rect -2063 -1517 -2040 -1469
rect -2120 -1528 -2040 -1517
rect -1820 -979 -1740 -968
rect -1820 -1027 -1797 -979
rect -1763 -1027 -1740 -979
rect -1820 -1051 -1740 -1027
rect -1820 -1095 -1797 -1051
rect -1763 -1095 -1740 -1051
rect -1820 -1123 -1740 -1095
rect -1820 -1163 -1797 -1123
rect -1763 -1163 -1740 -1123
rect -1820 -1195 -1740 -1163
rect -1820 -1231 -1797 -1195
rect -1763 -1231 -1740 -1195
rect -1820 -1265 -1740 -1231
rect -1820 -1301 -1797 -1265
rect -1763 -1301 -1740 -1265
rect -1820 -1333 -1740 -1301
rect -1820 -1373 -1797 -1333
rect -1763 -1373 -1740 -1333
rect -1820 -1401 -1740 -1373
rect -1820 -1445 -1797 -1401
rect -1763 -1445 -1740 -1401
rect -1820 -1469 -1740 -1445
rect -1820 -1517 -1797 -1469
rect -1763 -1517 -1740 -1469
rect -1820 -1528 -1740 -1517
rect -1569 -979 -1489 -968
rect -1569 -1027 -1546 -979
rect -1512 -1027 -1489 -979
rect -1569 -1051 -1489 -1027
rect -1569 -1095 -1546 -1051
rect -1512 -1095 -1489 -1051
rect -1569 -1123 -1489 -1095
rect -1569 -1163 -1546 -1123
rect -1512 -1163 -1489 -1123
rect -1569 -1195 -1489 -1163
rect -1569 -1231 -1546 -1195
rect -1512 -1231 -1489 -1195
rect -1569 -1265 -1489 -1231
rect -1569 -1301 -1546 -1265
rect -1512 -1301 -1489 -1265
rect -1569 -1333 -1489 -1301
rect -1569 -1373 -1546 -1333
rect -1512 -1373 -1489 -1333
rect -1569 -1401 -1489 -1373
rect -1569 -1445 -1546 -1401
rect -1512 -1445 -1489 -1401
rect -1569 -1469 -1489 -1445
rect -1569 -1517 -1546 -1469
rect -1512 -1517 -1489 -1469
rect -1569 -1528 -1489 -1517
rect -1419 -993 -1339 -968
rect -1419 -1027 -1396 -993
rect -1362 -1027 -1339 -993
rect -1419 -1061 -1339 -1027
rect -1419 -1095 -1396 -1061
rect -1362 -1095 -1339 -1061
rect -1419 -1129 -1339 -1095
rect -1419 -1163 -1396 -1129
rect -1362 -1163 -1339 -1129
rect -1419 -1197 -1339 -1163
rect -1419 -1231 -1396 -1197
rect -1362 -1231 -1339 -1197
rect -1419 -1265 -1339 -1231
rect -1419 -1299 -1396 -1265
rect -1362 -1299 -1339 -1265
rect -1419 -1333 -1339 -1299
rect -1419 -1367 -1396 -1333
rect -1362 -1367 -1339 -1333
rect -1419 -1401 -1339 -1367
rect -1419 -1435 -1396 -1401
rect -1362 -1435 -1339 -1401
rect -1419 -1469 -1339 -1435
rect -1419 -1503 -1396 -1469
rect -1362 -1503 -1339 -1469
rect -1419 -1528 -1339 -1503
rect -3654 -1563 -3631 -1529
rect -3597 -1563 -3574 -1529
rect -3654 -1598 -3574 -1563
rect -1920 -1598 -1840 -1578
rect -3654 -1601 -1840 -1598
rect -3654 -1635 -3631 -1601
rect -3597 -1635 -1897 -1601
rect -1863 -1635 -1840 -1601
rect -3654 -1638 -1840 -1635
rect -3654 -1673 -3574 -1638
rect -1920 -1658 -1840 -1638
rect -1481 -1594 -1329 -1574
rect -1295 -1594 -1255 -898
rect -897 -918 -817 -898
rect -747 -861 -277 -858
rect -747 -895 -334 -861
rect -300 -895 -277 -861
rect -747 -898 -277 -895
rect -747 -968 -707 -898
rect -357 -918 -277 -898
rect -207 -968 -167 -618
rect -81 -701 -1 -678
rect -81 -735 -58 -701
rect -24 -735 -1 -701
rect -81 -773 -1 -735
rect -81 -807 -58 -773
rect -24 -807 -1 -773
rect -81 -830 -1 -807
rect -61 -864 -21 -830
rect 315 -861 395 -838
rect 615 -858 655 -618
rect 855 -858 935 -838
rect 315 -864 338 -861
rect -61 -895 338 -864
rect 372 -895 395 -861
rect -61 -904 395 -895
rect 315 -918 395 -904
rect 465 -861 935 -858
rect 465 -895 878 -861
rect 912 -895 935 -861
rect 465 -898 935 -895
rect 465 -968 505 -898
rect 855 -918 935 -898
rect 1005 -968 1045 -618
rect -917 -979 -837 -968
rect -917 -1027 -894 -979
rect -860 -1027 -837 -979
rect -917 -1051 -837 -1027
rect -917 -1095 -894 -1051
rect -860 -1095 -837 -1051
rect -917 -1123 -837 -1095
rect -917 -1163 -894 -1123
rect -860 -1163 -837 -1123
rect -917 -1195 -837 -1163
rect -917 -1231 -894 -1195
rect -860 -1231 -837 -1195
rect -917 -1265 -837 -1231
rect -917 -1301 -894 -1265
rect -860 -1301 -837 -1265
rect -917 -1333 -837 -1301
rect -917 -1373 -894 -1333
rect -860 -1373 -837 -1333
rect -917 -1401 -837 -1373
rect -917 -1445 -894 -1401
rect -860 -1445 -837 -1401
rect -917 -1469 -837 -1445
rect -917 -1517 -894 -1469
rect -860 -1517 -837 -1469
rect -917 -1528 -837 -1517
rect -767 -993 -687 -968
rect -767 -1027 -744 -993
rect -710 -1027 -687 -993
rect -767 -1061 -687 -1027
rect -767 -1095 -744 -1061
rect -710 -1095 -687 -1061
rect -767 -1129 -687 -1095
rect -767 -1163 -744 -1129
rect -710 -1163 -687 -1129
rect -767 -1197 -687 -1163
rect -767 -1231 -744 -1197
rect -710 -1231 -687 -1197
rect -767 -1265 -687 -1231
rect -767 -1299 -744 -1265
rect -710 -1299 -687 -1265
rect -767 -1333 -687 -1299
rect -767 -1367 -744 -1333
rect -710 -1367 -687 -1333
rect -767 -1401 -687 -1367
rect -767 -1435 -744 -1401
rect -710 -1435 -687 -1401
rect -767 -1469 -687 -1435
rect -767 -1503 -744 -1469
rect -710 -1503 -687 -1469
rect -767 -1528 -687 -1503
rect -617 -979 -537 -968
rect -617 -1027 -594 -979
rect -560 -1027 -537 -979
rect -617 -1051 -537 -1027
rect -617 -1095 -594 -1051
rect -560 -1095 -537 -1051
rect -617 -1123 -537 -1095
rect -617 -1163 -594 -1123
rect -560 -1163 -537 -1123
rect -617 -1195 -537 -1163
rect -617 -1231 -594 -1195
rect -560 -1231 -537 -1195
rect -617 -1265 -537 -1231
rect -617 -1301 -594 -1265
rect -560 -1301 -537 -1265
rect -617 -1333 -537 -1301
rect -617 -1373 -594 -1333
rect -560 -1373 -537 -1333
rect -617 -1401 -537 -1373
rect -617 -1445 -594 -1401
rect -560 -1445 -537 -1401
rect -617 -1469 -537 -1445
rect -617 -1517 -594 -1469
rect -560 -1517 -537 -1469
rect -617 -1528 -537 -1517
rect -377 -979 -297 -968
rect -377 -1027 -354 -979
rect -320 -1027 -297 -979
rect -377 -1051 -297 -1027
rect -377 -1095 -354 -1051
rect -320 -1095 -297 -1051
rect -377 -1123 -297 -1095
rect -377 -1163 -354 -1123
rect -320 -1163 -297 -1123
rect -377 -1195 -297 -1163
rect -377 -1231 -354 -1195
rect -320 -1231 -297 -1195
rect -377 -1265 -297 -1231
rect -377 -1301 -354 -1265
rect -320 -1301 -297 -1265
rect -377 -1333 -297 -1301
rect -377 -1373 -354 -1333
rect -320 -1373 -297 -1333
rect -377 -1401 -297 -1373
rect -377 -1445 -354 -1401
rect -320 -1445 -297 -1401
rect -377 -1469 -297 -1445
rect -377 -1517 -354 -1469
rect -320 -1517 -297 -1469
rect -377 -1528 -297 -1517
rect -227 -993 -147 -968
rect -227 -1027 -204 -993
rect -170 -1027 -147 -993
rect -227 -1061 -147 -1027
rect -227 -1095 -204 -1061
rect -170 -1095 -147 -1061
rect -227 -1129 -147 -1095
rect -227 -1163 -204 -1129
rect -170 -1163 -147 -1129
rect -227 -1197 -147 -1163
rect -227 -1231 -204 -1197
rect -170 -1231 -147 -1197
rect -227 -1265 -147 -1231
rect -227 -1299 -204 -1265
rect -170 -1299 -147 -1265
rect -227 -1333 -147 -1299
rect -227 -1367 -204 -1333
rect -170 -1367 -147 -1333
rect -227 -1401 -147 -1367
rect -227 -1435 -204 -1401
rect -170 -1435 -147 -1401
rect -227 -1469 -147 -1435
rect -227 -1503 -204 -1469
rect -170 -1503 -147 -1469
rect -227 -1528 -147 -1503
rect 295 -979 375 -968
rect 295 -1027 318 -979
rect 352 -1027 375 -979
rect 295 -1051 375 -1027
rect 295 -1095 318 -1051
rect 352 -1095 375 -1051
rect 295 -1123 375 -1095
rect 295 -1163 318 -1123
rect 352 -1163 375 -1123
rect 295 -1195 375 -1163
rect 295 -1231 318 -1195
rect 352 -1231 375 -1195
rect 295 -1265 375 -1231
rect 295 -1301 318 -1265
rect 352 -1301 375 -1265
rect 295 -1333 375 -1301
rect 295 -1373 318 -1333
rect 352 -1373 375 -1333
rect 295 -1401 375 -1373
rect 295 -1445 318 -1401
rect 352 -1445 375 -1401
rect 295 -1469 375 -1445
rect 295 -1517 318 -1469
rect 352 -1517 375 -1469
rect 295 -1528 375 -1517
rect 445 -993 525 -968
rect 445 -1027 468 -993
rect 502 -1027 525 -993
rect 445 -1061 525 -1027
rect 445 -1095 468 -1061
rect 502 -1095 525 -1061
rect 445 -1129 525 -1095
rect 445 -1163 468 -1129
rect 502 -1163 525 -1129
rect 445 -1197 525 -1163
rect 445 -1231 468 -1197
rect 502 -1231 525 -1197
rect 445 -1265 525 -1231
rect 445 -1299 468 -1265
rect 502 -1299 525 -1265
rect 445 -1333 525 -1299
rect 445 -1367 468 -1333
rect 502 -1367 525 -1333
rect 445 -1401 525 -1367
rect 445 -1435 468 -1401
rect 502 -1435 525 -1401
rect 445 -1469 525 -1435
rect 445 -1503 468 -1469
rect 502 -1503 525 -1469
rect 445 -1528 525 -1503
rect 595 -979 675 -968
rect 595 -1027 618 -979
rect 652 -1027 675 -979
rect 595 -1051 675 -1027
rect 595 -1095 618 -1051
rect 652 -1095 675 -1051
rect 595 -1123 675 -1095
rect 595 -1163 618 -1123
rect 652 -1163 675 -1123
rect 595 -1195 675 -1163
rect 595 -1231 618 -1195
rect 652 -1231 675 -1195
rect 595 -1265 675 -1231
rect 595 -1301 618 -1265
rect 652 -1301 675 -1265
rect 595 -1333 675 -1301
rect 595 -1373 618 -1333
rect 652 -1373 675 -1333
rect 595 -1401 675 -1373
rect 595 -1445 618 -1401
rect 652 -1445 675 -1401
rect 595 -1469 675 -1445
rect 595 -1517 618 -1469
rect 652 -1517 675 -1469
rect 595 -1528 675 -1517
rect 835 -979 915 -968
rect 835 -1027 858 -979
rect 892 -1027 915 -979
rect 835 -1051 915 -1027
rect 835 -1095 858 -1051
rect 892 -1095 915 -1051
rect 835 -1123 915 -1095
rect 835 -1163 858 -1123
rect 892 -1163 915 -1123
rect 835 -1195 915 -1163
rect 835 -1231 858 -1195
rect 892 -1231 915 -1195
rect 835 -1265 915 -1231
rect 835 -1301 858 -1265
rect 892 -1301 915 -1265
rect 835 -1333 915 -1301
rect 835 -1373 858 -1333
rect 892 -1373 915 -1333
rect 835 -1401 915 -1373
rect 835 -1445 858 -1401
rect 892 -1445 915 -1401
rect 835 -1469 915 -1445
rect 835 -1517 858 -1469
rect 892 -1517 915 -1469
rect 835 -1528 915 -1517
rect 985 -993 1065 -968
rect 985 -1027 1008 -993
rect 1042 -1027 1065 -993
rect 985 -1061 1065 -1027
rect 985 -1095 1008 -1061
rect 1042 -1095 1065 -1061
rect 985 -1129 1065 -1095
rect 985 -1163 1008 -1129
rect 1042 -1163 1065 -1129
rect 985 -1197 1065 -1163
rect 985 -1231 1008 -1197
rect 1042 -1231 1065 -1197
rect 985 -1265 1065 -1231
rect 985 -1299 1008 -1265
rect 1042 -1299 1065 -1265
rect 985 -1333 1065 -1299
rect 985 -1367 1008 -1333
rect 1042 -1367 1065 -1333
rect 985 -1401 1065 -1367
rect 985 -1435 1008 -1401
rect 1042 -1435 1065 -1401
rect 985 -1469 1065 -1435
rect 985 -1503 1008 -1469
rect 1042 -1503 1065 -1469
rect 985 -1528 1065 -1503
rect -1481 -1597 -1255 -1594
rect -1481 -1631 -1458 -1597
rect -1424 -1631 -1386 -1597
rect -1352 -1631 -1255 -1597
rect -1481 -1634 -1255 -1631
rect -1481 -1654 -1329 -1634
rect -3654 -1707 -3631 -1673
rect -3597 -1707 -3574 -1673
rect -3654 -1730 -3574 -1707
rect -2520 -1715 -1294 -1692
rect -2520 -1749 -2497 -1715
rect -2463 -1749 -2425 -1715
rect -2391 -1749 -2353 -1715
rect -2319 -1749 -2281 -1715
rect -2247 -1749 -2209 -1715
rect -2175 -1749 -2137 -1715
rect -2103 -1749 -2065 -1715
rect -2031 -1749 -1993 -1715
rect -1959 -1749 -1921 -1715
rect -1887 -1749 -1849 -1715
rect -1815 -1749 -1777 -1715
rect -1743 -1749 -1705 -1715
rect -1671 -1749 -1633 -1715
rect -1599 -1749 -1561 -1715
rect -1527 -1749 -1489 -1715
rect -1455 -1749 -1417 -1715
rect -1383 -1749 -1345 -1715
rect -1311 -1749 -1294 -1715
rect -2520 -1772 -1294 -1749
rect -962 -1715 -82 -1692
rect -962 -1749 -939 -1715
rect -905 -1749 -867 -1715
rect -833 -1749 -795 -1715
rect -761 -1749 -723 -1715
rect -689 -1749 -651 -1715
rect -617 -1749 -579 -1715
rect -545 -1749 -507 -1715
rect -473 -1749 -435 -1715
rect -401 -1749 -363 -1715
rect -329 -1749 -291 -1715
rect -257 -1749 -219 -1715
rect -185 -1749 -147 -1715
rect -113 -1749 -82 -1715
rect -962 -1772 -82 -1749
rect 250 -1715 1130 -1692
rect 250 -1749 273 -1715
rect 307 -1749 345 -1715
rect 379 -1749 417 -1715
rect 451 -1749 489 -1715
rect 523 -1749 561 -1715
rect 595 -1749 633 -1715
rect 667 -1749 705 -1715
rect 739 -1749 777 -1715
rect 811 -1749 849 -1715
rect 883 -1749 921 -1715
rect 955 -1749 993 -1715
rect 1027 -1749 1065 -1715
rect 1099 -1749 1130 -1715
rect 250 -1772 1130 -1749
<< viali >>
rect -2947 1365 -2913 1399
rect -2497 1407 -2463 1441
rect -2425 1407 -2391 1441
rect -2353 1407 -2319 1441
rect -2281 1407 -2247 1441
rect -2209 1407 -2175 1441
rect -2137 1407 -2103 1441
rect -2065 1407 -2031 1441
rect -1993 1407 -1959 1441
rect -1921 1407 -1887 1441
rect -1849 1407 -1815 1441
rect -1777 1407 -1743 1441
rect -1705 1407 -1671 1441
rect -939 1407 -905 1441
rect -867 1407 -833 1441
rect -795 1407 -761 1441
rect -723 1407 -689 1441
rect -651 1407 -617 1441
rect -579 1407 -545 1441
rect -507 1407 -473 1441
rect -435 1407 -401 1441
rect -363 1407 -329 1441
rect -291 1407 -257 1441
rect -219 1407 -185 1441
rect -147 1407 -113 1441
rect 273 1407 307 1441
rect 345 1407 379 1441
rect 417 1407 451 1441
rect 489 1407 523 1441
rect 561 1407 595 1441
rect 633 1407 667 1441
rect 705 1407 739 1441
rect 777 1407 811 1441
rect 849 1407 883 1441
rect 921 1407 955 1441
rect 993 1407 1027 1441
rect 1065 1407 1099 1441
rect 1485 1407 1519 1441
rect 1557 1407 1591 1441
rect 1629 1407 1663 1441
rect 1701 1407 1735 1441
rect 1773 1407 1807 1441
rect 1845 1407 1879 1441
rect 1917 1407 1951 1441
rect 1989 1407 2023 1441
rect 2061 1407 2095 1441
rect 2133 1407 2167 1441
rect 2205 1407 2239 1441
rect 2277 1407 2311 1441
rect -2947 1293 -2913 1327
rect -1683 1289 -1649 1323
rect -1611 1289 -1577 1323
rect -2947 1221 -2913 1255
rect -2397 1195 -2363 1209
rect -2397 1175 -2363 1195
rect -2397 1127 -2363 1137
rect -2397 1103 -2363 1127
rect -2397 1059 -2363 1065
rect -2397 1031 -2363 1059
rect -2397 991 -2363 993
rect -2397 959 -2363 991
rect -2397 889 -2363 921
rect -2397 887 -2363 889
rect -2397 821 -2363 849
rect -2397 815 -2363 821
rect -2397 753 -2363 777
rect -2397 743 -2363 753
rect -2833 631 -2799 665
rect -2397 685 -2363 705
rect -2397 671 -2363 685
rect -2097 1195 -2063 1209
rect -2097 1175 -2063 1195
rect -2097 1127 -2063 1137
rect -2097 1103 -2063 1127
rect -2097 1059 -2063 1065
rect -2097 1031 -2063 1059
rect -2097 991 -2063 993
rect -2097 959 -2063 991
rect -2097 889 -2063 921
rect -2097 887 -2063 889
rect -2097 821 -2063 849
rect -2097 815 -2063 821
rect -2097 753 -2063 777
rect -2097 743 -2063 753
rect -2097 685 -2063 705
rect -2097 671 -2063 685
rect -1797 1195 -1763 1209
rect -1797 1175 -1763 1195
rect -1797 1127 -1763 1137
rect -1797 1103 -1763 1127
rect -1797 1059 -1763 1065
rect -1797 1031 -1763 1059
rect -1797 991 -1763 993
rect -1797 959 -1763 991
rect -1797 889 -1763 921
rect -1797 887 -1763 889
rect -1797 821 -1763 849
rect -1797 815 -1763 821
rect -1797 753 -1763 777
rect -1797 743 -1763 753
rect -1797 685 -1763 705
rect -1797 671 -1763 685
rect -2833 559 -2799 593
rect -3631 440 -3597 474
rect -2833 487 -2799 521
rect -1817 559 -1783 593
rect -894 1195 -860 1209
rect -894 1175 -860 1195
rect -894 1127 -860 1137
rect -894 1103 -860 1127
rect -894 1059 -860 1065
rect -894 1031 -860 1059
rect -894 991 -860 993
rect -894 959 -860 991
rect -894 889 -860 921
rect -894 887 -860 889
rect -894 821 -860 849
rect -894 815 -860 821
rect -894 753 -860 777
rect -894 743 -860 753
rect -894 685 -860 705
rect -894 671 -860 685
rect -354 1195 -320 1209
rect -354 1175 -320 1195
rect -354 1127 -320 1137
rect -354 1103 -320 1127
rect -354 1059 -320 1065
rect -354 1031 -320 1059
rect -354 991 -320 993
rect -354 959 -320 991
rect -354 889 -320 921
rect -354 887 -320 889
rect -354 821 -320 849
rect -354 815 -320 821
rect -354 753 -320 777
rect -354 743 -320 753
rect -354 685 -320 705
rect -354 671 -320 685
rect 318 1195 352 1209
rect 318 1175 352 1195
rect 318 1127 352 1137
rect 318 1103 352 1127
rect 318 1059 352 1065
rect 318 1031 352 1059
rect 318 991 352 993
rect 318 959 352 991
rect 318 889 352 921
rect 318 887 352 889
rect 318 821 352 849
rect 318 815 352 821
rect 318 753 352 777
rect 318 743 352 753
rect 318 685 352 705
rect 318 671 352 685
rect 618 1195 652 1209
rect 618 1175 652 1195
rect 618 1127 652 1137
rect 618 1103 652 1127
rect 618 1059 652 1065
rect 618 1031 652 1059
rect 618 991 652 993
rect 618 959 652 991
rect 618 889 652 921
rect 618 887 652 889
rect 618 821 652 849
rect 618 815 652 821
rect 618 753 652 777
rect 618 743 652 753
rect 618 685 652 705
rect 618 671 652 685
rect 858 1195 892 1209
rect 858 1175 892 1195
rect 858 1127 892 1137
rect 858 1103 892 1127
rect 858 1059 892 1065
rect 858 1031 892 1059
rect 858 991 892 993
rect 858 959 892 991
rect 858 889 892 921
rect 858 887 892 889
rect 858 821 892 849
rect 858 815 892 821
rect 858 753 892 777
rect 858 743 892 753
rect 858 685 892 705
rect 858 671 892 685
rect 1530 1195 1564 1209
rect 1530 1175 1564 1195
rect 1530 1127 1564 1137
rect 1530 1103 1564 1127
rect 1530 1059 1564 1065
rect 1530 1031 1564 1059
rect 1530 991 1564 993
rect 1530 959 1564 991
rect 1530 889 1564 921
rect 1530 887 1564 889
rect 1530 821 1564 849
rect 1530 815 1564 821
rect 1530 753 1564 777
rect 1530 743 1564 753
rect 1530 685 1564 705
rect 1530 671 1564 685
rect 2070 1195 2104 1209
rect 2070 1175 2104 1195
rect 2070 1127 2104 1137
rect 2070 1103 2104 1127
rect 2070 1059 2104 1065
rect 2070 1031 2104 1059
rect 2070 991 2104 993
rect 2070 959 2104 991
rect 2070 889 2104 921
rect 2070 887 2104 889
rect 2070 821 2104 849
rect 2070 815 2104 821
rect 2070 753 2104 777
rect 2070 743 2104 753
rect 2070 685 2104 705
rect 2070 671 2104 685
rect -3631 368 -3597 402
rect -2197 368 -2163 402
rect -3631 296 -3597 330
rect -58 465 -24 499
rect -2397 265 -2363 269
rect -2397 235 -2363 265
rect -2397 163 -2363 197
rect -2397 95 -2363 125
rect -2397 91 -2363 95
rect -2097 265 -2063 269
rect -2097 235 -2063 265
rect -2097 163 -2063 197
rect -2097 95 -2063 125
rect -2097 91 -2063 95
rect -1797 265 -1763 269
rect -1797 235 -1763 265
rect -1797 163 -1763 197
rect -1797 95 -1763 125
rect -1797 91 -1763 95
rect -894 265 -860 269
rect -894 235 -860 265
rect -894 163 -860 197
rect -894 95 -860 125
rect -894 91 -860 95
rect -594 265 -560 269
rect -594 235 -560 265
rect -594 163 -560 197
rect -594 95 -560 125
rect -594 91 -560 95
rect -354 265 -320 269
rect -354 235 -320 265
rect -354 163 -320 197
rect -354 95 -320 125
rect -354 91 -320 95
rect -3517 15 -3483 49
rect -3517 -57 -3483 -23
rect -3517 -129 -3483 -95
rect -2719 -99 -2685 -65
rect -1683 -53 -1649 -19
rect -1611 -53 -1577 -19
rect 2220 491 2254 525
rect 2220 419 2254 453
rect 318 265 352 269
rect 318 235 352 265
rect 318 163 352 197
rect 318 95 352 125
rect 318 91 352 95
rect 858 265 892 269
rect 858 235 892 265
rect 858 163 892 197
rect 858 95 892 125
rect 858 91 892 95
rect 1530 265 1564 269
rect 1530 235 1564 265
rect 1530 163 1564 197
rect 1530 95 1564 125
rect 1530 91 1564 95
rect 1830 265 1864 269
rect 1830 235 1864 265
rect 1830 163 1864 197
rect 1830 95 1864 125
rect 1830 91 1864 95
rect 2070 265 2104 269
rect 2070 235 2104 265
rect 2070 163 2104 197
rect 2070 95 2104 125
rect 2070 91 2104 95
rect -2833 -213 -2799 -179
rect -2833 -285 -2799 -251
rect -2719 -171 -2685 -137
rect -2497 -171 -2463 -137
rect -2425 -171 -2391 -137
rect -2353 -171 -2319 -137
rect -2281 -171 -2247 -137
rect -2209 -171 -2175 -137
rect -2137 -171 -2103 -137
rect -2065 -171 -2031 -137
rect -1993 -171 -1959 -137
rect -1921 -171 -1887 -137
rect -1849 -171 -1815 -137
rect -1777 -171 -1743 -137
rect -1705 -171 -1671 -137
rect -1633 -171 -1599 -137
rect -1561 -171 -1527 -137
rect -1489 -171 -1455 -137
rect -1417 -171 -1383 -137
rect -1345 -171 -1311 -137
rect -939 -171 -905 -137
rect -867 -171 -833 -137
rect -795 -171 -761 -137
rect -723 -171 -689 -137
rect -651 -171 -617 -137
rect -579 -171 -545 -137
rect -507 -171 -473 -137
rect -435 -171 -401 -137
rect -363 -171 -329 -137
rect -291 -171 -257 -137
rect -219 -171 -185 -137
rect -147 -171 -113 -137
rect 273 -171 307 -137
rect 345 -171 379 -137
rect 417 -171 451 -137
rect 489 -171 523 -137
rect 561 -171 595 -137
rect 633 -171 667 -137
rect 705 -171 739 -137
rect 777 -171 811 -137
rect 849 -171 883 -137
rect 921 -171 955 -137
rect 993 -171 1027 -137
rect 1065 -171 1099 -137
rect -2719 -243 -2685 -209
rect -1458 -289 -1424 -255
rect -1386 -289 -1352 -255
rect -2833 -357 -2799 -323
rect 1485 -171 1519 -137
rect 1557 -171 1591 -137
rect 1629 -171 1663 -137
rect 1701 -171 1735 -137
rect 1773 -171 1807 -137
rect 1845 -171 1879 -137
rect 1917 -171 1951 -137
rect 1989 -171 2023 -137
rect 2061 -171 2095 -137
rect 2133 -171 2167 -137
rect 2205 -171 2239 -137
rect 2277 -171 2311 -137
rect -2397 -403 -2363 -399
rect -2397 -433 -2363 -403
rect -2397 -505 -2363 -471
rect -2947 -638 -2913 -604
rect -2397 -573 -2363 -543
rect -2397 -577 -2363 -573
rect -2097 -403 -2063 -399
rect -2097 -433 -2063 -403
rect -2097 -505 -2063 -471
rect -2097 -573 -2063 -543
rect -2097 -577 -2063 -573
rect -1797 -403 -1763 -399
rect -1797 -433 -1763 -403
rect -1797 -505 -1763 -471
rect -1797 -573 -1763 -543
rect -1797 -577 -1763 -573
rect -1546 -403 -1512 -399
rect -1546 -433 -1512 -403
rect -1546 -505 -1512 -471
rect -1546 -573 -1512 -543
rect -1546 -577 -1512 -573
rect -894 -403 -860 -399
rect -894 -433 -860 -403
rect -894 -505 -860 -471
rect -894 -573 -860 -543
rect -894 -577 -860 -573
rect -354 -403 -320 -399
rect -354 -433 -320 -403
rect -354 -505 -320 -471
rect -354 -573 -320 -543
rect -354 -577 -320 -573
rect 318 -403 352 -399
rect 318 -433 352 -403
rect 318 -505 352 -471
rect 318 -573 352 -543
rect 318 -577 352 -573
rect 858 -403 892 -399
rect 858 -433 892 -403
rect 858 -505 892 -471
rect 858 -573 892 -543
rect 858 -577 892 -573
rect -2947 -710 -2913 -676
rect -2197 -710 -2163 -676
rect -3517 -829 -3483 -795
rect -2947 -782 -2913 -748
rect -1668 -789 -1634 -755
rect -3517 -901 -3483 -867
rect -1817 -901 -1783 -867
rect -1668 -861 -1634 -827
rect -1396 -735 -1362 -701
rect -1396 -807 -1362 -773
rect -3517 -973 -3483 -939
rect -2397 -993 -2363 -979
rect -2397 -1013 -2363 -993
rect -2397 -1061 -2363 -1051
rect -2397 -1085 -2363 -1061
rect -2397 -1129 -2363 -1123
rect -2397 -1157 -2363 -1129
rect -2397 -1197 -2363 -1195
rect -2397 -1229 -2363 -1197
rect -2397 -1299 -2363 -1267
rect -2397 -1301 -2363 -1299
rect -2397 -1367 -2363 -1339
rect -2397 -1373 -2363 -1367
rect -2397 -1435 -2363 -1411
rect -2397 -1445 -2363 -1435
rect -2397 -1503 -2363 -1483
rect -2397 -1517 -2363 -1503
rect -2097 -993 -2063 -979
rect -2097 -1013 -2063 -993
rect -2097 -1061 -2063 -1051
rect -2097 -1085 -2063 -1061
rect -2097 -1129 -2063 -1123
rect -2097 -1157 -2063 -1129
rect -2097 -1197 -2063 -1195
rect -2097 -1229 -2063 -1197
rect -2097 -1299 -2063 -1267
rect -2097 -1301 -2063 -1299
rect -2097 -1367 -2063 -1339
rect -2097 -1373 -2063 -1367
rect -2097 -1435 -2063 -1411
rect -2097 -1445 -2063 -1435
rect -2097 -1503 -2063 -1483
rect -2097 -1517 -2063 -1503
rect -1797 -993 -1763 -979
rect -1797 -1013 -1763 -993
rect -1797 -1061 -1763 -1051
rect -1797 -1085 -1763 -1061
rect -1797 -1129 -1763 -1123
rect -1797 -1157 -1763 -1129
rect -1797 -1197 -1763 -1195
rect -1797 -1229 -1763 -1197
rect -1797 -1299 -1763 -1267
rect -1797 -1301 -1763 -1299
rect -1797 -1367 -1763 -1339
rect -1797 -1373 -1763 -1367
rect -1797 -1435 -1763 -1411
rect -1797 -1445 -1763 -1435
rect -1797 -1503 -1763 -1483
rect -1797 -1517 -1763 -1503
rect -1546 -993 -1512 -979
rect -1546 -1013 -1512 -993
rect -1546 -1061 -1512 -1051
rect -1546 -1085 -1512 -1061
rect -1546 -1129 -1512 -1123
rect -1546 -1157 -1512 -1129
rect -1546 -1197 -1512 -1195
rect -1546 -1229 -1512 -1197
rect -1546 -1299 -1512 -1267
rect -1546 -1301 -1512 -1299
rect -1546 -1367 -1512 -1339
rect -1546 -1373 -1512 -1367
rect -1546 -1435 -1512 -1411
rect -1546 -1445 -1512 -1435
rect -1546 -1503 -1512 -1483
rect -1546 -1517 -1512 -1503
rect -3631 -1563 -3597 -1529
rect -3631 -1635 -3597 -1601
rect -58 -735 -24 -701
rect -58 -807 -24 -773
rect -894 -993 -860 -979
rect -894 -1013 -860 -993
rect -894 -1061 -860 -1051
rect -894 -1085 -860 -1061
rect -894 -1129 -860 -1123
rect -894 -1157 -860 -1129
rect -894 -1197 -860 -1195
rect -894 -1229 -860 -1197
rect -894 -1299 -860 -1267
rect -894 -1301 -860 -1299
rect -894 -1367 -860 -1339
rect -894 -1373 -860 -1367
rect -894 -1435 -860 -1411
rect -894 -1445 -860 -1435
rect -894 -1503 -860 -1483
rect -894 -1517 -860 -1503
rect -594 -993 -560 -979
rect -594 -1013 -560 -993
rect -594 -1061 -560 -1051
rect -594 -1085 -560 -1061
rect -594 -1129 -560 -1123
rect -594 -1157 -560 -1129
rect -594 -1197 -560 -1195
rect -594 -1229 -560 -1197
rect -594 -1299 -560 -1267
rect -594 -1301 -560 -1299
rect -594 -1367 -560 -1339
rect -594 -1373 -560 -1367
rect -594 -1435 -560 -1411
rect -594 -1445 -560 -1435
rect -594 -1503 -560 -1483
rect -594 -1517 -560 -1503
rect -354 -993 -320 -979
rect -354 -1013 -320 -993
rect -354 -1061 -320 -1051
rect -354 -1085 -320 -1061
rect -354 -1129 -320 -1123
rect -354 -1157 -320 -1129
rect -354 -1197 -320 -1195
rect -354 -1229 -320 -1197
rect -354 -1299 -320 -1267
rect -354 -1301 -320 -1299
rect -354 -1367 -320 -1339
rect -354 -1373 -320 -1367
rect -354 -1435 -320 -1411
rect -354 -1445 -320 -1435
rect -354 -1503 -320 -1483
rect -354 -1517 -320 -1503
rect 318 -993 352 -979
rect 318 -1013 352 -993
rect 318 -1061 352 -1051
rect 318 -1085 352 -1061
rect 318 -1129 352 -1123
rect 318 -1157 352 -1129
rect 318 -1197 352 -1195
rect 318 -1229 352 -1197
rect 318 -1299 352 -1267
rect 318 -1301 352 -1299
rect 318 -1367 352 -1339
rect 318 -1373 352 -1367
rect 318 -1435 352 -1411
rect 318 -1445 352 -1435
rect 318 -1503 352 -1483
rect 318 -1517 352 -1503
rect 618 -993 652 -979
rect 618 -1013 652 -993
rect 618 -1061 652 -1051
rect 618 -1085 652 -1061
rect 618 -1129 652 -1123
rect 618 -1157 652 -1129
rect 618 -1197 652 -1195
rect 618 -1229 652 -1197
rect 618 -1299 652 -1267
rect 618 -1301 652 -1299
rect 618 -1367 652 -1339
rect 618 -1373 652 -1367
rect 618 -1435 652 -1411
rect 618 -1445 652 -1435
rect 618 -1503 652 -1483
rect 618 -1517 652 -1503
rect 858 -993 892 -979
rect 858 -1013 892 -993
rect 858 -1061 892 -1051
rect 858 -1085 892 -1061
rect 858 -1129 892 -1123
rect 858 -1157 892 -1129
rect 858 -1197 892 -1195
rect 858 -1229 892 -1197
rect 858 -1299 892 -1267
rect 858 -1301 892 -1299
rect 858 -1367 892 -1339
rect 858 -1373 892 -1367
rect 858 -1435 892 -1411
rect 858 -1445 892 -1435
rect 858 -1503 892 -1483
rect 858 -1517 892 -1503
rect -1458 -1631 -1424 -1597
rect -1386 -1631 -1352 -1597
rect -3631 -1707 -3597 -1673
rect -2497 -1749 -2463 -1715
rect -2425 -1749 -2391 -1715
rect -2353 -1749 -2319 -1715
rect -2281 -1749 -2247 -1715
rect -2209 -1749 -2175 -1715
rect -2137 -1749 -2103 -1715
rect -2065 -1749 -2031 -1715
rect -1993 -1749 -1959 -1715
rect -1921 -1749 -1887 -1715
rect -1849 -1749 -1815 -1715
rect -1777 -1749 -1743 -1715
rect -1705 -1749 -1671 -1715
rect -1633 -1749 -1599 -1715
rect -1561 -1749 -1527 -1715
rect -1489 -1749 -1455 -1715
rect -1417 -1749 -1383 -1715
rect -1345 -1749 -1311 -1715
rect -939 -1749 -905 -1715
rect -867 -1749 -833 -1715
rect -795 -1749 -761 -1715
rect -723 -1749 -689 -1715
rect -651 -1749 -617 -1715
rect -579 -1749 -545 -1715
rect -507 -1749 -473 -1715
rect -435 -1749 -401 -1715
rect -363 -1749 -329 -1715
rect -291 -1749 -257 -1715
rect -219 -1749 -185 -1715
rect -147 -1749 -113 -1715
rect 273 -1749 307 -1715
rect 345 -1749 379 -1715
rect 417 -1749 451 -1715
rect 489 -1749 523 -1715
rect 561 -1749 595 -1715
rect 633 -1749 667 -1715
rect 705 -1749 739 -1715
rect 777 -1749 811 -1715
rect 849 -1749 883 -1715
rect 921 -1749 955 -1715
rect 993 -1749 1027 -1715
rect 1065 -1749 1099 -1715
<< metal1 >>
rect -3654 474 -3574 1474
rect -3654 440 -3631 474
rect -3597 440 -3574 474
rect -3654 402 -3574 440
rect -3654 368 -3631 402
rect -3597 368 -3574 402
rect -3654 330 -3574 368
rect -3654 296 -3631 330
rect -3597 296 -3574 330
rect -3654 -1529 -3574 296
rect -3654 -1563 -3631 -1529
rect -3597 -1563 -3574 -1529
rect -3654 -1601 -3574 -1563
rect -3654 -1635 -3631 -1601
rect -3597 -1635 -3574 -1601
rect -3654 -1673 -3574 -1635
rect -3654 -1707 -3631 -1673
rect -3597 -1707 -3574 -1673
rect -3654 -1783 -3574 -1707
rect -3540 49 -3460 1474
rect -3540 15 -3517 49
rect -3483 15 -3460 49
rect -3540 -23 -3460 15
rect -3540 -57 -3517 -23
rect -3483 -57 -3460 -23
rect -3540 -95 -3460 -57
rect -3540 -129 -3517 -95
rect -3483 -129 -3460 -95
rect -3540 -795 -3460 -129
rect -3540 -829 -3517 -795
rect -3483 -829 -3460 -795
rect -3540 -867 -3460 -829
rect -3540 -901 -3517 -867
rect -3483 -901 -3460 -867
rect -3540 -939 -3460 -901
rect -3540 -973 -3517 -939
rect -3483 -973 -3460 -939
rect -3540 -1783 -3460 -973
rect -3426 1400 -3346 1474
rect -3426 1348 -3412 1400
rect -3360 1348 -3346 1400
rect -3426 1332 -3346 1348
rect -3426 1280 -3412 1332
rect -3360 1280 -3346 1332
rect -3426 1264 -3346 1280
rect -3426 1212 -3412 1264
rect -3360 1212 -3346 1264
rect -3426 -1783 -3346 1212
rect -3312 -1524 -3232 1474
rect -3312 -1576 -3298 -1524
rect -3246 -1576 -3232 -1524
rect -3312 -1592 -3232 -1576
rect -3312 -1644 -3298 -1592
rect -3246 -1644 -3232 -1592
rect -3312 -1660 -3232 -1644
rect -3312 -1712 -3298 -1660
rect -3246 -1712 -3232 -1660
rect -3312 -1783 -3232 -1712
rect -3198 -178 -3118 1474
rect -3198 -230 -3184 -178
rect -3132 -230 -3118 -178
rect -3198 -246 -3118 -230
rect -3198 -298 -3184 -246
rect -3132 -298 -3118 -246
rect -3198 -314 -3118 -298
rect -3198 -366 -3184 -314
rect -3132 -366 -3118 -314
rect -3198 -1782 -3118 -366
rect -3084 58 -3004 1474
rect -3084 6 -3070 58
rect -3018 6 -3004 58
rect -3084 -10 -3004 6
rect -3084 -62 -3070 -10
rect -3018 -62 -3004 -10
rect -3084 -78 -3004 -62
rect -3084 -130 -3070 -78
rect -3018 -130 -3004 -78
rect -3084 -1783 -3004 -130
rect -2970 1399 -2890 1474
rect -2970 1365 -2947 1399
rect -2913 1365 -2890 1399
rect -2970 1327 -2890 1365
rect -2970 1293 -2947 1327
rect -2913 1293 -2890 1327
rect -2970 1255 -2890 1293
rect -2970 1221 -2947 1255
rect -2913 1221 -2890 1255
rect -2970 -604 -2890 1221
rect -2970 -638 -2947 -604
rect -2913 -638 -2890 -604
rect -2970 -676 -2890 -638
rect -2970 -710 -2947 -676
rect -2913 -710 -2890 -676
rect -2970 -748 -2890 -710
rect -2970 -782 -2947 -748
rect -2913 -782 -2890 -748
rect -2970 -1782 -2890 -782
rect -2856 665 -2776 1474
rect -2856 631 -2833 665
rect -2799 631 -2776 665
rect -2856 593 -2776 631
rect -2856 559 -2833 593
rect -2799 559 -2776 593
rect -2856 521 -2776 559
rect -2856 487 -2833 521
rect -2799 487 -2776 521
rect -2856 -179 -2776 487
rect -2856 -213 -2833 -179
rect -2799 -213 -2776 -179
rect -2856 -251 -2776 -213
rect -2856 -285 -2833 -251
rect -2799 -285 -2776 -251
rect -2856 -323 -2776 -285
rect -2856 -357 -2833 -323
rect -2799 -357 -2776 -323
rect -2856 -1782 -2776 -357
rect -2742 -65 -2662 1474
rect -2742 -99 -2719 -65
rect -2685 -99 -2662 -65
rect -2742 -137 -2662 -99
rect -2742 -171 -2719 -137
rect -2685 -171 -2662 -137
rect -2742 -209 -2662 -171
rect -2742 -243 -2719 -209
rect -2685 -243 -2662 -209
rect -2742 -1782 -2662 -243
rect -2628 1441 2342 1474
rect -2628 1407 -2497 1441
rect -2463 1407 -2425 1441
rect -2391 1407 -2353 1441
rect -2319 1407 -2281 1441
rect -2247 1407 -2209 1441
rect -2175 1407 -2137 1441
rect -2103 1407 -2065 1441
rect -2031 1407 -1993 1441
rect -1959 1407 -1921 1441
rect -1887 1407 -1849 1441
rect -1815 1407 -1777 1441
rect -1743 1407 -1705 1441
rect -1671 1407 -939 1441
rect -905 1407 -867 1441
rect -833 1407 -795 1441
rect -761 1407 -723 1441
rect -689 1407 -651 1441
rect -617 1407 -579 1441
rect -545 1407 -507 1441
rect -473 1407 -435 1441
rect -401 1407 -363 1441
rect -329 1407 -291 1441
rect -257 1407 -219 1441
rect -185 1407 -147 1441
rect -113 1407 273 1441
rect 307 1407 345 1441
rect 379 1407 417 1441
rect 451 1407 489 1441
rect 523 1407 561 1441
rect 595 1407 633 1441
rect 667 1407 705 1441
rect 739 1407 777 1441
rect 811 1407 849 1441
rect 883 1407 921 1441
rect 955 1407 993 1441
rect 1027 1407 1065 1441
rect 1099 1407 1485 1441
rect 1519 1407 1557 1441
rect 1591 1407 1629 1441
rect 1663 1407 1701 1441
rect 1735 1407 1773 1441
rect 1807 1407 1845 1441
rect 1879 1407 1917 1441
rect 1951 1407 1989 1441
rect 2023 1407 2061 1441
rect 2095 1407 2133 1441
rect 2167 1407 2205 1441
rect 2239 1407 2277 1441
rect 2311 1407 2342 1441
rect -2628 1374 2342 1407
rect -2628 -1682 -2548 1374
rect -2400 1220 -2360 1374
rect -1800 1220 -1760 1374
rect -1706 1332 -1554 1346
rect -1706 1280 -1692 1332
rect -1640 1280 -1620 1332
rect -1568 1280 -1554 1332
rect -1706 1266 -1554 1280
rect -897 1220 -857 1374
rect -357 1220 -317 1374
rect 315 1220 355 1374
rect 616 1220 656 1374
rect 855 1220 895 1374
rect 1527 1220 1567 1374
rect 2067 1220 2107 1374
rect -2420 1209 -2340 1220
rect -2420 1175 -2397 1209
rect -2363 1175 -2340 1209
rect -2420 1137 -2340 1175
rect -2420 1103 -2397 1137
rect -2363 1103 -2340 1137
rect -2420 1065 -2340 1103
rect -2420 1031 -2397 1065
rect -2363 1031 -2340 1065
rect -2420 993 -2340 1031
rect -2420 959 -2397 993
rect -2363 959 -2340 993
rect -2420 921 -2340 959
rect -2420 887 -2397 921
rect -2363 887 -2340 921
rect -2420 849 -2340 887
rect -2420 815 -2397 849
rect -2363 815 -2340 849
rect -2420 777 -2340 815
rect -2420 743 -2397 777
rect -2363 743 -2340 777
rect -2420 705 -2340 743
rect -2420 671 -2397 705
rect -2363 671 -2340 705
rect -2420 660 -2340 671
rect -2120 1218 -2040 1220
rect -2120 1166 -2106 1218
rect -2054 1166 -2040 1218
rect -2120 1146 -2040 1166
rect -2120 1094 -2106 1146
rect -2054 1094 -2040 1146
rect -2120 1074 -2040 1094
rect -2120 1022 -2106 1074
rect -2054 1022 -2040 1074
rect -2120 1002 -2040 1022
rect -2120 950 -2106 1002
rect -2054 950 -2040 1002
rect -2120 930 -2040 950
rect -2120 878 -2106 930
rect -2054 878 -2040 930
rect -2120 858 -2040 878
rect -2120 806 -2106 858
rect -2054 806 -2040 858
rect -2120 786 -2040 806
rect -2120 734 -2106 786
rect -2054 734 -2040 786
rect -2120 714 -2040 734
rect -2120 662 -2106 714
rect -2054 662 -2040 714
rect -2120 660 -2040 662
rect -1820 1209 -1740 1220
rect -1820 1175 -1797 1209
rect -1763 1175 -1740 1209
rect -1820 1137 -1740 1175
rect -1820 1103 -1797 1137
rect -1763 1103 -1740 1137
rect -1820 1065 -1740 1103
rect -1820 1031 -1797 1065
rect -1763 1031 -1740 1065
rect -1820 993 -1740 1031
rect -1820 959 -1797 993
rect -1763 959 -1740 993
rect -1820 921 -1740 959
rect -1820 887 -1797 921
rect -1763 887 -1740 921
rect -1820 849 -1740 887
rect -1820 815 -1797 849
rect -1763 815 -1740 849
rect -1820 777 -1740 815
rect -1820 743 -1797 777
rect -1763 743 -1740 777
rect -1820 705 -1740 743
rect -1820 671 -1797 705
rect -1763 671 -1740 705
rect -1820 660 -1740 671
rect -917 1209 -837 1220
rect -917 1175 -894 1209
rect -860 1175 -837 1209
rect -917 1137 -837 1175
rect -917 1103 -894 1137
rect -860 1103 -837 1137
rect -917 1065 -837 1103
rect -917 1031 -894 1065
rect -860 1031 -837 1065
rect -917 993 -837 1031
rect -917 959 -894 993
rect -860 959 -837 993
rect -917 921 -837 959
rect -917 887 -894 921
rect -860 887 -837 921
rect -917 849 -837 887
rect -917 815 -894 849
rect -860 815 -837 849
rect -917 777 -837 815
rect -917 743 -894 777
rect -860 743 -837 777
rect -917 705 -837 743
rect -917 671 -894 705
rect -860 671 -837 705
rect -917 660 -837 671
rect -377 1209 -297 1220
rect -377 1175 -354 1209
rect -320 1175 -297 1209
rect -377 1137 -297 1175
rect -377 1103 -354 1137
rect -320 1103 -297 1137
rect -377 1065 -297 1103
rect -377 1031 -354 1065
rect -320 1031 -297 1065
rect -377 993 -297 1031
rect -377 959 -354 993
rect -320 959 -297 993
rect -377 921 -297 959
rect -377 887 -354 921
rect -320 887 -297 921
rect -377 849 -297 887
rect -377 815 -354 849
rect -320 815 -297 849
rect -377 777 -297 815
rect -377 743 -354 777
rect -320 743 -297 777
rect -377 705 -297 743
rect -377 671 -354 705
rect -320 671 -297 705
rect -377 660 -297 671
rect 295 1209 375 1220
rect 295 1175 318 1209
rect 352 1175 375 1209
rect 295 1137 375 1175
rect 295 1103 318 1137
rect 352 1103 375 1137
rect 295 1065 375 1103
rect 295 1031 318 1065
rect 352 1031 375 1065
rect 295 993 375 1031
rect 295 959 318 993
rect 352 959 375 993
rect 295 921 375 959
rect 295 887 318 921
rect 352 887 375 921
rect 295 849 375 887
rect 295 815 318 849
rect 352 815 375 849
rect 295 777 375 815
rect 295 743 318 777
rect 352 743 375 777
rect 295 705 375 743
rect 295 671 318 705
rect 352 671 375 705
rect 295 660 375 671
rect 595 1209 675 1220
rect 595 1175 618 1209
rect 652 1175 675 1209
rect 595 1137 675 1175
rect 595 1103 618 1137
rect 652 1103 675 1137
rect 595 1065 675 1103
rect 595 1031 618 1065
rect 652 1031 675 1065
rect 595 993 675 1031
rect 595 959 618 993
rect 652 959 675 993
rect 595 921 675 959
rect 595 887 618 921
rect 652 887 675 921
rect 595 849 675 887
rect 595 815 618 849
rect 652 815 675 849
rect 595 777 675 815
rect 595 743 618 777
rect 652 743 675 777
rect 595 705 675 743
rect 595 671 618 705
rect 652 671 675 705
rect 595 660 675 671
rect 835 1209 915 1220
rect 835 1175 858 1209
rect 892 1175 915 1209
rect 835 1137 915 1175
rect 835 1103 858 1137
rect 892 1103 915 1137
rect 835 1065 915 1103
rect 835 1031 858 1065
rect 892 1031 915 1065
rect 835 993 915 1031
rect 835 959 858 993
rect 892 959 915 993
rect 835 921 915 959
rect 835 887 858 921
rect 892 887 915 921
rect 835 849 915 887
rect 835 815 858 849
rect 892 815 915 849
rect 835 777 915 815
rect 835 743 858 777
rect 892 743 915 777
rect 835 705 915 743
rect 835 671 858 705
rect 892 671 915 705
rect 835 660 915 671
rect 1507 1209 1587 1220
rect 1507 1175 1530 1209
rect 1564 1175 1587 1209
rect 1507 1137 1587 1175
rect 1507 1103 1530 1137
rect 1564 1103 1587 1137
rect 1507 1065 1587 1103
rect 1507 1031 1530 1065
rect 1564 1031 1587 1065
rect 1507 993 1587 1031
rect 1507 959 1530 993
rect 1564 959 1587 993
rect 1507 921 1587 959
rect 1507 887 1530 921
rect 1564 887 1587 921
rect 1507 849 1587 887
rect 1507 815 1530 849
rect 1564 815 1587 849
rect 1507 777 1587 815
rect 1507 743 1530 777
rect 1564 743 1587 777
rect 1507 705 1587 743
rect 1507 671 1530 705
rect 1564 671 1587 705
rect 1507 660 1587 671
rect 2047 1209 2127 1220
rect 2047 1175 2070 1209
rect 2104 1175 2127 1209
rect 2047 1137 2127 1175
rect 2047 1103 2070 1137
rect 2104 1103 2127 1137
rect 2047 1065 2127 1103
rect 2047 1031 2070 1065
rect 2104 1031 2127 1065
rect 2047 993 2127 1031
rect 2047 959 2070 993
rect 2104 959 2127 993
rect 2047 921 2127 959
rect 2047 887 2070 921
rect 2104 887 2127 921
rect 2047 849 2127 887
rect 2047 815 2070 849
rect 2104 815 2127 849
rect 2047 777 2127 815
rect 2047 743 2070 777
rect 2104 743 2127 777
rect 2047 705 2127 743
rect 2047 671 2070 705
rect 2104 671 2127 705
rect 2047 660 2127 671
rect -1840 593 -1760 616
rect -1840 559 -1817 593
rect -1783 559 -1760 593
rect -1840 536 -1760 559
rect -2220 405 -2140 425
rect -1820 405 -1781 536
rect 2197 534 2277 548
rect -1676 508 -1528 522
rect -1676 456 -1662 508
rect -1610 456 -1594 508
rect -1542 502 -1528 508
rect -81 502 -1 522
rect -1542 499 -1 502
rect -1542 465 -58 499
rect -24 465 -1 499
rect -1542 462 -1 465
rect -1542 456 -1528 462
rect -1676 442 -1528 456
rect -81 442 -1 462
rect 2197 482 2211 534
rect 2263 482 2277 534
rect 2197 462 2277 482
rect -2220 402 -1781 405
rect -2220 368 -2197 402
rect -2163 368 -1781 402
rect 2197 410 2211 462
rect 2263 410 2277 462
rect 2197 396 2277 410
rect -2220 365 -1781 368
rect -2220 345 -2140 365
rect -2420 269 -2340 310
rect -2420 235 -2397 269
rect -2363 235 -2340 269
rect -2420 197 -2340 235
rect -2420 163 -2397 197
rect -2363 163 -2340 197
rect -2420 125 -2340 163
rect -2420 91 -2397 125
rect -2363 91 -2340 125
rect -2420 50 -2340 91
rect -2120 278 -2040 310
rect -2120 226 -2106 278
rect -2054 226 -2040 278
rect -2120 206 -2040 226
rect -2120 154 -2106 206
rect -2054 154 -2040 206
rect -2120 134 -2040 154
rect -2120 82 -2106 134
rect -2054 82 -2040 134
rect -2120 50 -2040 82
rect -1820 269 -1740 310
rect -1820 235 -1797 269
rect -1763 235 -1740 269
rect -1820 197 -1740 235
rect -1820 163 -1797 197
rect -1763 163 -1740 197
rect -1820 125 -1740 163
rect -1820 91 -1797 125
rect -1763 91 -1740 125
rect -1820 50 -1740 91
rect -917 269 -837 310
rect -917 235 -894 269
rect -860 235 -837 269
rect -917 197 -837 235
rect -917 163 -894 197
rect -860 163 -837 197
rect -917 125 -837 163
rect -917 91 -894 125
rect -860 91 -837 125
rect -917 50 -837 91
rect -617 269 -537 310
rect -617 235 -594 269
rect -560 235 -537 269
rect -617 197 -537 235
rect -617 163 -594 197
rect -560 163 -537 197
rect -617 125 -537 163
rect -617 91 -594 125
rect -560 91 -537 125
rect -617 50 -537 91
rect -377 269 -297 310
rect -377 235 -354 269
rect -320 235 -297 269
rect -377 197 -297 235
rect -377 163 -354 197
rect -320 163 -297 197
rect -377 125 -297 163
rect -377 91 -354 125
rect -320 91 -297 125
rect -377 50 -297 91
rect 295 269 375 310
rect 295 235 318 269
rect 352 235 375 269
rect 295 197 375 235
rect 295 163 318 197
rect 352 163 375 197
rect 295 125 375 163
rect 295 91 318 125
rect 352 91 375 125
rect 295 50 375 91
rect 835 269 915 310
rect 835 235 858 269
rect 892 235 915 269
rect 835 197 915 235
rect 835 163 858 197
rect 892 163 915 197
rect 835 125 915 163
rect 835 91 858 125
rect 892 91 915 125
rect 835 50 915 91
rect 1507 269 1587 310
rect 1507 235 1530 269
rect 1564 235 1587 269
rect 1507 197 1587 235
rect 1507 163 1530 197
rect 1564 163 1587 197
rect 1507 125 1587 163
rect 1507 91 1530 125
rect 1564 91 1587 125
rect 1507 50 1587 91
rect 1807 269 1887 310
rect 1807 235 1830 269
rect 1864 235 1887 269
rect 1807 197 1887 235
rect 1807 163 1830 197
rect 1864 163 1887 197
rect 1807 125 1887 163
rect 1807 91 1830 125
rect 1864 91 1887 125
rect 1807 50 1887 91
rect 2047 269 2127 310
rect 2047 235 2070 269
rect 2104 235 2127 269
rect 2047 197 2127 235
rect 2047 163 2070 197
rect 2104 163 2127 197
rect 2047 125 2127 163
rect 2047 91 2070 125
rect 2104 91 2127 125
rect 2047 50 2127 91
rect -2400 -104 -2360 50
rect -1800 -104 -1760 50
rect -1706 -10 -1554 4
rect -1706 -62 -1692 -10
rect -1640 -62 -1620 -10
rect -1568 -62 -1554 -10
rect -1706 -76 -1554 -62
rect -897 -104 -857 50
rect -597 -104 -557 50
rect -357 -104 -317 50
rect 315 -104 355 50
rect 855 -104 895 50
rect 1527 -104 1567 50
rect 1827 -104 1867 50
rect 2067 -104 2107 50
rect -2520 -137 2342 -104
rect -2520 -171 -2497 -137
rect -2463 -171 -2425 -137
rect -2391 -171 -2353 -137
rect -2319 -171 -2281 -137
rect -2247 -171 -2209 -137
rect -2175 -171 -2137 -137
rect -2103 -171 -2065 -137
rect -2031 -171 -1993 -137
rect -1959 -171 -1921 -137
rect -1887 -171 -1849 -137
rect -1815 -171 -1777 -137
rect -1743 -171 -1705 -137
rect -1671 -171 -1633 -137
rect -1599 -171 -1561 -137
rect -1527 -171 -1489 -137
rect -1455 -171 -1417 -137
rect -1383 -171 -1345 -137
rect -1311 -171 -939 -137
rect -905 -171 -867 -137
rect -833 -171 -795 -137
rect -761 -171 -723 -137
rect -689 -171 -651 -137
rect -617 -171 -579 -137
rect -545 -171 -507 -137
rect -473 -171 -435 -137
rect -401 -171 -363 -137
rect -329 -171 -291 -137
rect -257 -171 -219 -137
rect -185 -171 -147 -137
rect -113 -171 273 -137
rect 307 -171 345 -137
rect 379 -171 417 -137
rect 451 -171 489 -137
rect 523 -171 561 -137
rect 595 -171 633 -137
rect 667 -171 705 -137
rect 739 -171 777 -137
rect 811 -171 849 -137
rect 883 -171 921 -137
rect 955 -171 993 -137
rect 1027 -171 1065 -137
rect 1099 -171 1485 -137
rect 1519 -171 1557 -137
rect 1591 -171 1629 -137
rect 1663 -171 1701 -137
rect 1735 -171 1773 -137
rect 1807 -171 1845 -137
rect 1879 -171 1917 -137
rect 1951 -171 1989 -137
rect 2023 -171 2061 -137
rect 2095 -171 2133 -137
rect 2167 -171 2205 -137
rect 2239 -171 2277 -137
rect 2311 -171 2342 -137
rect -2520 -204 2342 -171
rect -2400 -358 -2360 -204
rect -1800 -358 -1760 -204
rect -1549 -358 -1509 -204
rect -1481 -246 -1329 -232
rect -1481 -298 -1467 -246
rect -1415 -298 -1395 -246
rect -1343 -298 -1329 -246
rect -1481 -312 -1329 -298
rect -897 -358 -857 -204
rect -357 -358 -317 -204
rect 315 -358 355 -204
rect 855 -358 895 -204
rect -2420 -399 -2340 -358
rect -2420 -433 -2397 -399
rect -2363 -433 -2340 -399
rect -2420 -471 -2340 -433
rect -2420 -505 -2397 -471
rect -2363 -505 -2340 -471
rect -2420 -543 -2340 -505
rect -2420 -577 -2397 -543
rect -2363 -577 -2340 -543
rect -2420 -618 -2340 -577
rect -2120 -390 -2040 -358
rect -2120 -442 -2106 -390
rect -2054 -442 -2040 -390
rect -2120 -462 -2040 -442
rect -2120 -514 -2106 -462
rect -2054 -514 -2040 -462
rect -2120 -534 -2040 -514
rect -2120 -586 -2106 -534
rect -2054 -586 -2040 -534
rect -2120 -618 -2040 -586
rect -1820 -399 -1740 -358
rect -1820 -433 -1797 -399
rect -1763 -433 -1740 -399
rect -1820 -471 -1740 -433
rect -1820 -505 -1797 -471
rect -1763 -505 -1740 -471
rect -1820 -543 -1740 -505
rect -1820 -577 -1797 -543
rect -1763 -577 -1740 -543
rect -1820 -618 -1740 -577
rect -1569 -399 -1489 -358
rect -1569 -433 -1546 -399
rect -1512 -433 -1489 -399
rect -1569 -471 -1489 -433
rect -1569 -505 -1546 -471
rect -1512 -505 -1489 -471
rect -1569 -543 -1489 -505
rect -1569 -577 -1546 -543
rect -1512 -577 -1489 -543
rect -1569 -618 -1489 -577
rect -917 -399 -837 -358
rect -917 -433 -894 -399
rect -860 -433 -837 -399
rect -917 -471 -837 -433
rect -917 -505 -894 -471
rect -860 -505 -837 -471
rect -917 -543 -837 -505
rect -917 -577 -894 -543
rect -860 -577 -837 -543
rect -917 -618 -837 -577
rect -377 -399 -297 -358
rect -377 -433 -354 -399
rect -320 -433 -297 -399
rect -377 -471 -297 -433
rect -377 -505 -354 -471
rect -320 -505 -297 -471
rect -377 -543 -297 -505
rect -377 -577 -354 -543
rect -320 -577 -297 -543
rect -377 -618 -297 -577
rect 295 -399 375 -358
rect 295 -433 318 -399
rect 352 -433 375 -399
rect 295 -471 375 -433
rect 295 -505 318 -471
rect 352 -505 375 -471
rect 295 -543 375 -505
rect 295 -577 318 -543
rect 352 -577 375 -543
rect 295 -618 375 -577
rect 835 -399 915 -358
rect 835 -433 858 -399
rect 892 -433 915 -399
rect 835 -471 915 -433
rect 835 -505 858 -471
rect 892 -505 915 -471
rect 835 -543 915 -505
rect 835 -577 858 -543
rect 892 -577 915 -543
rect 835 -618 915 -577
rect -2220 -673 -2140 -653
rect -2220 -676 -1781 -673
rect -2220 -710 -2197 -676
rect -2163 -710 -1781 -676
rect -2220 -713 -1781 -710
rect -2220 -733 -2140 -713
rect -1820 -844 -1781 -713
rect -1419 -701 -1339 -678
rect -1691 -746 -1611 -732
rect -1691 -798 -1677 -746
rect -1625 -798 -1611 -746
rect -1691 -818 -1611 -798
rect -1840 -867 -1760 -844
rect -1840 -901 -1817 -867
rect -1783 -901 -1760 -867
rect -1691 -870 -1677 -818
rect -1625 -870 -1611 -818
rect -1419 -735 -1396 -701
rect -1362 -735 -1339 -701
rect -1419 -770 -1339 -735
rect -81 -701 -1 -678
rect -81 -735 -58 -701
rect -24 -735 -1 -701
rect -81 -770 -1 -735
rect -1419 -773 -1 -770
rect -1419 -807 -1396 -773
rect -1362 -807 -58 -773
rect -24 -807 -1 -773
rect -1419 -810 -1 -807
rect -1419 -830 -1339 -810
rect -81 -830 -1 -810
rect -1691 -884 -1611 -870
rect -1840 -924 -1760 -901
rect -2420 -979 -2340 -968
rect -2420 -1013 -2397 -979
rect -2363 -1013 -2340 -979
rect -2420 -1051 -2340 -1013
rect -2420 -1085 -2397 -1051
rect -2363 -1085 -2340 -1051
rect -2420 -1123 -2340 -1085
rect -2420 -1157 -2397 -1123
rect -2363 -1157 -2340 -1123
rect -2420 -1195 -2340 -1157
rect -2420 -1229 -2397 -1195
rect -2363 -1229 -2340 -1195
rect -2420 -1267 -2340 -1229
rect -2420 -1301 -2397 -1267
rect -2363 -1301 -2340 -1267
rect -2420 -1339 -2340 -1301
rect -2420 -1373 -2397 -1339
rect -2363 -1373 -2340 -1339
rect -2420 -1411 -2340 -1373
rect -2420 -1445 -2397 -1411
rect -2363 -1445 -2340 -1411
rect -2420 -1483 -2340 -1445
rect -2420 -1517 -2397 -1483
rect -2363 -1517 -2340 -1483
rect -2420 -1528 -2340 -1517
rect -2120 -970 -2040 -968
rect -2120 -1022 -2106 -970
rect -2054 -1022 -2040 -970
rect -2120 -1042 -2040 -1022
rect -2120 -1094 -2106 -1042
rect -2054 -1094 -2040 -1042
rect -2120 -1114 -2040 -1094
rect -2120 -1166 -2106 -1114
rect -2054 -1166 -2040 -1114
rect -2120 -1186 -2040 -1166
rect -2120 -1238 -2106 -1186
rect -2054 -1238 -2040 -1186
rect -2120 -1258 -2040 -1238
rect -2120 -1310 -2106 -1258
rect -2054 -1310 -2040 -1258
rect -2120 -1330 -2040 -1310
rect -2120 -1382 -2106 -1330
rect -2054 -1382 -2040 -1330
rect -2120 -1402 -2040 -1382
rect -2120 -1454 -2106 -1402
rect -2054 -1454 -2040 -1402
rect -2120 -1474 -2040 -1454
rect -2120 -1526 -2106 -1474
rect -2054 -1526 -2040 -1474
rect -2120 -1528 -2040 -1526
rect -1820 -979 -1740 -968
rect -1820 -1013 -1797 -979
rect -1763 -1013 -1740 -979
rect -1820 -1051 -1740 -1013
rect -1820 -1085 -1797 -1051
rect -1763 -1085 -1740 -1051
rect -1820 -1123 -1740 -1085
rect -1820 -1157 -1797 -1123
rect -1763 -1157 -1740 -1123
rect -1820 -1195 -1740 -1157
rect -1820 -1229 -1797 -1195
rect -1763 -1229 -1740 -1195
rect -1820 -1267 -1740 -1229
rect -1820 -1301 -1797 -1267
rect -1763 -1301 -1740 -1267
rect -1820 -1339 -1740 -1301
rect -1820 -1373 -1797 -1339
rect -1763 -1373 -1740 -1339
rect -1820 -1411 -1740 -1373
rect -1820 -1445 -1797 -1411
rect -1763 -1445 -1740 -1411
rect -1820 -1483 -1740 -1445
rect -1820 -1517 -1797 -1483
rect -1763 -1517 -1740 -1483
rect -1820 -1528 -1740 -1517
rect -1569 -979 -1489 -968
rect -1569 -1013 -1546 -979
rect -1512 -1013 -1489 -979
rect -1569 -1051 -1489 -1013
rect -1569 -1085 -1546 -1051
rect -1512 -1085 -1489 -1051
rect -1569 -1123 -1489 -1085
rect -1569 -1157 -1546 -1123
rect -1512 -1157 -1489 -1123
rect -1569 -1195 -1489 -1157
rect -1569 -1229 -1546 -1195
rect -1512 -1229 -1489 -1195
rect -1569 -1267 -1489 -1229
rect -1569 -1301 -1546 -1267
rect -1512 -1301 -1489 -1267
rect -1569 -1339 -1489 -1301
rect -1569 -1373 -1546 -1339
rect -1512 -1373 -1489 -1339
rect -1569 -1411 -1489 -1373
rect -1569 -1445 -1546 -1411
rect -1512 -1445 -1489 -1411
rect -1569 -1483 -1489 -1445
rect -1569 -1517 -1546 -1483
rect -1512 -1517 -1489 -1483
rect -1569 -1528 -1489 -1517
rect -917 -979 -837 -968
rect -917 -1013 -894 -979
rect -860 -1013 -837 -979
rect -917 -1051 -837 -1013
rect -917 -1085 -894 -1051
rect -860 -1085 -837 -1051
rect -917 -1123 -837 -1085
rect -917 -1157 -894 -1123
rect -860 -1157 -837 -1123
rect -917 -1195 -837 -1157
rect -917 -1229 -894 -1195
rect -860 -1229 -837 -1195
rect -917 -1267 -837 -1229
rect -917 -1301 -894 -1267
rect -860 -1301 -837 -1267
rect -917 -1339 -837 -1301
rect -917 -1373 -894 -1339
rect -860 -1373 -837 -1339
rect -917 -1411 -837 -1373
rect -917 -1445 -894 -1411
rect -860 -1445 -837 -1411
rect -917 -1483 -837 -1445
rect -917 -1517 -894 -1483
rect -860 -1517 -837 -1483
rect -917 -1528 -837 -1517
rect -617 -979 -537 -968
rect -617 -1013 -594 -979
rect -560 -1013 -537 -979
rect -617 -1051 -537 -1013
rect -617 -1085 -594 -1051
rect -560 -1085 -537 -1051
rect -617 -1123 -537 -1085
rect -617 -1157 -594 -1123
rect -560 -1157 -537 -1123
rect -617 -1195 -537 -1157
rect -617 -1229 -594 -1195
rect -560 -1229 -537 -1195
rect -617 -1267 -537 -1229
rect -617 -1301 -594 -1267
rect -560 -1301 -537 -1267
rect -617 -1339 -537 -1301
rect -617 -1373 -594 -1339
rect -560 -1373 -537 -1339
rect -617 -1411 -537 -1373
rect -617 -1445 -594 -1411
rect -560 -1445 -537 -1411
rect -617 -1483 -537 -1445
rect -617 -1517 -594 -1483
rect -560 -1517 -537 -1483
rect -617 -1528 -537 -1517
rect -377 -979 -297 -968
rect -377 -1013 -354 -979
rect -320 -1013 -297 -979
rect -377 -1051 -297 -1013
rect -377 -1085 -354 -1051
rect -320 -1085 -297 -1051
rect -377 -1123 -297 -1085
rect -377 -1157 -354 -1123
rect -320 -1157 -297 -1123
rect -377 -1195 -297 -1157
rect -377 -1229 -354 -1195
rect -320 -1229 -297 -1195
rect -377 -1267 -297 -1229
rect -377 -1301 -354 -1267
rect -320 -1301 -297 -1267
rect -377 -1339 -297 -1301
rect -377 -1373 -354 -1339
rect -320 -1373 -297 -1339
rect -377 -1411 -297 -1373
rect -377 -1445 -354 -1411
rect -320 -1445 -297 -1411
rect -377 -1483 -297 -1445
rect -377 -1517 -354 -1483
rect -320 -1517 -297 -1483
rect -377 -1528 -297 -1517
rect 295 -979 375 -968
rect 295 -1013 318 -979
rect 352 -1013 375 -979
rect 295 -1051 375 -1013
rect 295 -1085 318 -1051
rect 352 -1085 375 -1051
rect 295 -1123 375 -1085
rect 295 -1157 318 -1123
rect 352 -1157 375 -1123
rect 295 -1195 375 -1157
rect 295 -1229 318 -1195
rect 352 -1229 375 -1195
rect 295 -1267 375 -1229
rect 295 -1301 318 -1267
rect 352 -1301 375 -1267
rect 295 -1339 375 -1301
rect 295 -1373 318 -1339
rect 352 -1373 375 -1339
rect 295 -1411 375 -1373
rect 295 -1445 318 -1411
rect 352 -1445 375 -1411
rect 295 -1483 375 -1445
rect 295 -1517 318 -1483
rect 352 -1517 375 -1483
rect 295 -1528 375 -1517
rect 595 -979 675 -968
rect 595 -1013 618 -979
rect 652 -1013 675 -979
rect 595 -1051 675 -1013
rect 595 -1085 618 -1051
rect 652 -1085 675 -1051
rect 595 -1123 675 -1085
rect 595 -1157 618 -1123
rect 652 -1157 675 -1123
rect 595 -1195 675 -1157
rect 595 -1229 618 -1195
rect 652 -1229 675 -1195
rect 595 -1267 675 -1229
rect 595 -1301 618 -1267
rect 652 -1301 675 -1267
rect 595 -1339 675 -1301
rect 595 -1373 618 -1339
rect 652 -1373 675 -1339
rect 595 -1411 675 -1373
rect 595 -1445 618 -1411
rect 652 -1445 675 -1411
rect 595 -1483 675 -1445
rect 595 -1517 618 -1483
rect 652 -1517 675 -1483
rect 595 -1528 675 -1517
rect 835 -979 915 -968
rect 835 -1013 858 -979
rect 892 -1013 915 -979
rect 835 -1051 915 -1013
rect 835 -1085 858 -1051
rect 892 -1085 915 -1051
rect 835 -1123 915 -1085
rect 835 -1157 858 -1123
rect 892 -1157 915 -1123
rect 835 -1195 915 -1157
rect 835 -1229 858 -1195
rect 892 -1229 915 -1195
rect 835 -1267 915 -1229
rect 835 -1301 858 -1267
rect 892 -1301 915 -1267
rect 835 -1339 915 -1301
rect 835 -1373 858 -1339
rect 892 -1373 915 -1339
rect 835 -1411 915 -1373
rect 835 -1445 858 -1411
rect 892 -1445 915 -1411
rect 835 -1483 915 -1445
rect 835 -1517 858 -1483
rect 892 -1517 915 -1483
rect 835 -1528 915 -1517
rect -2400 -1682 -2360 -1528
rect -1800 -1682 -1760 -1528
rect -1549 -1682 -1509 -1528
rect -1481 -1588 -1329 -1574
rect -1481 -1640 -1467 -1588
rect -1415 -1640 -1395 -1588
rect -1343 -1640 -1329 -1588
rect -1481 -1654 -1329 -1640
rect -897 -1682 -857 -1528
rect -596 -1682 -556 -1528
rect -357 -1682 -317 -1528
rect 315 -1682 355 -1528
rect 616 -1682 656 -1528
rect 855 -1682 895 -1528
rect -2628 -1715 1130 -1682
rect -2628 -1749 -2497 -1715
rect -2463 -1749 -2425 -1715
rect -2391 -1749 -2353 -1715
rect -2319 -1749 -2281 -1715
rect -2247 -1749 -2209 -1715
rect -2175 -1749 -2137 -1715
rect -2103 -1749 -2065 -1715
rect -2031 -1749 -1993 -1715
rect -1959 -1749 -1921 -1715
rect -1887 -1749 -1849 -1715
rect -1815 -1749 -1777 -1715
rect -1743 -1749 -1705 -1715
rect -1671 -1749 -1633 -1715
rect -1599 -1749 -1561 -1715
rect -1527 -1749 -1489 -1715
rect -1455 -1749 -1417 -1715
rect -1383 -1749 -1345 -1715
rect -1311 -1749 -939 -1715
rect -905 -1749 -867 -1715
rect -833 -1749 -795 -1715
rect -761 -1749 -723 -1715
rect -689 -1749 -651 -1715
rect -617 -1749 -579 -1715
rect -545 -1749 -507 -1715
rect -473 -1749 -435 -1715
rect -401 -1749 -363 -1715
rect -329 -1749 -291 -1715
rect -257 -1749 -219 -1715
rect -185 -1749 -147 -1715
rect -113 -1749 273 -1715
rect 307 -1749 345 -1715
rect 379 -1749 417 -1715
rect 451 -1749 489 -1715
rect 523 -1749 561 -1715
rect 595 -1749 633 -1715
rect 667 -1749 705 -1715
rect 739 -1749 777 -1715
rect 811 -1749 849 -1715
rect 883 -1749 921 -1715
rect 955 -1749 993 -1715
rect 1027 -1749 1065 -1715
rect 1099 -1749 1130 -1715
rect -2628 -1782 1130 -1749
<< via1 >>
rect -3412 1348 -3360 1400
rect -3412 1280 -3360 1332
rect -3412 1212 -3360 1264
rect -3298 -1576 -3246 -1524
rect -3298 -1644 -3246 -1592
rect -3298 -1712 -3246 -1660
rect -3184 -230 -3132 -178
rect -3184 -298 -3132 -246
rect -3184 -366 -3132 -314
rect -3070 6 -3018 58
rect -3070 -62 -3018 -10
rect -3070 -130 -3018 -78
rect -1692 1323 -1640 1332
rect -1692 1289 -1683 1323
rect -1683 1289 -1649 1323
rect -1649 1289 -1640 1323
rect -1692 1280 -1640 1289
rect -1620 1323 -1568 1332
rect -1620 1289 -1611 1323
rect -1611 1289 -1577 1323
rect -1577 1289 -1568 1323
rect -1620 1280 -1568 1289
rect -2106 1209 -2054 1218
rect -2106 1175 -2097 1209
rect -2097 1175 -2063 1209
rect -2063 1175 -2054 1209
rect -2106 1166 -2054 1175
rect -2106 1137 -2054 1146
rect -2106 1103 -2097 1137
rect -2097 1103 -2063 1137
rect -2063 1103 -2054 1137
rect -2106 1094 -2054 1103
rect -2106 1065 -2054 1074
rect -2106 1031 -2097 1065
rect -2097 1031 -2063 1065
rect -2063 1031 -2054 1065
rect -2106 1022 -2054 1031
rect -2106 993 -2054 1002
rect -2106 959 -2097 993
rect -2097 959 -2063 993
rect -2063 959 -2054 993
rect -2106 950 -2054 959
rect -2106 921 -2054 930
rect -2106 887 -2097 921
rect -2097 887 -2063 921
rect -2063 887 -2054 921
rect -2106 878 -2054 887
rect -2106 849 -2054 858
rect -2106 815 -2097 849
rect -2097 815 -2063 849
rect -2063 815 -2054 849
rect -2106 806 -2054 815
rect -2106 777 -2054 786
rect -2106 743 -2097 777
rect -2097 743 -2063 777
rect -2063 743 -2054 777
rect -2106 734 -2054 743
rect -2106 705 -2054 714
rect -2106 671 -2097 705
rect -2097 671 -2063 705
rect -2063 671 -2054 705
rect -2106 662 -2054 671
rect -1662 456 -1610 508
rect -1594 456 -1542 508
rect 2211 525 2263 534
rect 2211 491 2220 525
rect 2220 491 2254 525
rect 2254 491 2263 525
rect 2211 482 2263 491
rect 2211 453 2263 462
rect 2211 419 2220 453
rect 2220 419 2254 453
rect 2254 419 2263 453
rect 2211 410 2263 419
rect -2106 269 -2054 278
rect -2106 235 -2097 269
rect -2097 235 -2063 269
rect -2063 235 -2054 269
rect -2106 226 -2054 235
rect -2106 197 -2054 206
rect -2106 163 -2097 197
rect -2097 163 -2063 197
rect -2063 163 -2054 197
rect -2106 154 -2054 163
rect -2106 125 -2054 134
rect -2106 91 -2097 125
rect -2097 91 -2063 125
rect -2063 91 -2054 125
rect -2106 82 -2054 91
rect -1692 -19 -1640 -10
rect -1692 -53 -1683 -19
rect -1683 -53 -1649 -19
rect -1649 -53 -1640 -19
rect -1692 -62 -1640 -53
rect -1620 -19 -1568 -10
rect -1620 -53 -1611 -19
rect -1611 -53 -1577 -19
rect -1577 -53 -1568 -19
rect -1620 -62 -1568 -53
rect -1467 -255 -1415 -246
rect -1467 -289 -1458 -255
rect -1458 -289 -1424 -255
rect -1424 -289 -1415 -255
rect -1467 -298 -1415 -289
rect -1395 -255 -1343 -246
rect -1395 -289 -1386 -255
rect -1386 -289 -1352 -255
rect -1352 -289 -1343 -255
rect -1395 -298 -1343 -289
rect -2106 -399 -2054 -390
rect -2106 -433 -2097 -399
rect -2097 -433 -2063 -399
rect -2063 -433 -2054 -399
rect -2106 -442 -2054 -433
rect -2106 -471 -2054 -462
rect -2106 -505 -2097 -471
rect -2097 -505 -2063 -471
rect -2063 -505 -2054 -471
rect -2106 -514 -2054 -505
rect -2106 -543 -2054 -534
rect -2106 -577 -2097 -543
rect -2097 -577 -2063 -543
rect -2063 -577 -2054 -543
rect -2106 -586 -2054 -577
rect -1677 -755 -1625 -746
rect -1677 -789 -1668 -755
rect -1668 -789 -1634 -755
rect -1634 -789 -1625 -755
rect -1677 -798 -1625 -789
rect -1677 -827 -1625 -818
rect -1677 -861 -1668 -827
rect -1668 -861 -1634 -827
rect -1634 -861 -1625 -827
rect -1677 -870 -1625 -861
rect -2106 -979 -2054 -970
rect -2106 -1013 -2097 -979
rect -2097 -1013 -2063 -979
rect -2063 -1013 -2054 -979
rect -2106 -1022 -2054 -1013
rect -2106 -1051 -2054 -1042
rect -2106 -1085 -2097 -1051
rect -2097 -1085 -2063 -1051
rect -2063 -1085 -2054 -1051
rect -2106 -1094 -2054 -1085
rect -2106 -1123 -2054 -1114
rect -2106 -1157 -2097 -1123
rect -2097 -1157 -2063 -1123
rect -2063 -1157 -2054 -1123
rect -2106 -1166 -2054 -1157
rect -2106 -1195 -2054 -1186
rect -2106 -1229 -2097 -1195
rect -2097 -1229 -2063 -1195
rect -2063 -1229 -2054 -1195
rect -2106 -1238 -2054 -1229
rect -2106 -1267 -2054 -1258
rect -2106 -1301 -2097 -1267
rect -2097 -1301 -2063 -1267
rect -2063 -1301 -2054 -1267
rect -2106 -1310 -2054 -1301
rect -2106 -1339 -2054 -1330
rect -2106 -1373 -2097 -1339
rect -2097 -1373 -2063 -1339
rect -2063 -1373 -2054 -1339
rect -2106 -1382 -2054 -1373
rect -2106 -1411 -2054 -1402
rect -2106 -1445 -2097 -1411
rect -2097 -1445 -2063 -1411
rect -2063 -1445 -2054 -1411
rect -2106 -1454 -2054 -1445
rect -2106 -1483 -2054 -1474
rect -2106 -1517 -2097 -1483
rect -2097 -1517 -2063 -1483
rect -2063 -1517 -2054 -1483
rect -2106 -1526 -2054 -1517
rect -1467 -1597 -1415 -1588
rect -1467 -1631 -1458 -1597
rect -1458 -1631 -1424 -1597
rect -1424 -1631 -1415 -1597
rect -1467 -1640 -1415 -1631
rect -1395 -1597 -1343 -1588
rect -1395 -1631 -1386 -1597
rect -1386 -1631 -1352 -1597
rect -1352 -1631 -1343 -1597
rect -1395 -1640 -1343 -1631
<< metal2 >>
rect -3426 1400 -3346 1414
rect -3426 1348 -3412 1400
rect -3360 1348 -3346 1400
rect -3426 1332 -3346 1348
rect -3426 1280 -3412 1332
rect -3360 1326 -3346 1332
rect -1706 1332 -1554 1346
rect -1706 1326 -1692 1332
rect -3360 1286 -1692 1326
rect -3360 1280 -3346 1286
rect -3426 1264 -3346 1280
rect -1706 1280 -1692 1286
rect -1640 1280 -1620 1332
rect -1568 1280 -1554 1332
rect -1706 1266 -1554 1280
rect -3426 1212 -3412 1264
rect -3360 1212 -3346 1264
rect -3426 1198 -3346 1212
rect -2120 1218 -2040 1220
rect -2120 1166 -2106 1218
rect -2054 1166 -2040 1218
rect -2120 1146 -2040 1166
rect -2120 1094 -2106 1146
rect -2054 1094 -2040 1146
rect -2120 1074 -2040 1094
rect -2120 1022 -2106 1074
rect -2054 1022 -2040 1074
rect -2120 1002 -2040 1022
rect -2120 950 -2106 1002
rect -2054 950 -2040 1002
rect -2120 930 -2040 950
rect -2120 878 -2106 930
rect -2054 878 -2040 930
rect -2120 858 -2040 878
rect -2120 806 -2106 858
rect -2054 806 -2040 858
rect -2120 786 -2040 806
rect -2120 734 -2106 786
rect -2054 734 -2040 786
rect -2120 714 -2040 734
rect -2120 662 -2106 714
rect -2054 662 -2040 714
rect -2120 660 -2040 662
rect -2100 504 -2060 660
rect 2197 534 2277 548
rect -1676 508 -1528 522
rect -1676 504 -1662 508
rect -2100 464 -1662 504
rect -2100 310 -2060 464
rect -1676 456 -1662 464
rect -1610 456 -1594 508
rect -1542 456 -1528 508
rect -1676 442 -1528 456
rect 2197 482 2211 534
rect 2263 492 2277 534
rect 2263 482 2322 492
rect 2197 462 2322 482
rect 2197 410 2211 462
rect 2263 452 2322 462
rect 2263 410 2277 452
rect 2197 396 2277 410
rect -2120 278 -2040 310
rect -2120 226 -2106 278
rect -2054 226 -2040 278
rect -2120 206 -2040 226
rect -2120 154 -2106 206
rect -2054 154 -2040 206
rect -2120 134 -2040 154
rect -2120 82 -2106 134
rect -2054 82 -2040 134
rect -3084 58 -3004 72
rect -3084 6 -3070 58
rect -3018 6 -3004 58
rect -2120 50 -2040 82
rect -3084 -10 -3004 6
rect -3084 -62 -3070 -10
rect -3018 -16 -3004 -10
rect -1706 -10 -1554 4
rect -1706 -16 -1692 -10
rect -3018 -56 -1692 -16
rect -3018 -62 -3004 -56
rect -3084 -78 -3004 -62
rect -1706 -62 -1692 -56
rect -1640 -62 -1620 -10
rect -1568 -62 -1554 -10
rect -1706 -76 -1554 -62
rect -3084 -130 -3070 -78
rect -3018 -130 -3004 -78
rect -3084 -144 -3004 -130
rect -3198 -178 -3118 -164
rect -3198 -230 -3184 -178
rect -3132 -230 -3118 -178
rect -3198 -246 -3118 -230
rect -3198 -298 -3184 -246
rect -3132 -252 -3118 -246
rect -1481 -246 -1329 -232
rect -1481 -252 -1467 -246
rect -3132 -292 -1467 -252
rect -3132 -298 -3118 -292
rect -3198 -314 -3118 -298
rect -1481 -298 -1467 -292
rect -1415 -298 -1395 -246
rect -1343 -298 -1329 -246
rect -1481 -312 -1329 -298
rect -3198 -366 -3184 -314
rect -3132 -366 -3118 -314
rect -3198 -380 -3118 -366
rect -2120 -390 -2040 -358
rect -2120 -442 -2106 -390
rect -2054 -442 -2040 -390
rect -2120 -462 -2040 -442
rect -2120 -514 -2106 -462
rect -2054 -514 -2040 -462
rect -2120 -534 -2040 -514
rect -2120 -586 -2106 -534
rect -2054 -586 -2040 -534
rect -2120 -618 -2040 -586
rect -2100 -772 -2060 -618
rect -1691 -746 -1611 -732
rect -1691 -772 -1677 -746
rect -2100 -798 -1677 -772
rect -1625 -798 -1611 -746
rect -2100 -812 -1611 -798
rect -2100 -968 -2060 -812
rect -1691 -818 -1611 -812
rect -1691 -870 -1677 -818
rect -1625 -870 -1611 -818
rect -1691 -884 -1611 -870
rect -2120 -970 -2040 -968
rect -2120 -1022 -2106 -970
rect -2054 -1022 -2040 -970
rect -2120 -1042 -2040 -1022
rect -2120 -1094 -2106 -1042
rect -2054 -1094 -2040 -1042
rect -2120 -1114 -2040 -1094
rect -2120 -1166 -2106 -1114
rect -2054 -1166 -2040 -1114
rect -2120 -1186 -2040 -1166
rect -2120 -1238 -2106 -1186
rect -2054 -1238 -2040 -1186
rect -2120 -1258 -2040 -1238
rect -2120 -1310 -2106 -1258
rect -2054 -1310 -2040 -1258
rect -2120 -1330 -2040 -1310
rect -2120 -1382 -2106 -1330
rect -2054 -1382 -2040 -1330
rect -2120 -1402 -2040 -1382
rect -2120 -1454 -2106 -1402
rect -2054 -1454 -2040 -1402
rect -2120 -1474 -2040 -1454
rect -3312 -1524 -3232 -1510
rect -3312 -1576 -3298 -1524
rect -3246 -1576 -3232 -1524
rect -2120 -1526 -2106 -1474
rect -2054 -1526 -2040 -1474
rect -2120 -1528 -2040 -1526
rect -3312 -1592 -3232 -1576
rect -3312 -1644 -3298 -1592
rect -3246 -1598 -3232 -1592
rect -1481 -1588 -1329 -1574
rect -1481 -1598 -1467 -1588
rect -3246 -1638 -1467 -1598
rect -3246 -1644 -3232 -1638
rect -3312 -1660 -3232 -1644
rect -1481 -1640 -1467 -1638
rect -1415 -1640 -1395 -1588
rect -1343 -1640 -1329 -1588
rect -1481 -1654 -1329 -1640
rect -3312 -1712 -3298 -1660
rect -3246 -1712 -3232 -1660
rect -3312 -1726 -3232 -1712
<< labels >>
flabel metal1 s -2719 -171 -2685 -137 2 FreeSans 2500 0 0 0 GND
port 1 nsew
flabel metal1 s -3644 1408 -3583 1468 2 FreeSans 3126 0 0 0 x0
port 2 nsew
flabel metal1 s -3531 1347 -3470 1407 2 FreeSans 3126 0 0 0 x0_bar
port 3 nsew
flabel metal1 s -3416 1408 -3355 1468 2 FreeSans 3126 0 0 0 x1
port 4 nsew
flabel metal1 s -3302 1347 -3241 1407 2 FreeSans 3126 0 0 0 x1_bar
port 5 nsew
flabel metal1 s -3188 1409 -3127 1469 2 FreeSans 3126 0 0 0 x2
port 6 nsew
flabel metal1 s -3075 1348 -3014 1408 2 FreeSans 3126 0 0 0 x2_bar
port 7 nsew
flabel metal1 s -2960 1409 -2899 1469 2 FreeSans 3126 0 0 0 x3
port 8 nsew
flabel metal1 s -2846 1348 -2785 1408 2 FreeSans 3126 0 0 0 x3_bar
port 9 nsew
flabel metal1 s -2610 1408 -2576 1442 2 FreeSans 2500 0 0 0 VDD
port 10 nsew
flabel metal2 s 2220 491 2254 525 2 FreeSans 2500 0 0 0 s0
port 11 nsew
rlabel metal1 -2140 -174 -2100 -134 2 CMOS_XNOR_0/GND!
rlabel metal1 -2140 -1752 -2100 -1712 2 CMOS_XNOR_0/VDD
flabel locali -1396 -800 -1362 -766 4 FreeSans 3126 0 0 0 CMOS_XNOR_0/XNOR
flabel locali -1897 -1635 -1863 -1601 4 FreeSans 3912 0 0 0 CMOS_XNOR_0/B
flabel locali -1897 -285 -1863 -251 4 FreeSans 3912 0 0 0 CMOS_XNOR_0/A_bar
flabel locali -2347 -710 -2313 -676 4 FreeSans 3912 0 0 0 CMOS_XNOR_0/A
rlabel locali -2383 -906 -2334 -859 2 CMOS_XNOR_0/B_bar
rlabel metal1 -582 -174 -542 -134 4 CMOS_OR_1/GND!
rlabel metal1 -582 1404 -542 1444 4 CMOS_OR_1/VDD
flabel locali -204 553 -170 587 2 FreeSans 2500 0 0 0 CMOS_OR_1/OR
flabel locali -694 -57 -660 -23 2 FreeSans 2500 0 0 0 CMOS_OR_1/B
flabel locali -874 553 -840 587 2 FreeSans 2500 0 0 0 CMOS_OR_1/A
rlabel metal1 1842 -174 1882 -134 4 CMOS_OR_0/GND!
rlabel metal1 1842 1404 1882 1444 4 CMOS_OR_0/VDD
flabel locali 2220 553 2254 587 2 FreeSans 2500 0 0 0 CMOS_OR_0/OR
flabel locali 1730 -57 1764 -23 2 FreeSans 2500 0 0 0 CMOS_OR_0/B
flabel locali 1550 553 1584 587 2 FreeSans 2500 0 0 0 CMOS_OR_0/A
rlabel metal1 -582 -174 -542 -134 2 CMOS_AND_2/GND!
rlabel metal1 -582 -1752 -542 -1712 2 CMOS_AND_2/VDD
flabel locali -204 -895 -170 -861 4 FreeSans 2500 0 0 0 CMOS_AND_2/AND
flabel locali -694 -285 -660 -251 4 FreeSans 2500 0 0 0 CMOS_AND_2/A
flabel locali -874 -895 -840 -861 4 FreeSans 2500 0 0 0 CMOS_AND_2/B
rlabel metal1 630 -174 670 -134 2 CMOS_AND_1/GND!
rlabel metal1 630 -1752 670 -1712 2 CMOS_AND_1/VDD
flabel locali 1008 -895 1042 -861 4 FreeSans 2500 0 0 0 CMOS_AND_1/AND
flabel locali 518 -285 552 -251 4 FreeSans 2500 0 0 0 CMOS_AND_1/A
flabel locali 338 -895 372 -861 4 FreeSans 2500 0 0 0 CMOS_AND_1/B
rlabel metal1 630 -174 670 -134 4 CMOS_AND_0/GND!
rlabel metal1 630 1404 670 1444 4 CMOS_AND_0/VDD
flabel locali 1008 553 1042 587 2 FreeSans 2500 0 0 0 CMOS_AND_0/AND
flabel locali 518 -57 552 -23 2 FreeSans 2500 0 0 0 CMOS_AND_0/A
flabel locali 338 553 372 587 2 FreeSans 2500 0 0 0 CMOS_AND_0/B
rlabel metal1 -2140 -174 -2100 -134 4 CMOS_XOR_0/GND!
rlabel metal1 -2140 1404 -2100 1444 4 CMOS_XOR_0/VDD
flabel locali -1897 1293 -1863 1327 2 FreeSans 3126 0 0 0 CMOS_XOR_0/B
flabel locali -1897 -57 -1863 -23 2 FreeSans 3126 0 0 0 CMOS_XOR_0/A_bar
flabel locali -2347 368 -2313 402 2 FreeSans 3126 0 0 0 CMOS_XOR_0/A
rlabel locali -2383 551 -2334 598 4 CMOS_XOR_0/B_bar
<< end >>
