* NGSPICE file created from EESPFAL_s2_flat.ext - technology: sky130A

.subckt EESPFAL_s2_flat GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar Dis1 Dis3 Dis2
+ s2_bar s2 CLK2 CLK1 CLK3
X0 GND.t18 EESPFAL_3in_NOR_v2_0/C.t5 EESPFAL_3in_NOR_v2_0/C_bar.t3 GND.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_385_214# x3.t0 CLK1.t31 GND.t55 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X2 EESPFAL_NAND_v3_1/A.t2 Dis1.t0 GND.t75 GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 EESPFAL_3in_NOR_v2_0/C.t2 EESPFAL_3in_NOR_v2_0/C_bar.t5 GND.t33 GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 CLK1.t38 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/A_bar CLK1.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X5 CLK2.t22 EESPFAL_NAND_v3_1/OUT_bar.t6 EESPFAL_NAND_v3_1/OUT CLK2.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X6 CLK1.t24 EESPFAL_NAND_v3_1/A.t6 EESPFAL_NAND_v3_1/A_bar.t2 CLK1.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 CLK2.t24 EESPFAL_INV4_2/A EESPFAL_3in_NOR_v2_0/C.t1 GND.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 EESPFAL_INV4_2/A EESPFAL_INV4_2/A_bar CLK1.t3 CLK1.t2 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X9 CLK1.t43 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/B CLK1.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X10 CLK1.t8 x1.t0 a_1645_n466# GND.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X11 a_1945_n466# x1_bar.t0 CLK1.t7 GND.t20 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X12 GND.t36 s2_bar.t5 s2.t5 GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 EESPFAL_INV4_2/A EESPFAL_INV4_2/A_bar GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X14 GND.t30 EESPFAL_3in_NOR_v2_0/B EESPFAL_3in_NOR_v2_0/B_bar GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X15 EESPFAL_3in_NOR_v2_0/B EESPFAL_3in_NOR_v2_0/B_bar GND.t46 GND.t45 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X16 CLK2.t14 EESPFAL_3in_NOR_v2_0/C_bar.t6 EESPFAL_3in_NOR_v2_0/C.t4 CLK2.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 CLK2.t26 EESPFAL_NAND_v3_0/B_bar EESPFAL_3in_NOR_v2_0/B_bar GND.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 s2_bar.t3 s2.t7 GND.t38 GND.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_1645_n2607# x2.t0 EESPFAL_INV4_2/A GND.t41 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X20 EESPFAL_NAND_v3_1/B_bar EESPFAL_NAND_v3_1/B CLK1.t36 CLK1.t35 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X21 GND.t66 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar GND.t59 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X22 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar.t7 GND.t76 GND.t45 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X23 CLK1.t44 x2_bar.t0 EESPFAL_INV4_2/A_bar GND.t78 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.6e+12p ps=1.68e+07u w=1.5e+06u l=150000u
X24 EESPFAL_NAND_v3_1/A_bar.t0 EESPFAL_NAND_v3_1/A.t7 GND.t87 GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X25 s2.t0 EESPFAL_3in_NOR_v2_0/C.t6 CLK3.t0 GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X26 CLK1.t20 EESPFAL_INV4_2/A EESPFAL_INV4_2/A_bar CLK1.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X27 EESPFAL_NAND_v3_0/B_bar Dis1.t1 GND.t63 GND.t62 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X28 EESPFAL_NAND_v3_0/A_bar Dis1.t2 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X29 a_5735_214# EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/OUT GND.t58 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X30 a_85_n466# x0_bar.t0 EESPFAL_NAND_v3_0/A_bar GND.t19 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X31 a_1645_214# x2_bar.t1 EESPFAL_NAND_v3_1/A_bar.t3 GND.t42 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X32 a_85_214# x2_bar.t2 EESPFAL_NAND_v3_1/A.t1 GND.t19 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X33 CLK3.t10 s2.t8 s2_bar.t0 CLK3.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X34 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar CLK1.t52 CLK1.t51 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X35 GND.t53 EESPFAL_INV4_2/A EESPFAL_INV4_2/A_bar GND.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X36 GND.t82 Dis1.t3 EESPFAL_NAND_v3_1/B GND.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X37 EESPFAL_3in_NOR_v2_0/C_bar.t1 Dis2.t0 GND.t14 GND.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X38 EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_3in_NOR_v2_0/B CLK2.t10 CLK2.t9 sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X39 CLK2.t27 EESPFAL_NAND_v3_1/B_bar EESPFAL_NAND_v3_1/OUT_bar.t2 GND.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X40 a_1945_214# x3_bar.t0 CLK1.t11 GND.t20 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X41 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/A CLK1.t37 CLK1.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X42 EESPFAL_NAND_v3_1/OUT_bar.t0 Dis2.t1 GND.t25 GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X43 CLK1.t28 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar CLK1.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X44 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar CLK1.t41 CLK1.t40 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X45 GND.t65 Dis2.t2 EESPFAL_3in_NOR_v2_0/B GND.t64 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X46 EESPFAL_3in_NOR_v2_0/C_bar.t0 EESPFAL_INV4_2/A_bar CLK2.t0 GND.t3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X47 EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_NAND_v3_0/A_bar CLK2.t1 GND.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X48 CLK2.t6 EESPFAL_3in_NOR_v2_0/C.t7 EESPFAL_3in_NOR_v2_0/C_bar.t4 CLK2.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X49 s2.t2 Dis3.t0 GND.t57 GND.t56 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X50 EESPFAL_NAND_v3_1/A.t4 EESPFAL_NAND_v3_1/A_bar.t6 CLK1.t48 CLK1.t47 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X51 GND.t86 EESPFAL_NAND_v3_1/A_bar.t7 EESPFAL_NAND_v3_1/A.t5 GND.t67 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X52 EESPFAL_3in_NOR_v2_0/C.t0 EESPFAL_3in_NOR_v2_0/C_bar.t7 CLK2.t12 CLK2.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X53 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/A_bar GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=0p ps=0u w=1.5e+06u l=150000u
X54 CLK3.t2 EESPFAL_NAND_v3_1/OUT_bar.t8 a_6065_n2606# GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X55 CLK1.t10 x3_bar.t1 a_1945_n2607# GND.t40 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X56 GND.t68 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/A_bar GND.t67 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X57 GND.t60 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar GND.t59 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X58 s2.t6 EESPFAL_NAND_v3_1/OUT CLK3.t11 GND.t85 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X59 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar GND.t73 GND.t72 sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=0p ps=0u w=1.5e+06u l=150000u
X60 EESPFAL_NAND_v3_0/B_bar x2.t1 CLK1.t22 GND.t47 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X61 EESPFAL_NAND_v3_1/A_bar.t4 x2.t2 a_1945_214# GND.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X62 CLK3.t1 EESPFAL_3in_NOR_v2_0/B s2.t1 GND.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X63 EESPFAL_INV4_2/A_bar EESPFAL_INV4_2/A CLK1.t18 CLK1.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X64 GND.t84 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar.t5 GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X65 a_5735_n466# EESPFAL_NAND_v3_0/B EESPFAL_3in_NOR_v2_0/B GND.t58 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X66 EESPFAL_3in_NOR_v2_0/B_bar Dis2.t3 GND.t77 GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X67 CLK3.t6 s2_bar.t6 s2.t3 CLK3.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X68 CLK1.t6 x1_bar.t1 EESPFAL_INV4_2/A_bar GND.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X69 CLK1.t5 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/A CLK1.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X70 CLK1.t32 x1_bar.t2 a_85_n466# GND.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X71 CLK1.t16 x3_bar.t2 a_85_214# GND.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X72 s2_bar.t4 s2.t9 CLK3.t8 CLK3.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X73 EESPFAL_INV4_2/A_bar Dis1.t4 GND.t89 GND.t88 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X74 EESPFAL_INV4_2/A_bar x3.t1 CLK1.t29 GND.t81 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X75 CLK1.t34 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar CLK1.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X76 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar.t9 CLK2.t20 CLK2.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X77 GND.t80 Dis2.t4 EESPFAL_NAND_v3_1/OUT GND.t64 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X78 CLK2.t18 EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_3in_NOR_v2_0/B CLK2.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X79 EESPFAL_NAND_v3_1/A_bar.t1 EESPFAL_NAND_v3_1/A.t8 CLK1.t15 CLK1.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X80 GND.t34 Dis1.t5 EESPFAL_NAND_v3_1/A_bar.t5 GND.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X81 CLK2.t2 EESPFAL_NAND_v3_1/A.t9 a_5735_214# GND.t61 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X82 CLK1.t30 x3.t2 a_1645_214# GND.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X83 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_0/B CLK1.t26 CLK1.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X84 EESPFAL_NAND_v3_1/B_bar x1.t1 CLK1.t12 GND.t47 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X85 EESPFAL_NAND_v3_1/A.t0 x2.t3 a_385_214# GND.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X86 EESPFAL_NAND_v3_0/A x0.t0 a_1945_n466# GND.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X87 CLK1.t50 EESPFAL_NAND_v3_1/B_bar EESPFAL_NAND_v3_1/B CLK1.t49 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X88 GND.t12 Dis1.t6 EESPFAL_NAND_v3_0/A GND.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X89 GND.t71 Dis2.t5 EESPFAL_3in_NOR_v2_0/C.t3 GND.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X90 EESPFAL_3in_NOR_v2_0/C_bar.t2 EESPFAL_3in_NOR_v2_0/C.t8 CLK2.t4 CLK2.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X91 CLK1.t1 EESPFAL_INV4_2/A_bar EESPFAL_INV4_2/A CLK1.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X92 GND.t49 Dis1.t7 EESPFAL_NAND_v3_0/B GND.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X93 EESPFAL_NAND_v3_1/OUT_bar.t1 EESPFAL_NAND_v3_1/A_bar.t8 CLK2.t23 GND.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X94 EESPFAL_NAND_v3_1/OUT_bar.t3 EESPFAL_NAND_v3_1/OUT CLK2.t31 CLK2.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X95 EESPFAL_NAND_v3_1/B_bar Dis1.t8 GND.t79 GND.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X96 a_6065_n2606# EESPFAL_3in_NOR_v2_0/B_bar a_5915_n2606# GND.t44 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X97 CLK2.t25 EESPFAL_NAND_v3_0/A a_5735_n466# GND.t61 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X98 a_385_n466# x1.t2 CLK1.t21 GND.t55 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X99 GND.t22 Dis1.t9 EESPFAL_INV4_2/A GND.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X100 a_1645_n466# x0_bar.t1 EESPFAL_NAND_v3_0/A GND.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X101 EESPFAL_NAND_v3_0/A_bar x0.t1 a_385_n466# GND.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X102 a_5915_n2606# EESPFAL_3in_NOR_v2_0/C_bar.t8 s2_bar.t2 GND.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X103 GND.t27 Dis3.t1 s2_bar.t1 GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X104 a_1795_n2607# x0.t2 a_1645_n2607# GND.t15 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X105 s2.t4 s2_bar.t7 CLK3.t4 CLK3.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X106 CLK1.t46 EESPFAL_NAND_v3_1/A_bar.t9 EESPFAL_NAND_v3_1/A.t3 CLK1.t45 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X107 EESPFAL_INV4_2/A_bar x0_bar.t2 CLK1.t39 GND.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X108 CLK1.t9 x2_bar.t3 EESPFAL_NAND_v3_0/B GND.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X109 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar GND.t83 GND.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X110 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/A_bar CLK1.t4 CLK1.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X111 CLK1.t13 x1_bar.t3 EESPFAL_NAND_v3_1/B GND.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X112 a_1945_n2607# x1.t3 a_1795_n2607# GND.t50 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X113 CLK2.t8 EESPFAL_3in_NOR_v2_0/B EESPFAL_3in_NOR_v2_0/B_bar CLK2.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X114 CLK2.t29 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar.t4 CLK2.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X115 EESPFAL_3in_NOR_v2_0/B EESPFAL_3in_NOR_v2_0/B_bar CLK2.t16 CLK2.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
R0 EESPFAL_3in_NOR_v2_0/C.t7 EESPFAL_3in_NOR_v2_0/C.t8 819.4
R1 EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_3in_NOR_v2_0/C.t6 775.706
R2 EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_3in_NOR_v2_0/C.t7 514.133
R3 EESPFAL_3in_NOR_v2_0/C.n2 EESPFAL_3in_NOR_v2_0/C.t5 305.266
R4 EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_3in_NOR_v2_0/C.n1 166.734
R5 EESPFAL_3in_NOR_v2_0/C EESPFAL_3in_NOR_v2_0/C.n7 163.511
R6 EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_3in_NOR_v2_0/C.n5 102.4
R7 EESPFAL_3in_NOR_v2_0/C.n7 EESPFAL_3in_NOR_v2_0/C.n6 88.292
R8 EESPFAL_3in_NOR_v2_0/C.n6 EESPFAL_3in_NOR_v2_0/C.t1 81.939
R9 EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_3in_NOR_v2_0/C.n2 76
R10 EESPFAL_3in_NOR_v2_0/C.n4 EESPFAL_3in_NOR_v2_0/C.n3 57.6
R11 EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_3in_NOR_v2_0/C.n0 51.537
R12 EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_3in_NOR_v2_0/C.t4 39.4
R13 EESPFAL_3in_NOR_v2_0/C.n1 EESPFAL_3in_NOR_v2_0/C.t0 39.4
R14 EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_3in_NOR_v2_0/C.t3 24
R15 EESPFAL_3in_NOR_v2_0/C.n0 EESPFAL_3in_NOR_v2_0/C.t2 24
R16 EESPFAL_3in_NOR_v2_0/C.n5 EESPFAL_3in_NOR_v2_0/C.n4 6.4
R17 EESPFAL_3in_NOR_v2_0/C.n3 EESPFAL_INV4_2/OUT_bar 3.2
R18 EESPFAL_3in_NOR_v2_0/C_bar.t7 EESPFAL_3in_NOR_v2_0/C_bar.t6 819.4
R19 EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_3in_NOR_v2_0/C_bar.t5 506.1
R20 EESPFAL_3in_NOR_v2_0/C_bar.n5 EESPFAL_3in_NOR_v2_0/C_bar.t7 313.3
R21 EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_3in_NOR_v2_0/C_bar.t8 305.997
R22 EESPFAL_INV4_2/OUT EESPFAL_3in_NOR_v2_0/C_bar.n0 210.945
R23 EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_3in_NOR_v2_0/C_bar.t0 187.539
R24 EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_3in_NOR_v2_0/C_bar.n1 128.334
R25 EESPFAL_3in_NOR_v2_0/C_bar.n0 EESPFAL_3in_NOR_v2_0/C_bar 115.2
R26 EESPFAL_3in_NOR_v2_0/C_bar.n3 EESPFAL_3in_NOR_v2_0/C_bar.n2 57.937
R27 EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_3in_NOR_v2_0/C_bar.n4 57.6
R28 EESPFAL_3in_NOR_v2_0/C_bar.n4 EESPFAL_3in_NOR_v2_0/C_bar.n3 41.6
R29 EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_3in_NOR_v2_0/C_bar.t4 39.4
R30 EESPFAL_3in_NOR_v2_0/C_bar.n1 EESPFAL_3in_NOR_v2_0/C_bar.t2 39.4
R31 EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_3in_NOR_v2_0/C_bar.t3 24
R32 EESPFAL_3in_NOR_v2_0/C_bar.n2 EESPFAL_3in_NOR_v2_0/C_bar.t1 24
R33 EESPFAL_3in_NOR_v2_0/C_bar.n6 EESPFAL_3in_NOR_v2_0/C_bar.n5 8.764
R34 EESPFAL_INV4_2/OUT EESPFAL_3in_NOR_v2_0/C_bar.n6 4.65
R35 GND.n413 GND.n412 341.085
R36 GND.n421 GND.n253 341.085
R37 GND.n423 GND.n422 341.085
R38 GND.n432 GND.n247 341.085
R39 GND.n433 GND.n432 341.085
R40 GND.n434 GND.n433 341.085
R41 GND.n445 GND.n241 341.085
R42 GND.n448 GND.n447 341.085
R43 GND.n458 GND.n457 341.085
R44 GND.n460 GND.n458 341.085
R45 GND.n460 GND.n459 341.085
R46 GND.n469 GND.n468 341.085
R47 GND.n471 GND.n470 341.085
R48 GND.n480 GND.n479 341.085
R49 GND.n319 GND.n318 341.085
R50 GND.n320 GND.n305 341.085
R51 GND.n329 GND.n305 341.085
R52 GND.n330 GND.n329 341.085
R53 GND.n332 GND.n331 341.085
R54 GND.n342 GND.n341 341.085
R55 GND.n351 GND.n292 341.085
R56 GND.n352 GND.n351 341.085
R57 GND.n353 GND.n352 341.085
R58 GND.n361 GND.n286 341.085
R59 GND.n373 GND.n372 341.085
R60 GND.n375 GND.n373 341.085
R61 GND.n375 GND.n374 341.085
R62 GND.n385 GND.n384 341.085
R63 GND.n395 GND.n268 341.085
R64 GND.n397 GND.n396 341.085
R65 GND.n397 GND.n262 341.085
R66 GND.n405 GND.n262 341.085
R67 GND.t42 GND.n247 319.767
R68 GND.n446 GND.t6 319.767
R69 GND.t67 GND.n446 319.767
R70 GND.n459 GND.t9 319.767
R71 GND.n320 GND.t58 319.767
R72 GND.n340 GND.t45 319.767
R73 GND.t29 GND.n340 319.767
R74 GND.n353 GND.t8 319.767
R75 GND.n372 GND.t39 319.767
R76 GND.n386 GND.t72 319.767
R77 GND.n386 GND.t59 319.767
R78 GND.t47 GND.n405 319.767
R79 GND.n422 GND.t23 277.131
R80 GND.t11 GND.n241 277.131
R81 GND.n447 GND.t0 277.131
R82 GND.t55 GND.n469 277.131
R83 GND.n318 GND.t61 277.131
R84 GND.n332 GND.t64 277.131
R85 GND.n342 GND.t24 277.131
R86 GND.t74 GND.n361 277.131
R87 GND.n384 GND.t48 277.131
R88 GND.t62 GND.n395 277.131
R89 GND.n167 GND.t40 267.309
R90 GND.n484 GND.t78 267.309
R91 GND.t20 GND.n253 234.496
R92 GND.n470 GND.t51 234.496
R93 GND.n93 GND.t85 192.984
R94 GND.n3 GND.t2 192.984
R95 GND.n412 GND.t43 191.86
R96 GND.t19 GND.n480 191.86
R97 GND.n175 GND.t50 185.81
R98 GND.n492 GND.t69 185.81
R99 GND.t43 GND.n411 158.378
R100 GND.n481 GND.t19 158.378
R101 GND.n411 GND.n258 157.6
R102 GND.n414 GND.n258 157.6
R103 GND.n414 GND.n254 157.6
R104 GND.n420 GND.n254 157.6
R105 GND.n420 GND.n252 157.6
R106 GND.n424 GND.n252 157.6
R107 GND.n424 GND.n248 157.6
R108 GND.n431 GND.n248 157.6
R109 GND.n431 GND.n246 157.6
R110 GND.n435 GND.n246 157.6
R111 GND.n435 GND.n242 157.6
R112 GND.n444 GND.n242 157.6
R113 GND.n444 GND.n240 157.6
R114 GND.n449 GND.n240 157.6
R115 GND.n449 GND.n237 157.6
R116 GND.n456 GND.n237 157.6
R117 GND.n456 GND.n236 157.6
R118 GND.n461 GND.n236 157.6
R119 GND.n461 GND.n232 157.6
R120 GND.n467 GND.n232 157.6
R121 GND.n467 GND.n231 157.6
R122 GND.n472 GND.n231 157.6
R123 GND.n472 GND.n226 157.6
R124 GND.n478 GND.n226 157.6
R125 GND.n478 GND.n225 157.6
R126 GND.n481 GND.n225 157.6
R127 GND.n317 GND.n311 157.6
R128 GND.n317 GND.n310 157.6
R129 GND.n321 GND.n310 157.6
R130 GND.n321 GND.n306 157.6
R131 GND.n328 GND.n306 157.6
R132 GND.n328 GND.n304 157.6
R133 GND.n333 GND.n304 157.6
R134 GND.n333 GND.n298 157.6
R135 GND.n339 GND.n298 157.6
R136 GND.n339 GND.n297 157.6
R137 GND.n343 GND.n297 157.6
R138 GND.n343 GND.n293 157.6
R139 GND.n350 GND.n293 157.6
R140 GND.n350 GND.n291 157.6
R141 GND.n354 GND.n291 157.6
R142 GND.n354 GND.n287 157.6
R143 GND.n360 GND.n287 157.6
R144 GND.n360 GND.n285 157.6
R145 GND.n371 GND.n281 157.6
R146 GND.n371 GND.n280 157.6
R147 GND.n376 GND.n280 157.6
R148 GND.n376 GND.n276 157.6
R149 GND.n383 GND.n276 157.6
R150 GND.n383 GND.n275 157.6
R151 GND.n387 GND.n275 157.6
R152 GND.n387 GND.n269 157.6
R153 GND.n394 GND.n269 157.6
R154 GND.n394 GND.n267 157.6
R155 GND.n398 GND.n267 157.6
R156 GND.n398 GND.n263 157.6
R157 GND.n404 GND.n263 157.6
R158 GND.n404 GND.n261 157.6
R159 GND.n314 GND.n313 118.661
R160 GND.n363 GND.n362 115.922
R161 GND.n366 GND.n365 115.922
R162 GND.n407 GND.n406 115.922
R163 GND.n118 GND.t70 111.486
R164 GND.n142 GND.t13 111.486
R165 GND.n11 GND.t44 111.486
R166 GND.n36 GND.t26 111.486
R167 GND.n60 GND.t56 111.486
R168 GND.n85 GND.t28 111.486
R169 GND.n183 GND.t15 111.486
R170 GND.n208 GND.t21 111.486
R171 GND.n525 GND.t88 111.486
R172 GND.n500 GND.t10 111.486
R173 GND.n413 GND.t20 106.589
R174 GND.n479 GND.t51 106.589
R175 GND.n313 GND.t61 70.155
R176 GND.n362 GND.t74 70.155
R177 GND.t23 GND.n421 63.953
R178 GND.n434 GND.t11 63.953
R179 GND.n457 GND.t0 63.953
R180 GND.n471 GND.t55 63.953
R181 GND.t64 GND.n330 63.953
R182 GND.t24 GND.n292 63.953
R183 GND.n374 GND.t48 63.953
R184 GND.n396 GND.t62 63.953
R185 GND.n159 GND.t3 44.336
R186 GND.n101 GND.t54 44.336
R187 GND GND.n482 37.956
R188 GND.n126 GND.t32 37.162
R189 GND.n134 GND.t17 37.162
R190 GND.n19 GND.t31 37.162
R191 GND.n44 GND.t37 37.162
R192 GND.n52 GND.t35 37.162
R193 GND.n77 GND.t16 37.162
R194 GND.n191 GND.t41 37.162
R195 GND.n216 GND.t4 37.162
R196 GND.n533 GND.t52 37.162
R197 GND.n508 GND.t81 37.162
R198 GND.n483 GND 29.511
R199 GND.n325 GND.t80 29.103
R200 GND.n347 GND.t25 29.103
R201 GND.n379 GND.t82 29.103
R202 GND.n265 GND.t79 29.103
R203 GND.n244 GND.t34 29.103
R204 GND.n453 GND.t75 29.103
R205 GND.n35 GND.t27 29.103
R206 GND.n64 GND.t57 29.103
R207 GND.n117 GND.t71 29.103
R208 GND.n146 GND.t14 29.103
R209 GND.n207 GND.t22 29.103
R210 GND.n524 GND.t89 29.103
R211 GND.n325 GND.t65 29.102
R212 GND.n347 GND.t77 29.102
R213 GND.n379 GND.t49 29.102
R214 GND.n265 GND.t63 29.102
R215 GND.n244 GND.t12 29.102
R216 GND.n453 GND.t1 29.102
R217 GND.n365 GND.t39 27.519
R218 GND.n406 GND.t47 27.519
R219 GND.n440 GND.t7 24
R220 GND.n440 GND.t68 24
R221 GND.n439 GND.t87 24
R222 GND.n439 GND.t86 24
R223 GND.n301 GND.t46 24
R224 GND.n301 GND.t30 24
R225 GND.n300 GND.t76 24
R226 GND.n300 GND.t84 24
R227 GND.n272 GND.t73 24
R228 GND.n272 GND.t60 24
R229 GND.n271 GND.t83 24
R230 GND.n271 GND.t66 24
R231 GND.n0 GND.t5 24
R232 GND.n0 GND.t53 24
R233 GND.n1 GND.t33 24
R234 GND.n1 GND.t18 24
R235 GND.n2 GND.t38 24
R236 GND.n2 GND.t36 24
R237 GND.n423 GND.t42 21.317
R238 GND.t6 GND.n445 21.317
R239 GND.n448 GND.t67 21.317
R240 GND.n468 GND.t9 21.317
R241 GND.t58 GND.n319 21.317
R242 GND.n331 GND.t45 21.317
R243 GND.n341 GND.t29 21.317
R244 GND.t8 GND.n286 21.317
R245 GND.t72 GND.n385 21.317
R246 GND.t59 GND.n268 21.317
R247 GND.n316 GND.n312 12.8
R248 GND.n316 GND.n309 12.8
R249 GND.n322 GND.n309 12.8
R250 GND.n322 GND.n307 12.8
R251 GND.n327 GND.n307 12.8
R252 GND.n327 GND.n303 12.8
R253 GND.n334 GND.n303 12.8
R254 GND.n334 GND.n299 12.8
R255 GND.n338 GND.n299 12.8
R256 GND.n338 GND.n296 12.8
R257 GND.n344 GND.n296 12.8
R258 GND.n344 GND.n294 12.8
R259 GND.n349 GND.n294 12.8
R260 GND.n349 GND.n290 12.8
R261 GND.n355 GND.n290 12.8
R262 GND.n355 GND.n288 12.8
R263 GND.n359 GND.n288 12.8
R264 GND.n359 GND.n284 12.8
R265 GND.n363 GND.n284 12.8
R266 GND.n366 GND.n282 12.8
R267 GND.n370 GND.n282 12.8
R268 GND.n370 GND.n279 12.8
R269 GND.n377 GND.n279 12.8
R270 GND.n377 GND.n277 12.8
R271 GND.n382 GND.n277 12.8
R272 GND.n382 GND.n274 12.8
R273 GND.n388 GND.n274 12.8
R274 GND.n388 GND.n270 12.8
R275 GND.n393 GND.n270 12.8
R276 GND.n393 GND.n266 12.8
R277 GND.n399 GND.n266 12.8
R278 GND.n399 GND.n264 12.8
R279 GND.n403 GND.n264 12.8
R280 GND.n403 GND.n260 12.8
R281 GND.n407 GND.n260 12.8
R282 GND.n410 GND.n257 12.8
R283 GND.n415 GND.n257 12.8
R284 GND.n415 GND.n255 12.8
R285 GND.n419 GND.n255 12.8
R286 GND.n419 GND.n251 12.8
R287 GND.n425 GND.n251 12.8
R288 GND.n425 GND.n249 12.8
R289 GND.n430 GND.n249 12.8
R290 GND.n430 GND.n245 12.8
R291 GND.n436 GND.n245 12.8
R292 GND.n436 GND.n243 12.8
R293 GND.n443 GND.n243 12.8
R294 GND.n443 GND.n239 12.8
R295 GND.n450 GND.n239 12.8
R296 GND.n450 GND.n238 12.8
R297 GND.n455 GND.n238 12.8
R298 GND.n455 GND.n235 12.8
R299 GND.n462 GND.n235 12.8
R300 GND.n462 GND.n233 12.8
R301 GND.n466 GND.n233 12.8
R302 GND.n466 GND.n230 12.8
R303 GND.n473 GND.n230 12.8
R304 GND.n473 GND.n227 12.8
R305 GND.n477 GND.n227 12.8
R306 GND.n477 GND.n228 12.8
R307 GND.n136 GND.n133 12.8
R308 GND.n54 GND.n51 12.8
R309 GND.n312 GND.n311 9.154
R310 GND.n282 GND.n281 9.154
R311 GND.n371 GND.n370 9.154
R312 GND.n372 GND.n371 9.154
R313 GND.n280 GND.n279 9.154
R314 GND.n373 GND.n280 9.154
R315 GND.n377 GND.n376 9.154
R316 GND.n376 GND.n375 9.154
R317 GND.n277 GND.n276 9.154
R318 GND.n374 GND.n276 9.154
R319 GND.n383 GND.n382 9.154
R320 GND.n384 GND.n383 9.154
R321 GND.n275 GND.n274 9.154
R322 GND.n385 GND.n275 9.154
R323 GND.n388 GND.n387 9.154
R324 GND.n387 GND.n386 9.154
R325 GND.n270 GND.n269 9.154
R326 GND.n269 GND.n268 9.154
R327 GND.n394 GND.n393 9.154
R328 GND.n395 GND.n394 9.154
R329 GND.n267 GND.n266 9.154
R330 GND.n396 GND.n267 9.154
R331 GND.n399 GND.n398 9.154
R332 GND.n398 GND.n397 9.154
R333 GND.n264 GND.n263 9.154
R334 GND.n263 GND.n262 9.154
R335 GND.n404 GND.n403 9.154
R336 GND.n405 GND.n404 9.154
R337 GND.n261 GND.n260 9.154
R338 GND.n317 GND.n316 9.154
R339 GND.n318 GND.n317 9.154
R340 GND.n310 GND.n309 9.154
R341 GND.n319 GND.n310 9.154
R342 GND.n322 GND.n321 9.154
R343 GND.n321 GND.n320 9.154
R344 GND.n307 GND.n306 9.154
R345 GND.n306 GND.n305 9.154
R346 GND.n328 GND.n327 9.154
R347 GND.n329 GND.n328 9.154
R348 GND.n304 GND.n303 9.154
R349 GND.n330 GND.n304 9.154
R350 GND.n334 GND.n333 9.154
R351 GND.n333 GND.n332 9.154
R352 GND.n299 GND.n298 9.154
R353 GND.n331 GND.n298 9.154
R354 GND.n339 GND.n338 9.154
R355 GND.n340 GND.n339 9.154
R356 GND.n297 GND.n296 9.154
R357 GND.n341 GND.n297 9.154
R358 GND.n344 GND.n343 9.154
R359 GND.n343 GND.n342 9.154
R360 GND.n294 GND.n293 9.154
R361 GND.n293 GND.n292 9.154
R362 GND.n350 GND.n349 9.154
R363 GND.n351 GND.n350 9.154
R364 GND.n291 GND.n290 9.154
R365 GND.n352 GND.n291 9.154
R366 GND.n355 GND.n354 9.154
R367 GND.n354 GND.n353 9.154
R368 GND.n288 GND.n287 9.154
R369 GND.n287 GND.n286 9.154
R370 GND.n360 GND.n359 9.154
R371 GND.n361 GND.n360 9.154
R372 GND.n285 GND.n284 9.154
R373 GND.n258 GND.n257 9.154
R374 GND.n412 GND.n258 9.154
R375 GND.n415 GND.n414 9.154
R376 GND.n414 GND.n413 9.154
R377 GND.n255 GND.n254 9.154
R378 GND.n254 GND.n253 9.154
R379 GND.n420 GND.n419 9.154
R380 GND.n421 GND.n420 9.154
R381 GND.n252 GND.n251 9.154
R382 GND.n422 GND.n252 9.154
R383 GND.n425 GND.n424 9.154
R384 GND.n424 GND.n423 9.154
R385 GND.n249 GND.n248 9.154
R386 GND.n248 GND.n247 9.154
R387 GND.n431 GND.n430 9.154
R388 GND.n432 GND.n431 9.154
R389 GND.n246 GND.n245 9.154
R390 GND.n433 GND.n246 9.154
R391 GND.n436 GND.n435 9.154
R392 GND.n435 GND.n434 9.154
R393 GND.n243 GND.n242 9.154
R394 GND.n242 GND.n241 9.154
R395 GND.n444 GND.n443 9.154
R396 GND.n445 GND.n444 9.154
R397 GND.n240 GND.n239 9.154
R398 GND.n446 GND.n240 9.154
R399 GND.n450 GND.n449 9.154
R400 GND.n449 GND.n448 9.154
R401 GND.n238 GND.n237 9.154
R402 GND.n447 GND.n237 9.154
R403 GND.n456 GND.n455 9.154
R404 GND.n457 GND.n456 9.154
R405 GND.n236 GND.n235 9.154
R406 GND.n458 GND.n236 9.154
R407 GND.n462 GND.n461 9.154
R408 GND.n461 GND.n460 9.154
R409 GND.n233 GND.n232 9.154
R410 GND.n459 GND.n232 9.154
R411 GND.n467 GND.n466 9.154
R412 GND.n468 GND.n467 9.154
R413 GND.n231 GND.n230 9.154
R414 GND.n469 GND.n231 9.154
R415 GND.n473 GND.n472 9.154
R416 GND.n472 GND.n471 9.154
R417 GND.n227 GND.n226 9.154
R418 GND.n470 GND.n226 9.154
R419 GND.n478 GND.n477 9.154
R420 GND.n479 GND.n478 9.154
R421 GND.n228 GND.n225 9.154
R422 GND.n480 GND.n225 9.154
R423 GND.n482 GND.n481 9.154
R424 GND.n411 GND.n410 9.154
R425 GND.n5 GND.n4 9.154
R426 GND.n9 GND.n8 9.154
R427 GND.n8 GND.n7 9.154
R428 GND.n13 GND.n12 9.154
R429 GND.n12 GND.n11 9.154
R430 GND.n17 GND.n16 9.154
R431 GND.n16 GND.n15 9.154
R432 GND.n21 GND.n20 9.154
R433 GND.n20 GND.n19 9.154
R434 GND.n25 GND.n24 9.154
R435 GND.n24 GND.n23 9.154
R436 GND.n29 GND.n28 9.154
R437 GND.n28 GND.n27 9.154
R438 GND.n33 GND.n32 9.154
R439 GND.n32 GND.n31 9.154
R440 GND.n38 GND.n37 9.154
R441 GND.n37 GND.n36 9.154
R442 GND.n42 GND.n41 9.154
R443 GND.n41 GND.n40 9.154
R444 GND.n46 GND.n45 9.154
R445 GND.n45 GND.n44 9.154
R446 GND.n51 GND.n50 9.154
R447 GND.n50 GND.n49 9.154
R448 GND.n54 GND.n53 9.154
R449 GND.n53 GND.n52 9.154
R450 GND.n58 GND.n57 9.154
R451 GND.n57 GND.n56 9.154
R452 GND.n62 GND.n61 9.154
R453 GND.n61 GND.n60 9.154
R454 GND.n67 GND.n66 9.154
R455 GND.n66 GND.n65 9.154
R456 GND.n71 GND.n70 9.154
R457 GND.n70 GND.n69 9.154
R458 GND.n75 GND.n74 9.154
R459 GND.n74 GND.n73 9.154
R460 GND.n79 GND.n78 9.154
R461 GND.n78 GND.n77 9.154
R462 GND.n83 GND.n82 9.154
R463 GND.n82 GND.n81 9.154
R464 GND.n87 GND.n86 9.154
R465 GND.n86 GND.n85 9.154
R466 GND.n91 GND.n90 9.154
R467 GND.n90 GND.n89 9.154
R468 GND.n95 GND.n94 9.154
R469 GND.n103 GND.n102 9.154
R470 GND.n107 GND.n106 9.154
R471 GND.n106 GND.n105 9.154
R472 GND.n111 GND.n110 9.154
R473 GND.n110 GND.n109 9.154
R474 GND.n115 GND.n114 9.154
R475 GND.n114 GND.n113 9.154
R476 GND.n120 GND.n119 9.154
R477 GND.n119 GND.n118 9.154
R478 GND.n124 GND.n123 9.154
R479 GND.n123 GND.n122 9.154
R480 GND.n128 GND.n127 9.154
R481 GND.n127 GND.n126 9.154
R482 GND.n133 GND.n132 9.154
R483 GND.n132 GND.n131 9.154
R484 GND.n136 GND.n135 9.154
R485 GND.n135 GND.n134 9.154
R486 GND.n140 GND.n139 9.154
R487 GND.n139 GND.n138 9.154
R488 GND.n144 GND.n143 9.154
R489 GND.n143 GND.n142 9.154
R490 GND.n149 GND.n148 9.154
R491 GND.n148 GND.n147 9.154
R492 GND.n153 GND.n152 9.154
R493 GND.n152 GND.n151 9.154
R494 GND.n157 GND.n156 9.154
R495 GND.n156 GND.n155 9.154
R496 GND.n161 GND.n160 9.154
R497 GND.n169 GND.n168 9.154
R498 GND.n173 GND.n172 9.154
R499 GND.n172 GND.n171 9.154
R500 GND.n177 GND.n176 9.154
R501 GND.n176 GND.n175 9.154
R502 GND.n181 GND.n180 9.154
R503 GND.n180 GND.n179 9.154
R504 GND.n185 GND.n184 9.154
R505 GND.n184 GND.n183 9.154
R506 GND.n189 GND.n188 9.154
R507 GND.n188 GND.n187 9.154
R508 GND.n193 GND.n192 9.154
R509 GND.n192 GND.n191 9.154
R510 GND.n197 GND.n196 9.154
R511 GND.n196 GND.n195 9.154
R512 GND.n201 GND.n200 9.154
R513 GND.n200 GND.n199 9.154
R514 GND.n205 GND.n204 9.154
R515 GND.n204 GND.n203 9.154
R516 GND.n210 GND.n209 9.154
R517 GND.n209 GND.n208 9.154
R518 GND.n214 GND.n213 9.154
R519 GND.n213 GND.n212 9.154
R520 GND.n218 GND.n217 9.154
R521 GND.n217 GND.n216 9.154
R522 GND.n222 GND.n221 9.154
R523 GND.n221 GND.n220 9.154
R524 GND.n535 GND.n534 9.154
R525 GND.n534 GND.n533 9.154
R526 GND.n531 GND.n530 9.154
R527 GND.n530 GND.n529 9.154
R528 GND.n527 GND.n526 9.154
R529 GND.n526 GND.n525 9.154
R530 GND.n522 GND.n521 9.154
R531 GND.n521 GND.n520 9.154
R532 GND.n518 GND.n517 9.154
R533 GND.n517 GND.n516 9.154
R534 GND.n514 GND.n513 9.154
R535 GND.n513 GND.n512 9.154
R536 GND.n510 GND.n509 9.154
R537 GND.n509 GND.n508 9.154
R538 GND.n506 GND.n505 9.154
R539 GND.n505 GND.n504 9.154
R540 GND.n502 GND.n501 9.154
R541 GND.n501 GND.n500 9.154
R542 GND.n498 GND.n497 9.154
R543 GND.n497 GND.n496 9.154
R544 GND.n494 GND.n493 9.154
R545 GND.n493 GND.n492 9.154
R546 GND.n490 GND.n489 9.154
R547 GND.n489 GND.n488 9.154
R548 GND.n486 GND.n485 9.154
R549 GND.n441 GND.n440 5.103
R550 GND.n441 GND.n439 5.103
R551 GND.n337 GND.n301 5.103
R552 GND.n337 GND.n300 5.103
R553 GND.n389 GND.n272 5.103
R554 GND.n389 GND.n271 5.103
R555 GND.n223 GND.n0 5.103
R556 GND.n130 GND.n1 5.103
R557 GND.n48 GND.n2 5.103
R558 GND.n408 GND.n407 4.65
R559 GND.n368 GND.n282 4.65
R560 GND.n370 GND.n369 4.65
R561 GND.n279 GND.n278 4.65
R562 GND.n378 GND.n377 4.65
R563 GND.n380 GND.n277 4.65
R564 GND.n382 GND.n381 4.65
R565 GND.n274 GND.n273 4.65
R566 GND.n389 GND.n388 4.65
R567 GND.n390 GND.n270 4.65
R568 GND.n393 GND.n392 4.65
R569 GND.n391 GND.n266 4.65
R570 GND.n400 GND.n399 4.65
R571 GND.n401 GND.n264 4.65
R572 GND.n403 GND.n402 4.65
R573 GND.n260 GND.n259 4.65
R574 GND.n367 GND.n366 4.65
R575 GND.n364 GND.n363 4.65
R576 GND.n316 GND.n315 4.65
R577 GND.n309 GND.n308 4.65
R578 GND.n323 GND.n322 4.65
R579 GND.n324 GND.n307 4.65
R580 GND.n327 GND.n326 4.65
R581 GND.n303 GND.n302 4.65
R582 GND.n335 GND.n334 4.65
R583 GND.n336 GND.n299 4.65
R584 GND.n338 GND.n337 4.65
R585 GND.n296 GND.n295 4.65
R586 GND.n345 GND.n344 4.65
R587 GND.n346 GND.n294 4.65
R588 GND.n349 GND.n348 4.65
R589 GND.n290 GND.n289 4.65
R590 GND.n356 GND.n355 4.65
R591 GND.n357 GND.n288 4.65
R592 GND.n359 GND.n358 4.65
R593 GND.n284 GND.n283 4.65
R594 GND.n257 GND.n256 4.65
R595 GND.n416 GND.n415 4.65
R596 GND.n417 GND.n255 4.65
R597 GND.n419 GND.n418 4.65
R598 GND.n251 GND.n250 4.65
R599 GND.n426 GND.n425 4.65
R600 GND.n427 GND.n249 4.65
R601 GND.n430 GND.n429 4.65
R602 GND.n428 GND.n245 4.65
R603 GND.n437 GND.n436 4.65
R604 GND.n438 GND.n243 4.65
R605 GND.n443 GND.n442 4.65
R606 GND.n441 GND.n239 4.65
R607 GND.n451 GND.n450 4.65
R608 GND.n452 GND.n238 4.65
R609 GND.n455 GND.n454 4.65
R610 GND.n235 GND.n234 4.65
R611 GND.n463 GND.n462 4.65
R612 GND.n464 GND.n233 4.65
R613 GND.n466 GND.n465 4.65
R614 GND.n230 GND.n229 4.65
R615 GND.n474 GND.n473 4.65
R616 GND.n475 GND.n227 4.65
R617 GND.n477 GND.n476 4.65
R618 GND.n410 GND.n409 4.65
R619 GND.n10 GND.n9 4.65
R620 GND.n14 GND.n13 4.65
R621 GND.n18 GND.n17 4.65
R622 GND.n22 GND.n21 4.65
R623 GND.n26 GND.n25 4.65
R624 GND.n30 GND.n29 4.65
R625 GND.n34 GND.n33 4.65
R626 GND.n39 GND.n38 4.65
R627 GND.n43 GND.n42 4.65
R628 GND.n47 GND.n46 4.65
R629 GND.n51 GND.n48 4.65
R630 GND.n55 GND.n54 4.65
R631 GND.n59 GND.n58 4.65
R632 GND.n63 GND.n62 4.65
R633 GND.n68 GND.n67 4.65
R634 GND.n72 GND.n71 4.65
R635 GND.n76 GND.n75 4.65
R636 GND.n80 GND.n79 4.65
R637 GND.n84 GND.n83 4.65
R638 GND.n88 GND.n87 4.65
R639 GND.n92 GND.n91 4.65
R640 GND.n96 GND.n95 4.65
R641 GND.n98 GND.n97 4.65
R642 GND.n100 GND.n99 4.65
R643 GND.n104 GND.n103 4.65
R644 GND.n108 GND.n107 4.65
R645 GND.n112 GND.n111 4.65
R646 GND.n116 GND.n115 4.65
R647 GND.n121 GND.n120 4.65
R648 GND.n125 GND.n124 4.65
R649 GND.n129 GND.n128 4.65
R650 GND.n133 GND.n130 4.65
R651 GND.n137 GND.n136 4.65
R652 GND.n141 GND.n140 4.65
R653 GND.n145 GND.n144 4.65
R654 GND.n150 GND.n149 4.65
R655 GND.n154 GND.n153 4.65
R656 GND.n158 GND.n157 4.65
R657 GND.n162 GND.n161 4.65
R658 GND.n164 GND.n163 4.65
R659 GND.n166 GND.n165 4.65
R660 GND.n170 GND.n169 4.65
R661 GND.n174 GND.n173 4.65
R662 GND.n178 GND.n177 4.65
R663 GND.n182 GND.n181 4.65
R664 GND.n186 GND.n185 4.65
R665 GND.n190 GND.n189 4.65
R666 GND.n194 GND.n193 4.65
R667 GND.n198 GND.n197 4.65
R668 GND.n202 GND.n201 4.65
R669 GND.n206 GND.n205 4.65
R670 GND.n211 GND.n210 4.65
R671 GND.n215 GND.n214 4.65
R672 GND.n219 GND.n218 4.65
R673 GND.n223 GND.n222 4.65
R674 GND.n536 GND.n535 4.65
R675 GND.n532 GND.n531 4.65
R676 GND.n528 GND.n527 4.65
R677 GND.n523 GND.n522 4.65
R678 GND.n519 GND.n518 4.65
R679 GND.n515 GND.n514 4.65
R680 GND.n511 GND.n510 4.65
R681 GND.n507 GND.n506 4.65
R682 GND.n503 GND.n502 4.65
R683 GND.n499 GND.n498 4.65
R684 GND.n495 GND.n494 4.65
R685 GND.n491 GND.n490 4.65
R686 GND.n313 GND.n311 2.791
R687 GND.n365 GND.n281 2.791
R688 GND.n406 GND.n261 2.791
R689 GND.n362 GND.n285 2.791
R690 GND.n482 GND.n224 2.739
R691 GND.n487 GND.n483 2.739
R692 GND.n6 GND.n5 2.682
R693 GND.n314 GND.n312 2.682
R694 GND.n228 GND.n224 2.682
R695 GND.n487 GND.n486 2.682
R696 GND.n4 GND.n3 1.873
R697 GND.n102 GND.n101 1.873
R698 GND.n485 GND.n484 1.873
R699 GND.n94 GND.n93 1.873
R700 GND.n160 GND.n159 1.873
R701 GND.n168 GND.n167 1.873
R702 GND.n10 GND.n6 1.096
R703 GND.n315 GND.n314 1.095
R704 GND.n476 GND.n224 1.095
R705 GND.n491 GND.n487 1.095
R706 GND.n409 GND.n408 0.662
R707 GND.n100 GND.n98 0.573
R708 GND.n166 GND.n164 0.563
R709 GND.n367 GND.n364 0.55
R710 GND.n315 GND.n308 0.1
R711 GND.n323 GND.n308 0.1
R712 GND.n324 GND.n323 0.1
R713 GND.n326 GND.n324 0.1
R714 GND.n335 GND.n302 0.1
R715 GND.n336 GND.n335 0.1
R716 GND.n337 GND.n336 0.1
R717 GND.n345 GND.n295 0.1
R718 GND.n346 GND.n345 0.1
R719 GND.n348 GND.n289 0.1
R720 GND.n356 GND.n289 0.1
R721 GND.n357 GND.n356 0.1
R722 GND.n358 GND.n357 0.1
R723 GND.n358 GND.n283 0.1
R724 GND.n364 GND.n283 0.1
R725 GND.n368 GND.n367 0.1
R726 GND.n369 GND.n368 0.1
R727 GND.n369 GND.n278 0.1
R728 GND.n378 GND.n278 0.1
R729 GND.n381 GND.n380 0.1
R730 GND.n381 GND.n273 0.1
R731 GND.n389 GND.n273 0.1
R732 GND.n392 GND.n390 0.1
R733 GND.n392 GND.n391 0.1
R734 GND.n401 GND.n400 0.1
R735 GND.n402 GND.n401 0.1
R736 GND.n402 GND.n259 0.1
R737 GND.n408 GND.n259 0.1
R738 GND.n409 GND.n256 0.1
R739 GND.n416 GND.n256 0.1
R740 GND.n417 GND.n416 0.1
R741 GND.n418 GND.n417 0.1
R742 GND.n418 GND.n250 0.1
R743 GND.n426 GND.n250 0.1
R744 GND.n427 GND.n426 0.1
R745 GND.n429 GND.n427 0.1
R746 GND.n429 GND.n428 0.1
R747 GND.n438 GND.n437 0.1
R748 GND.n442 GND.n438 0.1
R749 GND.n442 GND.n441 0.1
R750 GND.n452 GND.n451 0.1
R751 GND.n454 GND.n452 0.1
R752 GND.n463 GND.n234 0.1
R753 GND.n464 GND.n463 0.1
R754 GND.n465 GND.n464 0.1
R755 GND.n465 GND.n229 0.1
R756 GND.n474 GND.n229 0.1
R757 GND.n475 GND.n474 0.1
R758 GND.n476 GND.n475 0.1
R759 GND.n14 GND.n10 0.1
R760 GND.n18 GND.n14 0.1
R761 GND.n22 GND.n18 0.1
R762 GND.n26 GND.n22 0.1
R763 GND.n30 GND.n26 0.1
R764 GND.n34 GND.n30 0.1
R765 GND.n43 GND.n39 0.1
R766 GND.n47 GND.n43 0.1
R767 GND.n48 GND.n47 0.1
R768 GND.n59 GND.n55 0.1
R769 GND.n63 GND.n59 0.1
R770 GND.n72 GND.n68 0.1
R771 GND.n76 GND.n72 0.1
R772 GND.n80 GND.n76 0.1
R773 GND.n84 GND.n80 0.1
R774 GND.n88 GND.n84 0.1
R775 GND.n92 GND.n88 0.1
R776 GND.n96 GND.n92 0.1
R777 GND.n98 GND.n96 0.1
R778 GND.n104 GND.n100 0.1
R779 GND.n108 GND.n104 0.1
R780 GND.n112 GND.n108 0.1
R781 GND.n116 GND.n112 0.1
R782 GND.n125 GND.n121 0.1
R783 GND.n129 GND.n125 0.1
R784 GND.n130 GND.n129 0.1
R785 GND.n141 GND.n137 0.1
R786 GND.n145 GND.n141 0.1
R787 GND.n154 GND.n150 0.1
R788 GND.n158 GND.n154 0.1
R789 GND.n162 GND.n158 0.1
R790 GND.n164 GND.n162 0.1
R791 GND.n170 GND.n166 0.1
R792 GND.n174 GND.n170 0.1
R793 GND.n178 GND.n174 0.1
R794 GND.n182 GND.n178 0.1
R795 GND.n186 GND.n182 0.1
R796 GND.n190 GND.n186 0.1
R797 GND.n194 GND.n190 0.1
R798 GND.n198 GND.n194 0.1
R799 GND.n202 GND.n198 0.1
R800 GND.n206 GND.n202 0.1
R801 GND.n215 GND.n211 0.1
R802 GND.n219 GND.n215 0.1
R803 GND.n223 GND.n219 0.1
R804 GND.n536 GND.n532 0.1
R805 GND.n532 GND.n528 0.1
R806 GND.n523 GND.n519 0.1
R807 GND.n519 GND.n515 0.1
R808 GND.n515 GND.n511 0.1
R809 GND.n511 GND.n507 0.1
R810 GND.n507 GND.n503 0.1
R811 GND.n503 GND.n499 0.1
R812 GND.n499 GND.n495 0.1
R813 GND.n495 GND.n491 0.1
R814 GND.n325 GND.n302 0.075
R815 GND GND.n295 0.075
R816 GND.n347 GND.n346 0.075
R817 GND.n380 GND.n379 0.075
R818 GND.n390 EESPFAL_INV4_1/GND 0.075
R819 GND.n391 GND.n265 0.075
R820 GND.n437 GND.n244 0.075
R821 GND.n451 EESPFAL_XOR_v3_0/GND 0.075
R822 GND.n454 GND.n453 0.075
R823 GND.n39 GND.n35 0.075
R824 GND.n55 EESPFAL_3in_NOR_v2_0/GND 0.075
R825 GND.n64 GND.n63 0.075
R826 GND.n121 GND.n117 0.075
R827 GND.n137 EESPFAL_INV4_2/GND 0.075
R828 GND.n146 GND.n145 0.075
R829 GND.n211 GND.n207 0.075
R830 EESPFAL_4in_NAND_0/GND GND.n536 0.075
R831 GND.n528 GND.n524 0.075
R832 GND.n326 GND.n325 0.025
R833 GND.n337 GND 0.025
R834 GND.n348 GND.n347 0.025
R835 GND.n379 GND.n378 0.025
R836 EESPFAL_INV4_1/GND GND.n389 0.025
R837 GND.n400 GND.n265 0.025
R838 GND.n428 GND.n244 0.025
R839 GND.n441 EESPFAL_XOR_v3_0/GND 0.025
R840 GND.n453 GND.n234 0.025
R841 GND.n35 GND.n34 0.025
R842 GND.n48 EESPFAL_3in_NOR_v2_0/GND 0.025
R843 GND.n68 GND.n64 0.025
R844 GND.n117 GND.n116 0.025
R845 GND.n130 EESPFAL_INV4_2/GND 0.025
R846 GND.n150 GND.n146 0.025
R847 GND.n207 GND.n206 0.025
R848 EESPFAL_4in_NAND_0/GND GND.n223 0.025
R849 GND.n524 GND.n523 0.025
R850 x3.n0 x3.t0 1176.57
R851 x3.n0 x3.t2 1149.49
R852 EESPFAL_4in_NAND_0/A_bar x3.t1 1121.23
R853 x3 x3.n0 128
R854 EESPFAL_4in_NAND_0/A_bar x3 113.513
R855 CLK1.n26 CLK1.t43 44.338
R856 CLK1.n55 CLK1.t26 44.338
R857 CLK1.n171 CLK1.t5 44.338
R858 CLK1.n145 CLK1.t37 44.338
R859 CLK1.n369 CLK1.t48 44.337
R860 CLK1.n312 CLK1.t24 44.337
R861 CLK1.n171 CLK1.t1 44.337
R862 CLK1.n145 CLK1.t18 44.337
R863 CLK1.n253 CLK1.t36 44.337
R864 CLK1.n226 CLK1.t50 44.337
R865 CLK1.n0 CLK1.t15 39.4
R866 CLK1.n0 CLK1.t46 39.4
R867 CLK1.n207 CLK1.t52 39.4
R868 CLK1.n207 CLK1.t34 39.4
R869 CLK1.n95 CLK1.t3 39.4
R870 CLK1.n95 CLK1.t20 39.4
R871 CLK1.n94 CLK1.t4 39.4
R872 CLK1.n94 CLK1.t38 39.4
R873 CLK1.n7 CLK1.t41 39.4
R874 CLK1.n7 CLK1.t28 39.4
R875 CLK1.n77 CLK1.t10 31.775
R876 CLK1.n9 CLK1.t9 29.713
R877 CLK1.n72 CLK1.t22 29.713
R878 CLK1.n270 CLK1.t12 29.712
R879 CLK1.n209 CLK1.t13 29.712
R880 CLK1.n313 CLK1.t23 24.568
R881 CLK1.n370 CLK1.t47 24.568
R882 CLK1.n227 CLK1.t49 24.568
R883 CLK1.n249 CLK1.t35 24.568
R884 CLK1.n27 CLK1.t42 24.568
R885 CLK1.n51 CLK1.t25 24.568
R886 CLK1.n329 CLK1.t31 24
R887 CLK1.n329 CLK1.t16 24
R888 CLK1.n4 CLK1.t7 24
R889 CLK1.n4 CLK1.t8 24
R890 CLK1.n100 CLK1.t21 24
R891 CLK1.n100 CLK1.t32 24
R892 CLK1.n101 CLK1.t39 24
R893 CLK1.n101 CLK1.t44 24
R894 CLK1.n99 CLK1.t29 24
R895 CLK1.n99 CLK1.t6 24
R896 CLK1.n2 CLK1.t11 24
R897 CLK1.n2 CLK1.t30 24
R898 CLK1.n167 CLK1.t0 12.942
R899 CLK1.n146 CLK1.t17 12.942
R900 CLK1.n243 CLK1.n240 12.8
R901 CLK1.n45 CLK1.n42 12.8
R902 CLK1.n12 CLK1.n11 8.855
R903 CLK1.n16 CLK1.n15 8.855
R904 CLK1.n15 CLK1.n14 8.855
R905 CLK1.n20 CLK1.n19 8.855
R906 CLK1.n19 CLK1.n18 8.855
R907 CLK1.n24 CLK1.n23 8.855
R908 CLK1.n23 CLK1.n22 8.855
R909 CLK1.n29 CLK1.n28 8.855
R910 CLK1.n28 CLK1.n27 8.855
R911 CLK1.n33 CLK1.n32 8.855
R912 CLK1.n32 CLK1.n31 8.855
R913 CLK1.n37 CLK1.n36 8.855
R914 CLK1.n36 CLK1.n35 8.855
R915 CLK1.n42 CLK1.n41 8.855
R916 CLK1.n41 CLK1.n40 8.855
R917 CLK1.n45 CLK1.n44 8.855
R918 CLK1.n44 CLK1.n43 8.855
R919 CLK1.n49 CLK1.n48 8.855
R920 CLK1.n48 CLK1.n47 8.855
R921 CLK1.n53 CLK1.n52 8.855
R922 CLK1.n52 CLK1.n51 8.855
R923 CLK1.n58 CLK1.n57 8.855
R924 CLK1.n57 CLK1.n56 8.855
R925 CLK1.n62 CLK1.n61 8.855
R926 CLK1.n61 CLK1.n60 8.855
R927 CLK1.n66 CLK1.n65 8.855
R928 CLK1.n65 CLK1.n64 8.855
R929 CLK1.n70 CLK1.n69 8.855
R930 CLK1.n212 CLK1.n211 8.855
R931 CLK1.n216 CLK1.n215 8.855
R932 CLK1.n215 CLK1.n214 8.855
R933 CLK1.n220 CLK1.n219 8.855
R934 CLK1.n219 CLK1.n218 8.855
R935 CLK1.n224 CLK1.n223 8.855
R936 CLK1.n223 CLK1.n222 8.855
R937 CLK1.n229 CLK1.n228 8.855
R938 CLK1.n228 CLK1.n227 8.855
R939 CLK1.n233 CLK1.n232 8.855
R940 CLK1.n232 CLK1.n231 8.855
R941 CLK1.n237 CLK1.n236 8.855
R942 CLK1.n236 CLK1.n235 8.855
R943 CLK1.n240 CLK1.n206 8.855
R944 CLK1.n206 CLK1.n205 8.855
R945 CLK1.n243 CLK1.n242 8.855
R946 CLK1.n242 CLK1.n241 8.855
R947 CLK1.n247 CLK1.n246 8.855
R948 CLK1.n246 CLK1.n245 8.855
R949 CLK1.n251 CLK1.n250 8.855
R950 CLK1.n250 CLK1.n249 8.855
R951 CLK1.n256 CLK1.n255 8.855
R952 CLK1.n255 CLK1.n254 8.855
R953 CLK1.n260 CLK1.n259 8.855
R954 CLK1.n259 CLK1.n258 8.855
R955 CLK1.n264 CLK1.n263 8.855
R956 CLK1.n263 CLK1.n262 8.855
R957 CLK1.n268 CLK1.n267 8.855
R958 CLK1.n277 CLK1.n276 8.855
R959 CLK1.n281 CLK1.n280 8.855
R960 CLK1.n280 CLK1.n279 8.855
R961 CLK1.n285 CLK1.n284 8.855
R962 CLK1.n284 CLK1.n283 8.855
R963 CLK1.n290 CLK1.n289 8.855
R964 CLK1.n289 CLK1.n288 8.855
R965 CLK1.n294 CLK1.n293 8.855
R966 CLK1.n293 CLK1.n292 8.855
R967 CLK1.n298 CLK1.n297 8.855
R968 CLK1.n297 CLK1.n296 8.855
R969 CLK1.n302 CLK1.n301 8.855
R970 CLK1.n301 CLK1.n300 8.855
R971 CLK1.n306 CLK1.n305 8.855
R972 CLK1.n305 CLK1.n304 8.855
R973 CLK1.n310 CLK1.n309 8.855
R974 CLK1.n309 CLK1.n308 8.855
R975 CLK1.n315 CLK1.n314 8.855
R976 CLK1.n314 CLK1.n313 8.855
R977 CLK1.n319 CLK1.n318 8.855
R978 CLK1.n318 CLK1.n317 8.855
R979 CLK1.n323 CLK1.n322 8.855
R980 CLK1.n322 CLK1.n321 8.855
R981 CLK1.n327 CLK1.n326 8.855
R982 CLK1.n326 CLK1.n325 8.855
R983 CLK1.n380 CLK1.n379 8.855
R984 CLK1.n379 CLK1.n378 8.855
R985 CLK1.n376 CLK1.n375 8.855
R986 CLK1.n375 CLK1.n374 8.855
R987 CLK1.n372 CLK1.n371 8.855
R988 CLK1.n371 CLK1.n370 8.855
R989 CLK1.n367 CLK1.n366 8.855
R990 CLK1.n366 CLK1.n365 8.855
R991 CLK1.n363 CLK1.n362 8.855
R992 CLK1.n362 CLK1.n361 8.855
R993 CLK1.n359 CLK1.n358 8.855
R994 CLK1.n358 CLK1.n357 8.855
R995 CLK1.n355 CLK1.n354 8.855
R996 CLK1.n354 CLK1.n353 8.855
R997 CLK1.n351 CLK1.n350 8.855
R998 CLK1.n350 CLK1.n349 8.855
R999 CLK1.n347 CLK1.n346 8.855
R1000 CLK1.n346 CLK1.n345 8.855
R1001 CLK1.n342 CLK1.n341 8.855
R1002 CLK1.n341 CLK1.n340 8.855
R1003 CLK1.n338 CLK1.n337 8.855
R1004 CLK1.n337 CLK1.n336 8.855
R1005 CLK1.n334 CLK1.n333 8.855
R1006 CLK1.n321 CLK1.t14 8.189
R1007 CLK1.n378 CLK1.t45 8.189
R1008 CLK1.n235 CLK1.t51 8.189
R1009 CLK1.n241 CLK1.t33 8.189
R1010 CLK1.n35 CLK1.t40 8.189
R1011 CLK1.n43 CLK1.t27 8.189
R1012 CLK1.n110 CLK1.n101 7.776
R1013 CLK1.n128 CLK1.n99 7.776
R1014 CLK1.n344 CLK1.n329 6.776
R1015 CLK1.n119 CLK1.n100 6.776
R1016 CLK1.n201 CLK1.n3 6.754
R1017 CLK1.n328 CLK1.n0 4.938
R1018 CLK1.n239 CLK1.n207 4.938
R1019 CLK1.n158 CLK1.n94 4.938
R1020 CLK1.n158 CLK1.n95 4.938
R1021 CLK1.n39 CLK1.n7 4.938
R1022 CLK1.n9 CLK1.n8 4.662
R1023 CLK1.n209 CLK1.n208 4.662
R1024 CLK1.n74 CLK1.n73 4.65
R1025 CLK1.n13 CLK1.n12 4.65
R1026 CLK1.n17 CLK1.n16 4.65
R1027 CLK1.n21 CLK1.n20 4.65
R1028 CLK1.n25 CLK1.n24 4.65
R1029 CLK1.n30 CLK1.n29 4.65
R1030 CLK1.n34 CLK1.n33 4.65
R1031 CLK1.n38 CLK1.n37 4.65
R1032 CLK1.n42 CLK1.n39 4.65
R1033 CLK1.n46 CLK1.n45 4.65
R1034 CLK1.n50 CLK1.n49 4.65
R1035 CLK1.n54 CLK1.n53 4.65
R1036 CLK1.n59 CLK1.n58 4.65
R1037 CLK1.n63 CLK1.n62 4.65
R1038 CLK1.n67 CLK1.n66 4.65
R1039 CLK1.n71 CLK1.n70 4.65
R1040 CLK1.n198 CLK1.n6 4.65
R1041 CLK1.n204 CLK1.n1 4.65
R1042 CLK1.n203 CLK1.n202 4.65
R1043 CLK1.n213 CLK1.n212 4.65
R1044 CLK1.n217 CLK1.n216 4.65
R1045 CLK1.n221 CLK1.n220 4.65
R1046 CLK1.n225 CLK1.n224 4.65
R1047 CLK1.n230 CLK1.n229 4.65
R1048 CLK1.n234 CLK1.n233 4.65
R1049 CLK1.n238 CLK1.n237 4.65
R1050 CLK1.n240 CLK1.n239 4.65
R1051 CLK1.n244 CLK1.n243 4.65
R1052 CLK1.n248 CLK1.n247 4.65
R1053 CLK1.n252 CLK1.n251 4.65
R1054 CLK1.n257 CLK1.n256 4.65
R1055 CLK1.n261 CLK1.n260 4.65
R1056 CLK1.n265 CLK1.n264 4.65
R1057 CLK1.n269 CLK1.n268 4.65
R1058 CLK1.n272 CLK1.n271 4.65
R1059 CLK1.n274 CLK1.n273 4.65
R1060 CLK1.n278 CLK1.n277 4.65
R1061 CLK1.n282 CLK1.n281 4.65
R1062 CLK1.n286 CLK1.n285 4.65
R1063 CLK1.n291 CLK1.n290 4.65
R1064 CLK1.n295 CLK1.n294 4.65
R1065 CLK1.n299 CLK1.n298 4.65
R1066 CLK1.n303 CLK1.n302 4.65
R1067 CLK1.n307 CLK1.n306 4.65
R1068 CLK1.n311 CLK1.n310 4.65
R1069 CLK1.n316 CLK1.n315 4.65
R1070 CLK1.n320 CLK1.n319 4.65
R1071 CLK1.n324 CLK1.n323 4.65
R1072 CLK1.n328 CLK1.n327 4.65
R1073 CLK1.n381 CLK1.n380 4.65
R1074 CLK1.n377 CLK1.n376 4.65
R1075 CLK1.n373 CLK1.n372 4.65
R1076 CLK1.n368 CLK1.n367 4.65
R1077 CLK1.n364 CLK1.n363 4.65
R1078 CLK1.n360 CLK1.n359 4.65
R1079 CLK1.n356 CLK1.n355 4.65
R1080 CLK1.n352 CLK1.n351 4.65
R1081 CLK1.n348 CLK1.n347 4.65
R1082 CLK1.n343 CLK1.n342 4.65
R1083 CLK1.n339 CLK1.n338 4.65
R1084 CLK1.n335 CLK1.n334 4.65
R1085 CLK1.n157 CLK1.n154 4.633
R1086 CLK1.n154 CLK1.n98 4.633
R1087 CLK1.n80 CLK1.n79 4.427
R1088 CLK1.n84 CLK1.n83 4.427
R1089 CLK1.n83 CLK1.n82 4.427
R1090 CLK1.n88 CLK1.n87 4.427
R1091 CLK1.n87 CLK1.n86 4.427
R1092 CLK1.n92 CLK1.n91 4.427
R1093 CLK1.n91 CLK1.n90 4.427
R1094 CLK1.n194 CLK1.n193 4.427
R1095 CLK1.n193 CLK1.n192 4.427
R1096 CLK1.n190 CLK1.n189 4.427
R1097 CLK1.n189 CLK1.n188 4.427
R1098 CLK1.n186 CLK1.n185 4.427
R1099 CLK1.n185 CLK1.n184 4.427
R1100 CLK1.n182 CLK1.n181 4.427
R1101 CLK1.n181 CLK1.n180 4.427
R1102 CLK1.n178 CLK1.n177 4.427
R1103 CLK1.n174 CLK1.n173 4.427
R1104 CLK1.n169 CLK1.n168 4.427
R1105 CLK1.n165 CLK1.n164 4.427
R1106 CLK1.n161 CLK1.n160 4.427
R1107 CLK1.n157 CLK1.n156 4.427
R1108 CLK1.n154 CLK1.n153 4.427
R1109 CLK1.n98 CLK1.n97 4.427
R1110 CLK1.n148 CLK1.n147 4.427
R1111 CLK1.n143 CLK1.n142 4.427
R1112 CLK1.n139 CLK1.n138 4.427
R1113 CLK1.n135 CLK1.n134 4.427
R1114 CLK1.n134 CLK1.n133 4.427
R1115 CLK1.n131 CLK1.n130 4.427
R1116 CLK1.n130 CLK1.n129 4.427
R1117 CLK1.n126 CLK1.n125 4.427
R1118 CLK1.n125 CLK1.n124 4.427
R1119 CLK1.n122 CLK1.n121 4.427
R1120 CLK1.n121 CLK1.n120 4.427
R1121 CLK1.n117 CLK1.n116 4.427
R1122 CLK1.n116 CLK1.n115 4.427
R1123 CLK1.n113 CLK1.n112 4.427
R1124 CLK1.n112 CLK1.n111 4.427
R1125 CLK1.n108 CLK1.n107 4.427
R1126 CLK1.n107 CLK1.n106 4.427
R1127 CLK1.n104 CLK1.n103 4.427
R1128 CLK1.n177 CLK1.n176 4.427
R1129 CLK1.n173 CLK1.n172 4.427
R1130 CLK1.n168 CLK1.n167 4.427
R1131 CLK1.n164 CLK1.n163 4.427
R1132 CLK1.n160 CLK1.n159 4.427
R1133 CLK1.n156 CLK1.n155 4.427
R1134 CLK1.n153 CLK1.n152 4.427
R1135 CLK1.n97 CLK1.n96 4.427
R1136 CLK1.n147 CLK1.n146 4.427
R1137 CLK1.n142 CLK1.n141 4.427
R1138 CLK1.n138 CLK1.n137 4.427
R1139 CLK1.n159 CLK1.t2 4.314
R1140 CLK1.n152 CLK1.t19 4.314
R1141 CLK1.n6 CLK1.n5 3.715
R1142 CLK1.n200 CLK1.n199 3.039
R1143 CLK1.n331 CLK1.n330 3.038
R1144 CLK1.n201 CLK1.n200 2.849
R1145 CLK1.n5 CLK1.n4 2.57
R1146 CLK1.n3 CLK1.n2 2.57
R1147 CLK1.n81 CLK1.n80 2.325
R1148 CLK1.n85 CLK1.n84 2.325
R1149 CLK1.n89 CLK1.n88 2.325
R1150 CLK1.n93 CLK1.n92 2.325
R1151 CLK1.n195 CLK1.n194 2.325
R1152 CLK1.n191 CLK1.n190 2.325
R1153 CLK1.n187 CLK1.n186 2.325
R1154 CLK1.n183 CLK1.n182 2.325
R1155 CLK1.n179 CLK1.n178 2.325
R1156 CLK1.n175 CLK1.n174 2.325
R1157 CLK1.n170 CLK1.n169 2.325
R1158 CLK1.n166 CLK1.n165 2.325
R1159 CLK1.n162 CLK1.n161 2.325
R1160 CLK1.n158 CLK1.n157 2.325
R1161 CLK1.n154 CLK1.n151 2.325
R1162 CLK1.n149 CLK1.n148 2.325
R1163 CLK1.n144 CLK1.n143 2.325
R1164 CLK1.n140 CLK1.n139 2.325
R1165 CLK1.n136 CLK1.n135 2.325
R1166 CLK1.n132 CLK1.n131 2.325
R1167 CLK1.n127 CLK1.n126 2.325
R1168 CLK1.n123 CLK1.n122 2.325
R1169 CLK1.n118 CLK1.n117 2.325
R1170 CLK1.n114 CLK1.n113 2.325
R1171 CLK1.n109 CLK1.n108 2.325
R1172 CLK1.n76 CLK1.n75 2.325
R1173 CLK1.n197 CLK1.n196 2.203
R1174 CLK1.n287 CLK1.n204 2.203
R1175 CLK1.n211 CLK1.n210 1.655
R1176 CLK1.n276 CLK1.n275 1.655
R1177 CLK1.n11 CLK1.n10 1.655
R1178 CLK1.n69 CLK1.n68 1.655
R1179 CLK1.n267 CLK1.n266 1.655
R1180 CLK1.n333 CLK1.n332 1.655
R1181 CLK1.n105 CLK1.n104 1.156
R1182 CLK1.n331 CLK1 1.054
R1183 CLK1.n274 CLK1.n272 0.662
R1184 CLK1.n109 CLK1.n105 0.631
R1185 CLK1.n79 CLK1.n78 0.619
R1186 CLK1.n103 CLK1.n102 0.618
R1187 CLK1.n76 CLK1.n74 0.532
R1188 CLK1.n198 CLK1.n197 0.125
R1189 CLK1.n204 CLK1.n203 0.125
R1190 CLK1.n203 CLK1.n201 0.12
R1191 CLK1.n200 CLK1.n198 0.119
R1192 CLK1.n17 CLK1.n13 0.1
R1193 CLK1.n21 CLK1.n17 0.1
R1194 CLK1.n25 CLK1.n21 0.1
R1195 CLK1.n34 CLK1.n30 0.1
R1196 CLK1.n38 CLK1.n34 0.1
R1197 CLK1.n39 CLK1.n38 0.1
R1198 CLK1.n50 CLK1.n46 0.1
R1199 CLK1.n54 CLK1.n50 0.1
R1200 CLK1.n63 CLK1.n59 0.1
R1201 CLK1.n67 CLK1.n63 0.1
R1202 CLK1.n71 CLK1.n67 0.1
R1203 CLK1.n217 CLK1.n213 0.1
R1204 CLK1.n221 CLK1.n217 0.1
R1205 CLK1.n225 CLK1.n221 0.1
R1206 CLK1.n234 CLK1.n230 0.1
R1207 CLK1.n238 CLK1.n234 0.1
R1208 CLK1.n239 CLK1.n238 0.1
R1209 CLK1.n248 CLK1.n244 0.1
R1210 CLK1.n252 CLK1.n248 0.1
R1211 CLK1.n261 CLK1.n257 0.1
R1212 CLK1.n265 CLK1.n261 0.1
R1213 CLK1.n269 CLK1.n265 0.1
R1214 CLK1.n278 CLK1.n274 0.1
R1215 CLK1.n282 CLK1.n278 0.1
R1216 CLK1.n286 CLK1.n282 0.1
R1217 CLK1.n295 CLK1.n291 0.1
R1218 CLK1.n299 CLK1.n295 0.1
R1219 CLK1.n303 CLK1.n299 0.1
R1220 CLK1.n307 CLK1.n303 0.1
R1221 CLK1.n311 CLK1.n307 0.1
R1222 CLK1.n320 CLK1.n316 0.1
R1223 CLK1.n324 CLK1.n320 0.1
R1224 CLK1.n328 CLK1.n324 0.1
R1225 CLK1.n381 CLK1.n377 0.1
R1226 CLK1.n377 CLK1.n373 0.1
R1227 CLK1.n368 CLK1.n364 0.1
R1228 CLK1.n364 CLK1.n360 0.1
R1229 CLK1.n360 CLK1.n356 0.1
R1230 CLK1.n356 CLK1.n352 0.1
R1231 CLK1.n352 CLK1.n348 0.1
R1232 CLK1.n343 CLK1.n339 0.1
R1233 CLK1.n339 CLK1.n335 0.1
R1234 CLK1.n335 CLK1.n331 0.096
R1235 CLK1.n13 CLK1.n9 0.087
R1236 CLK1.n72 CLK1.n71 0.087
R1237 CLK1.n213 CLK1.n209 0.087
R1238 CLK1.n270 CLK1.n269 0.087
R1239 CLK1.n30 CLK1.n26 0.075
R1240 CLK1.n46 EESPFAL_INV4_0/CLK 0.075
R1241 CLK1.n55 CLK1.n54 0.075
R1242 CLK1.n230 CLK1.n226 0.075
R1243 CLK1.n244 CLK1 0.075
R1244 CLK1.n253 CLK1.n252 0.075
R1245 CLK1.n291 CLK1.n287 0.075
R1246 CLK1.n316 CLK1.n312 0.075
R1247 EESPFAL_XOR_v3_0/CLK CLK1.n381 0.075
R1248 CLK1.n373 CLK1.n369 0.075
R1249 CLK1.n348 CLK1.n344 0.075
R1250 CLK1.n85 CLK1.n81 0.041
R1251 CLK1.n89 CLK1.n85 0.041
R1252 CLK1.n93 CLK1.n89 0.041
R1253 CLK1.n195 CLK1.n191 0.041
R1254 CLK1.n191 CLK1.n187 0.041
R1255 CLK1.n187 CLK1.n183 0.041
R1256 CLK1.n183 CLK1.n179 0.041
R1257 CLK1.n179 CLK1.n175 0.041
R1258 CLK1.n170 CLK1.n166 0.041
R1259 CLK1.n166 CLK1.n162 0.041
R1260 CLK1.n162 CLK1.n158 0.041
R1261 CLK1.n151 CLK1.n150 0.041
R1262 CLK1.n150 CLK1.n149 0.041
R1263 CLK1.n144 CLK1.n140 0.041
R1264 CLK1.n140 CLK1.n136 0.041
R1265 CLK1.n136 CLK1.n132 0.041
R1266 CLK1.n127 CLK1.n123 0.041
R1267 CLK1.n118 CLK1.n114 0.041
R1268 CLK1.n132 CLK1.n128 0.036
R1269 CLK1.n196 CLK1.n195 0.031
R1270 CLK1.n171 CLK1.n170 0.031
R1271 CLK1.n151 EESPFAL_4in_NAND_0/CLK 0.031
R1272 CLK1.n149 CLK1.n145 0.031
R1273 CLK1.n123 CLK1.n119 0.031
R1274 CLK1.n26 CLK1.n25 0.025
R1275 CLK1.n39 EESPFAL_INV4_0/CLK 0.025
R1276 CLK1.n59 CLK1.n55 0.025
R1277 CLK1.n114 CLK1.n110 0.025
R1278 CLK1.n226 CLK1.n225 0.025
R1279 CLK1.n239 CLK1 0.025
R1280 CLK1.n257 CLK1.n253 0.025
R1281 CLK1.n287 CLK1.n286 0.025
R1282 CLK1.n312 CLK1.n311 0.025
R1283 EESPFAL_XOR_v3_0/CLK CLK1.n328 0.025
R1284 CLK1.n369 CLK1.n368 0.025
R1285 CLK1.n344 CLK1.n343 0.025
R1286 CLK1.n77 CLK1.n76 0.02
R1287 CLK1.n81 CLK1.n77 0.02
R1288 CLK1.n110 CLK1.n109 0.015
R1289 CLK1.n74 CLK1.n72 0.012
R1290 CLK1.n272 CLK1.n270 0.012
R1291 CLK1.n196 CLK1.n93 0.01
R1292 CLK1.n175 CLK1.n171 0.01
R1293 CLK1.n158 EESPFAL_4in_NAND_0/CLK 0.01
R1294 CLK1.n145 CLK1.n144 0.01
R1295 CLK1.n119 CLK1.n118 0.01
R1296 CLK1.n128 CLK1.n127 0.005
R1297 Dis1.n5 Dis1 563.2
R1298 Dis1.n2 EESPFAL_INV4_0/Dis 563.2
R1299 Dis1.n4 Dis1.t3 504.5
R1300 Dis1.n1 Dis1.t7 504.5
R1301 Dis1.n0 Dis1.t9 504.5
R1302 Dis1.n6 Dis1.t0 389.3
R1303 Dis1.n5 Dis1.t5 389.3
R1304 Dis1.n4 Dis1.t8 389.3
R1305 Dis1.n3 Dis1.t2 389.3
R1306 Dis1.n2 Dis1.t6 389.3
R1307 Dis1.n1 Dis1.t1 389.3
R1308 Dis1.n0 Dis1.t4 389.3
R1309 EESPFAL_4in_NAND_0/Dis Dis1.n8 290.754
R1310 Dis1.n7 EESPFAL_XOR_v3_0/Dis 137.537
R1311 Dis1.n8 EESPFAL_XOR_v3_1/Dis 137.536
R1312 Dis1.n6 Dis1.n5 115.2
R1313 Dis1.n3 Dis1.n2 115.2
R1314 Dis1.n7 Dis1 3.618
R1315 Dis1 Dis1.n4 3.2
R1316 EESPFAL_XOR_v3_0/Dis Dis1.n6 3.2
R1317 EESPFAL_INV4_0/Dis Dis1.n1 3.2
R1318 EESPFAL_XOR_v3_1/Dis Dis1.n3 3.2
R1319 EESPFAL_4in_NAND_0/Dis Dis1.n0 3.2
R1320 Dis1.n8 Dis1.n7 0.625
R1321 EESPFAL_NAND_v3_1/A.n0 EESPFAL_NAND_v3_1/A.t9 1071.62
R1322 EESPFAL_NAND_v3_1/A.t8 EESPFAL_NAND_v3_1/A.t6 819.4
R1323 EESPFAL_XOR_v3_0/OUT_bar EESPFAL_NAND_v3_1/A 526.587
R1324 EESPFAL_NAND_v3_1/A.n6 EESPFAL_NAND_v3_1/A.t7 506.1
R1325 EESPFAL_NAND_v3_1/A.n6 EESPFAL_NAND_v3_1/A.t8 313.3
R1326 EESPFAL_NAND_v3_1/A.n3 EESPFAL_NAND_v3_1/A.t1 273.936
R1327 EESPFAL_NAND_v3_1/A.n5 EESPFAL_NAND_v3_1/A.n1 128.334
R1328 EESPFAL_NAND_v3_1/A.n4 EESPFAL_NAND_v3_1/A.n3 105.6
R1329 EESPFAL_NAND_v3_1/A.n3 EESPFAL_NAND_v3_1/A.t0 81.939
R1330 EESPFAL_NAND_v3_1/A.n4 EESPFAL_NAND_v3_1/A.n2 57.937
R1331 EESPFAL_NAND_v3_1/A.n7 EESPFAL_NAND_v3_1/A.n5 57.6
R1332 EESPFAL_NAND_v3_1/A.n5 EESPFAL_NAND_v3_1/A.n4 41.6
R1333 EESPFAL_NAND_v3_1/A.n1 EESPFAL_NAND_v3_1/A.t3 39.4
R1334 EESPFAL_NAND_v3_1/A.n1 EESPFAL_NAND_v3_1/A.t4 39.4
R1335 EESPFAL_NAND_v3_1/A.n2 EESPFAL_NAND_v3_1/A.t5 24
R1336 EESPFAL_NAND_v3_1/A.n2 EESPFAL_NAND_v3_1/A.t2 24
R1337 EESPFAL_NAND_v3_1/A.n7 EESPFAL_NAND_v3_1/A.n6 8.764
R1338 EESPFAL_XOR_v3_0/OUT_bar EESPFAL_NAND_v3_1/A.n7 4.65
R1339 EESPFAL_NAND_v3_1/A.n0 EESPFAL_NAND_v3_1/A 3.2
R1340 EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/A.n0 2.37
R1341 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_3in_NOR_v2_0/A_bar 950.768
R1342 EESPFAL_NAND_v3_1/OUT_bar.t9 EESPFAL_NAND_v3_1/OUT_bar.t6 819.4
R1343 EESPFAL_3in_NOR_v2_0/A_bar EESPFAL_NAND_v3_1/OUT_bar.t8 684.833
R1344 EESPFAL_NAND_v3_1/OUT_bar.n5 EESPFAL_NAND_v3_1/OUT_bar.t7 506.1
R1345 EESPFAL_NAND_v3_1/OUT_bar.n5 EESPFAL_NAND_v3_1/OUT_bar.t9 313.3
R1346 EESPFAL_NAND_v3_1/OUT_bar.n1 EESPFAL_NAND_v3_1/OUT_bar.t2 177.936
R1347 EESPFAL_NAND_v3_1/OUT_bar.n4 EESPFAL_NAND_v3_1/OUT_bar.n0 128.334
R1348 EESPFAL_NAND_v3_1/OUT_bar.n3 EESPFAL_NAND_v3_1/OUT_bar.n1 105.6
R1349 EESPFAL_NAND_v3_1/OUT_bar.n1 EESPFAL_NAND_v3_1/OUT_bar.t1 81.937
R1350 EESPFAL_NAND_v3_1/OUT_bar.n3 EESPFAL_NAND_v3_1/OUT_bar.n2 58.267
R1351 EESPFAL_NAND_v3_1/OUT_bar.n6 EESPFAL_NAND_v3_1/OUT_bar.n4 57.6
R1352 EESPFAL_NAND_v3_1/OUT_bar.n4 EESPFAL_NAND_v3_1/OUT_bar.n3 41.6
R1353 EESPFAL_NAND_v3_1/OUT_bar.n0 EESPFAL_NAND_v3_1/OUT_bar.t4 39.4
R1354 EESPFAL_NAND_v3_1/OUT_bar.n0 EESPFAL_NAND_v3_1/OUT_bar.t3 39.4
R1355 EESPFAL_NAND_v3_1/OUT_bar.n2 EESPFAL_NAND_v3_1/OUT_bar.t5 24
R1356 EESPFAL_NAND_v3_1/OUT_bar.n2 EESPFAL_NAND_v3_1/OUT_bar.t0 24
R1357 EESPFAL_NAND_v3_1/OUT_bar.n6 EESPFAL_NAND_v3_1/OUT_bar.n5 8.764
R1358 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_1/OUT_bar.n6 4.65
R1359 CLK2.n132 CLK2.t18 44.338
R1360 CLK2.n103 CLK2.t10 44.338
R1361 CLK2.n241 CLK2.t31 44.337
R1362 CLK2.n194 CLK2.t22 44.337
R1363 CLK2.n34 CLK2.t4 44.337
R1364 CLK2.n63 CLK2.t14 44.337
R1365 CLK2.n0 CLK2.t20 39.4
R1366 CLK2.n0 CLK2.t29 39.4
R1367 CLK2.n6 CLK2.t16 39.4
R1368 CLK2.n6 CLK2.t8 39.4
R1369 CLK2.n15 CLK2.t12 39.4
R1370 CLK2.n15 CLK2.t6 39.4
R1371 CLK2.n17 CLK2.t0 29.712
R1372 CLK2.n10 CLK2.t24 29.712
R1373 CLK2.n195 CLK2.t21 24.568
R1374 CLK2.n242 CLK2.t30 24.568
R1375 CLK2.n128 CLK2.t17 24.568
R1376 CLK2.n104 CLK2.t9 24.568
R1377 CLK2.n59 CLK2.t13 24.568
R1378 CLK2.n35 CLK2.t3 24.568
R1379 CLK2.n216 CLK2.t23 24
R1380 CLK2.n216 CLK2.t27 24
R1381 CLK2.n161 CLK2.t25 24
R1382 CLK2.n7 CLK2.t1 24
R1383 CLK2.n7 CLK2.t26 24
R1384 CLK2.n1 CLK2.t2 24
R1385 CLK2.n118 CLK2.n115 12.8
R1386 CLK2.n49 CLK2.n46 12.8
R1387 CLK2.n155 CLK2.n154 8.855
R1388 CLK2.n13 CLK2.n12 8.855
R1389 CLK2.n74 CLK2.n73 8.855
R1390 CLK2.n73 CLK2.n72 8.855
R1391 CLK2.n70 CLK2.n69 8.855
R1392 CLK2.n69 CLK2.n68 8.855
R1393 CLK2.n66 CLK2.n65 8.855
R1394 CLK2.n65 CLK2.n64 8.855
R1395 CLK2.n61 CLK2.n60 8.855
R1396 CLK2.n60 CLK2.n59 8.855
R1397 CLK2.n57 CLK2.n56 8.855
R1398 CLK2.n56 CLK2.n55 8.855
R1399 CLK2.n53 CLK2.n52 8.855
R1400 CLK2.n52 CLK2.n51 8.855
R1401 CLK2.n49 CLK2.n48 8.855
R1402 CLK2.n48 CLK2.n47 8.855
R1403 CLK2.n46 CLK2.n45 8.855
R1404 CLK2.n45 CLK2.n44 8.855
R1405 CLK2.n41 CLK2.n40 8.855
R1406 CLK2.n40 CLK2.n39 8.855
R1407 CLK2.n37 CLK2.n36 8.855
R1408 CLK2.n36 CLK2.n35 8.855
R1409 CLK2.n32 CLK2.n31 8.855
R1410 CLK2.n31 CLK2.n30 8.855
R1411 CLK2.n28 CLK2.n27 8.855
R1412 CLK2.n27 CLK2.n26 8.855
R1413 CLK2.n24 CLK2.n23 8.855
R1414 CLK2.n23 CLK2.n22 8.855
R1415 CLK2.n20 CLK2.n19 8.855
R1416 CLK2.n151 CLK2.n150 8.855
R1417 CLK2.n150 CLK2.n149 8.855
R1418 CLK2.n147 CLK2.n146 8.855
R1419 CLK2.n146 CLK2.n145 8.855
R1420 CLK2.n143 CLK2.n142 8.855
R1421 CLK2.n142 CLK2.n141 8.855
R1422 CLK2.n139 CLK2.n138 8.855
R1423 CLK2.n138 CLK2.n137 8.855
R1424 CLK2.n135 CLK2.n134 8.855
R1425 CLK2.n134 CLK2.n133 8.855
R1426 CLK2.n130 CLK2.n129 8.855
R1427 CLK2.n129 CLK2.n128 8.855
R1428 CLK2.n126 CLK2.n125 8.855
R1429 CLK2.n125 CLK2.n124 8.855
R1430 CLK2.n122 CLK2.n121 8.855
R1431 CLK2.n121 CLK2.n120 8.855
R1432 CLK2.n118 CLK2.n117 8.855
R1433 CLK2.n117 CLK2.n116 8.855
R1434 CLK2.n115 CLK2.n114 8.855
R1435 CLK2.n114 CLK2.n113 8.855
R1436 CLK2.n110 CLK2.n109 8.855
R1437 CLK2.n109 CLK2.n108 8.855
R1438 CLK2.n106 CLK2.n105 8.855
R1439 CLK2.n105 CLK2.n104 8.855
R1440 CLK2.n101 CLK2.n100 8.855
R1441 CLK2.n100 CLK2.n99 8.855
R1442 CLK2.n97 CLK2.n96 8.855
R1443 CLK2.n96 CLK2.n95 8.855
R1444 CLK2.n93 CLK2.n92 8.855
R1445 CLK2.n92 CLK2.n91 8.855
R1446 CLK2.n89 CLK2.n88 8.855
R1447 CLK2.n88 CLK2.n87 8.855
R1448 CLK2.n84 CLK2.n83 8.855
R1449 CLK2.n83 CLK2.n82 8.855
R1450 CLK2.n80 CLK2.n79 8.855
R1451 CLK2.n172 CLK2.n171 8.855
R1452 CLK2.n176 CLK2.n175 8.855
R1453 CLK2.n175 CLK2.n174 8.855
R1454 CLK2.n180 CLK2.n179 8.855
R1455 CLK2.n179 CLK2.n178 8.855
R1456 CLK2.n184 CLK2.n183 8.855
R1457 CLK2.n183 CLK2.n182 8.855
R1458 CLK2.n188 CLK2.n187 8.855
R1459 CLK2.n187 CLK2.n186 8.855
R1460 CLK2.n192 CLK2.n191 8.855
R1461 CLK2.n191 CLK2.n190 8.855
R1462 CLK2.n197 CLK2.n196 8.855
R1463 CLK2.n196 CLK2.n195 8.855
R1464 CLK2.n201 CLK2.n200 8.855
R1465 CLK2.n200 CLK2.n199 8.855
R1466 CLK2.n205 CLK2.n204 8.855
R1467 CLK2.n204 CLK2.n203 8.855
R1468 CLK2.n209 CLK2.n208 8.855
R1469 CLK2.n208 CLK2.n207 8.855
R1470 CLK2.n252 CLK2.n251 8.855
R1471 CLK2.n251 CLK2.n250 8.855
R1472 CLK2.n248 CLK2.n247 8.855
R1473 CLK2.n247 CLK2.n246 8.855
R1474 CLK2.n244 CLK2.n243 8.855
R1475 CLK2.n243 CLK2.n242 8.855
R1476 CLK2.n239 CLK2.n238 8.855
R1477 CLK2.n238 CLK2.n237 8.855
R1478 CLK2.n235 CLK2.n234 8.855
R1479 CLK2.n234 CLK2.n233 8.855
R1480 CLK2.n231 CLK2.n230 8.855
R1481 CLK2.n230 CLK2.n229 8.855
R1482 CLK2.n215 CLK2.n214 8.855
R1483 CLK2.n214 CLK2.n213 8.855
R1484 CLK2.n223 CLK2.n222 8.855
R1485 CLK2.n222 CLK2.n221 8.855
R1486 CLK2.n219 CLK2.n218 8.855
R1487 CLK2.n167 CLK2.n2 8.365
R1488 CLK2.n203 CLK2.t19 8.189
R1489 CLK2.n250 CLK2.t28 8.189
R1490 CLK2.n120 CLK2.t15 8.189
R1491 CLK2.n113 CLK2.t7 8.189
R1492 CLK2.n51 CLK2.t11 8.189
R1493 CLK2.n44 CLK2.t5 8.189
R1494 CLK2.n225 CLK2.n216 6.776
R1495 CLK2.n86 CLK2.n7 6.776
R1496 CLK2.n163 CLK2.n162 6.754
R1497 CLK2.n210 CLK2.n0 4.938
R1498 CLK2.n119 CLK2.n6 4.938
R1499 CLK2.n50 CLK2.n15 4.938
R1500 CLK2.n157 CLK2.n5 4.675
R1501 CLK2.n169 CLK2.n168 4.675
R1502 CLK2.n10 CLK2.n9 4.662
R1503 CLK2.n17 CLK2.n16 4.662
R1504 CLK2.n14 CLK2.n13 4.65
R1505 CLK2.n75 CLK2.n74 4.65
R1506 CLK2.n71 CLK2.n70 4.65
R1507 CLK2.n67 CLK2.n66 4.65
R1508 CLK2.n62 CLK2.n61 4.65
R1509 CLK2.n58 CLK2.n57 4.65
R1510 CLK2.n54 CLK2.n53 4.65
R1511 CLK2.n50 CLK2.n49 4.65
R1512 CLK2.n46 CLK2.n43 4.65
R1513 CLK2.n42 CLK2.n41 4.65
R1514 CLK2.n38 CLK2.n37 4.65
R1515 CLK2.n33 CLK2.n32 4.65
R1516 CLK2.n29 CLK2.n28 4.65
R1517 CLK2.n25 CLK2.n24 4.65
R1518 CLK2.n21 CLK2.n20 4.65
R1519 CLK2.n77 CLK2.n8 4.65
R1520 CLK2.n156 CLK2.n155 4.65
R1521 CLK2.n152 CLK2.n151 4.65
R1522 CLK2.n148 CLK2.n147 4.65
R1523 CLK2.n144 CLK2.n143 4.65
R1524 CLK2.n140 CLK2.n139 4.65
R1525 CLK2.n136 CLK2.n135 4.65
R1526 CLK2.n131 CLK2.n130 4.65
R1527 CLK2.n127 CLK2.n126 4.65
R1528 CLK2.n123 CLK2.n122 4.65
R1529 CLK2.n119 CLK2.n118 4.65
R1530 CLK2.n115 CLK2.n112 4.65
R1531 CLK2.n111 CLK2.n110 4.65
R1532 CLK2.n107 CLK2.n106 4.65
R1533 CLK2.n102 CLK2.n101 4.65
R1534 CLK2.n98 CLK2.n97 4.65
R1535 CLK2.n94 CLK2.n93 4.65
R1536 CLK2.n90 CLK2.n89 4.65
R1537 CLK2.n85 CLK2.n84 4.65
R1538 CLK2.n81 CLK2.n80 4.65
R1539 CLK2.n160 CLK2.n4 4.65
R1540 CLK2.n159 CLK2.n158 4.65
R1541 CLK2.n166 CLK2.n165 4.65
R1542 CLK2.n173 CLK2.n172 4.65
R1543 CLK2.n177 CLK2.n176 4.65
R1544 CLK2.n181 CLK2.n180 4.65
R1545 CLK2.n185 CLK2.n184 4.65
R1546 CLK2.n189 CLK2.n188 4.65
R1547 CLK2.n193 CLK2.n192 4.65
R1548 CLK2.n198 CLK2.n197 4.65
R1549 CLK2.n202 CLK2.n201 4.65
R1550 CLK2.n206 CLK2.n205 4.65
R1551 CLK2.n210 CLK2.n209 4.65
R1552 CLK2.n253 CLK2.n252 4.65
R1553 CLK2.n249 CLK2.n248 4.65
R1554 CLK2.n245 CLK2.n244 4.65
R1555 CLK2.n240 CLK2.n239 4.65
R1556 CLK2.n236 CLK2.n235 4.65
R1557 CLK2.n232 CLK2.n231 4.65
R1558 CLK2.n224 CLK2.n223 4.65
R1559 CLK2.n164 CLK2.n3 3.039
R1560 CLK2.n227 CLK2.n215 3.033
R1561 CLK2.n220 CLK2.n219 2.682
R1562 CLK2.n162 CLK2.n161 2.57
R1563 CLK2.n2 CLK2.n1 2.57
R1564 CLK2.n164 CLK2.n163 2.224
R1565 CLK2.n159 CLK2.n157 2.203
R1566 CLK2.n169 CLK2.n167 2.203
R1567 CLK2.n171 CLK2.n170 1.655
R1568 CLK2.n154 CLK2.n153 1.655
R1569 CLK2.n12 CLK2.n11 1.655
R1570 CLK2.n19 CLK2.n18 1.655
R1571 CLK2.n79 CLK2.n78 1.655
R1572 CLK2.n218 CLK2.n217 1.655
R1573 CLK2.n228 CLK2.n212 1.495
R1574 CLK2.n224 CLK2.n220 1.095
R1575 CLK2.n77 CLK2.n76 1.047
R1576 CLK2.n211 CLK2 0.282
R1577 CLK2.n160 CLK2.n159 0.125
R1578 CLK2.n167 CLK2.n166 0.125
R1579 CLK2.n166 CLK2.n164 0.12
R1580 CLK2.n163 CLK2.n160 0.119
R1581 CLK2.n75 CLK2.n71 0.1
R1582 CLK2.n71 CLK2.n67 0.1
R1583 CLK2.n62 CLK2.n58 0.1
R1584 CLK2.n58 CLK2.n54 0.1
R1585 CLK2.n54 CLK2.n50 0.1
R1586 CLK2.n43 CLK2.n42 0.1
R1587 CLK2.n42 CLK2.n38 0.1
R1588 CLK2.n33 CLK2.n29 0.1
R1589 CLK2.n29 CLK2.n25 0.1
R1590 CLK2.n25 CLK2.n21 0.1
R1591 CLK2.n156 CLK2.n152 0.1
R1592 CLK2.n152 CLK2.n148 0.1
R1593 CLK2.n148 CLK2.n144 0.1
R1594 CLK2.n144 CLK2.n140 0.1
R1595 CLK2.n140 CLK2.n136 0.1
R1596 CLK2.n131 CLK2.n127 0.1
R1597 CLK2.n127 CLK2.n123 0.1
R1598 CLK2.n123 CLK2.n119 0.1
R1599 CLK2.n112 CLK2.n111 0.1
R1600 CLK2.n111 CLK2.n107 0.1
R1601 CLK2.n102 CLK2.n98 0.1
R1602 CLK2.n98 CLK2.n94 0.1
R1603 CLK2.n94 CLK2.n90 0.1
R1604 CLK2.n85 CLK2.n81 0.1
R1605 CLK2.n81 CLK2.n77 0.1
R1606 CLK2.n177 CLK2.n173 0.1
R1607 CLK2.n181 CLK2.n177 0.1
R1608 CLK2.n185 CLK2.n181 0.1
R1609 CLK2.n189 CLK2.n185 0.1
R1610 CLK2.n193 CLK2.n189 0.1
R1611 CLK2.n202 CLK2.n198 0.1
R1612 CLK2.n206 CLK2.n202 0.1
R1613 CLK2.n210 CLK2.n206 0.1
R1614 CLK2.n253 CLK2.n249 0.1
R1615 CLK2.n249 CLK2.n245 0.1
R1616 CLK2.n240 CLK2.n236 0.1
R1617 CLK2.n236 CLK2.n232 0.1
R1618 CLK2.n232 CLK2.n228 0.091
R1619 CLK2.n14 CLK2.n10 0.087
R1620 CLK2.n21 CLK2.n17 0.087
R1621 CLK2.n90 CLK2.n86 0.087
R1622 CLK2.n76 CLK2.n14 0.075
R1623 CLK2.n63 CLK2.n62 0.075
R1624 CLK2.n43 EESPFAL_INV4_2/CLK 0.075
R1625 CLK2.n38 CLK2.n34 0.075
R1626 CLK2.n157 CLK2.n156 0.075
R1627 CLK2.n132 CLK2.n131 0.075
R1628 CLK2.n112 EESPFAL_NAND_v3_0/CLK 0.075
R1629 CLK2.n107 CLK2.n103 0.075
R1630 CLK2.n173 CLK2.n169 0.075
R1631 CLK2.n198 CLK2.n194 0.075
R1632 CLK2 CLK2.n253 0.075
R1633 CLK2.n245 CLK2.n241 0.075
R1634 CLK2.n226 CLK2.n225 0.06
R1635 CLK2.n227 CLK2.n226 0.027
R1636 CLK2.n76 CLK2.n75 0.025
R1637 CLK2.n67 CLK2.n63 0.025
R1638 CLK2.n50 EESPFAL_INV4_2/CLK 0.025
R1639 CLK2.n34 CLK2.n33 0.025
R1640 CLK2.n136 CLK2.n132 0.025
R1641 CLK2.n119 EESPFAL_NAND_v3_0/CLK 0.025
R1642 CLK2.n103 CLK2.n102 0.025
R1643 CLK2.n194 CLK2.n193 0.025
R1644 CLK2 CLK2.n210 0.025
R1645 CLK2.n241 CLK2.n240 0.025
R1646 CLK2.n212 CLK2.n211 0.017
R1647 CLK2.n86 CLK2.n85 0.012
R1648 CLK2.n225 CLK2.n224 0.012
R1649 CLK2.n228 CLK2.n227 0.009
R1650 EESPFAL_NAND_v3_1/A_bar.t9 EESPFAL_NAND_v3_1/A_bar.t6 819.4
R1651 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/A_bar.t8 736.033
R1652 EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_NAND_v3_1/A_bar.t9 514.133
R1653 EESPFAL_NAND_v3_1/A_bar.n1 EESPFAL_NAND_v3_1/A_bar.t7 305.266
R1654 EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_NAND_v3_1/A_bar.n5 192
R1655 EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_NAND_v3_1/A_bar.n3 166.735
R1656 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/A_bar.n6 161.207
R1657 EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_NAND_v3_1/A_bar.n4 105.6
R1658 EESPFAL_NAND_v3_1/A_bar.n5 EESPFAL_NAND_v3_1/A_bar.t3 97.937
R1659 EESPFAL_NAND_v3_1/A_bar.n6 EESPFAL_NAND_v3_1/A_bar.t4 97.937
R1660 EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_NAND_v3_1/A_bar.n1 76
R1661 EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_NAND_v3_1/A_bar.n0 73.937
R1662 EESPFAL_NAND_v3_1/A_bar.n4 EESPFAL_NAND_v3_1/A_bar.n2 57.6
R1663 EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_NAND_v3_1/A_bar.t2 39.4
R1664 EESPFAL_NAND_v3_1/A_bar.n3 EESPFAL_NAND_v3_1/A_bar.t1 39.4
R1665 EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_NAND_v3_1/A_bar.t5 24
R1666 EESPFAL_NAND_v3_1/A_bar.n0 EESPFAL_NAND_v3_1/A_bar.t0 24
R1667 EESPFAL_NAND_v3_1/A_bar.n2 EESPFAL_XOR_v3_0/OUT 3.2
R1668 x1.n0 x1.t2 1176.57
R1669 x1.n0 x1.t0 1149.49
R1670 EESPFAL_4in_NAND_0/B x1.t3 446.232
R1671 x1 x1.t1 392.5
R1672 x1.n2 EESPFAL_4in_NAND_0/B 255.704
R1673 EESPFAL_XOR_v3_1/A x1.n2 254.89
R1674 x1.n1 x1 197.717
R1675 EESPFAL_XOR_v3_1/A x1.n0 128
R1676 x1.n2 x1.n1 2.168
R1677 x1.n1 x1 1.059
R1678 x1_bar.n0 x1_bar.t0 1069.04
R1679 x1_bar.n0 x1_bar.t2 1015.9
R1680 EESPFAL_4in_NAND_0/B_bar x1_bar.t1 912.566
R1681 x1_bar x1_bar.t3 778.1
R1682 x1_bar.n1 EESPFAL_4in_NAND_0/B_bar 220.027
R1683 EESPFAL_XOR_v3_1/A_bar x1_bar.n1 218.41
R1684 EESPFAL_XOR_v3_1/A_bar x1_bar.n0 89.6
R1685 x1_bar.n1 x1_bar 2.954
R1686 s2_bar.t6 s2_bar.t7 819.4
R1687 s2_bar.n4 s2_bar.t5 506.1
R1688 s2_bar.n4 s2_bar.t6 313.3
R1689 s2_bar.n2 s2_bar.t2 181.136
R1690 s2_bar.n3 s2_bar.n0 128.334
R1691 s2_bar.n2 s2_bar.n1 57.937
R1692 s2_bar.n5 s2_bar.n3 57.6
R1693 s2_bar.n3 s2_bar.n2 41.6
R1694 s2_bar.n0 s2_bar.t0 39.4
R1695 s2_bar.n0 s2_bar.t4 39.4
R1696 s2_bar.n1 s2_bar.t1 24
R1697 s2_bar.n1 s2_bar.t3 24
R1698 s2_bar.n5 s2_bar.n4 8.764
R1699 s2_bar s2_bar.n5 4.681
R1700 s2.t9 s2.t8 819.4
R1701 s2.n0 s2.t9 514.133
R1702 s2.n0 s2.t7 305.266
R1703 s2.n6 s2.n1 166.734
R1704 s2.n6 s2.n5 105.6
R1705 s2.n5 s2.t0 97.937
R1706 s2.n5 s2.n4 96
R1707 s2.n4 s2 83.813
R1708 s2 s2.n0 79.2
R1709 s2.n6 s2.n2 73.937
R1710 s2.n4 s2.n3 73.937
R1711 s2 s2.n6 54.4
R1712 s2.n1 s2.t3 39.4
R1713 s2.n1 s2.t4 39.4
R1714 s2.n2 s2.t5 24
R1715 s2.n2 s2.t2 24
R1716 s2.n3 s2.t1 24
R1717 s2.n3 s2.t6 24
R1718 x2.n0 x2.t2 800.452
R1719 x2.n0 x2.t3 787.997
R1720 EESPFAL_4in_NAND_0/D x2.t0 444.545
R1721 EESPFAL_INV4_0/A_bar x2.t1 392.5
R1722 EESPFAL_INV4_0/A_bar x2.n2 196.579
R1723 x2.n2 EESPFAL_4in_NAND_0/D 184.29
R1724 x2.n1 x2 181.93
R1725 x2 x2.n0 169.6
R1726 x2.n2 x2.n1 1.796
R1727 x2.n1 x2 0.26
R1728 x2_bar.n0 x2_bar.t1 810.772
R1729 EESPFAL_INV4_0/A x2_bar.t3 778.1
R1730 x2_bar.n0 x2_bar.t2 694.566
R1731 EESPFAL_4in_NAND_0/D_bar x2_bar.t0 495.233
R1732 x2_bar.n2 EESPFAL_4in_NAND_0/D_bar 147.293
R1733 x2_bar.n1 x2_bar 145.45
R1734 EESPFAL_INV4_0/A x2_bar.n2 41.057
R1735 x2_bar x2_bar.n0 25.6
R1736 x2_bar.n2 x2_bar.n1 2.782
R1737 x2_bar.n1 x2_bar 0.321
R1738 CLK3.n94 CLK3.t4 44.337
R1739 CLK3.n35 CLK3.t10 44.337
R1740 CLK3.n0 CLK3.t8 39.4
R1741 CLK3.n0 CLK3.t6 39.4
R1742 CLK3.n56 CLK3.t11 30.775
R1743 CLK3.n2 CLK3.t2 30.775
R1744 CLK3.n36 CLK3.t9 24.568
R1745 CLK3.n95 CLK3.t3 24.568
R1746 CLK3.n52 CLK3.t0 24
R1747 CLK3.n52 CLK3.t1 24
R1748 CLK3.n54 CLK3 9.095
R1749 CLK3.n5 CLK3.n4 8.855
R1750 CLK3.n9 CLK3.n8 8.855
R1751 CLK3.n8 CLK3.n7 8.855
R1752 CLK3.n13 CLK3.n12 8.855
R1753 CLK3.n12 CLK3.n11 8.855
R1754 CLK3.n17 CLK3.n16 8.855
R1755 CLK3.n16 CLK3.n15 8.855
R1756 CLK3.n21 CLK3.n20 8.855
R1757 CLK3.n20 CLK3.n19 8.855
R1758 CLK3.n25 CLK3.n24 8.855
R1759 CLK3.n24 CLK3.n23 8.855
R1760 CLK3.n29 CLK3.n28 8.855
R1761 CLK3.n28 CLK3.n27 8.855
R1762 CLK3.n33 CLK3.n32 8.855
R1763 CLK3.n32 CLK3.n31 8.855
R1764 CLK3.n38 CLK3.n37 8.855
R1765 CLK3.n37 CLK3.n36 8.855
R1766 CLK3.n42 CLK3.n41 8.855
R1767 CLK3.n41 CLK3.n40 8.855
R1768 CLK3.n46 CLK3.n45 8.855
R1769 CLK3.n45 CLK3.n44 8.855
R1770 CLK3.n50 CLK3.n49 8.855
R1771 CLK3.n49 CLK3.n48 8.855
R1772 CLK3.n105 CLK3.n104 8.855
R1773 CLK3.n104 CLK3.n103 8.855
R1774 CLK3.n101 CLK3.n100 8.855
R1775 CLK3.n100 CLK3.n99 8.855
R1776 CLK3.n97 CLK3.n96 8.855
R1777 CLK3.n96 CLK3.n95 8.855
R1778 CLK3.n92 CLK3.n91 8.855
R1779 CLK3.n91 CLK3.n90 8.855
R1780 CLK3.n88 CLK3.n87 8.855
R1781 CLK3.n87 CLK3.n86 8.855
R1782 CLK3.n84 CLK3.n83 8.855
R1783 CLK3.n83 CLK3.n82 8.855
R1784 CLK3.n80 CLK3.n79 8.855
R1785 CLK3.n79 CLK3.n78 8.855
R1786 CLK3.n75 CLK3.n74 8.855
R1787 CLK3.n74 CLK3.n73 8.855
R1788 CLK3.n71 CLK3.n70 8.855
R1789 CLK3.n70 CLK3.n69 8.855
R1790 CLK3.n67 CLK3.n66 8.855
R1791 CLK3.n66 CLK3.n65 8.855
R1792 CLK3.n62 CLK3.n61 8.855
R1793 CLK3.n44 CLK3.t7 8.189
R1794 CLK3.n103 CLK3.t5 8.189
R1795 CLK3.n77 CLK3.n52 6.776
R1796 CLK3.n51 CLK3.n0 4.938
R1797 CLK3.n56 CLK3.n55 4.687
R1798 CLK3.n2 CLK3.n1 4.687
R1799 CLK3.n6 CLK3.n5 4.65
R1800 CLK3.n10 CLK3.n9 4.65
R1801 CLK3.n14 CLK3.n13 4.65
R1802 CLK3.n18 CLK3.n17 4.65
R1803 CLK3.n22 CLK3.n21 4.65
R1804 CLK3.n26 CLK3.n25 4.65
R1805 CLK3.n30 CLK3.n29 4.65
R1806 CLK3.n34 CLK3.n33 4.65
R1807 CLK3.n39 CLK3.n38 4.65
R1808 CLK3.n43 CLK3.n42 4.65
R1809 CLK3.n47 CLK3.n46 4.65
R1810 CLK3.n51 CLK3.n50 4.65
R1811 CLK3.n106 CLK3.n105 4.65
R1812 CLK3.n102 CLK3.n101 4.65
R1813 CLK3.n98 CLK3.n97 4.65
R1814 CLK3.n93 CLK3.n92 4.65
R1815 CLK3.n89 CLK3.n88 4.65
R1816 CLK3.n85 CLK3.n84 4.65
R1817 CLK3.n81 CLK3.n80 4.65
R1818 CLK3.n76 CLK3.n75 4.65
R1819 CLK3.n72 CLK3.n71 4.65
R1820 CLK3.n68 CLK3.n67 4.65
R1821 CLK3.n63 CLK3.n62 3.033
R1822 CLK3.n58 CLK3.n54 2.251
R1823 CLK3.n59 CLK3.n53 2.249
R1824 CLK3.n4 CLK3.n3 1.655
R1825 CLK3.n61 CLK3.n60 1.655
R1826 CLK3.n10 CLK3.n6 0.1
R1827 CLK3.n14 CLK3.n10 0.1
R1828 CLK3.n18 CLK3.n14 0.1
R1829 CLK3.n22 CLK3.n18 0.1
R1830 CLK3.n26 CLK3.n22 0.1
R1831 CLK3.n30 CLK3.n26 0.1
R1832 CLK3.n34 CLK3.n30 0.1
R1833 CLK3.n43 CLK3.n39 0.1
R1834 CLK3.n47 CLK3.n43 0.1
R1835 CLK3.n51 CLK3.n47 0.1
R1836 CLK3.n106 CLK3.n102 0.1
R1837 CLK3.n102 CLK3.n98 0.1
R1838 CLK3.n93 CLK3.n89 0.1
R1839 CLK3.n89 CLK3.n85 0.1
R1840 CLK3.n85 CLK3.n81 0.1
R1841 CLK3.n76 CLK3.n72 0.1
R1842 CLK3.n72 CLK3.n68 0.1
R1843 CLK3.n81 CLK3.n77 0.087
R1844 CLK3.n68 CLK3.n64 0.076
R1845 CLK3.n39 CLK3.n35 0.075
R1846 CLK3 CLK3.n106 0.075
R1847 CLK3.n98 CLK3.n94 0.075
R1848 CLK3.n6 CLK3.n2 0.062
R1849 CLK3.n57 CLK3.n56 0.032
R1850 CLK3.n35 CLK3.n34 0.025
R1851 CLK3 CLK3.n51 0.025
R1852 CLK3.n94 CLK3.n93 0.025
R1853 CLK3.n58 CLK3.n57 0.025
R1854 CLK3.n64 CLK3.n63 0.023
R1855 CLK3.n77 CLK3.n76 0.012
R1856 CLK3.n59 CLK3.n58 0.003
R1857 CLK3.n63 CLK3.n59 0.003
R1858 x0_bar.n0 x0_bar.t1 810.772
R1859 x0_bar x0_bar.t2 703.9
R1860 x0_bar.n0 x0_bar.t0 694.566
R1861 x0_bar x0_bar.n1 293.496
R1862 x0_bar.n1 EESPFAL_XOR_v3_1/B_bar 291.37
R1863 EESPFAL_XOR_v3_1/B_bar x0_bar.n0 25.6
R1864 x0_bar.n1 x0_bar 2.601
R1865 Dis2.n1 Dis2.t4 504.5
R1866 Dis2.n0 Dis2.t2 504.5
R1867 Dis2.n4 Dis2.n3 408.185
R1868 Dis2.n1 Dis2.t1 389.3
R1869 Dis2.n0 Dis2.t3 389.3
R1870 Dis2.n4 Dis2.t5 389.3
R1871 Dis2.n5 Dis2.t0 389.3
R1872 Dis2.n2 Dis2 177.217
R1873 Dis2.n3 EESPFAL_NAND_v3_0/Dis 177.216
R1874 Dis2.n5 Dis2.n4 115.2
R1875 Dis2.n2 Dis2 3.612
R1876 Dis2 Dis2.n1 3.2
R1877 EESPFAL_NAND_v3_0/Dis Dis2.n0 3.2
R1878 EESPFAL_INV4_2/Dis Dis2.n5 3.2
R1879 Dis2.n3 Dis2.n2 0.625
R1880 x3_bar.n0 x3_bar.t0 1069.04
R1881 x3_bar.n0 x3_bar.t2 1015.9
R1882 EESPFAL_4in_NAND_0/A x3_bar.t1 447.076
R1883 x3_bar x3_bar.n0 89.6
R1884 EESPFAL_4in_NAND_0/A x3_bar 76.188
R1885 Dis3 Dis3.t1 392.5
R1886 Dis3.n0 Dis3.t0 389.3
R1887 Dis3.n0 Dis3 297.159
R1888 Dis3 Dis3.n0 112
R1889 x0.n0 x0.t0 800.452
R1890 x0.n0 x0.t1 787.997
R1891 x0 x0.t2 445.388
R1892 x0 x0.n1 329.196
R1893 x0.n1 EESPFAL_XOR_v3_1/B 327.85
R1894 EESPFAL_XOR_v3_1/B x0.n0 169.6
R1895 x0.n1 x0 2.882
C0 EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_0/B_bar 0.00fF
C1 Dis2 EESPFAL_NAND_v3_1/A_bar 0.01fF
C2 EESPFAL_NAND_v3_0/A x0_bar 0.08fF
C3 EESPFAL_INV4_2/A EESPFAL_3in_NOR_v2_0/B 0.00fF
C4 a_385_n466# x3_bar 0.00fF
C5 x0 a_85_214# 0.00fF
C6 x0 CLK1 0.95fF
C7 a_1945_214# EESPFAL_NAND_v3_1/B 0.00fF
C8 x1_bar Dis3 0.01fF
C9 EESPFAL_NAND_v3_0/A a_385_n466# 0.00fF
C10 Dis1 EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C11 a_85_214# EESPFAL_NAND_v3_0/A_bar 0.00fF
C12 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/B 1.00fF
C13 EESPFAL_NAND_v3_0/A_bar CLK1 1.92fF
C14 x2_bar EESPFAL_3in_NOR_v2_0/B_bar 0.01fF
C15 x1_bar a_1645_214# 0.00fF
C16 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/B 0.34fF
C17 Dis2 EESPFAL_3in_NOR_v2_0/B 0.10fF
C18 x1_bar EESPFAL_NAND_v3_1/B_bar 0.33fF
C19 x3 EESPFAL_NAND_v3_1/A_bar 0.04fF
C20 Dis3 EESPFAL_NAND_v3_0/B_bar 0.04fF
C21 x1_bar EESPFAL_NAND_v3_1/OUT 0.00fF
C22 s2_bar EESPFAL_NAND_v3_0/B_bar 0.00fF
C23 EESPFAL_NAND_v3_0/A_bar EESPFAL_3in_NOR_v2_0/B_bar 0.07fF
C24 EESPFAL_INV4_2/A Dis1 0.11fF
C25 a_5735_n466# CLK2 0.02fF
C26 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_1/B_bar 0.02fF
C27 EESPFAL_3in_NOR_v2_0/B EESPFAL_NAND_v3_1/B 0.02fF
C28 CLK1 CLK3 0.02fF
C29 x0 x2_bar 0.13fF
C30 EESPFAL_NAND_v3_0/A_bar x2_bar 0.24fF
C31 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_1/OUT_bar 0.02fF
C32 a_385_214# CLK1 0.01fF
C33 x1 x1_bar 5.84fF
C34 Dis2 Dis1 0.03fF
C35 EESPFAL_3in_NOR_v2_0/B_bar CLK3 0.58fF
C36 a_1945_n466# CLK1 0.02fF
C37 x0 EESPFAL_NAND_v3_0/A_bar 0.11fF
C38 EESPFAL_NAND_v3_0/A a_5735_n466# 0.01fF
C39 x1 EESPFAL_NAND_v3_0/B_bar 0.00fF
C40 Dis1 EESPFAL_NAND_v3_1/B 0.09fF
C41 CLK1 a_1795_n2607# 0.01fF
C42 x2 CLK2 0.02fF
C43 x2_bar CLK3 0.00fF
C44 Dis1 x3 0.26fF
C45 Dis2 a_5735_214# 0.00fF
C46 x3_bar CLK2 0.01fF
C47 a_385_214# x2_bar 0.00fF
C48 EESPFAL_NAND_v3_0/A CLK2 0.81fF
C49 a_1645_n466# x2 0.01fF
C50 EESPFAL_NAND_v3_0/A_bar CLK3 0.02fF
C51 a_1645_n466# x3_bar 0.00fF
C52 x3_bar x2 1.77fF
C53 a_1945_n466# x2_bar 0.00fF
C54 x0 a_385_214# 0.00fF
C55 a_5735_n466# EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C56 EESPFAL_NAND_v3_0/A x2 0.23fF
C57 EESPFAL_NAND_v3_0/A a_1645_n466# 0.01fF
C58 a_385_214# EESPFAL_NAND_v3_0/A_bar 0.00fF
C59 a_85_214# EESPFAL_NAND_v3_1/A 0.01fF
C60 EESPFAL_NAND_v3_0/A x3_bar 0.03fF
C61 EESPFAL_NAND_v3_1/A CLK1 1.43fF
C62 x0 a_1945_n466# 0.00fF
C63 a_1945_n466# EESPFAL_NAND_v3_0/A_bar 0.00fF
C64 x2_bar a_1795_n2607# 0.00fF
C65 EESPFAL_INV4_2/A_bar CLK1 1.83fF
C66 x1_bar a_1945_214# 0.00fF
C67 EESPFAL_NAND_v3_1/OUT_bar CLK2 1.18fF
C68 x0 a_1795_n2607# 0.00fF
C69 EESPFAL_NAND_v3_1/A EESPFAL_3in_NOR_v2_0/B_bar 0.00fF
C70 a_1645_n2607# x0_bar 0.00fF
C71 x1_bar EESPFAL_NAND_v3_1/A_bar 1.09fF
C72 EESPFAL_NAND_v3_0/B_bar EESPFAL_3in_NOR_v2_0/C 0.01fF
C73 Dis3 CLK1 0.25fF
C74 EESPFAL_NAND_v3_0/B EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C75 s2 EESPFAL_NAND_v3_0/B 0.00fF
C76 a_1645_214# CLK1 0.02fF
C77 EESPFAL_NAND_v3_1/A x2_bar 0.32fF
C78 CLK1 EESPFAL_NAND_v3_1/B_bar 0.89fF
C79 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_0/B_bar 0.01fF
C80 EESPFAL_INV4_2/A_bar x2_bar 0.19fF
C81 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/OUT_bar 0.01fF
C82 EESPFAL_NAND_v3_1/OUT CLK1 0.01fF
C83 Dis3 EESPFAL_3in_NOR_v2_0/B_bar 0.01fF
C84 s2_bar EESPFAL_3in_NOR_v2_0/B_bar 0.04fF
C85 EESPFAL_INV4_2/A x0_bar 0.01fF
C86 x0 EESPFAL_NAND_v3_1/A 0.01fF
C87 x0 EESPFAL_INV4_2/A_bar 0.06fF
C88 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_1/A 0.02fF
C89 CLK2 a_1945_n2607# 0.00fF
C90 EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_NAND_v3_1/B_bar 0.00fF
C91 EESPFAL_INV4_2/A EESPFAL_NAND_v3_0/B 0.01fF
C92 EESPFAL_INV4_2/A_bar EESPFAL_NAND_v3_0/A_bar 0.03fF
C93 EESPFAL_NAND_v3_0/B_bar EESPFAL_3in_NOR_v2_0/B 0.00fF
C94 x3 a_85_n466# 0.00fF
C95 EESPFAL_NAND_v3_1/OUT EESPFAL_3in_NOR_v2_0/B_bar 0.08fF
C96 Dis3 x2_bar 0.01fF
C97 x1 a_85_214# 0.01fF
C98 x1 CLK1 2.03fF
C99 a_1645_214# x2_bar 0.01fF
C100 Dis2 EESPFAL_NAND_v3_0/B 0.05fF
C101 x2_bar EESPFAL_NAND_v3_1/B_bar 0.02fF
C102 x3_bar a_1945_n2607# 0.01fF
C103 Dis1 x1_bar 0.23fF
C104 Dis3 EESPFAL_NAND_v3_0/A_bar 0.03fF
C105 s2_bar EESPFAL_NAND_v3_0/A_bar 0.00fF
C106 a_5735_n466# EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C107 EESPFAL_NAND_v3_1/A CLK3 0.02fF
C108 x0 a_1645_214# 0.00fF
C109 a_1645_214# EESPFAL_NAND_v3_0/A_bar 0.00fF
C110 x3 x0_bar 0.05fF
C111 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_1/B 0.03fF
C112 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_1/B_bar 0.04fF
C113 a_385_214# EESPFAL_NAND_v3_1/A 0.01fF
C114 Dis1 EESPFAL_NAND_v3_0/B_bar 0.16fF
C115 a_385_n466# x3 0.00fF
C116 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_1/OUT 0.00fF
C117 a_1945_n466# EESPFAL_NAND_v3_1/A 0.00fF
C118 EESPFAL_INV4_2/A_bar a_1945_n466# 0.00fF
C119 Dis3 CLK3 0.41fF
C120 a_1645_n2607# CLK2 0.00fF
C121 EESPFAL_NAND_v3_1/OUT_bar a_6065_n2606# 0.00fF
C122 x1 x2_bar 0.38fF
C123 CLK2 EESPFAL_3in_NOR_v2_0/C_bar 0.90fF
C124 s2 CLK2 0.12fF
C125 s2_bar CLK3 0.99fF
C126 CLK3 EESPFAL_NAND_v3_1/B_bar 0.02fF
C127 x0 x1 1.98fF
C128 CLK3 a_5915_n2606# 0.01fF
C129 x2 EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C130 EESPFAL_INV4_2/A_bar a_1795_n2607# 0.00fF
C131 x1 EESPFAL_NAND_v3_0/A_bar 0.11fF
C132 EESPFAL_NAND_v3_1/OUT CLK3 1.27fF
C133 Dis2 a_5735_n466# 0.00fF
C134 a_1645_n2607# x3_bar 0.00fF
C135 x3_bar EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C136 CLK1 EESPFAL_3in_NOR_v2_0/C 0.10fF
C137 EESPFAL_NAND_v3_0/A EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C138 EESPFAL_INV4_2/A CLK2 0.64fF
C139 EESPFAL_NAND_v3_0/A s2 0.01fF
C140 CLK1 a_1945_214# 0.02fF
C141 EESPFAL_NAND_v3_1/A_bar a_85_214# 0.00fF
C142 EESPFAL_INV4_2/A a_1645_n466# 0.00fF
C143 EESPFAL_INV4_2/A x2 0.14fF
C144 EESPFAL_NAND_v3_1/A_bar CLK1 1.28fF
C145 EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_3in_NOR_v2_0/C 0.06fF
C146 Dis2 CLK2 1.06fF
C147 EESPFAL_INV4_2/A x3_bar 0.07fF
C148 x1 a_385_214# 0.01fF
C149 EESPFAL_NAND_v3_0/A EESPFAL_INV4_2/A 0.07fF
C150 Dis2 x2 0.00fF
C151 EESPFAL_NAND_v3_1/A_bar EESPFAL_3in_NOR_v2_0/B_bar 0.00fF
C152 EESPFAL_3in_NOR_v2_0/B CLK1 0.01fF
C153 CLK2 EESPFAL_NAND_v3_1/B 0.42fF
C154 x1_bar a_85_n466# 0.00fF
C155 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C156 x2_bar EESPFAL_3in_NOR_v2_0/C 0.00fF
C157 x1 a_1945_n466# 0.00fF
C158 Dis2 x3_bar 0.00fF
C159 s2 EESPFAL_NAND_v3_1/OUT_bar 0.01fF
C160 x2_bar a_1945_214# 0.00fF
C161 EESPFAL_NAND_v3_0/A Dis2 0.03fF
C162 Dis3 EESPFAL_NAND_v3_1/A 0.02fF
C163 EESPFAL_INV4_2/A_bar Dis3 0.00fF
C164 x2 EESPFAL_NAND_v3_1/B 0.00fF
C165 x0 EESPFAL_3in_NOR_v2_0/C 0.00fF
C166 a_1645_214# EESPFAL_NAND_v3_1/A 0.00fF
C167 EESPFAL_3in_NOR_v2_0/B EESPFAL_3in_NOR_v2_0/B_bar 0.69fF
C168 x3 x2 0.61fF
C169 EESPFAL_NAND_v3_1/A_bar x2_bar 0.08fF
C170 EESPFAL_NAND_v3_0/A_bar EESPFAL_3in_NOR_v2_0/C 0.00fF
C171 a_1645_n466# x3 0.00fF
C172 x1 a_1795_n2607# 0.01fF
C173 x0 a_1945_214# 0.00fF
C174 x3_bar EESPFAL_NAND_v3_1/B 0.00fF
C175 EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/B_bar 0.03fF
C176 EESPFAL_NAND_v3_0/A_bar a_1945_214# 0.00fF
C177 x3 x3_bar 5.69fF
C178 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/A 0.04fF
C179 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/B 0.00fF
C180 x1_bar x0_bar 0.70fF
C181 a_6065_n2606# EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C182 EESPFAL_NAND_v3_0/A x3 0.00fF
C183 x0 EESPFAL_NAND_v3_1/A_bar 0.01fF
C184 s2 a_6065_n2606# 0.01fF
C185 Dis1 a_85_214# 0.01fF
C186 Dis1 CLK1 1.87fF
C187 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_0/A_bar 0.04fF
C188 a_385_n466# x1_bar 0.00fF
C189 x1_bar EESPFAL_NAND_v3_0/B 0.02fF
C190 s2_bar Dis3 0.28fF
C191 EESPFAL_3in_NOR_v2_0/B x2_bar 0.00fF
C192 a_1945_n2607# EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C193 Dis2 EESPFAL_NAND_v3_1/OUT_bar 0.27fF
C194 Dis3 EESPFAL_NAND_v3_1/B_bar 0.04fF
C195 CLK3 EESPFAL_3in_NOR_v2_0/C 0.50fF
C196 EESPFAL_NAND_v3_0/B_bar x0_bar 0.00fF
C197 Dis3 a_5915_n2606# 0.00fF
C198 s2_bar a_5915_n2606# 0.00fF
C199 Dis1 EESPFAL_3in_NOR_v2_0/B_bar 0.00fF
C200 Dis3 EESPFAL_NAND_v3_1/OUT 0.03fF
C201 EESPFAL_NAND_v3_0/A_bar EESPFAL_3in_NOR_v2_0/B 0.02fF
C202 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_0/B_bar 0.48fF
C203 x1 EESPFAL_NAND_v3_1/A 0.10fF
C204 a_1645_214# EESPFAL_NAND_v3_1/B_bar 0.00fF
C205 s2_bar EESPFAL_NAND_v3_1/OUT 0.07fF
C206 x1 EESPFAL_INV4_2/A_bar 0.06fF
C207 EESPFAL_NAND_v3_1/A_bar CLK3 0.01fF
C208 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/B_bar 0.00fF
C209 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_1/B 0.15fF
C210 EESPFAL_NAND_v3_1/OUT a_5915_n2606# 0.00fF
C211 EESPFAL_INV4_2/A a_1945_n2607# 0.01fF
C212 Dis1 x2_bar 0.28fF
C213 EESPFAL_NAND_v3_1/A_bar a_385_214# 0.00fF
C214 x1 Dis3 0.00fF
C215 EESPFAL_3in_NOR_v2_0/B_bar a_5735_214# 0.00fF
C216 EESPFAL_3in_NOR_v2_0/B CLK3 0.82fF
C217 a_1945_n466# EESPFAL_NAND_v3_1/A_bar 0.00fF
C218 a_1795_n2607# EESPFAL_3in_NOR_v2_0/C 0.00fF
C219 x0 Dis1 0.32fF
C220 x1 a_1645_214# 0.01fF
C221 Dis1 EESPFAL_NAND_v3_0/A_bar 0.38fF
C222 x1 EESPFAL_NAND_v3_1/B_bar 0.04fF
C223 a_1645_n2607# EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C224 s2 EESPFAL_3in_NOR_v2_0/C_bar 0.08fF
C225 x1_bar CLK2 0.02fF
C226 Dis1 CLK3 0.00fF
C227 EESPFAL_INV4_2/A a_1645_n2607# 0.01fF
C228 EESPFAL_INV4_2/A EESPFAL_3in_NOR_v2_0/C_bar 0.33fF
C229 EESPFAL_INV4_2/A_bar EESPFAL_3in_NOR_v2_0/C 0.01fF
C230 EESPFAL_NAND_v3_1/A a_1945_214# 0.00fF
C231 EESPFAL_INV4_2/A s2 0.00fF
C232 Dis1 a_385_214# 0.02fF
C233 CLK1 a_85_n466# 0.01fF
C234 a_1645_n466# x1_bar 0.00fF
C235 x1_bar x2 4.03fF
C236 EESPFAL_NAND_v3_0/B_bar CLK2 0.13fF
C237 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/A 2.86fF
C238 Dis2 EESPFAL_3in_NOR_v2_0/C_bar 0.23fF
C239 a_1945_n466# Dis1 0.00fF
C240 x1_bar x3_bar 0.13fF
C241 EESPFAL_INV4_2/A_bar EESPFAL_NAND_v3_1/A_bar 0.00fF
C242 Dis2 s2 0.01fF
C243 EESPFAL_NAND_v3_0/A x1_bar 0.08fF
C244 Dis3 EESPFAL_3in_NOR_v2_0/C 0.17fF
C245 a_5735_214# CLK3 0.00fF
C246 a_1645_n466# EESPFAL_NAND_v3_0/B_bar 0.00fF
C247 EESPFAL_NAND_v3_0/B_bar x2 0.04fF
C248 s2_bar EESPFAL_3in_NOR_v2_0/C 0.11fF
C249 EESPFAL_NAND_v3_1/A EESPFAL_3in_NOR_v2_0/B 0.00fF
C250 a_5915_n2606# EESPFAL_3in_NOR_v2_0/C 0.00fF
C251 a_85_214# x0_bar 0.00fF
C252 CLK1 x0_bar 0.34fF
C253 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/B_bar 0.08fF
C254 a_1945_214# EESPFAL_NAND_v3_1/B_bar 0.00fF
C255 EESPFAL_NAND_v3_1/A_bar Dis3 0.02fF
C256 EESPFAL_NAND_v3_1/OUT EESPFAL_3in_NOR_v2_0/C 0.10fF
C257 a_385_n466# CLK1 0.01fF
C258 EESPFAL_NAND_v3_0/B CLK1 1.04fF
C259 Dis2 EESPFAL_INV4_2/A 0.04fF
C260 x2_bar a_85_n466# 0.00fF
C261 EESPFAL_NAND_v3_1/A_bar a_1645_214# 0.01fF
C262 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/B_bar 0.42fF
C263 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/OUT 0.01fF
C264 Dis3 EESPFAL_3in_NOR_v2_0/B 0.02fF
C265 x1_bar EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C266 x0 a_85_n466# 0.00fF
C267 EESPFAL_NAND_v3_0/A_bar a_85_n466# 0.01fF
C268 EESPFAL_NAND_v3_0/B EESPFAL_3in_NOR_v2_0/B_bar 0.15fF
C269 s2_bar EESPFAL_3in_NOR_v2_0/B 0.10fF
C270 x1 EESPFAL_3in_NOR_v2_0/C 0.00fF
C271 Dis1 EESPFAL_NAND_v3_1/A 0.33fF
C272 EESPFAL_INV4_2/A x3 0.02fF
C273 EESPFAL_INV4_2/A_bar Dis1 0.37fF
C274 EESPFAL_3in_NOR_v2_0/B a_5915_n2606# 0.01fF
C275 x1 a_1945_214# 0.01fF
C276 x2_bar x0_bar 0.52fF
C277 EESPFAL_NAND_v3_1/OUT EESPFAL_3in_NOR_v2_0/B 1.75fF
C278 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_0/B_bar 0.00fF
C279 Dis2 EESPFAL_NAND_v3_1/B 0.04fF
C280 a_385_n466# x2_bar 0.00fF
C281 EESPFAL_NAND_v3_0/B x2_bar 0.06fF
C282 x1 EESPFAL_NAND_v3_1/A_bar 0.21fF
C283 x0 x0_bar 5.48fF
C284 EESPFAL_NAND_v3_0/A_bar x0_bar 0.31fF
C285 x0 a_385_n466# 0.01fF
C286 Dis1 Dis3 0.02fF
C287 x0 EESPFAL_NAND_v3_0/B 0.01fF
C288 a_385_n466# EESPFAL_NAND_v3_0/A_bar 0.01fF
C289 EESPFAL_NAND_v3_1/A a_5735_214# 0.01fF
C290 x1_bar a_1945_n2607# 0.00fF
C291 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/B 0.78fF
C292 Dis1 a_1645_214# 0.01fF
C293 x3 EESPFAL_NAND_v3_1/B 0.00fF
C294 Dis1 EESPFAL_NAND_v3_1/B_bar 0.16fF
C295 Dis1 EESPFAL_NAND_v3_1/OUT 0.00fF
C296 a_5735_n466# EESPFAL_3in_NOR_v2_0/B_bar 0.00fF
C297 Dis3 a_5735_214# 0.00fF
C298 CLK1 CLK2 1.21fF
C299 EESPFAL_NAND_v3_0/B CLK3 0.07fF
C300 a_385_214# x0_bar 0.00fF
C301 a_85_214# x2 0.00fF
C302 a_1645_n466# CLK1 0.02fF
C303 x2 CLK1 1.32fF
C304 x1 Dis1 0.52fF
C305 EESPFAL_NAND_v3_1/OUT a_5735_214# 0.01fF
C306 EESPFAL_3in_NOR_v2_0/B_bar CLK2 1.22fF
C307 a_85_214# x3_bar 0.00fF
C308 x3_bar CLK1 1.88fF
C309 a_1945_n466# EESPFAL_NAND_v3_0/B 0.00fF
C310 EESPFAL_NAND_v3_0/A CLK1 1.48fF
C311 x1_bar a_1645_n2607# 0.00fF
C312 EESPFAL_NAND_v3_1/A_bar a_1945_214# 0.01fF
C313 x2_bar CLK2 0.11fF
C314 EESPFAL_NAND_v3_1/A a_85_n466# 0.00fF
C315 EESPFAL_NAND_v3_0/A EESPFAL_3in_NOR_v2_0/B_bar 0.07fF
C316 EESPFAL_NAND_v3_0/B_bar EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C317 EESPFAL_3in_NOR_v2_0/B EESPFAL_3in_NOR_v2_0/C 1.44fF
C318 s2 EESPFAL_NAND_v3_0/B_bar 0.00fF
C319 x2_bar x2 5.04fF
C320 x0 CLK2 0.02fF
C321 a_1645_n466# x2_bar 0.01fF
C322 EESPFAL_NAND_v3_0/A_bar CLK2 0.18fF
C323 a_5735_n466# CLK3 0.01fF
C324 EESPFAL_INV4_2/A x1_bar 0.02fF
C325 x3_bar x2_bar 0.26fF
C326 EESPFAL_NAND_v3_1/OUT_bar CLK1 0.05fF
C327 EESPFAL_NAND_v3_0/A x2_bar 0.73fF
C328 x0 x2 1.60fF
C329 x0 a_1645_n466# 0.00fF
C330 EESPFAL_NAND_v3_1/A x0_bar 0.03fF
C331 a_1645_n466# EESPFAL_NAND_v3_0/A_bar 0.00fF
C332 EESPFAL_NAND_v3_0/A_bar x2 0.15fF
C333 EESPFAL_INV4_2/A_bar x0_bar 0.06fF
C334 x0 x3_bar 0.06fF
C335 Dis2 x1_bar 0.00fF
C336 EESPFAL_INV4_2/A EESPFAL_NAND_v3_0/B_bar 0.01fF
C337 a_385_n466# EESPFAL_NAND_v3_1/A 0.00fF
C338 EESPFAL_NAND_v3_0/A_bar x3_bar 0.04fF
C339 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_1/A 0.00fF
C340 x0 EESPFAL_NAND_v3_0/A 0.10fF
C341 Dis1 EESPFAL_3in_NOR_v2_0/C 0.00fF
C342 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_0/A_bar 1.17fF
C343 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_3in_NOR_v2_0/B_bar 0.81fF
C344 CLK2 CLK3 1.30fF
C345 Dis1 a_1945_214# 0.00fF
C346 Dis2 EESPFAL_NAND_v3_0/B_bar 0.02fF
C347 x1_bar EESPFAL_NAND_v3_1/B 0.07fF
C348 Dis1 EESPFAL_NAND_v3_1/A_bar 0.31fF
C349 x1_bar x3 0.79fF
C350 Dis3 EESPFAL_NAND_v3_0/B 0.06fF
C351 a_1645_214# x0_bar 0.00fF
C352 CLK1 a_1945_n2607# 0.01fF
C353 s2_bar EESPFAL_NAND_v3_0/B 0.00fF
C354 a_385_214# x2 0.01fF
C355 EESPFAL_NAND_v3_0/B_bar EESPFAL_NAND_v3_1/B 0.02fF
C356 x1 a_85_n466# 0.00fF
C357 EESPFAL_NAND_v3_0/A CLK3 0.20fF
C358 a_6065_n2606# EESPFAL_3in_NOR_v2_0/B_bar 0.00fF
C359 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_1/B_bar 0.02fF
C360 a_385_214# x3_bar 0.00fF
C361 Dis1 EESPFAL_3in_NOR_v2_0/B 0.00fF
C362 a_1945_n466# x2 0.01fF
C363 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C364 EESPFAL_NAND_v3_0/B EESPFAL_NAND_v3_1/OUT 0.03fF
C365 CLK2 a_1795_n2607# 0.00fF
C366 a_1945_n466# x3_bar 0.00fF
C367 a_5735_n466# EESPFAL_NAND_v3_1/A 0.00fF
C368 EESPFAL_NAND_v3_0/A a_1945_n466# 0.01fF
C369 x1 x0_bar 3.57fF
C370 x2_bar a_1945_n2607# 0.00fF
C371 x3_bar a_1795_n2607# 0.00fF
C372 x1 a_385_n466# 0.00fF
C373 EESPFAL_3in_NOR_v2_0/B a_5735_214# 0.00fF
C374 x1 EESPFAL_NAND_v3_0/B 0.00fF
C375 EESPFAL_NAND_v3_1/OUT_bar CLK3 0.20fF
C376 a_5735_n466# Dis3 0.00fF
C377 x0 a_1945_n2607# 0.00fF
C378 EESPFAL_NAND_v3_1/A CLK2 0.66fF
C379 a_1645_n2607# CLK1 0.01fF
C380 CLK1 EESPFAL_3in_NOR_v2_0/C_bar 0.15fF
C381 EESPFAL_INV4_2/A_bar CLK2 0.20fF
C382 EESPFAL_NAND_v3_1/A x2 0.18fF
C383 a_1645_n466# EESPFAL_NAND_v3_1/A 0.00fF
C384 EESPFAL_INV4_2/A_bar x2 0.13fF
C385 a_5735_n466# EESPFAL_NAND_v3_1/OUT 0.01fF
C386 EESPFAL_INV4_2/A_bar a_1645_n466# 0.00fF
C387 a_6065_n2606# CLK3 0.01fF
C388 EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_3in_NOR_v2_0/C_bar 0.22fF
C389 EESPFAL_NAND_v3_1/A x3_bar 0.09fF
C390 s2 EESPFAL_3in_NOR_v2_0/B_bar 0.02fF
C391 EESPFAL_INV4_2/A_bar x3_bar 0.05fF
C392 Dis3 CLK2 0.19fF
C393 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/A 0.02fF
C394 s2_bar CLK2 0.16fF
C395 EESPFAL_NAND_v3_0/A EESPFAL_INV4_2/A_bar 0.03fF
C396 EESPFAL_INV4_2/A CLK1 0.89fF
C397 CLK2 EESPFAL_NAND_v3_1/B_bar 0.03fF
C398 Dis3 x2 0.00fF
C399 a_1645_n2607# x2_bar 0.00fF
C400 CLK2 a_5915_n2606# 0.00fF
C401 x2_bar EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C402 EESPFAL_NAND_v3_1/OUT CLK2 0.96fF
C403 Dis2 CLK1 0.05fF
C404 a_1645_214# x2 0.01fF
C405 EESPFAL_NAND_v3_0/A Dis3 0.01fF
C406 x0 a_1645_n2607# 0.01fF
C407 x2 EESPFAL_NAND_v3_1/B_bar 0.01fF
C408 x0 EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C409 a_1645_214# x3_bar 0.00fF
C410 EESPFAL_NAND_v3_0/A s2_bar 0.02fF
C411 EESPFAL_NAND_v3_0/A_bar EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C412 EESPFAL_NAND_v3_0/B EESPFAL_3in_NOR_v2_0/C 0.01fF
C413 s2 EESPFAL_NAND_v3_0/A_bar 0.00fF
C414 x3_bar EESPFAL_NAND_v3_1/B_bar 0.00fF
C415 EESPFAL_NAND_v3_0/A a_1645_214# 0.00fF
C416 Dis2 EESPFAL_3in_NOR_v2_0/B_bar 0.26fF
C417 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_1/A 0.06fF
C418 EESPFAL_NAND_v3_1/A_bar x0_bar 0.02fF
C419 CLK1 EESPFAL_NAND_v3_1/B 0.83fF
C420 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/B_bar 0.00fF
C421 EESPFAL_INV4_2/A x2_bar 0.07fF
C422 x3 a_85_214# 0.00fF
C423 x1_bar EESPFAL_NAND_v3_0/B_bar 0.03fF
C424 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/OUT 0.08fF
C425 x3 CLK1 1.27fF
C426 x1 CLK2 0.02fF
C427 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_0/B 0.01fF
C428 x0 EESPFAL_INV4_2/A 0.09fF
C429 EESPFAL_3in_NOR_v2_0/B_bar EESPFAL_NAND_v3_1/B 0.02fF
C430 x1 a_1645_n466# 0.01fF
C431 Dis2 x2_bar 0.00fF
C432 x1 x2 0.50fF
C433 CLK3 EESPFAL_3in_NOR_v2_0/C_bar 0.32fF
C434 EESPFAL_INV4_2/A EESPFAL_NAND_v3_0/A_bar 0.02fF
C435 s2 CLK3 1.07fF
C436 Dis3 EESPFAL_NAND_v3_1/OUT_bar 0.01fF
C437 Dis1 a_85_n466# 0.01fF
C438 x1 x3_bar 1.88fF
C439 EESPFAL_NAND_v3_0/B EESPFAL_3in_NOR_v2_0/B 0.08fF
C440 s2_bar EESPFAL_NAND_v3_1/OUT_bar 0.10fF
C441 EESPFAL_NAND_v3_0/A x1 0.08fF
C442 x0 Dis2 0.00fF
C443 Dis2 EESPFAL_NAND_v3_0/A_bar 0.02fF
C444 x2_bar EESPFAL_NAND_v3_1/B 0.01fF
C445 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_NAND_v3_1/B_bar 0.09fF
C446 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/OUT_bar 0.80fF
C447 x3 x2_bar 3.12fF
C448 EESPFAL_INV4_2/A_bar a_1945_n2607# 0.00fF
C449 a_5735_n466# EESPFAL_3in_NOR_v2_0/C 0.00fF
C450 EESPFAL_INV4_2/A CLK3 0.01fF
C451 Dis3 a_6065_n2606# 0.00fF
C452 Dis1 x0_bar 0.15fF
C453 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_1/B 0.04fF
C454 s2_bar a_6065_n2606# 0.00fF
C455 x0 x3 0.04fF
C456 a_1795_n2607# EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C457 x3 EESPFAL_NAND_v3_0/A_bar 0.01fF
C458 a_385_n466# Dis1 0.02fF
C459 Dis1 EESPFAL_NAND_v3_0/B 0.09fF
C460 Dis2 CLK3 2.44fF
C461 EESPFAL_INV4_2/A a_1945_n466# 0.00fF
C462 EESPFAL_NAND_v3_1/OUT a_6065_n2606# 0.00fF
C463 CLK2 EESPFAL_3in_NOR_v2_0/C 1.06fF
C464 a_5735_n466# EESPFAL_3in_NOR_v2_0/B 0.01fF
C465 CLK3 EESPFAL_NAND_v3_1/B 0.03fF
C466 x2 EESPFAL_3in_NOR_v2_0/C 0.00fF
C467 EESPFAL_INV4_2/A a_1795_n2607# 0.01fF
C468 EESPFAL_NAND_v3_1/A_bar CLK2 0.07fF
C469 x2 a_1945_214# 0.01fF
C470 x3_bar EESPFAL_3in_NOR_v2_0/C 0.00fF
C471 EESPFAL_INV4_2/A_bar EESPFAL_3in_NOR_v2_0/C_bar 0.02fF
C472 EESPFAL_INV4_2/A_bar a_1645_n2607# 0.00fF
C473 x3_bar a_1945_214# 0.00fF
C474 EESPFAL_NAND_v3_0/A EESPFAL_3in_NOR_v2_0/C 0.03fF
C475 x3 a_385_214# 0.00fF
C476 EESPFAL_INV4_2/A_bar s2 0.00fF
C477 a_1645_n466# EESPFAL_NAND_v3_1/A_bar 0.00fF
C478 EESPFAL_NAND_v3_1/A_bar x2 0.13fF
C479 EESPFAL_NAND_v3_0/A a_1945_214# 0.00fF
C480 EESPFAL_3in_NOR_v2_0/B CLK2 0.94fF
C481 EESPFAL_NAND_v3_1/A_bar x3_bar 0.03fF
C482 EESPFAL_NAND_v3_0/A EESPFAL_NAND_v3_1/A_bar 0.02fF
C483 x1_bar a_85_214# 0.00fF
C484 x1_bar CLK1 1.99fF
C485 Dis3 EESPFAL_3in_NOR_v2_0/C_bar 0.18fF
C486 s2_bar EESPFAL_3in_NOR_v2_0/C_bar 1.69fF
C487 EESPFAL_INV4_2/A EESPFAL_NAND_v3_1/A 0.00fF
C488 s2 Dis3 0.41fF
C489 s2_bar s2 1.81fF
C490 EESPFAL_INV4_2/A EESPFAL_INV4_2/A_bar 0.97fF
C491 a_5915_n2606# EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C492 s2 a_5915_n2606# 0.01fF
C493 EESPFAL_NAND_v3_0/A EESPFAL_3in_NOR_v2_0/B 0.06fF
C494 EESPFAL_NAND_v3_0/B_bar CLK1 0.87fF
C495 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_3in_NOR_v2_0/C 0.10fF
C496 EESPFAL_NAND_v3_1/OUT EESPFAL_3in_NOR_v2_0/C_bar 0.01fF
C497 Dis2 EESPFAL_NAND_v3_1/A 0.01fF
C498 s2 EESPFAL_NAND_v3_1/OUT 0.04fF
C499 Dis2 EESPFAL_INV4_2/A_bar 0.01fF
C500 Dis1 CLK2 0.01fF
C501 EESPFAL_INV4_2/A Dis3 0.00fF
C502 EESPFAL_INV4_2/A s2_bar 0.00fF
C503 a_85_n466# x0_bar 0.00fF
C504 EESPFAL_NAND_v3_0/B_bar EESPFAL_3in_NOR_v2_0/B_bar 0.09fF
C505 EESPFAL_NAND_v3_1/A_bar EESPFAL_NAND_v3_1/OUT_bar 0.05fF
C506 x1_bar x2_bar 0.15fF
C507 Dis1 x2 0.56fF
C508 a_1645_n466# Dis1 0.01fF
C509 EESPFAL_NAND_v3_1/A EESPFAL_NAND_v3_1/B 0.97fF
C510 x3 EESPFAL_NAND_v3_1/A 0.07fF
C511 x1 EESPFAL_3in_NOR_v2_0/C_bar 0.00fF
C512 Dis2 Dis3 1.35fF
C513 x1 a_1645_n2607# 0.00fF
C514 Dis1 x3_bar 0.48fF
C515 EESPFAL_INV4_2/A_bar x3 0.05fF
C516 a_6065_n2606# EESPFAL_3in_NOR_v2_0/C 0.00fF
C517 EESPFAL_INV4_2/A EESPFAL_NAND_v3_1/OUT 0.01fF
C518 Dis2 s2_bar 0.01fF
C519 x0 x1_bar 1.94fF
C520 EESPFAL_NAND_v3_0/A Dis1 0.29fF
C521 EESPFAL_NAND_v3_1/OUT_bar EESPFAL_3in_NOR_v2_0/B 0.06fF
C522 EESPFAL_NAND_v3_0/B_bar x2_bar 0.30fF
C523 x1_bar EESPFAL_NAND_v3_0/A_bar 0.12fF
C524 a_5735_214# CLK2 0.02fF
C525 a_1945_n2607# EESPFAL_3in_NOR_v2_0/C 0.00fF
C526 Dis2 EESPFAL_NAND_v3_1/B_bar 0.02fF
C527 Dis2 EESPFAL_NAND_v3_1/OUT 0.11fF
C528 Dis3 EESPFAL_NAND_v3_1/B 0.05fF
C529 x0 EESPFAL_NAND_v3_0/B_bar 0.01fF
C530 a_385_n466# x0_bar 0.00fF
C531 EESPFAL_NAND_v3_0/B x0_bar 0.00fF
C532 EESPFAL_NAND_v3_0/A_bar EESPFAL_NAND_v3_0/B_bar 0.33fF
C533 x1 EESPFAL_INV4_2/A 0.09fF
C534 EESPFAL_NAND_v3_1/B EESPFAL_NAND_v3_1/B_bar 0.50fF
C535 x3 a_1645_214# 0.00fF
C536 EESPFAL_NAND_v3_0/A a_5735_214# 0.00fF
C537 x3 EESPFAL_NAND_v3_1/B_bar 0.00fF
C538 EESPFAL_NAND_v3_1/OUT EESPFAL_NAND_v3_1/B 0.07fF
C539 EESPFAL_3in_NOR_v2_0/B a_6065_n2606# 0.00fF
C540 x1_bar CLK3 0.00fF
C541 Dis1 EESPFAL_NAND_v3_1/OUT_bar 0.00fF
C542 x1 Dis2 0.00fF
C543 x1_bar a_385_214# 0.00fF
C544 EESPFAL_NAND_v3_0/B_bar CLK3 0.03fF
C545 a_1945_n466# x1_bar 0.00fF
C546 x1 EESPFAL_NAND_v3_1/B 0.01fF
C547 EESPFAL_3in_NOR_v2_0/C EESPFAL_3in_NOR_v2_0/C_bar 2.14fF
C548 x1 x3 0.11fF
C549 s2 EESPFAL_3in_NOR_v2_0/C 0.08fF
C550 EESPFAL_NAND_v3_1/OUT_bar a_5735_214# 0.00fF
C551 x1_bar a_1795_n2607# 0.00fF
C552 a_1945_n466# EESPFAL_NAND_v3_0/B_bar 0.00fF
C553 a_85_214# CLK1 0.01fF
C554 x2 a_85_n466# 0.01fF
C555 EESPFAL_INV4_2/A EESPFAL_3in_NOR_v2_0/C 0.07fF
C556 x3_bar a_85_n466# 0.00fF
C557 EESPFAL_NAND_v3_0/A a_85_n466# 0.00fF
C558 CLK1 EESPFAL_3in_NOR_v2_0/B_bar 0.04fF
C559 EESPFAL_3in_NOR_v2_0/B EESPFAL_3in_NOR_v2_0/C_bar 0.10fF
C560 s2 EESPFAL_3in_NOR_v2_0/B 0.05fF
C561 x1_bar EESPFAL_NAND_v3_1/A 0.27fF
C562 Dis2 EESPFAL_3in_NOR_v2_0/C 0.39fF
C563 EESPFAL_NAND_v3_0/B CLK2 0.50fF
C564 EESPFAL_INV4_2/A_bar x1_bar 0.06fF
C565 a_1645_n466# x0_bar 0.00fF
C566 x2 x0_bar 0.12fF
C567 a_85_214# x2_bar 0.00fF
C568 x2_bar CLK1 1.88fF
C569 a_385_n466# x2 0.01fF
C570 EESPFAL_NAND_v3_0/B x2 0.01fF
C571 x3_bar x0_bar 0.06fF
C572 a_6065_n2606# GND 0.02fF
C573 a_5915_n2606# GND 0.02fF
C574 a_1945_n2607# GND 0.02fF
C575 a_1795_n2607# GND 0.02fF
C576 a_1645_n2607# GND 0.02fF
C577 Dis3 GND 3.93fF
C578 s2 GND 1.26fF
C579 s2_bar GND 0.98fF
C580 EESPFAL_3in_NOR_v2_0/C_bar GND 1.25fF $ **FLOATING
C581 EESPFAL_3in_NOR_v2_0/C GND 1.26fF $ **FLOATING
C582 EESPFAL_INV4_2/A_bar GND 1.72fF
C583 EESPFAL_INV4_2/A GND 1.68fF
C584 a_5735_n466# GND 0.02fF
C585 a_1945_n466# GND 0.01fF
C586 a_1645_n466# GND 0.01fF
C587 a_385_n466# GND 0.02fF
C588 a_85_n466# GND 0.01fF
C589 EESPFAL_3in_NOR_v2_0/B_bar GND 1.53fF
C590 EESPFAL_3in_NOR_v2_0/B GND 1.16fF
C591 EESPFAL_NAND_v3_0/B_bar GND 1.09fF
C592 EESPFAL_NAND_v3_0/B GND 1.24fF
C593 EESPFAL_NAND_v3_0/A_bar GND 1.57fF
C594 EESPFAL_NAND_v3_0/A GND 1.41fF
C595 x0 GND 4.42fF
C596 x0_bar GND 3.37fF
C597 a_5735_214# GND 0.02fF
C598 a_1945_214# GND 0.01fF
C599 a_1645_214# GND 0.01fF
C600 a_385_214# GND 0.02fF
C601 a_85_214# GND 0.01fF
C602 Dis2 GND 5.04fF
C603 x1 GND 2.58fF
C604 x1_bar GND 7.60fF
C605 Dis1 GND 9.00fF
C606 EESPFAL_NAND_v3_1/OUT_bar GND 2.62fF $ **FLOATING
C607 EESPFAL_NAND_v3_1/OUT GND 1.72fF
C608 EESPFAL_NAND_v3_1/B_bar GND 1.18fF
C609 EESPFAL_NAND_v3_1/B GND 1.38fF
C610 x2 GND 2.17fF
C611 x2_bar GND 1.89fF
C612 x3_bar GND 9.41fF
C613 EESPFAL_NAND_v3_1/A GND 2.39fF $ **FLOATING
C614 EESPFAL_NAND_v3_1/A_bar GND 1.71fF $ **FLOATING
C615 x3 GND 6.66fF
C616 CLK3 GND 3.88fF
C617 CLK2 GND 9.51fF
C618 CLK1 GND 17.31fF
C619 x0.t2 GND 0.19fF
C620 x0.t1 GND 0.12fF
C621 x0.t0 GND 0.12fF
C622 x0.n0 GND 1.40fF $ **FLOATING
C623 EESPFAL_XOR_v3_1/B GND 0.33fF $ **FLOATING
C624 x0.n1 GND 2.97fF $ **FLOATING
C625 Dis3.t1 GND 0.08fF
C626 Dis3.t0 GND 0.08fF
C627 Dis3.n0 GND 0.39fF $ **FLOATING
C628 x3_bar.t1 GND 0.30fF
C629 x3_bar.t0 GND 0.36fF
C630 x3_bar.t2 GND 0.20fF
C631 x3_bar.n0 GND 1.90fF $ **FLOATING
C632 EESPFAL_4in_NAND_0/A GND 2.44fF $ **FLOATING
C633 Dis2.t2 GND 0.19fF
C634 Dis2.t3 GND 0.12fF
C635 Dis2.n0 GND 0.49fF $ **FLOATING
C636 EESPFAL_NAND_v3_0/Dis GND 0.20fF $ **FLOATING
C637 Dis2.t4 GND 0.19fF
C638 Dis2.t1 GND 0.12fF
C639 Dis2.n1 GND 0.49fF $ **FLOATING
C640 Dis2.n2 GND 0.80fF $ **FLOATING
C641 Dis2.n3 GND 2.24fF $ **FLOATING
C642 Dis2.t5 GND 0.12fF
C643 Dis2.n4 GND 1.26fF $ **FLOATING
C644 Dis2.t0 GND 0.12fF
C645 Dis2.n5 GND 0.26fF $ **FLOATING
C646 EESPFAL_INV4_2/Dis GND -0.23fF $ **FLOATING
C647 x0_bar.t2 GND 0.19fF
C648 x0_bar.t1 GND 0.49fF
C649 x0_bar.t0 GND 0.17fF
C650 x0_bar.n0 GND 1.62fF $ **FLOATING
C651 EESPFAL_XOR_v3_1/B_bar GND 0.32fF $ **FLOATING
C652 x0_bar.n1 GND 4.41fF $ **FLOATING
C653 CLK3.t8 GND 0.03fF
C654 CLK3.t6 GND 0.03fF
C655 CLK3.n0 GND 0.08fF $ **FLOATING
C656 CLK3.t10 GND 0.04fF
C657 CLK3.t2 GND 0.06fF
C658 CLK3.n1 GND 0.10fF $ **FLOATING
C659 CLK3.n2 GND 0.29fF $ **FLOATING
C660 CLK3.n3 GND 0.06fF $ **FLOATING
C661 CLK3.n4 GND 0.02fF $ **FLOATING
C662 CLK3.n5 GND 0.02fF $ **FLOATING
C663 CLK3.n6 GND 0.02fF $ **FLOATING
C664 CLK3.n7 GND 0.05fF $ **FLOATING
C665 CLK3.n8 GND 0.02fF $ **FLOATING
C666 CLK3.n9 GND 0.02fF $ **FLOATING
C667 CLK3.n10 GND 0.02fF $ **FLOATING
C668 CLK3.n11 GND 0.05fF $ **FLOATING
C669 CLK3.n12 GND 0.02fF $ **FLOATING
C670 CLK3.n13 GND 0.02fF $ **FLOATING
C671 CLK3.n14 GND 0.02fF $ **FLOATING
C672 CLK3.n15 GND 0.05fF $ **FLOATING
C673 CLK3.n16 GND 0.02fF $ **FLOATING
C674 CLK3.n17 GND 0.02fF $ **FLOATING
C675 CLK3.n18 GND 0.02fF $ **FLOATING
C676 CLK3.n19 GND 0.05fF $ **FLOATING
C677 CLK3.n20 GND 0.02fF $ **FLOATING
C678 CLK3.n21 GND 0.02fF $ **FLOATING
C679 CLK3.n22 GND 0.02fF $ **FLOATING
C680 CLK3.n23 GND 0.05fF $ **FLOATING
C681 CLK3.n24 GND 0.02fF $ **FLOATING
C682 CLK3.n25 GND 0.02fF $ **FLOATING
C683 CLK3.n26 GND 0.02fF $ **FLOATING
C684 CLK3.n27 GND 0.11fF $ **FLOATING
C685 CLK3.n28 GND 0.02fF $ **FLOATING
C686 CLK3.n29 GND 0.02fF $ **FLOATING
C687 CLK3.n30 GND 0.02fF $ **FLOATING
C688 CLK3.n31 GND 0.14fF $ **FLOATING
C689 CLK3.n32 GND 0.02fF $ **FLOATING
C690 CLK3.n33 GND 0.02fF $ **FLOATING
C691 CLK3.n34 GND 0.02fF $ **FLOATING
C692 CLK3.n35 GND 0.24fF $ **FLOATING
C693 CLK3.t9 GND 0.07fF
C694 CLK3.n36 GND 0.09fF $ **FLOATING
C695 CLK3.n37 GND 0.02fF $ **FLOATING
C696 CLK3.n38 GND 0.02fF $ **FLOATING
C697 CLK3.n39 GND 0.02fF $ **FLOATING
C698 CLK3.n40 GND 0.13fF $ **FLOATING
C699 CLK3.n41 GND 0.02fF $ **FLOATING
C700 CLK3.n42 GND 0.02fF $ **FLOATING
C701 CLK3.n43 GND 0.02fF $ **FLOATING
C702 CLK3.t7 GND 0.07fF
C703 CLK3.n44 GND 0.08fF $ **FLOATING
C704 CLK3.n45 GND 0.02fF $ **FLOATING
C705 CLK3.n46 GND 0.02fF $ **FLOATING
C706 CLK3.n47 GND 0.02fF $ **FLOATING
C707 CLK3.n48 GND 0.14fF $ **FLOATING
C708 CLK3.n49 GND 0.02fF $ **FLOATING
C709 CLK3.n50 GND 0.02fF $ **FLOATING
C710 CLK3.n51 GND 0.14fF $ **FLOATING
C711 CLK3.t4 GND 0.04fF
C712 CLK3.t0 GND 0.03fF
C713 CLK3.t1 GND 0.03fF
C714 CLK3.n52 GND 0.13fF $ **FLOATING
C715 CLK3.n53 GND 0.01fF $ **FLOATING
C716 CLK3.n54 GND 0.19fF $ **FLOATING
C717 CLK3.t11 GND 0.06fF
C718 CLK3.n55 GND 0.10fF $ **FLOATING
C719 CLK3.n56 GND 0.29fF $ **FLOATING
C720 CLK3.n57 GND 0.01fF $ **FLOATING
C721 CLK3.n58 GND 0.00fF $ **FLOATING
C722 CLK3.n60 GND 0.06fF $ **FLOATING
C723 CLK3.n61 GND 0.02fF $ **FLOATING
C724 CLK3.n62 GND 0.02fF $ **FLOATING
C725 CLK3.n63 GND 0.00fF $ **FLOATING
C726 CLK3.n64 GND 0.01fF $ **FLOATING
C727 CLK3.n65 GND 0.05fF $ **FLOATING
C728 CLK3.n66 GND 0.02fF $ **FLOATING
C729 CLK3.n67 GND 0.02fF $ **FLOATING
C730 CLK3.n68 GND 0.02fF $ **FLOATING
C731 CLK3.n69 GND 0.05fF $ **FLOATING
C732 CLK3.n70 GND 0.02fF $ **FLOATING
C733 CLK3.n71 GND 0.02fF $ **FLOATING
C734 CLK3.n72 GND 0.02fF $ **FLOATING
C735 CLK3.n73 GND 0.05fF $ **FLOATING
C736 CLK3.n74 GND 0.02fF $ **FLOATING
C737 CLK3.n75 GND 0.02fF $ **FLOATING
C738 CLK3.n76 GND 0.01fF $ **FLOATING
C739 CLK3.n77 GND 0.15fF $ **FLOATING
C740 CLK3.n78 GND 0.05fF $ **FLOATING
C741 CLK3.n79 GND 0.02fF $ **FLOATING
C742 CLK3.n80 GND 0.02fF $ **FLOATING
C743 CLK3.n81 GND 0.02fF $ **FLOATING
C744 CLK3.n82 GND 0.05fF $ **FLOATING
C745 CLK3.n83 GND 0.02fF $ **FLOATING
C746 CLK3.n84 GND 0.02fF $ **FLOATING
C747 CLK3.n85 GND 0.02fF $ **FLOATING
C748 CLK3.n86 GND 0.11fF $ **FLOATING
C749 CLK3.n87 GND 0.02fF $ **FLOATING
C750 CLK3.n88 GND 0.02fF $ **FLOATING
C751 CLK3.n89 GND 0.02fF $ **FLOATING
C752 CLK3.n90 GND 0.14fF $ **FLOATING
C753 CLK3.n91 GND 0.02fF $ **FLOATING
C754 CLK3.n92 GND 0.02fF $ **FLOATING
C755 CLK3.n93 GND 0.02fF $ **FLOATING
C756 CLK3.n94 GND 0.24fF $ **FLOATING
C757 CLK3.t3 GND 0.07fF
C758 CLK3.n95 GND 0.09fF $ **FLOATING
C759 CLK3.n96 GND 0.02fF $ **FLOATING
C760 CLK3.n97 GND 0.02fF $ **FLOATING
C761 CLK3.n98 GND 0.02fF $ **FLOATING
C762 CLK3.n99 GND 0.13fF $ **FLOATING
C763 CLK3.n100 GND 0.02fF $ **FLOATING
C764 CLK3.n101 GND 0.02fF $ **FLOATING
C765 CLK3.n102 GND 0.02fF $ **FLOATING
C766 CLK3.t5 GND 0.07fF
C767 CLK3.n103 GND 0.08fF $ **FLOATING
C768 CLK3.n104 GND 0.02fF $ **FLOATING
C769 CLK3.n105 GND 0.02fF $ **FLOATING
C770 CLK3.n106 GND 0.02fF $ **FLOATING
C771 x2_bar.t3 GND 0.11fF
C772 x2_bar.t1 GND 0.29fF
C773 x2_bar.t2 GND 0.10fF
C774 x2_bar.n0 GND 0.97fF $ **FLOATING
C775 x2_bar.n1 GND 0.88fF $ **FLOATING
C776 x2_bar.t0 GND 0.09fF
C777 EESPFAL_4in_NAND_0/D_bar GND 0.25fF $ **FLOATING
C778 x2_bar.n2 GND 4.63fF $ **FLOATING
C779 EESPFAL_INV4_0/A GND 0.56fF $ **FLOATING
C780 x2.t1 GND 0.08fF
C781 x2.t3 GND 0.11fF
C782 x2.t2 GND 0.11fF
C783 x2.n0 GND 1.31fF $ **FLOATING
C784 x2.n1 GND 0.67fF $ **FLOATING
C785 x2.t0 GND 0.17fF
C786 EESPFAL_4in_NAND_0/D GND 1.29fF $ **FLOATING
C787 x2.n2 GND 4.70fF $ **FLOATING
C788 EESPFAL_INV4_0/A_bar GND 0.30fF $ **FLOATING
C789 x1_bar.t0 GND 0.31fF
C790 x1_bar.t2 GND 0.17fF
C791 x1_bar.n0 GND 1.63fF $ **FLOATING
C792 x1_bar.t3 GND 0.15fF
C793 x1_bar.t1 GND 0.19fF
C794 EESPFAL_4in_NAND_0/B_bar GND 0.56fF $ **FLOATING
C795 x1_bar.n1 GND 3.37fF $ **FLOATING
C796 EESPFAL_XOR_v3_1/A_bar GND 0.25fF $ **FLOATING
C797 x1.t0 GND 0.20fF
C798 x1.t2 GND 0.17fF
C799 x1.n0 GND 1.50fF $ **FLOATING
C800 x1.t1 GND 0.10fF
C801 x1.n1 GND 3.66fF $ **FLOATING
C802 x1.t3 GND 0.22fF
C803 EESPFAL_4in_NAND_0/B GND 1.80fF $ **FLOATING
C804 x1.n2 GND 2.78fF $ **FLOATING
C805 EESPFAL_XOR_v3_1/A GND 0.28fF $ **FLOATING
C806 EESPFAL_NAND_v3_1/A_bar.t8 GND 0.07fF
C807 EESPFAL_NAND_v3_1/A_bar.t4 GND 0.21fF
C808 EESPFAL_NAND_v3_1/A_bar.t3 GND 0.21fF
C809 EESPFAL_NAND_v3_1/A_bar.t5 GND 0.05fF
C810 EESPFAL_NAND_v3_1/A_bar.t0 GND 0.05fF
C811 EESPFAL_NAND_v3_1/A_bar.n0 GND 0.17fF $ **FLOATING
C812 EESPFAL_NAND_v3_1/A_bar.t6 GND 0.07fF
C813 EESPFAL_NAND_v3_1/A_bar.t9 GND 0.07fF
C814 EESPFAL_NAND_v3_1/A_bar.t7 GND 0.04fF
C815 EESPFAL_NAND_v3_1/A_bar.n1 GND 0.07fF $ **FLOATING
C816 EESPFAL_XOR_v3_0/OUT GND 0.01fF $ **FLOATING
C817 EESPFAL_NAND_v3_1/A_bar.n2 GND 0.04fF $ **FLOATING
C818 EESPFAL_NAND_v3_1/A_bar.t2 GND 0.05fF
C819 EESPFAL_NAND_v3_1/A_bar.t1 GND 0.05fF
C820 EESPFAL_NAND_v3_1/A_bar.n3 GND 0.15fF $ **FLOATING
C821 EESPFAL_NAND_v3_1/A_bar.n4 GND 0.22fF $ **FLOATING
C822 EESPFAL_NAND_v3_1/A_bar.n5 GND 0.22fF $ **FLOATING
C823 EESPFAL_NAND_v3_1/A_bar.n6 GND 0.76fF $ **FLOATING
C824 CLK2.t20 GND 0.02fF
C825 CLK2.t29 GND 0.02fF
C826 CLK2.n0 GND 0.05fF $ **FLOATING
C827 CLK2.t22 GND 0.03fF
C828 CLK2.t2 GND 0.02fF
C829 CLK2.n1 GND 0.05fF $ **FLOATING
C830 CLK2.n2 GND 0.01fF $ **FLOATING
C831 CLK2.n3 GND 0.01fF $ **FLOATING
C832 CLK2.n4 GND 0.01fF $ **FLOATING
C833 CLK2.n5 GND 0.07fF $ **FLOATING
C834 CLK2.t18 GND 0.03fF
C835 CLK2.t16 GND 0.02fF
C836 CLK2.t8 GND 0.02fF
C837 CLK2.n6 GND 0.05fF $ **FLOATING
C838 EESPFAL_NAND_v3_0/CLK GND 0.01fF $ **FLOATING
C839 CLK2.t10 GND 0.03fF
C840 CLK2.t1 GND 0.02fF
C841 CLK2.t26 GND 0.02fF
C842 CLK2.n7 GND 0.08fF $ **FLOATING
C843 CLK2.n8 GND 0.07fF $ **FLOATING
C844 CLK2.t24 GND 0.04fF
C845 CLK2.n9 GND 0.08fF $ **FLOATING
C846 CLK2.n10 GND 0.24fF $ **FLOATING
C847 CLK2.n11 GND 0.04fF $ **FLOATING
C848 CLK2.n12 GND 0.02fF $ **FLOATING
C849 CLK2.n13 GND 0.01fF $ **FLOATING
C850 CLK2.n14 GND 0.01fF $ **FLOATING
C851 CLK2.t14 GND 0.03fF
C852 CLK2.t12 GND 0.02fF
C853 CLK2.t6 GND 0.02fF
C854 CLK2.n15 GND 0.05fF $ **FLOATING
C855 EESPFAL_INV4_2/CLK GND 0.01fF $ **FLOATING
C856 CLK2.t4 GND 0.03fF
C857 CLK2.t0 GND 0.04fF
C858 CLK2.n16 GND 0.08fF $ **FLOATING
C859 CLK2.n17 GND 0.24fF $ **FLOATING
C860 CLK2.n18 GND 0.04fF $ **FLOATING
C861 CLK2.n19 GND 0.02fF $ **FLOATING
C862 CLK2.n20 GND 0.01fF $ **FLOATING
C863 CLK2.n21 GND 0.01fF $ **FLOATING
C864 CLK2.n22 GND 0.03fF $ **FLOATING
C865 CLK2.n23 GND 0.02fF $ **FLOATING
C866 CLK2.n24 GND 0.01fF $ **FLOATING
C867 CLK2.n25 GND 0.02fF $ **FLOATING
C868 CLK2.n26 GND 0.07fF $ **FLOATING
C869 CLK2.n27 GND 0.02fF $ **FLOATING
C870 CLK2.n28 GND 0.01fF $ **FLOATING
C871 CLK2.n29 GND 0.02fF $ **FLOATING
C872 CLK2.n30 GND 0.09fF $ **FLOATING
C873 CLK2.n31 GND 0.02fF $ **FLOATING
C874 CLK2.n32 GND 0.01fF $ **FLOATING
C875 CLK2.n33 GND 0.01fF $ **FLOATING
C876 CLK2.n34 GND 0.15fF $ **FLOATING
C877 CLK2.t3 GND 0.05fF
C878 CLK2.n35 GND 0.05fF $ **FLOATING
C879 CLK2.n36 GND 0.02fF $ **FLOATING
C880 CLK2.n37 GND 0.01fF $ **FLOATING
C881 CLK2.n38 GND 0.01fF $ **FLOATING
C882 CLK2.n39 GND 0.08fF $ **FLOATING
C883 CLK2.n40 GND 0.02fF $ **FLOATING
C884 CLK2.n41 GND 0.01fF $ **FLOATING
C885 CLK2.n42 GND 0.02fF $ **FLOATING
C886 CLK2.n43 GND 0.01fF $ **FLOATING
C887 CLK2.t5 GND 0.05fF
C888 CLK2.n44 GND 0.05fF $ **FLOATING
C889 CLK2.n45 GND 0.02fF $ **FLOATING
C890 CLK2.n46 GND 0.01fF $ **FLOATING
C891 CLK2.n47 GND 0.09fF $ **FLOATING
C892 CLK2.n48 GND 0.02fF $ **FLOATING
C893 CLK2.n49 GND 0.01fF $ **FLOATING
C894 CLK2.n50 GND 0.09fF $ **FLOATING
C895 CLK2.t11 GND 0.05fF
C896 CLK2.n51 GND 0.05fF $ **FLOATING
C897 CLK2.n52 GND 0.02fF $ **FLOATING
C898 CLK2.n53 GND 0.01fF $ **FLOATING
C899 CLK2.n54 GND 0.02fF $ **FLOATING
C900 CLK2.n55 GND 0.08fF $ **FLOATING
C901 CLK2.n56 GND 0.02fF $ **FLOATING
C902 CLK2.n57 GND 0.01fF $ **FLOATING
C903 CLK2.n58 GND 0.02fF $ **FLOATING
C904 CLK2.t13 GND 0.05fF
C905 CLK2.n59 GND 0.05fF $ **FLOATING
C906 CLK2.n60 GND 0.02fF $ **FLOATING
C907 CLK2.n61 GND 0.01fF $ **FLOATING
C908 CLK2.n62 GND 0.01fF $ **FLOATING
C909 CLK2.n63 GND 0.15fF $ **FLOATING
C910 CLK2.n64 GND 0.09fF $ **FLOATING
C911 CLK2.n65 GND 0.02fF $ **FLOATING
C912 CLK2.n66 GND 0.01fF $ **FLOATING
C913 CLK2.n67 GND 0.01fF $ **FLOATING
C914 CLK2.n68 GND 0.07fF $ **FLOATING
C915 CLK2.n69 GND 0.02fF $ **FLOATING
C916 CLK2.n70 GND 0.01fF $ **FLOATING
C917 CLK2.n71 GND 0.02fF $ **FLOATING
C918 CLK2.n72 GND 0.03fF $ **FLOATING
C919 CLK2.n73 GND 0.02fF $ **FLOATING
C920 CLK2.n74 GND 0.01fF $ **FLOATING
C921 CLK2.n75 GND 0.01fF $ **FLOATING
C922 CLK2.n76 GND 0.11fF $ **FLOATING
C923 CLK2.n77 GND 0.11fF $ **FLOATING
C924 CLK2.n78 GND 0.04fF $ **FLOATING
C925 CLK2.n79 GND 0.02fF $ **FLOATING
C926 CLK2.n80 GND 0.01fF $ **FLOATING
C927 CLK2.n81 GND 0.02fF $ **FLOATING
C928 CLK2.n82 GND 0.03fF $ **FLOATING
C929 CLK2.n83 GND 0.02fF $ **FLOATING
C930 CLK2.n84 GND 0.01fF $ **FLOATING
C931 CLK2.n85 GND 0.01fF $ **FLOATING
C932 CLK2.n86 GND 0.10fF $ **FLOATING
C933 CLK2.n87 GND 0.03fF $ **FLOATING
C934 CLK2.n88 GND 0.02fF $ **FLOATING
C935 CLK2.n89 GND 0.01fF $ **FLOATING
C936 CLK2.n90 GND 0.01fF $ **FLOATING
C937 CLK2.n91 GND 0.03fF $ **FLOATING
C938 CLK2.n92 GND 0.02fF $ **FLOATING
C939 CLK2.n93 GND 0.01fF $ **FLOATING
C940 CLK2.n94 GND 0.02fF $ **FLOATING
C941 CLK2.n95 GND 0.07fF $ **FLOATING
C942 CLK2.n96 GND 0.02fF $ **FLOATING
C943 CLK2.n97 GND 0.01fF $ **FLOATING
C944 CLK2.n98 GND 0.02fF $ **FLOATING
C945 CLK2.n99 GND 0.09fF $ **FLOATING
C946 CLK2.n100 GND 0.02fF $ **FLOATING
C947 CLK2.n101 GND 0.01fF $ **FLOATING
C948 CLK2.n102 GND 0.01fF $ **FLOATING
C949 CLK2.n103 GND 0.15fF $ **FLOATING
C950 CLK2.t9 GND 0.05fF
C951 CLK2.n104 GND 0.05fF $ **FLOATING
C952 CLK2.n105 GND 0.02fF $ **FLOATING
C953 CLK2.n106 GND 0.01fF $ **FLOATING
C954 CLK2.n107 GND 0.01fF $ **FLOATING
C955 CLK2.n108 GND 0.08fF $ **FLOATING
C956 CLK2.n109 GND 0.02fF $ **FLOATING
C957 CLK2.n110 GND 0.01fF $ **FLOATING
C958 CLK2.n111 GND 0.02fF $ **FLOATING
C959 CLK2.n112 GND 0.01fF $ **FLOATING
C960 CLK2.t7 GND 0.05fF
C961 CLK2.n113 GND 0.05fF $ **FLOATING
C962 CLK2.n114 GND 0.02fF $ **FLOATING
C963 CLK2.n115 GND 0.01fF $ **FLOATING
C964 CLK2.n116 GND 0.09fF $ **FLOATING
C965 CLK2.n117 GND 0.02fF $ **FLOATING
C966 CLK2.n118 GND 0.01fF $ **FLOATING
C967 CLK2.n119 GND 0.09fF $ **FLOATING
C968 CLK2.t15 GND 0.05fF
C969 CLK2.n120 GND 0.05fF $ **FLOATING
C970 CLK2.n121 GND 0.02fF $ **FLOATING
C971 CLK2.n122 GND 0.01fF $ **FLOATING
C972 CLK2.n123 GND 0.02fF $ **FLOATING
C973 CLK2.n124 GND 0.08fF $ **FLOATING
C974 CLK2.n125 GND 0.02fF $ **FLOATING
C975 CLK2.n126 GND 0.01fF $ **FLOATING
C976 CLK2.n127 GND 0.02fF $ **FLOATING
C977 CLK2.t17 GND 0.05fF
C978 CLK2.n128 GND 0.05fF $ **FLOATING
C979 CLK2.n129 GND 0.02fF $ **FLOATING
C980 CLK2.n130 GND 0.01fF $ **FLOATING
C981 CLK2.n131 GND 0.01fF $ **FLOATING
C982 CLK2.n132 GND 0.15fF $ **FLOATING
C983 CLK2.n133 GND 0.09fF $ **FLOATING
C984 CLK2.n134 GND 0.02fF $ **FLOATING
C985 CLK2.n135 GND 0.01fF $ **FLOATING
C986 CLK2.n136 GND 0.01fF $ **FLOATING
C987 CLK2.n137 GND 0.07fF $ **FLOATING
C988 CLK2.n138 GND 0.02fF $ **FLOATING
C989 CLK2.n139 GND 0.01fF $ **FLOATING
C990 CLK2.n140 GND 0.02fF $ **FLOATING
C991 CLK2.n141 GND 0.03fF $ **FLOATING
C992 CLK2.n142 GND 0.02fF $ **FLOATING
C993 CLK2.n143 GND 0.01fF $ **FLOATING
C994 CLK2.n144 GND 0.02fF $ **FLOATING
C995 CLK2.n145 GND 0.03fF $ **FLOATING
C996 CLK2.n146 GND 0.02fF $ **FLOATING
C997 CLK2.n147 GND 0.01fF $ **FLOATING
C998 CLK2.n148 GND 0.02fF $ **FLOATING
C999 CLK2.n149 GND 0.03fF $ **FLOATING
C1000 CLK2.n150 GND 0.02fF $ **FLOATING
C1001 CLK2.n151 GND 0.01fF $ **FLOATING
C1002 CLK2.n152 GND 0.02fF $ **FLOATING
C1003 CLK2.n153 GND 0.04fF $ **FLOATING
C1004 CLK2.n154 GND 0.02fF $ **FLOATING
C1005 CLK2.n155 GND 0.01fF $ **FLOATING
C1006 CLK2.n156 GND 0.01fF $ **FLOATING
C1007 CLK2.n157 GND 0.05fF $ **FLOATING
C1008 CLK2.n158 GND 0.01fF $ **FLOATING
C1009 CLK2.n159 GND 0.04fF $ **FLOATING
C1010 CLK2.n160 GND 0.01fF $ **FLOATING
C1011 CLK2.t25 GND 0.02fF
C1012 CLK2.n161 GND 0.05fF $ **FLOATING
C1013 CLK2.n162 GND 0.01fF $ **FLOATING
C1014 CLK2.n163 GND 0.06fF $ **FLOATING
C1015 CLK2.n164 GND 0.06fF $ **FLOATING
C1016 CLK2.n165 GND 0.01fF $ **FLOATING
C1017 CLK2.n166 GND 0.01fF $ **FLOATING
C1018 CLK2.n167 GND 0.05fF $ **FLOATING
C1019 CLK2.n168 GND 0.07fF $ **FLOATING
C1020 CLK2.n169 GND 0.05fF $ **FLOATING
C1021 CLK2.n170 GND 0.04fF $ **FLOATING
C1022 CLK2.n171 GND 0.02fF $ **FLOATING
C1023 CLK2.n172 GND 0.01fF $ **FLOATING
C1024 CLK2.n173 GND 0.01fF $ **FLOATING
C1025 CLK2.n174 GND 0.03fF $ **FLOATING
C1026 CLK2.n175 GND 0.02fF $ **FLOATING
C1027 CLK2.n176 GND 0.01fF $ **FLOATING
C1028 CLK2.n177 GND 0.02fF $ **FLOATING
C1029 CLK2.n178 GND 0.03fF $ **FLOATING
C1030 CLK2.n179 GND 0.02fF $ **FLOATING
C1031 CLK2.n180 GND 0.01fF $ **FLOATING
C1032 CLK2.n181 GND 0.02fF $ **FLOATING
C1033 CLK2.n182 GND 0.03fF $ **FLOATING
C1034 CLK2.n183 GND 0.02fF $ **FLOATING
C1035 CLK2.n184 GND 0.01fF $ **FLOATING
C1036 CLK2.n185 GND 0.02fF $ **FLOATING
C1037 CLK2.n186 GND 0.07fF $ **FLOATING
C1038 CLK2.n187 GND 0.02fF $ **FLOATING
C1039 CLK2.n188 GND 0.01fF $ **FLOATING
C1040 CLK2.n189 GND 0.02fF $ **FLOATING
C1041 CLK2.n190 GND 0.09fF $ **FLOATING
C1042 CLK2.n191 GND 0.02fF $ **FLOATING
C1043 CLK2.n192 GND 0.01fF $ **FLOATING
C1044 CLK2.n193 GND 0.01fF $ **FLOATING
C1045 CLK2.n194 GND 0.15fF $ **FLOATING
C1046 CLK2.t21 GND 0.05fF
C1047 CLK2.n195 GND 0.05fF $ **FLOATING
C1048 CLK2.n196 GND 0.02fF $ **FLOATING
C1049 CLK2.n197 GND 0.01fF $ **FLOATING
C1050 CLK2.n198 GND 0.01fF $ **FLOATING
C1051 CLK2.n199 GND 0.08fF $ **FLOATING
C1052 CLK2.n200 GND 0.02fF $ **FLOATING
C1053 CLK2.n201 GND 0.01fF $ **FLOATING
C1054 CLK2.n202 GND 0.02fF $ **FLOATING
C1055 CLK2.t19 GND 0.05fF
C1056 CLK2.n203 GND 0.05fF $ **FLOATING
C1057 CLK2.n204 GND 0.02fF $ **FLOATING
C1058 CLK2.n205 GND 0.01fF $ **FLOATING
C1059 CLK2.n206 GND 0.02fF $ **FLOATING
C1060 CLK2.n207 GND 0.09fF $ **FLOATING
C1061 CLK2.n208 GND 0.02fF $ **FLOATING
C1062 CLK2.n209 GND 0.01fF $ **FLOATING
C1063 CLK2.n210 GND 0.09fF $ **FLOATING
C1064 CLK2.t31 GND 0.03fF
C1065 CLK2.n211 GND 0.01fF $ **FLOATING
C1066 CLK2.n212 GND 0.01fF $ **FLOATING
C1067 CLK2.n213 GND 0.03fF $ **FLOATING
C1068 CLK2.n214 GND 0.02fF $ **FLOATING
C1069 CLK2.n215 GND 0.01fF $ **FLOATING
C1070 CLK2.t23 GND 0.02fF
C1071 CLK2.t27 GND 0.02fF
C1072 CLK2.n216 GND 0.08fF $ **FLOATING
C1073 CLK2.n217 GND 0.04fF $ **FLOATING
C1074 CLK2.n218 GND 0.02fF $ **FLOATING
C1075 CLK2.n219 GND 0.01fF $ **FLOATING
C1076 CLK2.n220 GND 0.07fF $ **FLOATING
C1077 CLK2.n221 GND 0.03fF $ **FLOATING
C1078 CLK2.n222 GND 0.02fF $ **FLOATING
C1079 CLK2.n223 GND 0.01fF $ **FLOATING
C1080 CLK2.n224 GND 0.04fF $ **FLOATING
C1081 CLK2.n225 GND 0.09fF $ **FLOATING
C1082 CLK2.n226 GND 0.01fF $ **FLOATING
C1083 CLK2.n227 GND 0.00fF $ **FLOATING
C1084 CLK2.n228 GND 0.01fF $ **FLOATING
C1085 CLK2.n229 GND 0.03fF $ **FLOATING
C1086 CLK2.n230 GND 0.02fF $ **FLOATING
C1087 CLK2.n231 GND 0.01fF $ **FLOATING
C1088 CLK2.n232 GND 0.02fF $ **FLOATING
C1089 CLK2.n233 GND 0.07fF $ **FLOATING
C1090 CLK2.n234 GND 0.02fF $ **FLOATING
C1091 CLK2.n235 GND 0.01fF $ **FLOATING
C1092 CLK2.n236 GND 0.02fF $ **FLOATING
C1093 CLK2.n237 GND 0.09fF $ **FLOATING
C1094 CLK2.n238 GND 0.02fF $ **FLOATING
C1095 CLK2.n239 GND 0.01fF $ **FLOATING
C1096 CLK2.n240 GND 0.01fF $ **FLOATING
C1097 CLK2.n241 GND 0.15fF $ **FLOATING
C1098 CLK2.t30 GND 0.05fF
C1099 CLK2.n242 GND 0.05fF $ **FLOATING
C1100 CLK2.n243 GND 0.02fF $ **FLOATING
C1101 CLK2.n244 GND 0.01fF $ **FLOATING
C1102 CLK2.n245 GND 0.01fF $ **FLOATING
C1103 CLK2.n246 GND 0.08fF $ **FLOATING
C1104 CLK2.n247 GND 0.02fF $ **FLOATING
C1105 CLK2.n248 GND 0.01fF $ **FLOATING
C1106 CLK2.n249 GND 0.02fF $ **FLOATING
C1107 CLK2.t28 GND 0.05fF
C1108 CLK2.n250 GND 0.05fF $ **FLOATING
C1109 CLK2.n251 GND 0.02fF $ **FLOATING
C1110 CLK2.n252 GND 0.01fF $ **FLOATING
C1111 CLK2.n253 GND 0.01fF $ **FLOATING
C1112 EESPFAL_NAND_v3_1/OUT_bar.t8 GND 0.04fF
C1113 EESPFAL_3in_NOR_v2_0/A_bar GND 0.53fF $ **FLOATING
C1114 EESPFAL_NAND_v3_1/OUT_bar.t4 GND 0.04fF
C1115 EESPFAL_NAND_v3_1/OUT_bar.t3 GND 0.04fF
C1116 EESPFAL_NAND_v3_1/OUT_bar.n0 GND 0.09fF $ **FLOATING
C1117 EESPFAL_NAND_v3_1/OUT_bar.t1 GND 0.14fF
C1118 EESPFAL_NAND_v3_1/OUT_bar.t2 GND 0.20fF
C1119 EESPFAL_NAND_v3_1/OUT_bar.n1 GND 0.20fF $ **FLOATING
C1120 EESPFAL_NAND_v3_1/OUT_bar.t5 GND 0.04fF
C1121 EESPFAL_NAND_v3_1/OUT_bar.t0 GND 0.04fF
C1122 EESPFAL_NAND_v3_1/OUT_bar.n2 GND 0.11fF $ **FLOATING
C1123 EESPFAL_NAND_v3_1/OUT_bar.n3 GND 0.09fF $ **FLOATING
C1124 EESPFAL_NAND_v3_1/OUT_bar.n4 GND 0.10fF $ **FLOATING
C1125 EESPFAL_NAND_v3_1/OUT_bar.t6 GND 0.05fF
C1126 EESPFAL_NAND_v3_1/OUT_bar.t9 GND 0.05fF
C1127 EESPFAL_NAND_v3_1/OUT_bar.t7 GND 0.03fF
C1128 EESPFAL_NAND_v3_1/OUT_bar.n5 GND 0.05fF $ **FLOATING
C1129 EESPFAL_NAND_v3_1/OUT_bar.n6 GND 0.04fF $ **FLOATING
C1130 EESPFAL_XOR_v3_0/OUT_bar GND 0.35fF $ **FLOATING
C1131 EESPFAL_NAND_v3_1/A.t9 GND 0.11fF
C1132 EESPFAL_NAND_v3_1/A.n0 GND 0.43fF $ **FLOATING
C1133 EESPFAL_NAND_v3_1/A.t3 GND 0.04fF
C1134 EESPFAL_NAND_v3_1/A.t4 GND 0.04fF
C1135 EESPFAL_NAND_v3_1/A.n1 GND 0.10fF $ **FLOATING
C1136 EESPFAL_NAND_v3_1/A.t5 GND 0.04fF
C1137 EESPFAL_NAND_v3_1/A.t2 GND 0.04fF
C1138 EESPFAL_NAND_v3_1/A.n2 GND 0.12fF $ **FLOATING
C1139 EESPFAL_NAND_v3_1/A.t1 GND 0.27fF
C1140 EESPFAL_NAND_v3_1/A.t0 GND 0.15fF
C1141 EESPFAL_NAND_v3_1/A.n3 GND 0.23fF $ **FLOATING
C1142 EESPFAL_NAND_v3_1/A.n4 GND 0.10fF $ **FLOATING
C1143 EESPFAL_NAND_v3_1/A.n5 GND 0.11fF $ **FLOATING
C1144 EESPFAL_NAND_v3_1/A.t6 GND 0.05fF
C1145 EESPFAL_NAND_v3_1/A.t8 GND 0.05fF
C1146 EESPFAL_NAND_v3_1/A.t7 GND 0.04fF
C1147 EESPFAL_NAND_v3_1/A.n6 GND 0.06fF $ **FLOATING
C1148 EESPFAL_NAND_v3_1/A.n7 GND 0.04fF $ **FLOATING
C1149 Dis1.t9 GND 0.16fF
C1150 Dis1.t4 GND 0.10fF
C1151 Dis1.n0 GND 0.40fF $ **FLOATING
C1152 Dis1.t7 GND 0.16fF
C1153 Dis1.t1 GND 0.10fF
C1154 Dis1.n1 GND 0.40fF $ **FLOATING
C1155 EESPFAL_INV4_0/Dis GND 0.45fF $ **FLOATING
C1156 Dis1.t6 GND 0.10fF
C1157 Dis1.n2 GND 0.66fF $ **FLOATING
C1158 Dis1.t2 GND 0.10fF
C1159 Dis1.n3 GND 0.21fF $ **FLOATING
C1160 EESPFAL_XOR_v3_1/Dis GND 0.13fF $ **FLOATING
C1161 Dis1.t3 GND 0.16fF
C1162 Dis1.t8 GND 0.10fF
C1163 Dis1.n4 GND 0.40fF $ **FLOATING
C1164 Dis1.t5 GND 0.10fF
C1165 Dis1.n5 GND 0.66fF $ **FLOATING
C1166 Dis1.t0 GND 0.10fF
C1167 Dis1.n6 GND 0.21fF $ **FLOATING
C1168 EESPFAL_XOR_v3_0/Dis GND 0.13fF $ **FLOATING
C1169 Dis1.n7 GND 0.43fF $ **FLOATING
C1170 Dis1.n8 GND 1.98fF $ **FLOATING
C1171 EESPFAL_4in_NAND_0/Dis GND 0.28fF $ **FLOATING
C1172 CLK1.t15 GND 0.02fF
C1173 CLK1.t46 GND 0.02fF
C1174 CLK1.n0 GND 0.06fF $ **FLOATING
C1175 CLK1.t24 GND 0.03fF
C1176 CLK1.n1 GND 0.02fF $ **FLOATING
C1177 CLK1.t11 GND 0.02fF
C1178 CLK1.t30 GND 0.02fF
C1179 CLK1.n2 GND 0.04fF $ **FLOATING
C1180 CLK1.n3 GND 0.01fF $ **FLOATING
C1181 CLK1.t7 GND 0.02fF
C1182 CLK1.t8 GND 0.02fF
C1183 CLK1.n4 GND 0.04fF $ **FLOATING
C1184 CLK1.n5 GND 0.01fF $ **FLOATING
C1185 CLK1.n6 GND 0.01fF $ **FLOATING
C1186 CLK1.t10 GND 0.05fF
C1187 CLK1.t22 GND 0.04fF
C1188 CLK1.t26 GND 0.03fF
C1189 EESPFAL_INV4_0/CLK GND 0.01fF $ **FLOATING
C1190 CLK1.t41 GND 0.02fF
C1191 CLK1.t28 GND 0.02fF
C1192 CLK1.n7 GND 0.06fF $ **FLOATING
C1193 CLK1.t43 GND 0.03fF
C1194 CLK1.t9 GND 0.04fF
C1195 CLK1.n8 GND 0.08fF $ **FLOATING
C1196 CLK1.n9 GND 0.26fF $ **FLOATING
C1197 CLK1.n10 GND 0.04fF $ **FLOATING
C1198 CLK1.n11 GND 0.02fF $ **FLOATING
C1199 CLK1.n12 GND 0.01fF $ **FLOATING
C1200 CLK1.n13 GND 0.02fF $ **FLOATING
C1201 CLK1.n14 GND 0.03fF $ **FLOATING
C1202 CLK1.n15 GND 0.02fF $ **FLOATING
C1203 CLK1.n16 GND 0.01fF $ **FLOATING
C1204 CLK1.n17 GND 0.02fF $ **FLOATING
C1205 CLK1.n18 GND 0.07fF $ **FLOATING
C1206 CLK1.n19 GND 0.02fF $ **FLOATING
C1207 CLK1.n20 GND 0.01fF $ **FLOATING
C1208 CLK1.n21 GND 0.02fF $ **FLOATING
C1209 CLK1.n22 GND 0.10fF $ **FLOATING
C1210 CLK1.n23 GND 0.02fF $ **FLOATING
C1211 CLK1.n24 GND 0.01fF $ **FLOATING
C1212 CLK1.n25 GND 0.01fF $ **FLOATING
C1213 CLK1.n26 GND 0.16fF $ **FLOATING
C1214 CLK1.t42 GND 0.05fF
C1215 CLK1.n27 GND 0.06fF $ **FLOATING
C1216 CLK1.n28 GND 0.02fF $ **FLOATING
C1217 CLK1.n29 GND 0.01fF $ **FLOATING
C1218 CLK1.n30 GND 0.01fF $ **FLOATING
C1219 CLK1.n31 GND 0.09fF $ **FLOATING
C1220 CLK1.n32 GND 0.02fF $ **FLOATING
C1221 CLK1.n33 GND 0.01fF $ **FLOATING
C1222 CLK1.n34 GND 0.02fF $ **FLOATING
C1223 CLK1.t40 GND 0.05fF
C1224 CLK1.n35 GND 0.05fF $ **FLOATING
C1225 CLK1.n36 GND 0.02fF $ **FLOATING
C1226 CLK1.n37 GND 0.01fF $ **FLOATING
C1227 CLK1.n38 GND 0.02fF $ **FLOATING
C1228 CLK1.n39 GND 0.10fF $ **FLOATING
C1229 CLK1.n40 GND 0.09fF $ **FLOATING
C1230 CLK1.n41 GND 0.02fF $ **FLOATING
C1231 CLK1.n42 GND 0.01fF $ **FLOATING
C1232 CLK1.t27 GND 0.05fF
C1233 CLK1.n43 GND 0.05fF $ **FLOATING
C1234 CLK1.n44 GND 0.02fF $ **FLOATING
C1235 CLK1.n45 GND 0.01fF $ **FLOATING
C1236 CLK1.n46 GND 0.01fF $ **FLOATING
C1237 CLK1.n47 GND 0.09fF $ **FLOATING
C1238 CLK1.n48 GND 0.02fF $ **FLOATING
C1239 CLK1.n49 GND 0.01fF $ **FLOATING
C1240 CLK1.n50 GND 0.02fF $ **FLOATING
C1241 CLK1.t25 GND 0.05fF
C1242 CLK1.n51 GND 0.06fF $ **FLOATING
C1243 CLK1.n52 GND 0.02fF $ **FLOATING
C1244 CLK1.n53 GND 0.01fF $ **FLOATING
C1245 CLK1.n54 GND 0.01fF $ **FLOATING
C1246 CLK1.n55 GND 0.16fF $ **FLOATING
C1247 CLK1.n56 GND 0.10fF $ **FLOATING
C1248 CLK1.n57 GND 0.02fF $ **FLOATING
C1249 CLK1.n58 GND 0.01fF $ **FLOATING
C1250 CLK1.n59 GND 0.01fF $ **FLOATING
C1251 CLK1.n60 GND 0.07fF $ **FLOATING
C1252 CLK1.n61 GND 0.02fF $ **FLOATING
C1253 CLK1.n62 GND 0.01fF $ **FLOATING
C1254 CLK1.n63 GND 0.02fF $ **FLOATING
C1255 CLK1.n64 GND 0.03fF $ **FLOATING
C1256 CLK1.n65 GND 0.02fF $ **FLOATING
C1257 CLK1.n66 GND 0.01fF $ **FLOATING
C1258 CLK1.n67 GND 0.02fF $ **FLOATING
C1259 CLK1.n68 GND 0.04fF $ **FLOATING
C1260 CLK1.n69 GND 0.02fF $ **FLOATING
C1261 CLK1.n70 GND 0.01fF $ **FLOATING
C1262 CLK1.n71 GND 0.02fF $ **FLOATING
C1263 CLK1.n72 GND 0.25fF $ **FLOATING
C1264 CLK1.n73 GND 0.09fF $ **FLOATING
C1265 CLK1.n74 GND 0.05fF $ **FLOATING
C1266 CLK1.n75 GND 0.14fF $ **FLOATING
C1267 CLK1.n76 GND 0.07fF $ **FLOATING
C1268 CLK1.n77 GND 0.22fF $ **FLOATING
C1269 CLK1.n78 GND 0.07fF $ **FLOATING
C1270 CLK1.n79 GND 0.04fF $ **FLOATING
C1271 CLK1.n80 GND 0.04fF $ **FLOATING
C1272 CLK1.n81 GND 0.03fF $ **FLOATING
C1273 CLK1.n82 GND 0.06fF $ **FLOATING
C1274 CLK1.n83 GND 0.04fF $ **FLOATING
C1275 CLK1.n84 GND 0.04fF $ **FLOATING
C1276 CLK1.n85 GND 0.04fF $ **FLOATING
C1277 CLK1.n86 GND 0.05fF $ **FLOATING
C1278 CLK1.n87 GND 0.04fF $ **FLOATING
C1279 CLK1.n88 GND 0.04fF $ **FLOATING
C1280 CLK1.n89 GND 0.04fF $ **FLOATING
C1281 CLK1.n90 GND 0.05fF $ **FLOATING
C1282 CLK1.n91 GND 0.04fF $ **FLOATING
C1283 CLK1.n92 GND 0.04fF $ **FLOATING
C1284 CLK1.n93 GND 0.03fF $ **FLOATING
C1285 CLK1.t5 GND 0.03fF
C1286 CLK1.t1 GND 0.03fF
C1287 CLK1.t4 GND 0.02fF
C1288 CLK1.t38 GND 0.02fF
C1289 CLK1.n94 GND 0.06fF $ **FLOATING
C1290 CLK1.t3 GND 0.02fF
C1291 CLK1.t20 GND 0.02fF
C1292 CLK1.n95 GND 0.06fF $ **FLOATING
C1293 EESPFAL_4in_NAND_0/CLK GND 0.02fF $ **FLOATING
C1294 CLK1.n96 GND 0.17fF $ **FLOATING
C1295 CLK1.n97 GND 0.04fF $ **FLOATING
C1296 CLK1.n98 GND 0.04fF $ **FLOATING
C1297 CLK1.t37 GND 0.03fF
C1298 CLK1.t18 GND 0.03fF
C1299 CLK1.t29 GND 0.02fF
C1300 CLK1.t6 GND 0.02fF
C1301 CLK1.n99 GND 0.10fF $ **FLOATING
C1302 CLK1.t21 GND 0.02fF
C1303 CLK1.t32 GND 0.02fF
C1304 CLK1.n100 GND 0.09fF $ **FLOATING
C1305 CLK1.t39 GND 0.02fF
C1306 CLK1.t44 GND 0.02fF
C1307 CLK1.n101 GND 0.10fF $ **FLOATING
C1308 CLK1.n102 GND 0.08fF $ **FLOATING
C1309 CLK1.n103 GND 0.04fF $ **FLOATING
C1310 CLK1.n104 GND 0.04fF $ **FLOATING
C1311 CLK1.n105 GND 0.16fF $ **FLOATING
C1312 CLK1.n106 GND 0.06fF $ **FLOATING
C1313 CLK1.n107 GND 0.04fF $ **FLOATING
C1314 CLK1.n108 GND 0.04fF $ **FLOATING
C1315 CLK1.n109 GND 0.10fF $ **FLOATING
C1316 CLK1.n110 GND 0.13fF $ **FLOATING
C1317 CLK1.n111 GND 0.05fF $ **FLOATING
C1318 CLK1.n112 GND 0.04fF $ **FLOATING
C1319 CLK1.n113 GND 0.04fF $ **FLOATING
C1320 CLK1.n114 GND 0.03fF $ **FLOATING
C1321 CLK1.n115 GND 0.05fF $ **FLOATING
C1322 CLK1.n116 GND 0.04fF $ **FLOATING
C1323 CLK1.n117 GND 0.04fF $ **FLOATING
C1324 CLK1.n118 GND 0.03fF $ **FLOATING
C1325 CLK1.n119 GND 0.12fF $ **FLOATING
C1326 CLK1.n120 GND 0.05fF $ **FLOATING
C1327 CLK1.n121 GND 0.04fF $ **FLOATING
C1328 CLK1.n122 GND 0.04fF $ **FLOATING
C1329 CLK1.n123 GND 0.04fF $ **FLOATING
C1330 CLK1.n124 GND 0.05fF $ **FLOATING
C1331 CLK1.n125 GND 0.04fF $ **FLOATING
C1332 CLK1.n126 GND 0.04fF $ **FLOATING
C1333 CLK1.n127 GND 0.02fF $ **FLOATING
C1334 CLK1.n128 GND 0.13fF $ **FLOATING
C1335 CLK1.n129 GND 0.05fF $ **FLOATING
C1336 CLK1.n130 GND 0.04fF $ **FLOATING
C1337 CLK1.n131 GND 0.04fF $ **FLOATING
C1338 CLK1.n132 GND 0.04fF $ **FLOATING
C1339 CLK1.n133 GND 0.05fF $ **FLOATING
C1340 CLK1.n134 GND 0.04fF $ **FLOATING
C1341 CLK1.n135 GND 0.04fF $ **FLOATING
C1342 CLK1.n136 GND 0.04fF $ **FLOATING
C1343 CLK1.n137 GND 0.14fF $ **FLOATING
C1344 CLK1.n138 GND 0.04fF $ **FLOATING
C1345 CLK1.n139 GND 0.04fF $ **FLOATING
C1346 CLK1.n140 GND 0.04fF $ **FLOATING
C1347 CLK1.n141 GND 0.19fF $ **FLOATING
C1348 CLK1.n142 GND 0.04fF $ **FLOATING
C1349 CLK1.n143 GND 0.04fF $ **FLOATING
C1350 CLK1.n144 GND 0.03fF $ **FLOATING
C1351 CLK1.n145 GND 0.33fF $ **FLOATING
C1352 CLK1.t17 GND 0.09fF
C1353 CLK1.n146 GND 0.11fF $ **FLOATING
C1354 CLK1.n147 GND 0.04fF $ **FLOATING
C1355 CLK1.n148 GND 0.04fF $ **FLOATING
C1356 CLK1.n149 GND 0.04fF $ **FLOATING
C1357 CLK1.n150 GND 0.04fF $ **FLOATING
C1358 CLK1.n151 GND 0.04fF $ **FLOATING
C1359 CLK1.t19 GND 0.09fF
C1360 CLK1.n152 GND 0.10fF $ **FLOATING
C1361 CLK1.n153 GND 0.04fF $ **FLOATING
C1362 CLK1.n154 GND 0.04fF $ **FLOATING
C1363 CLK1.n155 GND 0.17fF $ **FLOATING
C1364 CLK1.n156 GND 0.04fF $ **FLOATING
C1365 CLK1.n157 GND 0.04fF $ **FLOATING
C1366 CLK1.n158 GND 0.20fF $ **FLOATING
C1367 CLK1.t2 GND 0.09fF
C1368 CLK1.n159 GND 0.10fF $ **FLOATING
C1369 CLK1.n160 GND 0.04fF $ **FLOATING
C1370 CLK1.n161 GND 0.04fF $ **FLOATING
C1371 CLK1.n162 GND 0.04fF $ **FLOATING
C1372 CLK1.n163 GND 0.17fF $ **FLOATING
C1373 CLK1.n164 GND 0.04fF $ **FLOATING
C1374 CLK1.n165 GND 0.04fF $ **FLOATING
C1375 CLK1.n166 GND 0.04fF $ **FLOATING
C1376 CLK1.t0 GND 0.09fF
C1377 CLK1.n167 GND 0.11fF $ **FLOATING
C1378 CLK1.n168 GND 0.04fF $ **FLOATING
C1379 CLK1.n169 GND 0.04fF $ **FLOATING
C1380 CLK1.n170 GND 0.04fF $ **FLOATING
C1381 CLK1.n171 GND 0.33fF $ **FLOATING
C1382 CLK1.n172 GND 0.19fF $ **FLOATING
C1383 CLK1.n173 GND 0.04fF $ **FLOATING
C1384 CLK1.n174 GND 0.04fF $ **FLOATING
C1385 CLK1.n175 GND 0.03fF $ **FLOATING
C1386 CLK1.n176 GND 0.14fF $ **FLOATING
C1387 CLK1.n177 GND 0.04fF $ **FLOATING
C1388 CLK1.n178 GND 0.04fF $ **FLOATING
C1389 CLK1.n179 GND 0.04fF $ **FLOATING
C1390 CLK1.n180 GND 0.05fF $ **FLOATING
C1391 CLK1.n181 GND 0.04fF $ **FLOATING
C1392 CLK1.n182 GND 0.04fF $ **FLOATING
C1393 CLK1.n183 GND 0.04fF $ **FLOATING
C1394 CLK1.n184 GND 0.05fF $ **FLOATING
C1395 CLK1.n185 GND 0.04fF $ **FLOATING
C1396 CLK1.n186 GND 0.04fF $ **FLOATING
C1397 CLK1.n187 GND 0.04fF $ **FLOATING
C1398 CLK1.n188 GND 0.05fF $ **FLOATING
C1399 CLK1.n189 GND 0.04fF $ **FLOATING
C1400 CLK1.n190 GND 0.04fF $ **FLOATING
C1401 CLK1.n191 GND 0.04fF $ **FLOATING
C1402 CLK1.n192 GND 0.05fF $ **FLOATING
C1403 CLK1.n193 GND 0.04fF $ **FLOATING
C1404 CLK1.n194 GND 0.04fF $ **FLOATING
C1405 CLK1.n195 GND 0.04fF $ **FLOATING
C1406 CLK1.n196 GND 0.05fF $ **FLOATING
C1407 CLK1.n197 GND 0.05fF $ **FLOATING
C1408 CLK1.n198 GND 0.01fF $ **FLOATING
C1409 CLK1.n199 GND 0.01fF $ **FLOATING
C1410 CLK1.n200 GND 0.04fF $ **FLOATING
C1411 CLK1.n201 GND 0.05fF $ **FLOATING
C1412 CLK1.n202 GND 0.01fF $ **FLOATING
C1413 CLK1.n203 GND 0.01fF $ **FLOATING
C1414 CLK1.n204 GND 0.04fF $ **FLOATING
C1415 CLK1.t12 GND 0.04fF
C1416 CLK1.t36 GND 0.03fF
C1417 CLK1.n205 GND 0.09fF $ **FLOATING
C1418 CLK1.n206 GND 0.02fF $ **FLOATING
C1419 CLK1.t52 GND 0.02fF
C1420 CLK1.t34 GND 0.02fF
C1421 CLK1.n207 GND 0.06fF $ **FLOATING
C1422 CLK1.t50 GND 0.03fF
C1423 CLK1.t13 GND 0.04fF
C1424 CLK1.n208 GND 0.08fF $ **FLOATING
C1425 CLK1.n209 GND 0.26fF $ **FLOATING
C1426 CLK1.n210 GND 0.04fF $ **FLOATING
C1427 CLK1.n211 GND 0.02fF $ **FLOATING
C1428 CLK1.n212 GND 0.01fF $ **FLOATING
C1429 CLK1.n213 GND 0.02fF $ **FLOATING
C1430 CLK1.n214 GND 0.03fF $ **FLOATING
C1431 CLK1.n215 GND 0.02fF $ **FLOATING
C1432 CLK1.n216 GND 0.01fF $ **FLOATING
C1433 CLK1.n217 GND 0.02fF $ **FLOATING
C1434 CLK1.n218 GND 0.07fF $ **FLOATING
C1435 CLK1.n219 GND 0.02fF $ **FLOATING
C1436 CLK1.n220 GND 0.01fF $ **FLOATING
C1437 CLK1.n221 GND 0.02fF $ **FLOATING
C1438 CLK1.n222 GND 0.10fF $ **FLOATING
C1439 CLK1.n223 GND 0.02fF $ **FLOATING
C1440 CLK1.n224 GND 0.01fF $ **FLOATING
C1441 CLK1.n225 GND 0.01fF $ **FLOATING
C1442 CLK1.n226 GND 0.16fF $ **FLOATING
C1443 CLK1.t49 GND 0.05fF
C1444 CLK1.n227 GND 0.06fF $ **FLOATING
C1445 CLK1.n228 GND 0.02fF $ **FLOATING
C1446 CLK1.n229 GND 0.01fF $ **FLOATING
C1447 CLK1.n230 GND 0.01fF $ **FLOATING
C1448 CLK1.n231 GND 0.09fF $ **FLOATING
C1449 CLK1.n232 GND 0.02fF $ **FLOATING
C1450 CLK1.n233 GND 0.01fF $ **FLOATING
C1451 CLK1.n234 GND 0.02fF $ **FLOATING
C1452 CLK1.t51 GND 0.05fF
C1453 CLK1.n235 GND 0.05fF $ **FLOATING
C1454 CLK1.n236 GND 0.02fF $ **FLOATING
C1455 CLK1.n237 GND 0.01fF $ **FLOATING
C1456 CLK1.n238 GND 0.02fF $ **FLOATING
C1457 CLK1.n239 GND 0.10fF $ **FLOATING
C1458 CLK1.n240 GND 0.01fF $ **FLOATING
C1459 CLK1.t33 GND 0.05fF
C1460 CLK1.n241 GND 0.05fF $ **FLOATING
C1461 CLK1.n242 GND 0.02fF $ **FLOATING
C1462 CLK1.n243 GND 0.01fF $ **FLOATING
C1463 CLK1.n244 GND 0.01fF $ **FLOATING
C1464 CLK1.n245 GND 0.09fF $ **FLOATING
C1465 CLK1.n246 GND 0.02fF $ **FLOATING
C1466 CLK1.n247 GND 0.01fF $ **FLOATING
C1467 CLK1.n248 GND 0.02fF $ **FLOATING
C1468 CLK1.t35 GND 0.05fF
C1469 CLK1.n249 GND 0.06fF $ **FLOATING
C1470 CLK1.n250 GND 0.02fF $ **FLOATING
C1471 CLK1.n251 GND 0.01fF $ **FLOATING
C1472 CLK1.n252 GND 0.01fF $ **FLOATING
C1473 CLK1.n253 GND 0.16fF $ **FLOATING
C1474 CLK1.n254 GND 0.10fF $ **FLOATING
C1475 CLK1.n255 GND 0.02fF $ **FLOATING
C1476 CLK1.n256 GND 0.01fF $ **FLOATING
C1477 CLK1.n257 GND 0.01fF $ **FLOATING
C1478 CLK1.n258 GND 0.07fF $ **FLOATING
C1479 CLK1.n259 GND 0.02fF $ **FLOATING
C1480 CLK1.n260 GND 0.01fF $ **FLOATING
C1481 CLK1.n261 GND 0.02fF $ **FLOATING
C1482 CLK1.n262 GND 0.03fF $ **FLOATING
C1483 CLK1.n263 GND 0.02fF $ **FLOATING
C1484 CLK1.n264 GND 0.01fF $ **FLOATING
C1485 CLK1.n265 GND 0.02fF $ **FLOATING
C1486 CLK1.n266 GND 0.04fF $ **FLOATING
C1487 CLK1.n267 GND 0.02fF $ **FLOATING
C1488 CLK1.n268 GND 0.01fF $ **FLOATING
C1489 CLK1.n269 GND 0.02fF $ **FLOATING
C1490 CLK1.n270 GND 0.25fF $ **FLOATING
C1491 CLK1.n271 GND 0.09fF $ **FLOATING
C1492 CLK1.n272 GND 0.06fF $ **FLOATING
C1493 CLK1.n273 GND 0.11fF $ **FLOATING
C1494 CLK1.n274 GND 0.06fF $ **FLOATING
C1495 CLK1.n275 GND 0.04fF $ **FLOATING
C1496 CLK1.n276 GND 0.02fF $ **FLOATING
C1497 CLK1.n277 GND 0.01fF $ **FLOATING
C1498 CLK1.n278 GND 0.02fF $ **FLOATING
C1499 CLK1.n279 GND 0.03fF $ **FLOATING
C1500 CLK1.n280 GND 0.02fF $ **FLOATING
C1501 CLK1.n281 GND 0.01fF $ **FLOATING
C1502 CLK1.n282 GND 0.02fF $ **FLOATING
C1503 CLK1.n283 GND 0.03fF $ **FLOATING
C1504 CLK1.n284 GND 0.02fF $ **FLOATING
C1505 CLK1.n285 GND 0.01fF $ **FLOATING
C1506 CLK1.n286 GND 0.01fF $ **FLOATING
C1507 CLK1.n287 GND 0.04fF $ **FLOATING
C1508 CLK1.n288 GND 0.03fF $ **FLOATING
C1509 CLK1.n289 GND 0.02fF $ **FLOATING
C1510 CLK1.n290 GND 0.01fF $ **FLOATING
C1511 CLK1.n291 GND 0.01fF $ **FLOATING
C1512 CLK1.n292 GND 0.03fF $ **FLOATING
C1513 CLK1.n293 GND 0.02fF $ **FLOATING
C1514 CLK1.n294 GND 0.01fF $ **FLOATING
C1515 CLK1.n295 GND 0.02fF $ **FLOATING
C1516 CLK1.n296 GND 0.03fF $ **FLOATING
C1517 CLK1.n297 GND 0.02fF $ **FLOATING
C1518 CLK1.n298 GND 0.01fF $ **FLOATING
C1519 CLK1.n299 GND 0.02fF $ **FLOATING
C1520 CLK1.n300 GND 0.03fF $ **FLOATING
C1521 CLK1.n301 GND 0.02fF $ **FLOATING
C1522 CLK1.n302 GND 0.01fF $ **FLOATING
C1523 CLK1.n303 GND 0.02fF $ **FLOATING
C1524 CLK1.n304 GND 0.07fF $ **FLOATING
C1525 CLK1.n305 GND 0.02fF $ **FLOATING
C1526 CLK1.n306 GND 0.01fF $ **FLOATING
C1527 CLK1.n307 GND 0.02fF $ **FLOATING
C1528 CLK1.n308 GND 0.10fF $ **FLOATING
C1529 CLK1.n309 GND 0.02fF $ **FLOATING
C1530 CLK1.n310 GND 0.01fF $ **FLOATING
C1531 CLK1.n311 GND 0.01fF $ **FLOATING
C1532 CLK1.n312 GND 0.16fF $ **FLOATING
C1533 CLK1.t23 GND 0.05fF
C1534 CLK1.n313 GND 0.06fF $ **FLOATING
C1535 CLK1.n314 GND 0.02fF $ **FLOATING
C1536 CLK1.n315 GND 0.01fF $ **FLOATING
C1537 CLK1.n316 GND 0.01fF $ **FLOATING
C1538 CLK1.n317 GND 0.09fF $ **FLOATING
C1539 CLK1.n318 GND 0.02fF $ **FLOATING
C1540 CLK1.n319 GND 0.01fF $ **FLOATING
C1541 CLK1.n320 GND 0.02fF $ **FLOATING
C1542 CLK1.t14 GND 0.05fF
C1543 CLK1.n321 GND 0.05fF $ **FLOATING
C1544 CLK1.n322 GND 0.02fF $ **FLOATING
C1545 CLK1.n323 GND 0.01fF $ **FLOATING
C1546 CLK1.n324 GND 0.02fF $ **FLOATING
C1547 CLK1.n325 GND 0.09fF $ **FLOATING
C1548 CLK1.n326 GND 0.02fF $ **FLOATING
C1549 CLK1.n327 GND 0.01fF $ **FLOATING
C1550 CLK1.n328 GND 0.10fF $ **FLOATING
C1551 CLK1.t48 GND 0.03fF
C1552 CLK1.t31 GND 0.02fF
C1553 CLK1.t16 GND 0.02fF
C1554 CLK1.n329 GND 0.09fF $ **FLOATING
C1555 CLK1.n330 GND 0.11fF $ **FLOATING
C1556 CLK1.n331 GND 0.03fF $ **FLOATING
C1557 CLK1.n332 GND 0.04fF $ **FLOATING
C1558 CLK1.n333 GND 0.02fF $ **FLOATING
C1559 CLK1.n334 GND 0.01fF $ **FLOATING
C1560 CLK1.n335 GND 0.02fF $ **FLOATING
C1561 CLK1.n336 GND 0.03fF $ **FLOATING
C1562 CLK1.n337 GND 0.02fF $ **FLOATING
C1563 CLK1.n338 GND 0.01fF $ **FLOATING
C1564 CLK1.n339 GND 0.02fF $ **FLOATING
C1565 CLK1.n340 GND 0.03fF $ **FLOATING
C1566 CLK1.n341 GND 0.02fF $ **FLOATING
C1567 CLK1.n342 GND 0.01fF $ **FLOATING
C1568 CLK1.n343 GND 0.01fF $ **FLOATING
C1569 CLK1.n344 GND 0.10fF $ **FLOATING
C1570 CLK1.n345 GND 0.03fF $ **FLOATING
C1571 CLK1.n346 GND 0.02fF $ **FLOATING
C1572 CLK1.n347 GND 0.01fF $ **FLOATING
C1573 CLK1.n348 GND 0.01fF $ **FLOATING
C1574 CLK1.n349 GND 0.03fF $ **FLOATING
C1575 CLK1.n350 GND 0.02fF $ **FLOATING
C1576 CLK1.n351 GND 0.01fF $ **FLOATING
C1577 CLK1.n352 GND 0.02fF $ **FLOATING
C1578 CLK1.n353 GND 0.03fF $ **FLOATING
C1579 CLK1.n354 GND 0.02fF $ **FLOATING
C1580 CLK1.n355 GND 0.01fF $ **FLOATING
C1581 CLK1.n356 GND 0.02fF $ **FLOATING
C1582 CLK1.n357 GND 0.03fF $ **FLOATING
C1583 CLK1.n358 GND 0.02fF $ **FLOATING
C1584 CLK1.n359 GND 0.01fF $ **FLOATING
C1585 CLK1.n360 GND 0.02fF $ **FLOATING
C1586 CLK1.n361 GND 0.07fF $ **FLOATING
C1587 CLK1.n362 GND 0.02fF $ **FLOATING
C1588 CLK1.n363 GND 0.01fF $ **FLOATING
C1589 CLK1.n364 GND 0.02fF $ **FLOATING
C1590 CLK1.n365 GND 0.10fF $ **FLOATING
C1591 CLK1.n366 GND 0.02fF $ **FLOATING
C1592 CLK1.n367 GND 0.01fF $ **FLOATING
C1593 CLK1.n368 GND 0.01fF $ **FLOATING
C1594 CLK1.n369 GND 0.16fF $ **FLOATING
C1595 CLK1.t47 GND 0.05fF
C1596 CLK1.n370 GND 0.06fF $ **FLOATING
C1597 CLK1.n371 GND 0.02fF $ **FLOATING
C1598 CLK1.n372 GND 0.01fF $ **FLOATING
C1599 CLK1.n373 GND 0.01fF $ **FLOATING
C1600 CLK1.n374 GND 0.09fF $ **FLOATING
C1601 CLK1.n375 GND 0.02fF $ **FLOATING
C1602 CLK1.n376 GND 0.01fF $ **FLOATING
C1603 CLK1.n377 GND 0.02fF $ **FLOATING
C1604 CLK1.t45 GND 0.05fF
C1605 CLK1.n378 GND 0.05fF $ **FLOATING
C1606 CLK1.n379 GND 0.02fF $ **FLOATING
C1607 CLK1.n380 GND 0.01fF $ **FLOATING
C1608 CLK1.n381 GND 0.01fF $ **FLOATING
C1609 EESPFAL_XOR_v3_0/CLK GND 0.01fF $ **FLOATING
C1610 x3.t1 GND 0.27fF
C1611 x3.t2 GND 0.26fF
C1612 x3.t0 GND 0.23fF
C1613 x3.n0 GND 1.98fF $ **FLOATING
C1614 EESPFAL_4in_NAND_0/A_bar GND 0.78fF $ **FLOATING
C1615 EESPFAL_INV4_2/OUT GND 0.23fF $ **FLOATING
C1616 EESPFAL_3in_NOR_v2_0/C_bar.t8 GND 0.03fF
C1617 EESPFAL_3in_NOR_v2_0/C_bar.n0 GND 0.63fF $ **FLOATING
C1618 EESPFAL_3in_NOR_v2_0/C_bar.t4 GND 0.04fF
C1619 EESPFAL_3in_NOR_v2_0/C_bar.t2 GND 0.04fF
C1620 EESPFAL_3in_NOR_v2_0/C_bar.n1 GND 0.11fF $ **FLOATING
C1621 EESPFAL_3in_NOR_v2_0/C_bar.t3 GND 0.04fF
C1622 EESPFAL_3in_NOR_v2_0/C_bar.t1 GND 0.04fF
C1623 EESPFAL_3in_NOR_v2_0/C_bar.n2 GND 0.13fF $ **FLOATING
C1624 EESPFAL_3in_NOR_v2_0/C_bar.t0 GND 0.25fF
C1625 EESPFAL_3in_NOR_v2_0/C_bar.n3 GND 0.17fF $ **FLOATING
C1626 EESPFAL_3in_NOR_v2_0/C_bar.n4 GND 0.12fF $ **FLOATING
C1627 EESPFAL_3in_NOR_v2_0/C_bar.t6 GND 0.06fF
C1628 EESPFAL_3in_NOR_v2_0/C_bar.t7 GND 0.05fF
C1629 EESPFAL_3in_NOR_v2_0/C_bar.t5 GND 0.04fF
C1630 EESPFAL_3in_NOR_v2_0/C_bar.n5 GND 0.06fF $ **FLOATING
C1631 EESPFAL_3in_NOR_v2_0/C_bar.n6 GND 0.04fF $ **FLOATING
C1632 EESPFAL_3in_NOR_v2_0/C.t6 GND 0.05fF
C1633 EESPFAL_3in_NOR_v2_0/C.t3 GND 0.04fF
C1634 EESPFAL_3in_NOR_v2_0/C.t2 GND 0.04fF
C1635 EESPFAL_3in_NOR_v2_0/C.n0 GND 0.12fF $ **FLOATING
C1636 EESPFAL_3in_NOR_v2_0/C.t4 GND 0.04fF
C1637 EESPFAL_3in_NOR_v2_0/C.t0 GND 0.04fF
C1638 EESPFAL_3in_NOR_v2_0/C.n1 GND 0.13fF $ **FLOATING
C1639 EESPFAL_3in_NOR_v2_0/C.t8 GND 0.06fF
C1640 EESPFAL_3in_NOR_v2_0/C.t7 GND 0.06fF
C1641 EESPFAL_3in_NOR_v2_0/C.t5 GND 0.03fF
C1642 EESPFAL_3in_NOR_v2_0/C.n2 GND 0.06fF $ **FLOATING
C1643 EESPFAL_INV4_2/OUT_bar GND 0.01fF $ **FLOATING
C1644 EESPFAL_3in_NOR_v2_0/C.n3 GND 0.03fF $ **FLOATING
C1645 EESPFAL_3in_NOR_v2_0/C.n4 GND 0.11fF $ **FLOATING
C1646 EESPFAL_3in_NOR_v2_0/C.n5 GND 0.11fF $ **FLOATING
C1647 EESPFAL_3in_NOR_v2_0/C.t1 GND 0.17fF
C1648 EESPFAL_3in_NOR_v2_0/C.n6 GND 0.18fF $ **FLOATING
C1649 EESPFAL_3in_NOR_v2_0/C.n7 GND 0.78fF $ **FLOATING
.ends

