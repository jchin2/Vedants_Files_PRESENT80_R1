magic
tech sky130A
timestamp 1667077063
<< nwell >>
rect -1240 645 -200 740
rect -925 450 -515 645
<< nmos >>
rect -1155 30 -1140 180
rect -1080 30 -1065 180
rect -1005 30 -990 180
rect -840 30 -825 180
rect -765 30 -750 180
rect -690 30 -675 180
rect -615 30 -600 180
rect -450 30 -435 180
rect -375 30 -360 180
rect -300 30 -285 180
<< pmos >>
rect -840 475 -825 625
rect -765 475 -750 625
rect -690 475 -675 625
rect -615 475 -600 625
<< ndiff >>
rect -1215 145 -1155 180
rect -1215 125 -1195 145
rect -1175 125 -1155 145
rect -1215 105 -1155 125
rect -1215 85 -1195 105
rect -1175 85 -1155 105
rect -1215 65 -1155 85
rect -1215 45 -1195 65
rect -1175 45 -1155 65
rect -1215 30 -1155 45
rect -1140 145 -1080 180
rect -1140 125 -1120 145
rect -1100 125 -1080 145
rect -1140 105 -1080 125
rect -1140 85 -1120 105
rect -1100 85 -1080 105
rect -1140 65 -1080 85
rect -1140 45 -1120 65
rect -1100 45 -1080 65
rect -1140 30 -1080 45
rect -1065 145 -1005 180
rect -1065 125 -1045 145
rect -1025 125 -1005 145
rect -1065 105 -1005 125
rect -1065 85 -1045 105
rect -1025 85 -1005 105
rect -1065 65 -1005 85
rect -1065 45 -1045 65
rect -1025 45 -1005 65
rect -1065 30 -1005 45
rect -990 145 -930 180
rect -990 125 -970 145
rect -950 125 -930 145
rect -990 105 -930 125
rect -990 85 -970 105
rect -950 85 -930 105
rect -990 65 -930 85
rect -990 45 -970 65
rect -950 45 -930 65
rect -990 30 -930 45
rect -900 145 -840 180
rect -900 125 -880 145
rect -860 125 -840 145
rect -900 105 -840 125
rect -900 85 -880 105
rect -860 85 -840 105
rect -900 65 -840 85
rect -900 45 -880 65
rect -860 45 -840 65
rect -900 30 -840 45
rect -825 145 -765 180
rect -825 125 -805 145
rect -785 125 -765 145
rect -825 105 -765 125
rect -825 85 -805 105
rect -785 85 -765 105
rect -825 65 -765 85
rect -825 45 -805 65
rect -785 45 -765 65
rect -825 30 -765 45
rect -750 145 -690 180
rect -750 125 -730 145
rect -710 125 -690 145
rect -750 105 -690 125
rect -750 85 -730 105
rect -710 85 -690 105
rect -750 65 -690 85
rect -750 45 -730 65
rect -710 45 -690 65
rect -750 30 -690 45
rect -675 145 -615 180
rect -675 125 -655 145
rect -635 125 -615 145
rect -675 105 -615 125
rect -675 85 -655 105
rect -635 85 -615 105
rect -675 65 -615 85
rect -675 45 -655 65
rect -635 45 -615 65
rect -675 30 -615 45
rect -600 145 -540 180
rect -600 125 -580 145
rect -560 125 -540 145
rect -600 105 -540 125
rect -600 85 -580 105
rect -560 85 -540 105
rect -600 65 -540 85
rect -600 45 -580 65
rect -560 45 -540 65
rect -600 30 -540 45
rect -510 145 -450 180
rect -510 125 -490 145
rect -470 125 -450 145
rect -510 105 -450 125
rect -510 85 -490 105
rect -470 85 -450 105
rect -510 65 -450 85
rect -510 45 -490 65
rect -470 45 -450 65
rect -510 30 -450 45
rect -435 30 -375 180
rect -360 30 -300 180
rect -285 145 -225 180
rect -285 125 -265 145
rect -245 125 -225 145
rect -285 105 -225 125
rect -285 85 -265 105
rect -245 85 -225 105
rect -285 65 -225 85
rect -285 45 -265 65
rect -245 45 -225 65
rect -285 30 -225 45
<< pdiff >>
rect -900 590 -840 625
rect -900 570 -880 590
rect -860 570 -840 590
rect -900 550 -840 570
rect -900 530 -880 550
rect -860 530 -840 550
rect -900 510 -840 530
rect -900 490 -880 510
rect -860 490 -840 510
rect -900 475 -840 490
rect -825 590 -765 625
rect -825 570 -805 590
rect -785 570 -765 590
rect -825 550 -765 570
rect -825 530 -805 550
rect -785 530 -765 550
rect -825 510 -765 530
rect -825 490 -805 510
rect -785 490 -765 510
rect -825 475 -765 490
rect -750 590 -690 625
rect -750 570 -730 590
rect -710 570 -690 590
rect -750 550 -690 570
rect -750 530 -730 550
rect -710 530 -690 550
rect -750 510 -690 530
rect -750 490 -730 510
rect -710 490 -690 510
rect -750 475 -690 490
rect -675 590 -615 625
rect -675 570 -655 590
rect -635 570 -615 590
rect -675 550 -615 570
rect -675 530 -655 550
rect -635 530 -615 550
rect -675 510 -615 530
rect -675 490 -655 510
rect -635 490 -615 510
rect -675 475 -615 490
rect -600 590 -540 625
rect -600 570 -580 590
rect -560 570 -540 590
rect -600 550 -540 570
rect -600 530 -580 550
rect -560 530 -540 550
rect -600 510 -540 530
rect -600 490 -580 510
rect -560 490 -540 510
rect -600 475 -540 490
<< ndiffc >>
rect -1195 125 -1175 145
rect -1195 85 -1175 105
rect -1195 45 -1175 65
rect -1120 125 -1100 145
rect -1120 85 -1100 105
rect -1120 45 -1100 65
rect -1045 125 -1025 145
rect -1045 85 -1025 105
rect -1045 45 -1025 65
rect -970 125 -950 145
rect -970 85 -950 105
rect -970 45 -950 65
rect -880 125 -860 145
rect -880 85 -860 105
rect -880 45 -860 65
rect -805 125 -785 145
rect -805 85 -785 105
rect -805 45 -785 65
rect -730 125 -710 145
rect -730 85 -710 105
rect -730 45 -710 65
rect -655 125 -635 145
rect -655 85 -635 105
rect -655 45 -635 65
rect -580 125 -560 145
rect -580 85 -560 105
rect -580 45 -560 65
rect -490 125 -470 145
rect -490 85 -470 105
rect -490 45 -470 65
rect -265 125 -245 145
rect -265 85 -245 105
rect -265 45 -245 65
<< pdiffc >>
rect -880 570 -860 590
rect -880 530 -860 550
rect -880 490 -860 510
rect -805 570 -785 590
rect -805 530 -785 550
rect -805 490 -785 510
rect -730 570 -710 590
rect -730 530 -710 550
rect -730 490 -710 510
rect -655 570 -635 590
rect -655 530 -635 550
rect -655 490 -635 510
rect -580 570 -560 590
rect -580 530 -560 550
rect -580 490 -560 510
<< psubdiff >>
rect -1220 -55 -220 -40
rect -1220 -75 -1210 -55
rect -1190 -75 -1170 -55
rect -1150 -75 -1130 -55
rect -1110 -75 -1090 -55
rect -1070 -75 -1050 -55
rect -1030 -75 -1010 -55
rect -990 -75 -970 -55
rect -950 -75 -930 -55
rect -910 -75 -890 -55
rect -870 -75 -850 -55
rect -830 -75 -810 -55
rect -790 -75 -770 -55
rect -750 -75 -730 -55
rect -710 -75 -690 -55
rect -670 -75 -650 -55
rect -630 -75 -610 -55
rect -590 -75 -570 -55
rect -550 -75 -530 -55
rect -510 -75 -490 -55
rect -470 -75 -450 -55
rect -430 -75 -410 -55
rect -390 -75 -370 -55
rect -350 -75 -330 -55
rect -310 -75 -290 -55
rect -270 -75 -250 -55
rect -230 -75 -220 -55
rect -1220 -90 -220 -75
<< nsubdiff >>
rect -1220 700 -220 715
rect -1220 680 -1210 700
rect -1190 680 -1170 700
rect -1150 680 -1130 700
rect -1110 680 -1090 700
rect -1070 680 -1050 700
rect -1030 680 -1010 700
rect -990 680 -970 700
rect -950 680 -930 700
rect -910 680 -890 700
rect -870 680 -850 700
rect -830 680 -810 700
rect -790 680 -770 700
rect -750 680 -730 700
rect -710 680 -690 700
rect -670 680 -650 700
rect -630 680 -610 700
rect -590 680 -570 700
rect -550 680 -530 700
rect -510 680 -490 700
rect -470 680 -450 700
rect -430 680 -410 700
rect -390 680 -370 700
rect -350 680 -330 700
rect -310 680 -290 700
rect -270 680 -250 700
rect -230 680 -220 700
rect -1220 665 -220 680
<< psubdiffcont >>
rect -1210 -75 -1190 -55
rect -1170 -75 -1150 -55
rect -1130 -75 -1110 -55
rect -1090 -75 -1070 -55
rect -1050 -75 -1030 -55
rect -1010 -75 -990 -55
rect -970 -75 -950 -55
rect -930 -75 -910 -55
rect -890 -75 -870 -55
rect -850 -75 -830 -55
rect -810 -75 -790 -55
rect -770 -75 -750 -55
rect -730 -75 -710 -55
rect -690 -75 -670 -55
rect -650 -75 -630 -55
rect -610 -75 -590 -55
rect -570 -75 -550 -55
rect -530 -75 -510 -55
rect -490 -75 -470 -55
rect -450 -75 -430 -55
rect -410 -75 -390 -55
rect -370 -75 -350 -55
rect -330 -75 -310 -55
rect -290 -75 -270 -55
rect -250 -75 -230 -55
<< nsubdiffcont >>
rect -1210 680 -1190 700
rect -1170 680 -1150 700
rect -1130 680 -1110 700
rect -1090 680 -1070 700
rect -1050 680 -1030 700
rect -1010 680 -990 700
rect -970 680 -950 700
rect -930 680 -910 700
rect -890 680 -870 700
rect -850 680 -830 700
rect -810 680 -790 700
rect -770 680 -750 700
rect -730 680 -710 700
rect -690 680 -670 700
rect -650 680 -630 700
rect -610 680 -590 700
rect -570 680 -550 700
rect -530 680 -510 700
rect -490 680 -470 700
rect -450 680 -430 700
rect -410 680 -390 700
rect -370 680 -350 700
rect -330 680 -310 700
rect -290 680 -270 700
rect -250 680 -230 700
<< poly >>
rect -840 640 -750 655
rect -840 625 -825 640
rect -765 625 -750 640
rect -690 640 -600 655
rect -690 625 -675 640
rect -615 625 -600 640
rect -840 460 -825 475
rect -765 400 -750 475
rect -690 460 -675 475
rect -615 460 -600 475
rect -715 450 -675 460
rect -715 430 -705 450
rect -685 430 -675 450
rect -715 420 -675 430
rect -765 390 -725 400
rect -765 370 -755 390
rect -735 370 -725 390
rect -765 360 -725 370
rect -1030 280 -990 290
rect -1115 270 -1065 280
rect -1115 250 -1105 270
rect -1085 250 -1065 270
rect -1030 260 -1020 280
rect -1000 260 -990 280
rect -1030 250 -990 260
rect -1115 240 -1065 250
rect -1180 230 -1140 240
rect -1180 210 -1170 230
rect -1150 210 -1140 230
rect -1180 200 -1140 210
rect -1155 180 -1140 200
rect -1080 180 -1065 240
rect -1005 180 -990 250
rect -840 180 -825 195
rect -765 180 -750 360
rect -690 180 -675 420
rect -325 340 -285 350
rect -325 320 -315 340
rect -295 320 -285 340
rect -325 310 -285 320
rect -400 290 -360 300
rect -400 270 -390 290
rect -370 270 -360 290
rect -400 260 -360 270
rect -465 240 -425 250
rect -465 220 -455 240
rect -435 220 -425 240
rect -465 210 -425 220
rect -615 180 -600 195
rect -450 180 -435 210
rect -375 180 -360 260
rect -300 180 -285 310
rect -1155 15 -1140 30
rect -1080 15 -1065 30
rect -1005 15 -990 30
rect -840 15 -825 30
rect -765 15 -750 30
rect -690 15 -675 30
rect -615 15 -600 30
rect -450 15 -435 30
rect -375 15 -360 30
rect -300 15 -285 30
rect -840 5 -800 15
rect -840 -15 -830 5
rect -810 -15 -800 5
rect -840 -25 -800 -15
rect -640 5 -600 15
rect -640 -15 -630 5
rect -610 -15 -600 5
rect -640 -25 -600 -15
<< polycont >>
rect -705 430 -685 450
rect -755 370 -735 390
rect -1105 250 -1085 270
rect -1020 260 -1000 280
rect -1170 210 -1150 230
rect -315 320 -295 340
rect -390 270 -370 290
rect -455 220 -435 240
rect -830 -15 -810 5
rect -630 -15 -610 5
<< locali >>
rect -1220 700 -220 710
rect -1220 680 -1210 700
rect -1190 680 -1170 700
rect -1150 680 -1130 700
rect -1110 680 -1090 700
rect -1070 680 -1050 700
rect -1030 680 -1010 700
rect -990 680 -970 700
rect -950 680 -930 700
rect -910 680 -890 700
rect -870 680 -850 700
rect -830 680 -810 700
rect -790 680 -770 700
rect -750 680 -730 700
rect -710 680 -690 700
rect -670 680 -650 700
rect -630 680 -610 700
rect -590 680 -570 700
rect -550 680 -530 700
rect -510 680 -490 700
rect -470 680 -450 700
rect -430 680 -410 700
rect -390 680 -370 700
rect -350 680 -330 700
rect -310 680 -290 700
rect -270 680 -250 700
rect -230 680 -220 700
rect -1220 670 -220 680
rect -890 590 -850 605
rect -890 570 -880 590
rect -860 570 -850 590
rect -890 550 -850 570
rect -890 530 -880 550
rect -860 530 -850 550
rect -890 510 -850 530
rect -890 490 -880 510
rect -860 490 -850 510
rect -890 480 -850 490
rect -815 590 -775 605
rect -815 570 -805 590
rect -785 570 -775 590
rect -815 550 -775 570
rect -815 530 -805 550
rect -785 530 -775 550
rect -815 510 -775 530
rect -815 490 -805 510
rect -785 490 -775 510
rect -815 475 -775 490
rect -740 590 -700 605
rect -740 570 -730 590
rect -710 570 -700 590
rect -740 550 -700 570
rect -740 530 -730 550
rect -710 530 -700 550
rect -740 510 -700 530
rect -740 490 -730 510
rect -710 490 -700 510
rect -740 480 -700 490
rect -665 590 -625 605
rect -665 570 -655 590
rect -635 570 -625 590
rect -665 550 -625 570
rect -665 530 -655 550
rect -635 530 -625 550
rect -665 510 -625 530
rect -665 490 -655 510
rect -635 490 -625 510
rect -665 475 -625 490
rect -590 590 -550 605
rect -590 570 -580 590
rect -560 570 -550 590
rect -590 550 -550 570
rect -590 530 -580 550
rect -560 530 -550 550
rect -590 510 -550 530
rect -590 490 -580 510
rect -560 490 -550 510
rect -590 480 -550 490
rect -805 450 -785 475
rect -715 450 -675 460
rect -1215 430 -825 450
rect -865 420 -825 430
rect -925 400 -885 410
rect -1215 380 -915 400
rect -895 380 -885 400
rect -865 400 -855 420
rect -835 400 -825 420
rect -865 390 -825 400
rect -805 430 -705 450
rect -685 430 -675 450
rect -925 370 -885 380
rect -1215 350 -940 360
rect -1215 340 -970 350
rect -980 330 -970 340
rect -950 330 -940 350
rect -980 320 -940 330
rect -1215 300 -1000 320
rect -1030 290 -1000 300
rect -1030 280 -990 290
rect -1215 270 -1075 280
rect -1215 260 -1105 270
rect -1115 250 -1105 260
rect -1085 250 -1075 270
rect -1030 260 -1020 280
rect -1000 260 -990 280
rect -1030 250 -990 260
rect -1115 240 -1075 250
rect -1180 230 -1140 240
rect -1215 210 -1170 230
rect -1150 210 -1140 230
rect -1180 200 -1140 210
rect -805 200 -785 430
rect -715 420 -675 430
rect -765 390 -725 400
rect -655 390 -635 475
rect -515 450 -475 460
rect -515 430 -505 450
rect -485 430 -225 450
rect -515 420 -475 430
rect -765 370 -755 390
rect -735 370 -225 390
rect -765 360 -725 370
rect -655 200 -635 370
rect -325 340 -285 350
rect -325 320 -315 340
rect -295 320 -285 340
rect -325 310 -285 320
rect -400 290 -360 300
rect -400 270 -390 290
rect -370 270 -360 290
rect -400 260 -360 270
rect -465 240 -425 250
rect -465 220 -455 240
rect -435 220 -425 240
rect -465 210 -425 220
rect -1120 180 -775 200
rect -1120 160 -1100 180
rect -970 160 -950 180
rect -1205 145 -1165 160
rect -1205 125 -1195 145
rect -1175 125 -1165 145
rect -1205 105 -1165 125
rect -1205 85 -1195 105
rect -1175 85 -1165 105
rect -1205 65 -1165 85
rect -1205 45 -1195 65
rect -1175 45 -1165 65
rect -1205 35 -1165 45
rect -1130 145 -1090 160
rect -1130 125 -1120 145
rect -1100 125 -1090 145
rect -1130 105 -1090 125
rect -1130 85 -1120 105
rect -1100 85 -1090 105
rect -1130 65 -1090 85
rect -1130 45 -1120 65
rect -1100 45 -1090 65
rect -1130 35 -1090 45
rect -1055 145 -1015 160
rect -1055 125 -1045 145
rect -1025 125 -1015 145
rect -1055 105 -1015 125
rect -1055 85 -1045 105
rect -1025 85 -1015 105
rect -1055 65 -1015 85
rect -1055 45 -1045 65
rect -1025 45 -1015 65
rect -1055 35 -1015 45
rect -980 145 -940 160
rect -980 125 -970 145
rect -950 125 -940 145
rect -980 105 -940 125
rect -980 85 -970 105
rect -950 85 -940 105
rect -980 65 -940 85
rect -980 45 -970 65
rect -950 45 -940 65
rect -980 35 -940 45
rect -890 145 -850 160
rect -890 125 -880 145
rect -860 125 -850 145
rect -890 105 -850 125
rect -890 85 -880 105
rect -860 85 -850 105
rect -890 65 -850 85
rect -890 45 -880 65
rect -860 45 -850 65
rect -890 35 -850 45
rect -815 145 -775 180
rect -665 180 -480 200
rect -815 125 -805 145
rect -785 125 -775 145
rect -815 105 -775 125
rect -815 85 -805 105
rect -785 85 -775 105
rect -815 65 -775 85
rect -815 45 -805 65
rect -785 45 -775 65
rect -815 35 -775 45
rect -740 145 -700 160
rect -740 125 -730 145
rect -710 125 -700 145
rect -740 105 -700 125
rect -740 85 -730 105
rect -710 85 -700 105
rect -740 65 -700 85
rect -740 45 -730 65
rect -710 45 -700 65
rect -740 35 -700 45
rect -665 145 -625 180
rect -500 160 -480 180
rect -665 125 -655 145
rect -635 125 -625 145
rect -665 105 -625 125
rect -665 85 -655 105
rect -635 85 -625 105
rect -665 65 -625 85
rect -665 45 -655 65
rect -635 45 -625 65
rect -665 35 -625 45
rect -590 145 -550 160
rect -590 125 -580 145
rect -560 125 -550 145
rect -590 105 -550 125
rect -590 85 -580 105
rect -560 85 -550 105
rect -590 65 -550 85
rect -590 45 -580 65
rect -560 45 -550 65
rect -590 35 -550 45
rect -500 145 -460 160
rect -500 125 -490 145
rect -470 125 -460 145
rect -500 105 -460 125
rect -500 85 -490 105
rect -470 85 -460 105
rect -500 65 -460 85
rect -500 45 -490 65
rect -470 45 -460 65
rect -500 35 -460 45
rect -275 145 -235 160
rect -275 125 -265 145
rect -245 125 -235 145
rect -275 105 -235 125
rect -275 85 -265 105
rect -245 85 -235 105
rect -275 65 -235 85
rect -275 45 -265 65
rect -245 45 -235 65
rect -275 35 -235 45
rect -840 5 -800 15
rect -640 5 -600 15
rect -1215 -15 -830 5
rect -810 -15 -630 5
rect -610 -15 -600 5
rect -840 -25 -800 -15
rect -640 -25 -600 -15
rect -1220 -55 -220 -45
rect -1220 -75 -1210 -55
rect -1190 -75 -1170 -55
rect -1150 -75 -1130 -55
rect -1110 -75 -1090 -55
rect -1070 -75 -1050 -55
rect -1030 -75 -1010 -55
rect -990 -75 -970 -55
rect -950 -75 -930 -55
rect -910 -75 -890 -55
rect -870 -75 -850 -55
rect -830 -75 -810 -55
rect -790 -75 -770 -55
rect -750 -75 -730 -55
rect -710 -75 -690 -55
rect -670 -75 -650 -55
rect -630 -75 -610 -55
rect -590 -75 -570 -55
rect -550 -75 -530 -55
rect -510 -75 -490 -55
rect -470 -75 -450 -55
rect -430 -75 -410 -55
rect -390 -75 -370 -55
rect -350 -75 -330 -55
rect -310 -75 -290 -55
rect -270 -75 -250 -55
rect -230 -75 -220 -55
rect -1220 -85 -220 -75
<< viali >>
rect -1210 680 -1190 700
rect -1170 680 -1150 700
rect -1130 680 -1110 700
rect -1090 680 -1070 700
rect -1050 680 -1030 700
rect -1010 680 -990 700
rect -970 680 -950 700
rect -930 680 -910 700
rect -890 680 -870 700
rect -850 680 -830 700
rect -810 680 -790 700
rect -770 680 -750 700
rect -730 680 -710 700
rect -690 680 -670 700
rect -650 680 -630 700
rect -610 680 -590 700
rect -570 680 -550 700
rect -530 680 -510 700
rect -490 680 -470 700
rect -450 680 -430 700
rect -410 680 -390 700
rect -370 680 -350 700
rect -330 680 -310 700
rect -290 680 -270 700
rect -250 680 -230 700
rect -880 570 -860 590
rect -880 530 -860 550
rect -880 490 -860 510
rect -730 570 -710 590
rect -730 530 -710 550
rect -730 490 -710 510
rect -580 570 -560 590
rect -580 530 -560 550
rect -580 490 -560 510
rect -915 380 -895 400
rect -855 400 -835 420
rect -705 430 -685 450
rect -970 330 -950 350
rect -505 430 -485 450
rect -315 320 -295 340
rect -390 270 -370 290
rect -455 220 -435 240
rect -1195 125 -1175 145
rect -1195 85 -1175 105
rect -1195 45 -1175 65
rect -1045 125 -1025 145
rect -1045 85 -1025 105
rect -1045 45 -1025 65
rect -880 125 -860 145
rect -880 85 -860 105
rect -880 45 -860 65
rect -730 125 -710 145
rect -730 85 -710 105
rect -730 45 -710 65
rect -580 125 -560 145
rect -580 85 -560 105
rect -580 45 -560 65
rect -265 125 -245 145
rect -265 85 -245 105
rect -265 45 -245 65
rect -1210 -75 -1190 -55
rect -1170 -75 -1150 -55
rect -1130 -75 -1110 -55
rect -1090 -75 -1070 -55
rect -1050 -75 -1030 -55
rect -1010 -75 -990 -55
rect -970 -75 -950 -55
rect -930 -75 -910 -55
rect -890 -75 -870 -55
rect -850 -75 -830 -55
rect -810 -75 -790 -55
rect -770 -75 -750 -55
rect -730 -75 -710 -55
rect -690 -75 -670 -55
rect -650 -75 -630 -55
rect -610 -75 -590 -55
rect -570 -75 -550 -55
rect -530 -75 -510 -55
rect -490 -75 -470 -55
rect -450 -75 -430 -55
rect -410 -75 -390 -55
rect -370 -75 -350 -55
rect -330 -75 -310 -55
rect -290 -75 -270 -55
rect -250 -75 -230 -55
<< metal1 >>
rect -1220 700 -220 715
rect -1220 680 -1210 700
rect -1190 680 -1170 700
rect -1150 680 -1130 700
rect -1110 680 -1090 700
rect -1070 680 -1050 700
rect -1030 680 -1010 700
rect -990 680 -970 700
rect -950 680 -930 700
rect -910 680 -890 700
rect -870 680 -850 700
rect -830 680 -810 700
rect -790 680 -770 700
rect -750 680 -730 700
rect -710 680 -690 700
rect -670 680 -650 700
rect -630 680 -610 700
rect -590 680 -570 700
rect -550 680 -530 700
rect -510 680 -490 700
rect -470 680 -450 700
rect -430 680 -410 700
rect -390 680 -370 700
rect -350 680 -330 700
rect -310 680 -290 700
rect -270 680 -250 700
rect -230 680 -220 700
rect -1220 665 -220 680
rect -1195 160 -1175 665
rect -1045 160 -1025 665
rect -890 590 -850 665
rect -890 570 -880 590
rect -860 570 -850 590
rect -890 550 -850 570
rect -890 530 -880 550
rect -860 530 -850 550
rect -890 510 -850 530
rect -890 490 -880 510
rect -860 490 -850 510
rect -890 480 -850 490
rect -740 590 -700 665
rect -740 570 -730 590
rect -710 570 -700 590
rect -740 550 -700 570
rect -740 530 -730 550
rect -710 530 -700 550
rect -740 510 -700 530
rect -740 490 -730 510
rect -710 490 -700 510
rect -740 480 -700 490
rect -590 590 -550 665
rect -590 570 -580 590
rect -560 570 -550 590
rect -590 550 -550 570
rect -590 530 -580 550
rect -560 530 -550 550
rect -590 510 -550 530
rect -590 490 -580 510
rect -560 490 -550 510
rect -590 480 -550 490
rect -715 450 -675 460
rect -515 450 -475 460
rect -715 430 -705 450
rect -685 430 -505 450
rect -485 430 -475 450
rect -865 420 -825 430
rect -715 420 -675 430
rect -515 420 -475 430
rect -925 400 -885 410
rect -925 380 -915 400
rect -895 380 -885 400
rect -865 400 -855 420
rect -835 400 -825 420
rect -865 390 -825 400
rect -925 370 -885 380
rect -980 350 -940 360
rect -980 330 -970 350
rect -950 330 -940 350
rect -980 320 -940 330
rect -970 240 -950 320
rect -915 290 -895 370
rect -855 340 -835 390
rect -325 340 -285 350
rect -855 320 -315 340
rect -295 320 -285 340
rect -325 310 -285 320
rect -400 290 -360 300
rect -915 270 -390 290
rect -370 270 -360 290
rect -400 260 -360 270
rect -465 240 -425 250
rect -970 220 -455 240
rect -435 220 -425 240
rect -465 210 -425 220
rect -265 160 -245 665
rect -1205 145 -1165 160
rect -1205 125 -1195 145
rect -1175 125 -1165 145
rect -1205 105 -1165 125
rect -1205 85 -1195 105
rect -1175 85 -1165 105
rect -1205 65 -1165 85
rect -1205 45 -1195 65
rect -1175 45 -1165 65
rect -1205 35 -1165 45
rect -1055 145 -1015 160
rect -1055 125 -1045 145
rect -1025 125 -1015 145
rect -1055 105 -1015 125
rect -1055 85 -1045 105
rect -1025 85 -1015 105
rect -1055 65 -1015 85
rect -1055 45 -1045 65
rect -1025 45 -1015 65
rect -1055 35 -1015 45
rect -890 145 -850 160
rect -890 125 -880 145
rect -860 125 -850 145
rect -890 105 -850 125
rect -890 85 -880 105
rect -860 85 -850 105
rect -890 65 -850 85
rect -890 45 -880 65
rect -860 45 -850 65
rect -890 35 -850 45
rect -740 145 -700 160
rect -740 125 -730 145
rect -710 125 -700 145
rect -740 105 -700 125
rect -740 85 -730 105
rect -710 85 -700 105
rect -740 65 -700 85
rect -740 45 -730 65
rect -710 45 -700 65
rect -740 35 -700 45
rect -590 145 -550 160
rect -590 125 -580 145
rect -560 125 -550 145
rect -590 105 -550 125
rect -590 85 -580 105
rect -560 85 -550 105
rect -590 65 -550 85
rect -590 45 -580 65
rect -560 45 -550 65
rect -590 35 -550 45
rect -275 145 -235 160
rect -275 125 -265 145
rect -245 125 -235 145
rect -275 105 -235 125
rect -275 85 -265 105
rect -245 85 -235 105
rect -275 65 -235 85
rect -275 45 -265 65
rect -245 45 -235 65
rect -275 35 -235 45
rect -880 -40 -860 35
rect -730 -40 -710 35
rect -580 -40 -560 35
rect -1220 -55 -220 -40
rect -1220 -75 -1210 -55
rect -1190 -75 -1170 -55
rect -1150 -75 -1130 -55
rect -1110 -75 -1090 -55
rect -1070 -75 -1050 -55
rect -1030 -75 -1010 -55
rect -990 -75 -970 -55
rect -950 -75 -930 -55
rect -910 -75 -890 -55
rect -870 -75 -850 -55
rect -830 -75 -810 -55
rect -790 -75 -770 -55
rect -750 -75 -730 -55
rect -710 -75 -690 -55
rect -670 -75 -650 -55
rect -630 -75 -610 -55
rect -590 -75 -570 -55
rect -550 -75 -530 -55
rect -510 -75 -490 -55
rect -470 -75 -450 -55
rect -430 -75 -410 -55
rect -390 -75 -370 -55
rect -350 -75 -330 -55
rect -310 -75 -290 -55
rect -270 -75 -250 -55
rect -230 -75 -220 -55
rect -1220 -90 -220 -75
<< labels >>
rlabel viali -705 430 -685 450 7 OUT_bar
port 8 w
rlabel locali -755 370 -735 390 7 OUT
port 7 w
rlabel metal1 -730 680 -710 700 7 CLK
port 11 w
rlabel locali -1210 435 -1200 445 7 A
port 1 w
rlabel locali -1210 385 -1200 395 7 B
port 3 w
rlabel locali -830 -15 -810 5 7 Dis
port 9 w
rlabel locali -1210 265 -1200 275 7 B_bar
port 4 w
rlabel locali -1210 305 -1200 315 7 A_bar
port 2 w
rlabel locali -1210 345 -1200 355 7 C
port 5 w
rlabel locali -1210 215 -1200 225 7 C_bar
port 6 w
rlabel metal1 -730 -75 -710 -55 7 GND!
port 10 w
<< end >>
