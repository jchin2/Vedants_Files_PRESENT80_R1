magic
tech sky130A
magscale 1 2
timestamp 1671306811
<< metal4 >>
rect -1231 918 1231 1000
rect -1231 682 975 918
rect 1211 682 1231 918
rect -1231 598 1231 682
rect -1231 362 975 598
rect 1211 362 1231 598
rect -1231 278 1231 362
rect -1231 42 975 278
rect 1211 42 1231 278
rect -1231 -42 1231 42
rect -1231 -278 975 -42
rect 1211 -278 1231 -42
rect -1231 -362 1231 -278
rect -1231 -598 975 -362
rect 1211 -598 1231 -362
rect -1231 -682 1231 -598
rect -1231 -918 975 -682
rect 1211 -918 1231 -682
rect -1231 -1000 1231 -918
<< via4 >>
rect 975 682 1211 918
rect 975 362 1211 598
rect 975 42 1211 278
rect 975 -278 1211 -42
rect 975 -598 1211 -362
rect 975 -918 1211 -682
<< mimcap2 >>
rect -1131 758 629 900
rect -1131 -758 -1009 758
rect 507 -758 629 758
rect -1131 -900 629 -758
<< mimcap2contact >>
rect -1009 -758 507 758
<< metal5 >>
rect 933 918 1253 1001
rect -1115 758 613 884
rect -1115 -758 -1009 758
rect 507 -758 613 758
rect -1115 -884 613 -758
rect 933 682 975 918
rect 1211 682 1253 918
rect 933 598 1253 682
rect 933 362 975 598
rect 1211 362 1253 598
rect 933 278 1253 362
rect 933 42 975 278
rect 1211 42 1253 278
rect 933 -42 1253 42
rect 933 -278 975 -42
rect 1211 -278 1253 -42
rect 933 -362 1253 -278
rect 933 -598 975 -362
rect 1211 -598 1253 -362
rect 933 -682 1253 -598
rect 933 -918 975 -682
rect 1211 -918 1253 -682
rect 933 -1001 1253 -918
<< properties >>
string FIXED_BBOX -1231 -1000 729 1000
<< end >>
