**.subckt untitled-21
Vx0 __UNCONNECTED_PIN__0 __UNCONNECTED_PIN__1 3
Vx0_bar __UNCONNECTED_PIN__2 __UNCONNECTED_PIN__3 3
Vk0 __UNCONNECTED_PIN__4 __UNCONNECTED_PIN__5 3
Vk0_bar __UNCONNECTED_PIN__6 __UNCONNECTED_PIN__7 3
Vx1 __UNCONNECTED_PIN__8 __UNCONNECTED_PIN__9 3
Vx1_bar __UNCONNECTED_PIN__10 __UNCONNECTED_PIN__11 3
Vk1 __UNCONNECTED_PIN__12 __UNCONNECTED_PIN__13 3
Vk1_bar __UNCONNECTED_PIN__14 __UNCONNECTED_PIN__15 3
Vx2 __UNCONNECTED_PIN__16 __UNCONNECTED_PIN__17 3
Vx2_bar __UNCONNECTED_PIN__18 __UNCONNECTED_PIN__19 3
Vk2 __UNCONNECTED_PIN__20 __UNCONNECTED_PIN__21 3
Vk2_bar __UNCONNECTED_PIN__22 __UNCONNECTED_PIN__23 3
Vx3 __UNCONNECTED_PIN__24 __UNCONNECTED_PIN__25 3
Vx3_bar __UNCONNECTED_PIN__26 __UNCONNECTED_PIN__27 3
Vk3 __UNCONNECTED_PIN__28 __UNCONNECTED_PIN__29 3
Vk3_bar __UNCONNECTED_PIN__30 __UNCONNECTED_PIN__31 3
Vx4 __UNCONNECTED_PIN__32 __UNCONNECTED_PIN__33 3
Vx4_bar __UNCONNECTED_PIN__34 __UNCONNECTED_PIN__35 3
Vk4 __UNCONNECTED_PIN__36 __UNCONNECTED_PIN__37 3
Vk4_bar __UNCONNECTED_PIN__38 __UNCONNECTED_PIN__39 3
Vx5 __UNCONNECTED_PIN__40 __UNCONNECTED_PIN__41 3
Vx5_bar __UNCONNECTED_PIN__42 __UNCONNECTED_PIN__43 3
Vk5 __UNCONNECTED_PIN__44 __UNCONNECTED_PIN__45 3
Vk5_bar __UNCONNECTED_PIN__46 __UNCONNECTED_PIN__47 3
Vx6 __UNCONNECTED_PIN__48 __UNCONNECTED_PIN__49 3
Vx6_bar __UNCONNECTED_PIN__50 __UNCONNECTED_PIN__51 3
Vk6 __UNCONNECTED_PIN__52 __UNCONNECTED_PIN__53 3
Vk6_bar __UNCONNECTED_PIN__54 __UNCONNECTED_PIN__55 3
Vx7 __UNCONNECTED_PIN__56 __UNCONNECTED_PIN__57 3
Vx7_bar __UNCONNECTED_PIN__58 __UNCONNECTED_PIN__59 3
Vk7 __UNCONNECTED_PIN__60 __UNCONNECTED_PIN__61 3
Vk7_bar __UNCONNECTED_PIN__62 __UNCONNECTED_PIN__63 3
Vx8 __UNCONNECTED_PIN__64 __UNCONNECTED_PIN__65 3
Vx8_bar __UNCONNECTED_PIN__66 __UNCONNECTED_PIN__67 3
Vk8 __UNCONNECTED_PIN__68 __UNCONNECTED_PIN__69 3
Vk8_bar __UNCONNECTED_PIN__70 __UNCONNECTED_PIN__71 3
Vx9 __UNCONNECTED_PIN__72 __UNCONNECTED_PIN__73 3
Vx9_bar __UNCONNECTED_PIN__74 __UNCONNECTED_PIN__75 3
Vk9 __UNCONNECTED_PIN__76 __UNCONNECTED_PIN__77 3
Vk9_bar __UNCONNECTED_PIN__78 __UNCONNECTED_PIN__79 3
Vx10 __UNCONNECTED_PIN__80 __UNCONNECTED_PIN__81 3
Vx10_bar __UNCONNECTED_PIN__82 __UNCONNECTED_PIN__83 3
Vk10 __UNCONNECTED_PIN__84 __UNCONNECTED_PIN__85 3
Vk10_bar __UNCONNECTED_PIN__86 __UNCONNECTED_PIN__87 3
Vx11 __UNCONNECTED_PIN__88 __UNCONNECTED_PIN__89 3
Vx11_bar __UNCONNECTED_PIN__90 __UNCONNECTED_PIN__91 3
Vk11 __UNCONNECTED_PIN__92 __UNCONNECTED_PIN__93 3
Vk11_bar __UNCONNECTED_PIN__94 __UNCONNECTED_PIN__95 3
Vx12 __UNCONNECTED_PIN__96 __UNCONNECTED_PIN__97 3
Vx12_bar __UNCONNECTED_PIN__98 __UNCONNECTED_PIN__99 3
Vk12 __UNCONNECTED_PIN__100 __UNCONNECTED_PIN__101 3
Vk12_bar __UNCONNECTED_PIN__102 __UNCONNECTED_PIN__103 3
Vx13 __UNCONNECTED_PIN__104 __UNCONNECTED_PIN__105 3
Vx13_bar __UNCONNECTED_PIN__106 __UNCONNECTED_PIN__107 3
Vk13 __UNCONNECTED_PIN__108 __UNCONNECTED_PIN__109 3
Vk13_bar __UNCONNECTED_PIN__110 __UNCONNECTED_PIN__111 3
Vx14 __UNCONNECTED_PIN__112 __UNCONNECTED_PIN__113 3
Vx14_bar __UNCONNECTED_PIN__114 __UNCONNECTED_PIN__115 3
Vk14 __UNCONNECTED_PIN__116 __UNCONNECTED_PIN__117 3
Vk14_bar __UNCONNECTED_PIN__118 __UNCONNECTED_PIN__119 3
Vx15 __UNCONNECTED_PIN__120 __UNCONNECTED_PIN__121 3
Vx15_bar __UNCONNECTED_PIN__122 __UNCONNECTED_PIN__123 3
Vk15 __UNCONNECTED_PIN__124 __UNCONNECTED_PIN__125 3
Vk15_bar __UNCONNECTED_PIN__126 __UNCONNECTED_PIN__127 3
Vx16 __UNCONNECTED_PIN__128 __UNCONNECTED_PIN__129 3
Vx16_bar __UNCONNECTED_PIN__130 __UNCONNECTED_PIN__131 3
Vk16 __UNCONNECTED_PIN__132 __UNCONNECTED_PIN__133 3
Vk16_bar __UNCONNECTED_PIN__134 __UNCONNECTED_PIN__135 3
Vx17 __UNCONNECTED_PIN__136 __UNCONNECTED_PIN__137 3
Vx17_bar __UNCONNECTED_PIN__138 __UNCONNECTED_PIN__139 3
Vk17 __UNCONNECTED_PIN__140 __UNCONNECTED_PIN__141 3
Vk17_bar __UNCONNECTED_PIN__142 __UNCONNECTED_PIN__143 3
Vx18 __UNCONNECTED_PIN__144 __UNCONNECTED_PIN__145 3
Vx18_bar __UNCONNECTED_PIN__146 __UNCONNECTED_PIN__147 3
Vk18 __UNCONNECTED_PIN__148 __UNCONNECTED_PIN__149 3
Vk18_bar __UNCONNECTED_PIN__150 __UNCONNECTED_PIN__151 3
Vx19 __UNCONNECTED_PIN__152 __UNCONNECTED_PIN__153 3
Vx19_bar __UNCONNECTED_PIN__154 __UNCONNECTED_PIN__155 3
Vk19 __UNCONNECTED_PIN__156 __UNCONNECTED_PIN__157 3
Vk19_bar __UNCONNECTED_PIN__158 __UNCONNECTED_PIN__159 3
Vx20 __UNCONNECTED_PIN__160 __UNCONNECTED_PIN__161 3
Vx20_bar __UNCONNECTED_PIN__162 __UNCONNECTED_PIN__163 3
Vk20 __UNCONNECTED_PIN__164 __UNCONNECTED_PIN__165 3
Vk20_bar __UNCONNECTED_PIN__166 __UNCONNECTED_PIN__167 3
Vx21 __UNCONNECTED_PIN__168 __UNCONNECTED_PIN__169 3
Vx21_bar __UNCONNECTED_PIN__170 __UNCONNECTED_PIN__171 3
Vk21 __UNCONNECTED_PIN__172 __UNCONNECTED_PIN__173 3
Vk21_bar __UNCONNECTED_PIN__174 __UNCONNECTED_PIN__175 3
Vx22 __UNCONNECTED_PIN__176 __UNCONNECTED_PIN__177 3
Vx22_bar __UNCONNECTED_PIN__178 __UNCONNECTED_PIN__179 3
Vk22 __UNCONNECTED_PIN__180 __UNCONNECTED_PIN__181 3
Vk22_bar __UNCONNECTED_PIN__182 __UNCONNECTED_PIN__183 3
Vx23 __UNCONNECTED_PIN__184 __UNCONNECTED_PIN__185 3
Vx23_bar __UNCONNECTED_PIN__186 __UNCONNECTED_PIN__187 3
Vk23 __UNCONNECTED_PIN__188 __UNCONNECTED_PIN__189 3
Vk23_bar __UNCONNECTED_PIN__190 __UNCONNECTED_PIN__191 3
Vx24 __UNCONNECTED_PIN__192 __UNCONNECTED_PIN__193 3
Vx24_bar __UNCONNECTED_PIN__194 __UNCONNECTED_PIN__195 3
Vk24 __UNCONNECTED_PIN__196 __UNCONNECTED_PIN__197 3
Vk24_bar __UNCONNECTED_PIN__198 __UNCONNECTED_PIN__199 3
Vx25 __UNCONNECTED_PIN__200 __UNCONNECTED_PIN__201 3
Vx25_bar __UNCONNECTED_PIN__202 __UNCONNECTED_PIN__203 3
Vk25 __UNCONNECTED_PIN__204 __UNCONNECTED_PIN__205 3
Vk25_bar __UNCONNECTED_PIN__206 __UNCONNECTED_PIN__207 3
Vx26 __UNCONNECTED_PIN__208 __UNCONNECTED_PIN__209 3
Vx26_bar __UNCONNECTED_PIN__210 __UNCONNECTED_PIN__211 3
Vk26 __UNCONNECTED_PIN__212 __UNCONNECTED_PIN__213 3
Vk26_bar __UNCONNECTED_PIN__214 __UNCONNECTED_PIN__215 3
Vx27 __UNCONNECTED_PIN__216 __UNCONNECTED_PIN__217 3
Vx27_bar __UNCONNECTED_PIN__218 __UNCONNECTED_PIN__219 3
Vk27 __UNCONNECTED_PIN__220 __UNCONNECTED_PIN__221 3
Vk27_bar __UNCONNECTED_PIN__222 __UNCONNECTED_PIN__223 3
Vx28 __UNCONNECTED_PIN__224 __UNCONNECTED_PIN__225 3
Vx28_bar __UNCONNECTED_PIN__226 __UNCONNECTED_PIN__227 3
Vk28 __UNCONNECTED_PIN__228 __UNCONNECTED_PIN__229 3
Vk28_bar __UNCONNECTED_PIN__230 __UNCONNECTED_PIN__231 3
Vx29 __UNCONNECTED_PIN__232 __UNCONNECTED_PIN__233 3
Vx29_bar __UNCONNECTED_PIN__234 __UNCONNECTED_PIN__235 3
Vk29 __UNCONNECTED_PIN__236 __UNCONNECTED_PIN__237 3
Vk29_bar __UNCONNECTED_PIN__238 __UNCONNECTED_PIN__239 3
Vx30 __UNCONNECTED_PIN__240 __UNCONNECTED_PIN__241 3
Vx30_bar __UNCONNECTED_PIN__242 __UNCONNECTED_PIN__243 3
Vk30 __UNCONNECTED_PIN__244 __UNCONNECTED_PIN__245 3
Vk30_bar __UNCONNECTED_PIN__246 __UNCONNECTED_PIN__247 3
Vx31 __UNCONNECTED_PIN__248 __UNCONNECTED_PIN__249 3
Vx31_bar __UNCONNECTED_PIN__250 __UNCONNECTED_PIN__251 3
Vk31 __UNCONNECTED_PIN__252 __UNCONNECTED_PIN__253 3
Vk31_bar __UNCONNECTED_PIN__254 __UNCONNECTED_PIN__255 3
Vx32 __UNCONNECTED_PIN__256 __UNCONNECTED_PIN__257 3
Vx32_bar __UNCONNECTED_PIN__258 __UNCONNECTED_PIN__259 3
Vk32 __UNCONNECTED_PIN__260 __UNCONNECTED_PIN__261 3
Vk32_bar __UNCONNECTED_PIN__262 __UNCONNECTED_PIN__263 3
Vx33 __UNCONNECTED_PIN__264 __UNCONNECTED_PIN__265 3
Vx33_bar __UNCONNECTED_PIN__266 __UNCONNECTED_PIN__267 3
Vk33 __UNCONNECTED_PIN__268 __UNCONNECTED_PIN__269 3
Vk33_bar __UNCONNECTED_PIN__270 __UNCONNECTED_PIN__271 3
Vx34 __UNCONNECTED_PIN__272 __UNCONNECTED_PIN__273 3
Vx34_bar __UNCONNECTED_PIN__274 __UNCONNECTED_PIN__275 3
Vk34 __UNCONNECTED_PIN__276 __UNCONNECTED_PIN__277 3
Vk34_bar __UNCONNECTED_PIN__278 __UNCONNECTED_PIN__279 3
Vx35 __UNCONNECTED_PIN__280 __UNCONNECTED_PIN__281 3
Vx35_bar __UNCONNECTED_PIN__282 __UNCONNECTED_PIN__283 3
Vk35 __UNCONNECTED_PIN__284 __UNCONNECTED_PIN__285 3
Vk35_bar __UNCONNECTED_PIN__286 __UNCONNECTED_PIN__287 3
Vx36 __UNCONNECTED_PIN__288 __UNCONNECTED_PIN__289 3
Vx36_bar __UNCONNECTED_PIN__290 __UNCONNECTED_PIN__291 3
Vk36 __UNCONNECTED_PIN__292 __UNCONNECTED_PIN__293 3
Vk36_bar __UNCONNECTED_PIN__294 __UNCONNECTED_PIN__295 3
Vx37 __UNCONNECTED_PIN__296 __UNCONNECTED_PIN__297 3
Vx37_bar __UNCONNECTED_PIN__298 __UNCONNECTED_PIN__299 3
Vk37 __UNCONNECTED_PIN__300 __UNCONNECTED_PIN__301 3
Vk37_bar __UNCONNECTED_PIN__302 __UNCONNECTED_PIN__303 3
Vx38 __UNCONNECTED_PIN__304 __UNCONNECTED_PIN__305 3
Vx38_bar __UNCONNECTED_PIN__306 __UNCONNECTED_PIN__307 3
Vk38 __UNCONNECTED_PIN__308 __UNCONNECTED_PIN__309 3
Vk38_bar __UNCONNECTED_PIN__310 __UNCONNECTED_PIN__311 3
Vx39 __UNCONNECTED_PIN__312 __UNCONNECTED_PIN__313 3
Vx39_bar __UNCONNECTED_PIN__314 __UNCONNECTED_PIN__315 3
Vk39 __UNCONNECTED_PIN__316 __UNCONNECTED_PIN__317 3
Vk39_bar __UNCONNECTED_PIN__318 __UNCONNECTED_PIN__319 3
Vx40 __UNCONNECTED_PIN__320 __UNCONNECTED_PIN__321 3
Vx40_bar __UNCONNECTED_PIN__322 __UNCONNECTED_PIN__323 3
Vk40 __UNCONNECTED_PIN__324 __UNCONNECTED_PIN__325 3
Vk40_bar __UNCONNECTED_PIN__326 __UNCONNECTED_PIN__327 3
Vx41 __UNCONNECTED_PIN__328 __UNCONNECTED_PIN__329 3
Vx41_bar __UNCONNECTED_PIN__330 __UNCONNECTED_PIN__331 3
Vk41 __UNCONNECTED_PIN__332 __UNCONNECTED_PIN__333 3
Vk41_bar __UNCONNECTED_PIN__334 __UNCONNECTED_PIN__335 3
Vx42 __UNCONNECTED_PIN__336 __UNCONNECTED_PIN__337 3
Vx42_bar __UNCONNECTED_PIN__338 __UNCONNECTED_PIN__339 3
Vk42 __UNCONNECTED_PIN__340 __UNCONNECTED_PIN__341 3
Vk42_bar __UNCONNECTED_PIN__342 __UNCONNECTED_PIN__343 3
Vx43 __UNCONNECTED_PIN__344 __UNCONNECTED_PIN__345 3
Vx43_bar __UNCONNECTED_PIN__346 __UNCONNECTED_PIN__347 3
Vk43 __UNCONNECTED_PIN__348 __UNCONNECTED_PIN__349 3
Vk43_bar __UNCONNECTED_PIN__350 __UNCONNECTED_PIN__351 3
Vx44 __UNCONNECTED_PIN__352 __UNCONNECTED_PIN__353 3
Vx44_bar __UNCONNECTED_PIN__354 __UNCONNECTED_PIN__355 3
Vk44 __UNCONNECTED_PIN__356 __UNCONNECTED_PIN__357 3
Vk44_bar __UNCONNECTED_PIN__358 __UNCONNECTED_PIN__359 3
Vx45 __UNCONNECTED_PIN__360 __UNCONNECTED_PIN__361 3
Vx45_bar __UNCONNECTED_PIN__362 __UNCONNECTED_PIN__363 3
Vk45 __UNCONNECTED_PIN__364 __UNCONNECTED_PIN__365 3
Vk45_bar __UNCONNECTED_PIN__366 __UNCONNECTED_PIN__367 3
Vx46 __UNCONNECTED_PIN__368 __UNCONNECTED_PIN__369 3
Vx46_bar __UNCONNECTED_PIN__370 __UNCONNECTED_PIN__371 3
Vk46 __UNCONNECTED_PIN__372 __UNCONNECTED_PIN__373 3
Vk46_bar __UNCONNECTED_PIN__374 __UNCONNECTED_PIN__375 3
Vx47 __UNCONNECTED_PIN__376 __UNCONNECTED_PIN__377 3
Vx47_bar __UNCONNECTED_PIN__378 __UNCONNECTED_PIN__379 3
Vk47 __UNCONNECTED_PIN__380 __UNCONNECTED_PIN__381 3
Vk47_bar __UNCONNECTED_PIN__382 __UNCONNECTED_PIN__383 3
Vx48 __UNCONNECTED_PIN__384 __UNCONNECTED_PIN__385 3
Vx48_bar __UNCONNECTED_PIN__386 __UNCONNECTED_PIN__387 3
Vk48 __UNCONNECTED_PIN__388 __UNCONNECTED_PIN__389 3
Vk48_bar __UNCONNECTED_PIN__390 __UNCONNECTED_PIN__391 3
Vx49 __UNCONNECTED_PIN__392 __UNCONNECTED_PIN__393 3
Vx49_bar __UNCONNECTED_PIN__394 __UNCONNECTED_PIN__395 3
Vk49 __UNCONNECTED_PIN__396 __UNCONNECTED_PIN__397 3
Vk49_bar __UNCONNECTED_PIN__398 __UNCONNECTED_PIN__399 3
Vx50 __UNCONNECTED_PIN__400 __UNCONNECTED_PIN__401 3
Vx50_bar __UNCONNECTED_PIN__402 __UNCONNECTED_PIN__403 3
Vk50 __UNCONNECTED_PIN__404 __UNCONNECTED_PIN__405 3
Vk50_bar __UNCONNECTED_PIN__406 __UNCONNECTED_PIN__407 3
Vx51 __UNCONNECTED_PIN__408 __UNCONNECTED_PIN__409 3
Vx51_bar __UNCONNECTED_PIN__410 __UNCONNECTED_PIN__411 3
Vk51 __UNCONNECTED_PIN__412 __UNCONNECTED_PIN__413 3
Vk51_bar __UNCONNECTED_PIN__414 __UNCONNECTED_PIN__415 3
Vx52 __UNCONNECTED_PIN__416 __UNCONNECTED_PIN__417 3
Vx52_bar __UNCONNECTED_PIN__418 __UNCONNECTED_PIN__419 3
Vk52 __UNCONNECTED_PIN__420 __UNCONNECTED_PIN__421 3
Vk52_bar __UNCONNECTED_PIN__422 __UNCONNECTED_PIN__423 3
Vx53 __UNCONNECTED_PIN__424 __UNCONNECTED_PIN__425 3
Vx53_bar __UNCONNECTED_PIN__426 __UNCONNECTED_PIN__427 3
Vk53 __UNCONNECTED_PIN__428 __UNCONNECTED_PIN__429 3
Vk53_bar __UNCONNECTED_PIN__430 __UNCONNECTED_PIN__431 3
Vx54 __UNCONNECTED_PIN__432 __UNCONNECTED_PIN__433 3
Vx54_bar __UNCONNECTED_PIN__434 __UNCONNECTED_PIN__435 3
Vk54 __UNCONNECTED_PIN__436 __UNCONNECTED_PIN__437 3
Vk54_bar __UNCONNECTED_PIN__438 __UNCONNECTED_PIN__439 3
Vx55 __UNCONNECTED_PIN__440 __UNCONNECTED_PIN__441 3
Vx55_bar __UNCONNECTED_PIN__442 __UNCONNECTED_PIN__443 3
Vk55 __UNCONNECTED_PIN__444 __UNCONNECTED_PIN__445 3
Vk55_bar __UNCONNECTED_PIN__446 __UNCONNECTED_PIN__447 3
Vx56 __UNCONNECTED_PIN__448 __UNCONNECTED_PIN__449 3
Vx56_bar __UNCONNECTED_PIN__450 __UNCONNECTED_PIN__451 3
Vk56 __UNCONNECTED_PIN__452 __UNCONNECTED_PIN__453 3
Vk56_bar __UNCONNECTED_PIN__454 __UNCONNECTED_PIN__455 3
Vx57 __UNCONNECTED_PIN__456 __UNCONNECTED_PIN__457 3
Vx57_bar __UNCONNECTED_PIN__458 __UNCONNECTED_PIN__459 3
Vk57 __UNCONNECTED_PIN__460 __UNCONNECTED_PIN__461 3
Vk57_bar __UNCONNECTED_PIN__462 __UNCONNECTED_PIN__463 3
Vx58 __UNCONNECTED_PIN__464 __UNCONNECTED_PIN__465 3
Vx58_bar __UNCONNECTED_PIN__466 __UNCONNECTED_PIN__467 3
Vk58 __UNCONNECTED_PIN__468 __UNCONNECTED_PIN__469 3
Vk58_bar __UNCONNECTED_PIN__470 __UNCONNECTED_PIN__471 3
Vx59 __UNCONNECTED_PIN__472 __UNCONNECTED_PIN__473 3
Vx59_bar __UNCONNECTED_PIN__474 __UNCONNECTED_PIN__475 3
Vk59 __UNCONNECTED_PIN__476 __UNCONNECTED_PIN__477 3
Vk59_bar __UNCONNECTED_PIN__478 __UNCONNECTED_PIN__479 3
Vx60 __UNCONNECTED_PIN__480 __UNCONNECTED_PIN__481 3
Vx60_bar __UNCONNECTED_PIN__482 __UNCONNECTED_PIN__483 3
Vk60 __UNCONNECTED_PIN__484 __UNCONNECTED_PIN__485 3
Vk60_bar __UNCONNECTED_PIN__486 __UNCONNECTED_PIN__487 3
Vx61 __UNCONNECTED_PIN__488 __UNCONNECTED_PIN__489 3
Vx61_bar __UNCONNECTED_PIN__490 __UNCONNECTED_PIN__491 3
Vk61 __UNCONNECTED_PIN__492 __UNCONNECTED_PIN__493 3
Vk61_bar __UNCONNECTED_PIN__494 __UNCONNECTED_PIN__495 3
Vx62 __UNCONNECTED_PIN__496 __UNCONNECTED_PIN__497 3
Vx62_bar __UNCONNECTED_PIN__498 __UNCONNECTED_PIN__499 3
Vk62 __UNCONNECTED_PIN__500 __UNCONNECTED_PIN__501 3
Vk62_bar __UNCONNECTED_PIN__502 __UNCONNECTED_PIN__503 3
Vx63 __UNCONNECTED_PIN__504 __UNCONNECTED_PIN__505 3
Vx63_bar __UNCONNECTED_PIN__506 __UNCONNECTED_PIN__507 3
Vk63 __UNCONNECTED_PIN__508 __UNCONNECTED_PIN__509 3
Vk63_bar __UNCONNECTED_PIN__510 __UNCONNECTED_PIN__511 3
**.ends
** flattened .save nodes
.end
