magic
tech sky130A
magscale 1 2
timestamp 1671306811
<< pwell >>
rect -1316 -6 536 1038
<< nmoslvt >>
rect -990 20 -960 1012
rect -840 20 -810 1012
rect -690 20 -660 1012
rect -540 20 -510 1012
rect -390 20 -360 1012
rect -240 20 -210 1012
rect -90 20 -60 1012
rect 60 20 90 1012
rect 210 20 240 1012
rect 360 20 390 1012
<< ndiff >>
rect -1110 984 -990 1012
rect -1110 950 -1067 984
rect -1033 950 -990 984
rect -1110 916 -990 950
rect -1110 882 -1067 916
rect -1033 882 -990 916
rect -1110 848 -990 882
rect -1110 814 -1067 848
rect -1033 814 -990 848
rect -1110 780 -990 814
rect -1110 746 -1067 780
rect -1033 746 -990 780
rect -1110 712 -990 746
rect -1110 678 -1067 712
rect -1033 678 -990 712
rect -1110 644 -990 678
rect -1110 610 -1067 644
rect -1033 610 -990 644
rect -1110 576 -990 610
rect -1110 542 -1067 576
rect -1033 542 -990 576
rect -1110 508 -990 542
rect -1110 474 -1067 508
rect -1033 474 -990 508
rect -1110 440 -990 474
rect -1110 406 -1067 440
rect -1033 406 -990 440
rect -1110 372 -990 406
rect -1110 338 -1067 372
rect -1033 338 -990 372
rect -1110 304 -990 338
rect -1110 270 -1067 304
rect -1033 270 -990 304
rect -1110 236 -990 270
rect -1110 202 -1067 236
rect -1033 202 -990 236
rect -1110 168 -990 202
rect -1110 134 -1067 168
rect -1033 134 -990 168
rect -1110 100 -990 134
rect -1110 66 -1067 100
rect -1033 66 -990 100
rect -1110 20 -990 66
rect -960 984 -840 1012
rect -960 950 -917 984
rect -883 950 -840 984
rect -960 916 -840 950
rect -960 882 -917 916
rect -883 882 -840 916
rect -960 848 -840 882
rect -960 814 -917 848
rect -883 814 -840 848
rect -960 780 -840 814
rect -960 746 -917 780
rect -883 746 -840 780
rect -960 712 -840 746
rect -960 678 -917 712
rect -883 678 -840 712
rect -960 644 -840 678
rect -960 610 -917 644
rect -883 610 -840 644
rect -960 576 -840 610
rect -960 542 -917 576
rect -883 542 -840 576
rect -960 508 -840 542
rect -960 474 -917 508
rect -883 474 -840 508
rect -960 440 -840 474
rect -960 406 -917 440
rect -883 406 -840 440
rect -960 372 -840 406
rect -960 338 -917 372
rect -883 338 -840 372
rect -960 304 -840 338
rect -960 270 -917 304
rect -883 270 -840 304
rect -960 236 -840 270
rect -960 202 -917 236
rect -883 202 -840 236
rect -960 168 -840 202
rect -960 134 -917 168
rect -883 134 -840 168
rect -960 100 -840 134
rect -960 66 -917 100
rect -883 66 -840 100
rect -960 20 -840 66
rect -810 984 -690 1012
rect -810 950 -767 984
rect -733 950 -690 984
rect -810 916 -690 950
rect -810 882 -767 916
rect -733 882 -690 916
rect -810 848 -690 882
rect -810 814 -767 848
rect -733 814 -690 848
rect -810 780 -690 814
rect -810 746 -767 780
rect -733 746 -690 780
rect -810 712 -690 746
rect -810 678 -767 712
rect -733 678 -690 712
rect -810 644 -690 678
rect -810 610 -767 644
rect -733 610 -690 644
rect -810 576 -690 610
rect -810 542 -767 576
rect -733 542 -690 576
rect -810 508 -690 542
rect -810 474 -767 508
rect -733 474 -690 508
rect -810 440 -690 474
rect -810 406 -767 440
rect -733 406 -690 440
rect -810 372 -690 406
rect -810 338 -767 372
rect -733 338 -690 372
rect -810 304 -690 338
rect -810 270 -767 304
rect -733 270 -690 304
rect -810 236 -690 270
rect -810 202 -767 236
rect -733 202 -690 236
rect -810 168 -690 202
rect -810 134 -767 168
rect -733 134 -690 168
rect -810 100 -690 134
rect -810 66 -767 100
rect -733 66 -690 100
rect -810 20 -690 66
rect -660 984 -540 1012
rect -660 950 -617 984
rect -583 950 -540 984
rect -660 916 -540 950
rect -660 882 -617 916
rect -583 882 -540 916
rect -660 848 -540 882
rect -660 814 -617 848
rect -583 814 -540 848
rect -660 780 -540 814
rect -660 746 -617 780
rect -583 746 -540 780
rect -660 712 -540 746
rect -660 678 -617 712
rect -583 678 -540 712
rect -660 644 -540 678
rect -660 610 -617 644
rect -583 610 -540 644
rect -660 576 -540 610
rect -660 542 -617 576
rect -583 542 -540 576
rect -660 508 -540 542
rect -660 474 -617 508
rect -583 474 -540 508
rect -660 440 -540 474
rect -660 406 -617 440
rect -583 406 -540 440
rect -660 372 -540 406
rect -660 338 -617 372
rect -583 338 -540 372
rect -660 304 -540 338
rect -660 270 -617 304
rect -583 270 -540 304
rect -660 236 -540 270
rect -660 202 -617 236
rect -583 202 -540 236
rect -660 168 -540 202
rect -660 134 -617 168
rect -583 134 -540 168
rect -660 100 -540 134
rect -660 66 -617 100
rect -583 66 -540 100
rect -660 20 -540 66
rect -510 984 -390 1012
rect -510 950 -467 984
rect -433 950 -390 984
rect -510 916 -390 950
rect -510 882 -467 916
rect -433 882 -390 916
rect -510 848 -390 882
rect -510 814 -467 848
rect -433 814 -390 848
rect -510 780 -390 814
rect -510 746 -467 780
rect -433 746 -390 780
rect -510 712 -390 746
rect -510 678 -467 712
rect -433 678 -390 712
rect -510 644 -390 678
rect -510 610 -467 644
rect -433 610 -390 644
rect -510 576 -390 610
rect -510 542 -467 576
rect -433 542 -390 576
rect -510 508 -390 542
rect -510 474 -467 508
rect -433 474 -390 508
rect -510 440 -390 474
rect -510 406 -467 440
rect -433 406 -390 440
rect -510 372 -390 406
rect -510 338 -467 372
rect -433 338 -390 372
rect -510 304 -390 338
rect -510 270 -467 304
rect -433 270 -390 304
rect -510 236 -390 270
rect -510 202 -467 236
rect -433 202 -390 236
rect -510 168 -390 202
rect -510 134 -467 168
rect -433 134 -390 168
rect -510 100 -390 134
rect -510 66 -467 100
rect -433 66 -390 100
rect -510 20 -390 66
rect -360 984 -240 1012
rect -360 950 -317 984
rect -283 950 -240 984
rect -360 916 -240 950
rect -360 882 -317 916
rect -283 882 -240 916
rect -360 848 -240 882
rect -360 814 -317 848
rect -283 814 -240 848
rect -360 780 -240 814
rect -360 746 -317 780
rect -283 746 -240 780
rect -360 712 -240 746
rect -360 678 -317 712
rect -283 678 -240 712
rect -360 644 -240 678
rect -360 610 -317 644
rect -283 610 -240 644
rect -360 576 -240 610
rect -360 542 -317 576
rect -283 542 -240 576
rect -360 508 -240 542
rect -360 474 -317 508
rect -283 474 -240 508
rect -360 440 -240 474
rect -360 406 -317 440
rect -283 406 -240 440
rect -360 372 -240 406
rect -360 338 -317 372
rect -283 338 -240 372
rect -360 304 -240 338
rect -360 270 -317 304
rect -283 270 -240 304
rect -360 236 -240 270
rect -360 202 -317 236
rect -283 202 -240 236
rect -360 168 -240 202
rect -360 134 -317 168
rect -283 134 -240 168
rect -360 100 -240 134
rect -360 66 -317 100
rect -283 66 -240 100
rect -360 20 -240 66
rect -210 984 -90 1012
rect -210 950 -167 984
rect -133 950 -90 984
rect -210 916 -90 950
rect -210 882 -167 916
rect -133 882 -90 916
rect -210 848 -90 882
rect -210 814 -167 848
rect -133 814 -90 848
rect -210 780 -90 814
rect -210 746 -167 780
rect -133 746 -90 780
rect -210 712 -90 746
rect -210 678 -167 712
rect -133 678 -90 712
rect -210 644 -90 678
rect -210 610 -167 644
rect -133 610 -90 644
rect -210 576 -90 610
rect -210 542 -167 576
rect -133 542 -90 576
rect -210 508 -90 542
rect -210 474 -167 508
rect -133 474 -90 508
rect -210 440 -90 474
rect -210 406 -167 440
rect -133 406 -90 440
rect -210 372 -90 406
rect -210 338 -167 372
rect -133 338 -90 372
rect -210 304 -90 338
rect -210 270 -167 304
rect -133 270 -90 304
rect -210 236 -90 270
rect -210 202 -167 236
rect -133 202 -90 236
rect -210 168 -90 202
rect -210 134 -167 168
rect -133 134 -90 168
rect -210 100 -90 134
rect -210 66 -167 100
rect -133 66 -90 100
rect -210 20 -90 66
rect -60 984 60 1012
rect -60 950 -17 984
rect 17 950 60 984
rect -60 916 60 950
rect -60 882 -17 916
rect 17 882 60 916
rect -60 848 60 882
rect -60 814 -17 848
rect 17 814 60 848
rect -60 780 60 814
rect -60 746 -17 780
rect 17 746 60 780
rect -60 712 60 746
rect -60 678 -17 712
rect 17 678 60 712
rect -60 644 60 678
rect -60 610 -17 644
rect 17 610 60 644
rect -60 576 60 610
rect -60 542 -17 576
rect 17 542 60 576
rect -60 508 60 542
rect -60 474 -17 508
rect 17 474 60 508
rect -60 440 60 474
rect -60 406 -17 440
rect 17 406 60 440
rect -60 372 60 406
rect -60 338 -17 372
rect 17 338 60 372
rect -60 304 60 338
rect -60 270 -17 304
rect 17 270 60 304
rect -60 236 60 270
rect -60 202 -17 236
rect 17 202 60 236
rect -60 168 60 202
rect -60 134 -17 168
rect 17 134 60 168
rect -60 100 60 134
rect -60 66 -17 100
rect 17 66 60 100
rect -60 20 60 66
rect 90 984 210 1012
rect 90 950 133 984
rect 167 950 210 984
rect 90 916 210 950
rect 90 882 133 916
rect 167 882 210 916
rect 90 848 210 882
rect 90 814 133 848
rect 167 814 210 848
rect 90 780 210 814
rect 90 746 133 780
rect 167 746 210 780
rect 90 712 210 746
rect 90 678 133 712
rect 167 678 210 712
rect 90 644 210 678
rect 90 610 133 644
rect 167 610 210 644
rect 90 576 210 610
rect 90 542 133 576
rect 167 542 210 576
rect 90 508 210 542
rect 90 474 133 508
rect 167 474 210 508
rect 90 440 210 474
rect 90 406 133 440
rect 167 406 210 440
rect 90 372 210 406
rect 90 338 133 372
rect 167 338 210 372
rect 90 304 210 338
rect 90 270 133 304
rect 167 270 210 304
rect 90 236 210 270
rect 90 202 133 236
rect 167 202 210 236
rect 90 168 210 202
rect 90 134 133 168
rect 167 134 210 168
rect 90 100 210 134
rect 90 66 133 100
rect 167 66 210 100
rect 90 20 210 66
rect 240 984 360 1012
rect 240 950 283 984
rect 317 950 360 984
rect 240 916 360 950
rect 240 882 283 916
rect 317 882 360 916
rect 240 848 360 882
rect 240 814 283 848
rect 317 814 360 848
rect 240 780 360 814
rect 240 746 283 780
rect 317 746 360 780
rect 240 712 360 746
rect 240 678 283 712
rect 317 678 360 712
rect 240 644 360 678
rect 240 610 283 644
rect 317 610 360 644
rect 240 576 360 610
rect 240 542 283 576
rect 317 542 360 576
rect 240 508 360 542
rect 240 474 283 508
rect 317 474 360 508
rect 240 440 360 474
rect 240 406 283 440
rect 317 406 360 440
rect 240 372 360 406
rect 240 338 283 372
rect 317 338 360 372
rect 240 304 360 338
rect 240 270 283 304
rect 317 270 360 304
rect 240 236 360 270
rect 240 202 283 236
rect 317 202 360 236
rect 240 168 360 202
rect 240 134 283 168
rect 317 134 360 168
rect 240 100 360 134
rect 240 66 283 100
rect 317 66 360 100
rect 240 20 360 66
rect 390 984 510 1012
rect 390 950 433 984
rect 467 950 510 984
rect 390 916 510 950
rect 390 882 433 916
rect 467 882 510 916
rect 390 848 510 882
rect 390 814 433 848
rect 467 814 510 848
rect 390 780 510 814
rect 390 746 433 780
rect 467 746 510 780
rect 390 712 510 746
rect 390 678 433 712
rect 467 678 510 712
rect 390 644 510 678
rect 390 610 433 644
rect 467 610 510 644
rect 390 576 510 610
rect 390 542 433 576
rect 467 542 510 576
rect 390 508 510 542
rect 390 474 433 508
rect 467 474 510 508
rect 390 440 510 474
rect 390 406 433 440
rect 467 406 510 440
rect 390 372 510 406
rect 390 338 433 372
rect 467 338 510 372
rect 390 304 510 338
rect 390 270 433 304
rect 467 270 510 304
rect 390 236 510 270
rect 390 202 433 236
rect 467 202 510 236
rect 390 168 510 202
rect 390 134 433 168
rect 467 134 510 168
rect 390 100 510 134
rect 390 66 433 100
rect 467 66 510 100
rect 390 20 510 66
<< ndiffc >>
rect -1067 950 -1033 984
rect -1067 882 -1033 916
rect -1067 814 -1033 848
rect -1067 746 -1033 780
rect -1067 678 -1033 712
rect -1067 610 -1033 644
rect -1067 542 -1033 576
rect -1067 474 -1033 508
rect -1067 406 -1033 440
rect -1067 338 -1033 372
rect -1067 270 -1033 304
rect -1067 202 -1033 236
rect -1067 134 -1033 168
rect -1067 66 -1033 100
rect -917 950 -883 984
rect -917 882 -883 916
rect -917 814 -883 848
rect -917 746 -883 780
rect -917 678 -883 712
rect -917 610 -883 644
rect -917 542 -883 576
rect -917 474 -883 508
rect -917 406 -883 440
rect -917 338 -883 372
rect -917 270 -883 304
rect -917 202 -883 236
rect -917 134 -883 168
rect -917 66 -883 100
rect -767 950 -733 984
rect -767 882 -733 916
rect -767 814 -733 848
rect -767 746 -733 780
rect -767 678 -733 712
rect -767 610 -733 644
rect -767 542 -733 576
rect -767 474 -733 508
rect -767 406 -733 440
rect -767 338 -733 372
rect -767 270 -733 304
rect -767 202 -733 236
rect -767 134 -733 168
rect -767 66 -733 100
rect -617 950 -583 984
rect -617 882 -583 916
rect -617 814 -583 848
rect -617 746 -583 780
rect -617 678 -583 712
rect -617 610 -583 644
rect -617 542 -583 576
rect -617 474 -583 508
rect -617 406 -583 440
rect -617 338 -583 372
rect -617 270 -583 304
rect -617 202 -583 236
rect -617 134 -583 168
rect -617 66 -583 100
rect -467 950 -433 984
rect -467 882 -433 916
rect -467 814 -433 848
rect -467 746 -433 780
rect -467 678 -433 712
rect -467 610 -433 644
rect -467 542 -433 576
rect -467 474 -433 508
rect -467 406 -433 440
rect -467 338 -433 372
rect -467 270 -433 304
rect -467 202 -433 236
rect -467 134 -433 168
rect -467 66 -433 100
rect -317 950 -283 984
rect -317 882 -283 916
rect -317 814 -283 848
rect -317 746 -283 780
rect -317 678 -283 712
rect -317 610 -283 644
rect -317 542 -283 576
rect -317 474 -283 508
rect -317 406 -283 440
rect -317 338 -283 372
rect -317 270 -283 304
rect -317 202 -283 236
rect -317 134 -283 168
rect -317 66 -283 100
rect -167 950 -133 984
rect -167 882 -133 916
rect -167 814 -133 848
rect -167 746 -133 780
rect -167 678 -133 712
rect -167 610 -133 644
rect -167 542 -133 576
rect -167 474 -133 508
rect -167 406 -133 440
rect -167 338 -133 372
rect -167 270 -133 304
rect -167 202 -133 236
rect -167 134 -133 168
rect -167 66 -133 100
rect -17 950 17 984
rect -17 882 17 916
rect -17 814 17 848
rect -17 746 17 780
rect -17 678 17 712
rect -17 610 17 644
rect -17 542 17 576
rect -17 474 17 508
rect -17 406 17 440
rect -17 338 17 372
rect -17 270 17 304
rect -17 202 17 236
rect -17 134 17 168
rect -17 66 17 100
rect 133 950 167 984
rect 133 882 167 916
rect 133 814 167 848
rect 133 746 167 780
rect 133 678 167 712
rect 133 610 167 644
rect 133 542 167 576
rect 133 474 167 508
rect 133 406 167 440
rect 133 338 167 372
rect 133 270 167 304
rect 133 202 167 236
rect 133 134 167 168
rect 133 66 167 100
rect 283 950 317 984
rect 283 882 317 916
rect 283 814 317 848
rect 283 746 317 780
rect 283 678 317 712
rect 283 610 317 644
rect 283 542 317 576
rect 283 474 317 508
rect 283 406 317 440
rect 283 338 317 372
rect 283 270 317 304
rect 283 202 317 236
rect 283 134 317 168
rect 283 66 317 100
rect 433 950 467 984
rect 433 882 467 916
rect 433 814 467 848
rect 433 746 467 780
rect 433 678 467 712
rect 433 610 467 644
rect 433 542 467 576
rect 433 474 467 508
rect 433 406 467 440
rect 433 338 467 372
rect 433 270 467 304
rect 433 202 467 236
rect 433 134 467 168
rect 433 66 467 100
<< psubdiff >>
rect -1290 984 -1170 1012
rect -1290 950 -1247 984
rect -1213 950 -1170 984
rect -1290 916 -1170 950
rect -1290 882 -1247 916
rect -1213 882 -1170 916
rect -1290 848 -1170 882
rect -1290 814 -1247 848
rect -1213 814 -1170 848
rect -1290 780 -1170 814
rect -1290 746 -1247 780
rect -1213 746 -1170 780
rect -1290 712 -1170 746
rect -1290 678 -1247 712
rect -1213 678 -1170 712
rect -1290 644 -1170 678
rect -1290 610 -1247 644
rect -1213 610 -1170 644
rect -1290 576 -1170 610
rect -1290 542 -1247 576
rect -1213 542 -1170 576
rect -1290 508 -1170 542
rect -1290 474 -1247 508
rect -1213 474 -1170 508
rect -1290 440 -1170 474
rect -1290 406 -1247 440
rect -1213 406 -1170 440
rect -1290 372 -1170 406
rect -1290 338 -1247 372
rect -1213 338 -1170 372
rect -1290 304 -1170 338
rect -1290 270 -1247 304
rect -1213 270 -1170 304
rect -1290 236 -1170 270
rect -1290 202 -1247 236
rect -1213 202 -1170 236
rect -1290 168 -1170 202
rect -1290 134 -1247 168
rect -1213 134 -1170 168
rect -1290 100 -1170 134
rect -1290 66 -1247 100
rect -1213 66 -1170 100
rect -1290 20 -1170 66
<< psubdiffcont >>
rect -1247 950 -1213 984
rect -1247 882 -1213 916
rect -1247 814 -1213 848
rect -1247 746 -1213 780
rect -1247 678 -1213 712
rect -1247 610 -1213 644
rect -1247 542 -1213 576
rect -1247 474 -1213 508
rect -1247 406 -1213 440
rect -1247 338 -1213 372
rect -1247 270 -1213 304
rect -1247 202 -1213 236
rect -1247 134 -1213 168
rect -1247 66 -1213 100
<< poly >>
rect -990 1012 -960 1042
rect -840 1012 -810 1042
rect -690 1012 -660 1043
rect -540 1012 -510 1043
rect -390 1012 -360 1040
rect -240 1012 -210 1043
rect -90 1012 -60 1043
rect 60 1012 90 1042
rect 210 1012 240 1042
rect 360 1012 390 1042
rect -990 -10 -960 20
rect -840 -10 -810 20
rect -690 -10 -660 20
rect -540 -10 -510 20
rect -390 -10 -360 20
rect -240 -10 -210 20
rect -90 -10 -60 20
rect 60 -10 90 20
rect 210 -10 240 20
rect 360 -10 390 20
<< locali >>
rect -1270 984 -1190 990
rect -1270 950 -1247 984
rect -1213 950 -1190 984
rect -1270 916 -1190 950
rect -1270 882 -1247 916
rect -1213 882 -1190 916
rect -1270 848 -1190 882
rect -1270 814 -1247 848
rect -1213 814 -1190 848
rect -1270 780 -1190 814
rect -1270 746 -1247 780
rect -1213 746 -1190 780
rect -1270 712 -1190 746
rect -1270 678 -1247 712
rect -1213 678 -1190 712
rect -1270 644 -1190 678
rect -1270 610 -1247 644
rect -1213 610 -1190 644
rect -1270 576 -1190 610
rect -1270 542 -1247 576
rect -1213 542 -1190 576
rect -1270 508 -1190 542
rect -1270 474 -1247 508
rect -1213 474 -1190 508
rect -1270 440 -1190 474
rect -1270 406 -1247 440
rect -1213 406 -1190 440
rect -1270 372 -1190 406
rect -1270 338 -1247 372
rect -1213 338 -1190 372
rect -1270 304 -1190 338
rect -1270 270 -1247 304
rect -1213 270 -1190 304
rect -1270 236 -1190 270
rect -1270 202 -1247 236
rect -1213 202 -1190 236
rect -1270 168 -1190 202
rect -1270 134 -1247 168
rect -1213 134 -1190 168
rect -1270 100 -1190 134
rect -1270 66 -1247 100
rect -1213 66 -1190 100
rect -1270 40 -1190 66
rect -1090 984 -1010 990
rect -1090 950 -1067 984
rect -1033 950 -1010 984
rect -1090 916 -1010 950
rect -1090 882 -1067 916
rect -1033 882 -1010 916
rect -1090 848 -1010 882
rect -1090 814 -1067 848
rect -1033 814 -1010 848
rect -1090 780 -1010 814
rect -1090 746 -1067 780
rect -1033 746 -1010 780
rect -1090 712 -1010 746
rect -1090 678 -1067 712
rect -1033 678 -1010 712
rect -1090 644 -1010 678
rect -1090 610 -1067 644
rect -1033 610 -1010 644
rect -1090 576 -1010 610
rect -1090 542 -1067 576
rect -1033 542 -1010 576
rect -1090 508 -1010 542
rect -1090 474 -1067 508
rect -1033 474 -1010 508
rect -1090 440 -1010 474
rect -1090 406 -1067 440
rect -1033 406 -1010 440
rect -1090 372 -1010 406
rect -1090 338 -1067 372
rect -1033 338 -1010 372
rect -1090 304 -1010 338
rect -1090 270 -1067 304
rect -1033 270 -1010 304
rect -1090 236 -1010 270
rect -1090 202 -1067 236
rect -1033 202 -1010 236
rect -1090 168 -1010 202
rect -1090 134 -1067 168
rect -1033 134 -1010 168
rect -1090 100 -1010 134
rect -1090 66 -1067 100
rect -1033 66 -1010 100
rect -1090 40 -1010 66
rect -940 984 -860 990
rect -940 950 -917 984
rect -883 950 -860 984
rect -940 916 -860 950
rect -940 882 -917 916
rect -883 882 -860 916
rect -940 848 -860 882
rect -940 814 -917 848
rect -883 814 -860 848
rect -940 780 -860 814
rect -940 746 -917 780
rect -883 746 -860 780
rect -940 712 -860 746
rect -940 678 -917 712
rect -883 678 -860 712
rect -940 644 -860 678
rect -940 610 -917 644
rect -883 610 -860 644
rect -940 576 -860 610
rect -940 542 -917 576
rect -883 542 -860 576
rect -940 508 -860 542
rect -940 474 -917 508
rect -883 474 -860 508
rect -940 440 -860 474
rect -940 406 -917 440
rect -883 406 -860 440
rect -940 372 -860 406
rect -940 338 -917 372
rect -883 338 -860 372
rect -940 304 -860 338
rect -940 270 -917 304
rect -883 270 -860 304
rect -940 236 -860 270
rect -940 202 -917 236
rect -883 202 -860 236
rect -940 168 -860 202
rect -940 134 -917 168
rect -883 134 -860 168
rect -940 100 -860 134
rect -940 66 -917 100
rect -883 66 -860 100
rect -940 40 -860 66
rect -790 984 -710 990
rect -790 950 -767 984
rect -733 950 -710 984
rect -790 916 -710 950
rect -790 882 -767 916
rect -733 882 -710 916
rect -790 848 -710 882
rect -790 814 -767 848
rect -733 814 -710 848
rect -790 780 -710 814
rect -790 746 -767 780
rect -733 746 -710 780
rect -790 712 -710 746
rect -790 678 -767 712
rect -733 678 -710 712
rect -790 644 -710 678
rect -790 610 -767 644
rect -733 610 -710 644
rect -790 576 -710 610
rect -790 542 -767 576
rect -733 542 -710 576
rect -790 508 -710 542
rect -790 474 -767 508
rect -733 474 -710 508
rect -790 440 -710 474
rect -790 406 -767 440
rect -733 406 -710 440
rect -790 372 -710 406
rect -790 338 -767 372
rect -733 338 -710 372
rect -790 304 -710 338
rect -790 270 -767 304
rect -733 270 -710 304
rect -790 236 -710 270
rect -790 202 -767 236
rect -733 202 -710 236
rect -790 168 -710 202
rect -790 134 -767 168
rect -733 134 -710 168
rect -790 100 -710 134
rect -790 66 -767 100
rect -733 66 -710 100
rect -790 40 -710 66
rect -640 984 -560 990
rect -640 950 -617 984
rect -583 950 -560 984
rect -640 916 -560 950
rect -640 882 -617 916
rect -583 882 -560 916
rect -640 848 -560 882
rect -640 814 -617 848
rect -583 814 -560 848
rect -640 780 -560 814
rect -640 746 -617 780
rect -583 746 -560 780
rect -640 712 -560 746
rect -640 678 -617 712
rect -583 678 -560 712
rect -640 644 -560 678
rect -640 610 -617 644
rect -583 610 -560 644
rect -640 576 -560 610
rect -640 542 -617 576
rect -583 542 -560 576
rect -640 508 -560 542
rect -640 474 -617 508
rect -583 474 -560 508
rect -640 440 -560 474
rect -640 406 -617 440
rect -583 406 -560 440
rect -640 372 -560 406
rect -640 338 -617 372
rect -583 338 -560 372
rect -640 304 -560 338
rect -640 270 -617 304
rect -583 270 -560 304
rect -640 236 -560 270
rect -640 202 -617 236
rect -583 202 -560 236
rect -640 168 -560 202
rect -640 134 -617 168
rect -583 134 -560 168
rect -640 100 -560 134
rect -640 66 -617 100
rect -583 66 -560 100
rect -640 40 -560 66
rect -490 984 -410 990
rect -490 950 -467 984
rect -433 950 -410 984
rect -490 916 -410 950
rect -490 882 -467 916
rect -433 882 -410 916
rect -490 848 -410 882
rect -490 814 -467 848
rect -433 814 -410 848
rect -490 780 -410 814
rect -490 746 -467 780
rect -433 746 -410 780
rect -490 712 -410 746
rect -490 678 -467 712
rect -433 678 -410 712
rect -490 644 -410 678
rect -490 610 -467 644
rect -433 610 -410 644
rect -490 576 -410 610
rect -490 542 -467 576
rect -433 542 -410 576
rect -490 508 -410 542
rect -490 474 -467 508
rect -433 474 -410 508
rect -490 440 -410 474
rect -490 406 -467 440
rect -433 406 -410 440
rect -490 372 -410 406
rect -490 338 -467 372
rect -433 338 -410 372
rect -490 304 -410 338
rect -490 270 -467 304
rect -433 270 -410 304
rect -490 236 -410 270
rect -490 202 -467 236
rect -433 202 -410 236
rect -490 168 -410 202
rect -490 134 -467 168
rect -433 134 -410 168
rect -490 100 -410 134
rect -490 66 -467 100
rect -433 66 -410 100
rect -490 40 -410 66
rect -340 984 -260 990
rect -340 950 -317 984
rect -283 950 -260 984
rect -340 916 -260 950
rect -340 882 -317 916
rect -283 882 -260 916
rect -340 848 -260 882
rect -340 814 -317 848
rect -283 814 -260 848
rect -340 780 -260 814
rect -340 746 -317 780
rect -283 746 -260 780
rect -340 712 -260 746
rect -340 678 -317 712
rect -283 678 -260 712
rect -340 644 -260 678
rect -340 610 -317 644
rect -283 610 -260 644
rect -340 576 -260 610
rect -340 542 -317 576
rect -283 542 -260 576
rect -340 508 -260 542
rect -340 474 -317 508
rect -283 474 -260 508
rect -340 440 -260 474
rect -340 406 -317 440
rect -283 406 -260 440
rect -340 372 -260 406
rect -340 338 -317 372
rect -283 338 -260 372
rect -340 304 -260 338
rect -340 270 -317 304
rect -283 270 -260 304
rect -340 236 -260 270
rect -340 202 -317 236
rect -283 202 -260 236
rect -340 168 -260 202
rect -340 134 -317 168
rect -283 134 -260 168
rect -340 100 -260 134
rect -340 66 -317 100
rect -283 66 -260 100
rect -340 40 -260 66
rect -190 984 -110 990
rect -190 950 -167 984
rect -133 950 -110 984
rect -190 916 -110 950
rect -190 882 -167 916
rect -133 882 -110 916
rect -190 848 -110 882
rect -190 814 -167 848
rect -133 814 -110 848
rect -190 780 -110 814
rect -190 746 -167 780
rect -133 746 -110 780
rect -190 712 -110 746
rect -190 678 -167 712
rect -133 678 -110 712
rect -190 644 -110 678
rect -190 610 -167 644
rect -133 610 -110 644
rect -190 576 -110 610
rect -190 542 -167 576
rect -133 542 -110 576
rect -190 508 -110 542
rect -190 474 -167 508
rect -133 474 -110 508
rect -190 440 -110 474
rect -190 406 -167 440
rect -133 406 -110 440
rect -190 372 -110 406
rect -190 338 -167 372
rect -133 338 -110 372
rect -190 304 -110 338
rect -190 270 -167 304
rect -133 270 -110 304
rect -190 236 -110 270
rect -190 202 -167 236
rect -133 202 -110 236
rect -190 168 -110 202
rect -190 134 -167 168
rect -133 134 -110 168
rect -190 100 -110 134
rect -190 66 -167 100
rect -133 66 -110 100
rect -190 40 -110 66
rect -40 984 40 990
rect -40 950 -17 984
rect 17 950 40 984
rect -40 916 40 950
rect -40 882 -17 916
rect 17 882 40 916
rect -40 848 40 882
rect -40 814 -17 848
rect 17 814 40 848
rect -40 780 40 814
rect -40 746 -17 780
rect 17 746 40 780
rect -40 712 40 746
rect -40 678 -17 712
rect 17 678 40 712
rect -40 644 40 678
rect -40 610 -17 644
rect 17 610 40 644
rect -40 576 40 610
rect -40 542 -17 576
rect 17 542 40 576
rect -40 508 40 542
rect -40 474 -17 508
rect 17 474 40 508
rect -40 440 40 474
rect -40 406 -17 440
rect 17 406 40 440
rect -40 372 40 406
rect -40 338 -17 372
rect 17 338 40 372
rect -40 304 40 338
rect -40 270 -17 304
rect 17 270 40 304
rect -40 236 40 270
rect -40 202 -17 236
rect 17 202 40 236
rect -40 168 40 202
rect -40 134 -17 168
rect 17 134 40 168
rect -40 100 40 134
rect -40 66 -17 100
rect 17 66 40 100
rect -40 40 40 66
rect 110 984 190 990
rect 110 950 133 984
rect 167 950 190 984
rect 110 916 190 950
rect 110 882 133 916
rect 167 882 190 916
rect 110 848 190 882
rect 110 814 133 848
rect 167 814 190 848
rect 110 780 190 814
rect 110 746 133 780
rect 167 746 190 780
rect 110 712 190 746
rect 110 678 133 712
rect 167 678 190 712
rect 110 644 190 678
rect 110 610 133 644
rect 167 610 190 644
rect 110 576 190 610
rect 110 542 133 576
rect 167 542 190 576
rect 110 508 190 542
rect 110 474 133 508
rect 167 474 190 508
rect 110 440 190 474
rect 110 406 133 440
rect 167 406 190 440
rect 110 372 190 406
rect 110 338 133 372
rect 167 338 190 372
rect 110 304 190 338
rect 110 270 133 304
rect 167 270 190 304
rect 110 236 190 270
rect 110 202 133 236
rect 167 202 190 236
rect 110 168 190 202
rect 110 134 133 168
rect 167 134 190 168
rect 110 100 190 134
rect 110 66 133 100
rect 167 66 190 100
rect 110 40 190 66
rect 260 984 340 990
rect 260 950 283 984
rect 317 950 340 984
rect 260 916 340 950
rect 260 882 283 916
rect 317 882 340 916
rect 260 848 340 882
rect 260 814 283 848
rect 317 814 340 848
rect 260 780 340 814
rect 260 746 283 780
rect 317 746 340 780
rect 260 712 340 746
rect 260 678 283 712
rect 317 678 340 712
rect 260 644 340 678
rect 260 610 283 644
rect 317 610 340 644
rect 260 576 340 610
rect 260 542 283 576
rect 317 542 340 576
rect 260 508 340 542
rect 260 474 283 508
rect 317 474 340 508
rect 260 440 340 474
rect 260 406 283 440
rect 317 406 340 440
rect 260 372 340 406
rect 260 338 283 372
rect 317 338 340 372
rect 260 304 340 338
rect 260 270 283 304
rect 317 270 340 304
rect 260 236 340 270
rect 260 202 283 236
rect 317 202 340 236
rect 260 168 340 202
rect 260 134 283 168
rect 317 134 340 168
rect 260 100 340 134
rect 260 66 283 100
rect 317 66 340 100
rect 260 40 340 66
rect 410 984 490 990
rect 410 950 433 984
rect 467 950 490 984
rect 410 916 490 950
rect 410 882 433 916
rect 467 882 490 916
rect 410 848 490 882
rect 410 814 433 848
rect 467 814 490 848
rect 410 780 490 814
rect 410 746 433 780
rect 467 746 490 780
rect 410 712 490 746
rect 410 678 433 712
rect 467 678 490 712
rect 410 644 490 678
rect 410 610 433 644
rect 467 610 490 644
rect 410 576 490 610
rect 410 542 433 576
rect 467 542 490 576
rect 410 508 490 542
rect 410 474 433 508
rect 467 474 490 508
rect 410 440 490 474
rect 410 406 433 440
rect 467 406 490 440
rect 410 372 490 406
rect 410 338 433 372
rect 467 338 490 372
rect 410 304 490 338
rect 410 270 433 304
rect 467 270 490 304
rect 410 236 490 270
rect 410 202 433 236
rect 467 202 490 236
rect 410 168 490 202
rect 410 134 433 168
rect 467 134 490 168
rect 410 100 490 134
rect 410 66 433 100
rect 467 66 490 100
rect 410 40 490 66
<< end >>
