magic
tech sky130A
magscale 1 2
timestamp 1680667442
<< locali >>
rect 929 8898 949 8917
rect 930 8800 950 8819
rect 931 8696 951 8715
rect 928 8599 948 8618
rect 928 7103 948 7122
rect 927 7000 947 7019
rect 926 6897 946 6916
rect 933 6795 953 6815
rect 929 6538 949 6558
rect 928 6440 948 6459
rect 932 6338 952 6357
rect 927 6239 947 6258
rect 927 4737 947 4756
rect 928 4639 948 4658
rect 928 4538 948 4557
rect 928 4438 948 4458
rect 951 -17102 971 -17082
rect 954 -17203 974 -17184
rect 952 -17300 972 -17281
rect 954 -17404 974 -17385
rect 932 -18903 952 -18884
rect 948 -19006 968 -18987
rect 952 -19104 972 -19085
rect 929 -19207 949 -19187
rect 945 -19465 965 -19445
rect 948 -19564 968 -19545
rect 952 -19662 972 -19643
rect 943 -19763 963 -19744
rect 949 -21266 969 -21247
rect 950 -21362 970 -21343
rect 949 -21464 969 -21445
rect 953 -21564 973 -21544
rect 946 -21902 966 -21882
rect 950 -22004 970 -21985
rect 953 -22101 973 -22082
rect 950 -22200 970 -22181
rect 949 -23704 969 -23685
rect 951 -23801 971 -23782
rect 950 -23899 970 -23880
rect 948 -24003 968 -23983
rect 949 -24269 969 -24249
rect 955 -24361 975 -24342
rect 948 -24462 968 -24443
rect 951 -24565 971 -24546
rect 949 -26063 969 -26044
rect 953 -26165 973 -26146
rect 956 -26263 976 -26244
rect 951 -26365 971 -26345
rect 949 -47903 969 -47883
rect 946 -48003 966 -47984
rect 947 -48104 967 -48085
rect 947 -48202 967 -48183
rect 947 -49707 967 -49688
rect 947 -49804 967 -49785
rect 948 -49905 968 -49886
rect 947 -50007 967 -49987
rect 948 -50266 968 -50246
rect 948 -50365 968 -50346
rect 947 -50465 967 -50446
rect 947 -50568 967 -50549
rect 949 -52066 969 -52047
rect 953 -52164 973 -52145
rect 948 -52266 968 -52247
rect 950 -52364 970 -52344
rect 943 -52708 963 -52688
rect 947 -52807 967 -52788
rect 943 -52907 963 -52888
rect 944 -53007 964 -52988
rect 945 -54506 965 -54487
rect 950 -54604 970 -54585
rect 948 -54702 968 -54683
rect 949 -54806 969 -54786
rect 952 -55066 972 -55046
rect 954 -55162 974 -55143
rect 951 -55262 971 -55243
rect 950 -55362 970 -55343
rect 948 -56866 968 -56847
rect 949 -56968 969 -56949
rect 946 -57064 966 -57045
rect 949 -57165 969 -57145
rect 950 -78707 970 -78687
rect 950 -78807 970 -78788
rect 943 -78909 963 -78890
rect 945 -79009 965 -78990
rect 945 -80509 965 -80490
rect 949 -80606 969 -80587
rect 947 -80706 967 -80687
rect 954 -80810 974 -80790
rect 949 -81067 969 -81047
rect 948 -81166 968 -81147
rect 951 -81266 971 -81247
rect 948 -81369 968 -81350
rect 952 -82867 972 -82848
rect 950 -82965 970 -82946
rect 953 -83068 973 -83048
rect 951 -83168 971 -83149
rect 949 -83510 969 -83491
rect 945 -83609 965 -83589
rect 947 -83703 967 -83684
rect 948 -83809 968 -83790
rect 949 -85303 969 -85284
rect 946 -85407 966 -85388
rect 946 -85508 966 -85488
rect 946 -85606 966 -85587
rect 946 -85865 966 -85846
rect 943 -85967 963 -85947
rect 946 -86066 966 -86047
rect 946 -86164 966 -86145
rect 952 -87667 972 -87648
rect 948 -87770 968 -87751
rect 949 -87867 969 -87847
rect 948 -87968 968 -87949
rect 950 -109508 970 -109489
rect 947 -109610 967 -109590
rect 947 -109710 967 -109691
rect 947 -109804 967 -109785
rect 955 -111312 975 -111293
rect 949 -111410 969 -111391
rect 951 -111507 971 -111487
rect 950 -111607 970 -111588
rect 956 -111870 976 -111850
rect 955 -111968 975 -111949
rect 948 -112070 968 -112051
rect 945 -112171 965 -112152
rect 954 -113670 974 -113651
rect 955 -113772 975 -113753
rect 954 -113868 974 -113848
rect 949 -113969 969 -113950
rect 951 -114308 971 -114288
rect 947 -114409 967 -114390
rect 949 -114510 969 -114491
rect 950 -114608 970 -114589
rect 952 -116107 972 -116088
rect 948 -116210 968 -116191
rect 944 -116309 964 -116290
rect 951 -116410 971 -116390
rect 946 -116670 966 -116650
rect 949 -116765 969 -116746
rect 953 -116867 973 -116848
rect 951 -116969 971 -116950
rect 950 -118472 970 -118453
rect 948 -118567 968 -118548
rect 946 -118668 966 -118648
rect 951 -118769 971 -118750
rect 953 -140310 973 -140291
rect 944 -140411 964 -140391
rect 949 -140508 969 -140489
rect 945 -140608 965 -140589
rect 957 -142113 977 -142094
rect 946 -142215 966 -142196
rect 945 -142310 965 -142290
rect 943 -142412 963 -142393
rect 950 -142673 970 -142654
rect 950 -142773 970 -142753
rect 951 -142874 971 -142855
rect 948 -142972 968 -142953
rect 947 -144473 967 -144454
rect 949 -144572 969 -144553
rect 949 -144675 969 -144655
rect 949 -144773 969 -144754
rect 950 -145112 970 -145093
rect 951 -145210 971 -145190
rect 945 -145311 965 -145292
rect 945 -145411 965 -145392
rect 949 -146910 969 -146891
rect 954 -147006 974 -146987
rect 948 -147110 968 -147090
rect 950 -147213 970 -147194
rect 947 -147474 967 -147455
rect 946 -147571 966 -147551
rect 943 -147672 963 -147653
rect 946 -147770 966 -147751
rect 948 -149271 968 -149252
rect 949 -149370 969 -149351
rect 946 -149474 966 -149455
rect 947 -149571 967 -149551
rect 948 -171113 968 -171093
rect 948 -171213 968 -171194
rect 948 -171314 968 -171295
rect 944 -171413 964 -171394
rect 946 -172913 966 -172894
rect 948 -173013 968 -172994
rect 947 -173115 967 -173096
rect 949 -173213 969 -173193
rect 945 -173474 965 -173454
rect 949 -173574 969 -173555
rect 946 -173676 966 -173657
rect 946 -173773 966 -173754
rect 949 -175272 969 -175253
rect 953 -175371 973 -175352
rect 948 -175474 968 -175455
rect 947 -175576 967 -175556
rect 951 -175911 971 -175892
rect 947 -176014 967 -175994
rect 950 -176112 970 -176093
rect 943 -176210 963 -176191
rect 951 -177713 971 -177694
rect 949 -177814 969 -177795
rect 945 -177912 965 -177893
rect 951 -178013 971 -177993
rect 944 -178274 964 -178254
rect 946 -178372 966 -178353
rect 948 -178477 968 -178458
rect 943 -178570 963 -178551
rect 944 -180073 964 -180054
rect 950 -180170 970 -180151
rect 950 -180276 970 -180256
rect 947 -180374 967 -180355
rect 945 -201915 965 -201895
rect 949 -202015 969 -201996
rect 947 -202115 967 -202096
rect 948 -202215 968 -202196
rect 947 -203716 967 -203697
rect 948 -203815 968 -203796
rect 946 -203916 966 -203897
rect 947 -204015 967 -203995
rect 950 -204274 970 -204254
rect 948 -204375 968 -204356
rect 947 -204475 967 -204456
rect 952 -204576 972 -204557
rect 949 -206074 969 -206055
rect 947 -206178 967 -206159
rect 949 -206276 969 -206256
rect 947 -206376 967 -206357
rect 955 -206715 975 -206695
rect 950 -206815 970 -206796
rect 952 -206914 972 -206895
rect 946 -207015 966 -206996
rect 945 -208513 965 -208494
rect 950 -208614 970 -208595
rect 951 -208714 971 -208695
rect 948 -208814 968 -208794
rect 948 -209074 968 -209054
rect 946 -209173 966 -209154
rect 947 -209273 967 -209254
rect 946 -209373 966 -209354
rect 948 -210875 968 -210856
rect 954 -210973 974 -210954
rect 949 -211076 969 -211056
rect 948 -211174 968 -211155
rect 950 -232718 970 -232699
rect 948 -232817 968 -232797
rect 949 -232917 969 -232898
rect 948 -233016 968 -232997
rect 948 -234519 968 -234500
rect 947 -234617 967 -234598
rect 948 -234718 968 -234699
rect 948 -234818 968 -234798
rect 949 -235076 969 -235056
rect 948 -235179 968 -235160
rect 947 -235278 967 -235259
rect 948 -235379 968 -235360
rect 945 -236876 965 -236857
rect 948 -236979 968 -236960
rect 950 -237079 970 -237060
rect 949 -237179 969 -237159
<< metal1 >>
rect 945 7841 979 7875
<< via1 >>
rect 2864 4292 2916 4344
rect 2944 4292 2996 4344
rect 3024 4292 3076 4344
rect 8221 -5949 8273 -5897
rect 8701 -5949 8753 -5897
rect 8221 -6029 8273 -5977
rect 8701 -6029 8753 -5977
rect 8221 -6109 8273 -6057
rect 8701 -6109 8753 -6057
rect 8221 -6589 8273 -6537
rect 8701 -6589 8753 -6537
rect 8221 -6669 8273 -6617
rect 8701 -6669 8753 -6617
rect 8221 -6749 8273 -6697
rect 8701 -6749 8753 -6697
rect 2864 -16990 2916 -16938
rect 2944 -16990 2996 -16938
rect 3024 -16990 3076 -16938
rect 2864 -26510 2916 -26458
rect 2944 -26510 2996 -26458
rect 3024 -26510 3076 -26458
rect 8221 -36751 8273 -36699
rect 8701 -36751 8753 -36699
rect 8221 -36831 8273 -36779
rect 8701 -36831 8753 -36779
rect 8221 -36911 8273 -36859
rect 8701 -36911 8753 -36859
rect 8221 -37391 8273 -37339
rect 8701 -37391 8753 -37339
rect 8221 -37471 8273 -37419
rect 8701 -37471 8753 -37419
rect 8221 -37551 8273 -37499
rect 8701 -37551 8753 -37499
rect 2864 -47792 2916 -47740
rect 2944 -47792 2996 -47740
rect 3024 -47792 3076 -47740
rect 2864 -57312 2916 -57260
rect 2944 -57312 2996 -57260
rect 3024 -57312 3076 -57260
rect 8221 -67553 8273 -67501
rect 8701 -67553 8753 -67501
rect 8221 -67633 8273 -67581
rect 8701 -67633 8753 -67581
rect 8221 -67713 8273 -67661
rect 8701 -67713 8753 -67661
rect 8221 -68193 8273 -68141
rect 8701 -68193 8753 -68141
rect 8221 -68273 8273 -68221
rect 8701 -68273 8753 -68221
rect 8221 -68353 8273 -68301
rect 8701 -68353 8753 -68301
rect 2864 -78594 2916 -78542
rect 2944 -78594 2996 -78542
rect 3024 -78594 3076 -78542
rect 2864 -88114 2916 -88062
rect 2944 -88114 2996 -88062
rect 3024 -88114 3076 -88062
rect 8221 -98355 8273 -98303
rect 8701 -98355 8753 -98303
rect 8221 -98435 8273 -98383
rect 8701 -98435 8753 -98383
rect 8221 -98515 8273 -98463
rect 8701 -98515 8753 -98463
rect 8221 -98995 8273 -98943
rect 8701 -98995 8753 -98943
rect 8221 -99075 8273 -99023
rect 8701 -99075 8753 -99023
rect 8221 -99155 8273 -99103
rect 8701 -99155 8753 -99103
rect 2864 -109396 2916 -109344
rect 2944 -109396 2996 -109344
rect 3024 -109396 3076 -109344
rect 2864 -118916 2916 -118864
rect 2944 -118916 2996 -118864
rect 3024 -118916 3076 -118864
rect 8221 -129157 8273 -129105
rect 8701 -129157 8753 -129105
rect 8221 -129237 8273 -129185
rect 8701 -129237 8753 -129185
rect 8221 -129317 8273 -129265
rect 8701 -129317 8753 -129265
rect 8221 -129797 8273 -129745
rect 8701 -129797 8753 -129745
rect 8221 -129877 8273 -129825
rect 8701 -129877 8753 -129825
rect 8221 -129957 8273 -129905
rect 8701 -129957 8753 -129905
rect 2864 -140198 2916 -140146
rect 2944 -140198 2996 -140146
rect 3024 -140198 3076 -140146
rect 2864 -149718 2916 -149666
rect 2944 -149718 2996 -149666
rect 3024 -149718 3076 -149666
rect 8221 -159959 8273 -159907
rect 8701 -159959 8753 -159907
rect 8221 -160039 8273 -159987
rect 8701 -160039 8753 -159987
rect 8221 -160119 8273 -160067
rect 8701 -160119 8753 -160067
rect 8221 -160599 8273 -160547
rect 8701 -160599 8753 -160547
rect 8221 -160679 8273 -160627
rect 8701 -160679 8753 -160627
rect 8221 -160759 8273 -160707
rect 8701 -160759 8753 -160707
rect 2864 -171000 2916 -170948
rect 2944 -171000 2996 -170948
rect 3024 -171000 3076 -170948
rect 2864 -180520 2916 -180468
rect 2944 -180520 2996 -180468
rect 3024 -180520 3076 -180468
rect 8221 -190761 8273 -190709
rect 8701 -190761 8753 -190709
rect 8221 -190841 8273 -190789
rect 8701 -190841 8753 -190789
rect 8221 -190921 8273 -190869
rect 8701 -190921 8753 -190869
rect 8221 -191401 8273 -191349
rect 8701 -191401 8753 -191349
rect 8221 -191481 8273 -191429
rect 8701 -191481 8753 -191429
rect 8221 -191561 8273 -191509
rect 8701 -191561 8753 -191509
rect 2864 -201802 2916 -201750
rect 2944 -201802 2996 -201750
rect 3024 -201802 3076 -201750
rect 2864 -211322 2916 -211270
rect 2944 -211322 2996 -211270
rect 3024 -211322 3076 -211270
rect 8221 -221563 8273 -221511
rect 8701 -221563 8753 -221511
rect 8221 -221643 8273 -221591
rect 8701 -221643 8753 -221591
rect 8221 -221723 8273 -221671
rect 8701 -221723 8753 -221671
rect 8221 -222203 8273 -222151
rect 8701 -222203 8753 -222151
rect 8221 -222283 8273 -222231
rect 8701 -222283 8753 -222231
rect 8221 -222363 8273 -222311
rect 8701 -222363 8753 -222311
rect 2864 -232604 2916 -232552
rect 2944 -232604 2996 -232552
rect 3024 -232604 3076 -232552
<< metal2 >>
rect 1113 9021 1147 9055
rect 1231 9022 1261 9054
rect 4444 9020 4485 9062
rect 4566 9027 4586 9048
rect 8892 9025 8917 9053
rect 9172 9021 9203 9055
rect 9255 9021 9296 9064
rect 9355 9028 9383 9058
rect 10877 7287 10898 7309
rect 10876 7167 10897 7189
rect 1206 -17974 1286 5328
rect 2840 4344 3090 4358
rect 2840 4292 2864 4344
rect 2916 4292 2944 4344
rect 2996 4292 3024 4344
rect 3076 4292 3090 4344
rect 2840 -16938 3090 4292
rect 10653 2870 10674 2892
rect 10652 2766 10673 2788
rect 10913 1586 10934 1608
rect 10919 1459 10940 1481
rect 4461 -7462 4541 -5184
rect 10652 -5670 10674 -5650
rect 10652 -5672 10673 -5670
rect 10653 -5776 10674 -5754
rect 8207 -5897 8287 -5873
rect 8207 -5949 8221 -5897
rect 8273 -5949 8287 -5897
rect 8207 -5977 8287 -5949
rect 8207 -6029 8221 -5977
rect 8273 -6029 8287 -5977
rect 8207 -6057 8287 -6029
rect 8207 -6109 8221 -6057
rect 8273 -6109 8287 -6057
rect 4577 -6403 4657 -6243
rect 8207 -6537 8287 -6109
rect 8207 -6589 8221 -6537
rect 8273 -6589 8287 -6537
rect 8207 -6617 8287 -6589
rect 8207 -6669 8221 -6617
rect 8273 -6669 8287 -6617
rect 8207 -6697 8287 -6669
rect 8207 -6749 8221 -6697
rect 8273 -6749 8287 -6697
rect 8207 -6773 8287 -6749
rect 8390 -5967 8404 -5887
rect 8687 -5897 8767 -5873
rect 8687 -5949 8701 -5897
rect 8753 -5949 8767 -5897
rect 8390 -6679 8470 -5967
rect 8687 -5977 8767 -5949
rect 8687 -6029 8701 -5977
rect 8753 -6029 8767 -5977
rect 8687 -6057 8767 -6029
rect 8687 -6109 8701 -6057
rect 8753 -6109 8767 -6057
rect 8498 -6401 8578 -6245
rect 8687 -6537 8767 -6109
rect 8687 -6589 8701 -6537
rect 8753 -6589 8767 -6537
rect 8687 -6617 8767 -6589
rect 8687 -6669 8701 -6617
rect 8753 -6669 8767 -6617
rect 8390 -6759 8404 -6679
rect 8687 -6697 8767 -6669
rect 8687 -6749 8701 -6697
rect 8753 -6749 8767 -6697
rect 8687 -6773 8767 -6749
rect 10637 -6873 10658 -6869
rect 10637 -6891 10676 -6873
rect 10656 -6892 10676 -6891
rect 10636 -6976 10657 -6974
rect 10636 -6996 10674 -6976
rect 10882 -14127 10903 -14105
rect 10878 -14256 10899 -14234
rect 10610 -15434 10631 -15412
rect 10610 -15538 10631 -15516
rect 2840 -16990 2864 -16938
rect 2916 -16990 2944 -16938
rect 2996 -16990 3024 -16938
rect 3076 -16990 3090 -16938
rect 2840 -17004 3090 -16990
rect 10844 -19834 10865 -19812
rect 10838 -19954 10859 -19932
rect 10838 -23515 10859 -23493
rect 10841 -23636 10862 -23614
rect 1206 -48776 1286 -25474
rect 2840 -26458 3090 -26444
rect 2840 -26510 2864 -26458
rect 2916 -26510 2944 -26458
rect 2996 -26510 3024 -26458
rect 3076 -26510 3090 -26458
rect 2840 -47740 3090 -26510
rect 10610 -27931 10631 -27909
rect 10613 -28036 10634 -28014
rect 10877 -29215 10898 -29193
rect 10880 -29340 10901 -29318
rect 4461 -38264 4541 -35986
rect 10616 -36470 10637 -36448
rect 10617 -36578 10638 -36556
rect 8207 -36699 8287 -36675
rect 8207 -36751 8221 -36699
rect 8273 -36751 8287 -36699
rect 8207 -36779 8287 -36751
rect 8207 -36831 8221 -36779
rect 8273 -36831 8287 -36779
rect 8207 -36859 8287 -36831
rect 8207 -36911 8221 -36859
rect 8273 -36911 8287 -36859
rect 4577 -37205 4657 -37045
rect 8207 -37339 8287 -36911
rect 8207 -37391 8221 -37339
rect 8273 -37391 8287 -37339
rect 8207 -37419 8287 -37391
rect 8207 -37471 8221 -37419
rect 8273 -37471 8287 -37419
rect 8207 -37499 8287 -37471
rect 8207 -37551 8221 -37499
rect 8273 -37551 8287 -37499
rect 8207 -37575 8287 -37551
rect 8390 -36769 8404 -36689
rect 8687 -36699 8767 -36675
rect 8687 -36751 8701 -36699
rect 8753 -36751 8767 -36699
rect 8390 -37481 8470 -36769
rect 8687 -36779 8767 -36751
rect 8687 -36831 8701 -36779
rect 8753 -36831 8767 -36779
rect 8687 -36859 8767 -36831
rect 8687 -36911 8701 -36859
rect 8753 -36911 8767 -36859
rect 8498 -37203 8578 -37047
rect 8687 -37339 8767 -36911
rect 8687 -37391 8701 -37339
rect 8753 -37391 8767 -37339
rect 8687 -37419 8767 -37391
rect 8687 -37471 8701 -37419
rect 8753 -37471 8767 -37419
rect 8390 -37561 8404 -37481
rect 8687 -37499 8767 -37471
rect 8687 -37551 8701 -37499
rect 8753 -37551 8767 -37499
rect 8687 -37575 8767 -37551
rect 10653 -37695 10674 -37673
rect 10651 -37799 10672 -37777
rect 10879 -44933 10900 -44911
rect 10878 -45058 10899 -45036
rect 10612 -46234 10633 -46212
rect 10611 -46340 10632 -46318
rect 2840 -47792 2864 -47740
rect 2916 -47792 2944 -47740
rect 2996 -47792 3024 -47740
rect 3076 -47792 3090 -47740
rect 2840 -47806 3090 -47792
rect 10843 -50635 10864 -50613
rect 10842 -50758 10863 -50736
rect 10840 -54315 10861 -54293
rect 10839 -54440 10860 -54418
rect 1206 -79578 1286 -56276
rect 2840 -57260 3090 -57246
rect 2840 -57312 2864 -57260
rect 2916 -57312 2944 -57260
rect 2996 -57312 3024 -57260
rect 3076 -57312 3090 -57260
rect 2840 -78542 3090 -57312
rect 10610 -58733 10631 -58711
rect 10613 -58839 10634 -58817
rect 10879 -60014 10900 -59992
rect 10883 -60143 10904 -60121
rect 4461 -69066 4541 -66788
rect 10612 -67274 10633 -67252
rect 10615 -67379 10636 -67357
rect 8207 -67501 8287 -67477
rect 8207 -67553 8221 -67501
rect 8273 -67553 8287 -67501
rect 8207 -67581 8287 -67553
rect 8207 -67633 8221 -67581
rect 8273 -67633 8287 -67581
rect 8207 -67661 8287 -67633
rect 8207 -67713 8221 -67661
rect 8273 -67713 8287 -67661
rect 4577 -68007 4657 -67847
rect 8207 -68141 8287 -67713
rect 8207 -68193 8221 -68141
rect 8273 -68193 8287 -68141
rect 8207 -68221 8287 -68193
rect 8207 -68273 8221 -68221
rect 8273 -68273 8287 -68221
rect 8207 -68301 8287 -68273
rect 8207 -68353 8221 -68301
rect 8273 -68353 8287 -68301
rect 8207 -68377 8287 -68353
rect 8390 -67571 8404 -67491
rect 8687 -67501 8767 -67477
rect 8687 -67553 8701 -67501
rect 8753 -67553 8767 -67501
rect 8390 -68283 8470 -67571
rect 8687 -67581 8767 -67553
rect 8687 -67633 8701 -67581
rect 8753 -67633 8767 -67581
rect 8687 -67661 8767 -67633
rect 8687 -67713 8701 -67661
rect 8753 -67713 8767 -67661
rect 8498 -68005 8578 -67849
rect 8687 -68141 8767 -67713
rect 8687 -68193 8701 -68141
rect 8753 -68193 8767 -68141
rect 8687 -68221 8767 -68193
rect 8687 -68273 8701 -68221
rect 8753 -68273 8767 -68221
rect 8390 -68363 8404 -68283
rect 8687 -68301 8767 -68273
rect 8687 -68353 8701 -68301
rect 8753 -68353 8767 -68301
rect 8687 -68377 8767 -68353
rect 10614 -68497 10635 -68475
rect 10615 -68600 10636 -68578
rect 10882 -75732 10903 -75710
rect 10875 -75858 10896 -75836
rect 10611 -77023 10631 -77017
rect 10611 -77036 10639 -77023
rect 10618 -77045 10639 -77036
rect 10611 -77129 10630 -77122
rect 10611 -77141 10638 -77129
rect 10617 -77151 10638 -77141
rect 2840 -78594 2864 -78542
rect 2916 -78594 2944 -78542
rect 2996 -78594 3024 -78542
rect 3076 -78594 3090 -78542
rect 2840 -78608 3090 -78594
rect 10843 -81438 10864 -81416
rect 10840 -81559 10861 -81537
rect 10842 -85118 10863 -85096
rect 10841 -85239 10862 -85217
rect 1206 -110380 1286 -87078
rect 2840 -88062 3090 -88048
rect 2840 -88114 2864 -88062
rect 2916 -88114 2944 -88062
rect 2996 -88114 3024 -88062
rect 3076 -88114 3090 -88062
rect 2840 -109344 3090 -88114
rect 10606 -89535 10627 -89513
rect 10613 -89621 10634 -89618
rect 10611 -89640 10634 -89621
rect 10880 -90799 10901 -90796
rect 10876 -90818 10901 -90799
rect 10876 -90819 10896 -90818
rect 10883 -90944 10904 -90922
rect 4461 -99868 4541 -97590
rect 10614 -98074 10637 -98054
rect 10616 -98076 10637 -98074
rect 10618 -98181 10639 -98159
rect 8207 -98303 8287 -98279
rect 8207 -98355 8221 -98303
rect 8273 -98355 8287 -98303
rect 8207 -98383 8287 -98355
rect 8207 -98435 8221 -98383
rect 8273 -98435 8287 -98383
rect 8207 -98463 8287 -98435
rect 8207 -98515 8221 -98463
rect 8273 -98515 8287 -98463
rect 4577 -98809 4657 -98649
rect 8207 -98943 8287 -98515
rect 8207 -98995 8221 -98943
rect 8273 -98995 8287 -98943
rect 8207 -99023 8287 -98995
rect 8207 -99075 8221 -99023
rect 8273 -99075 8287 -99023
rect 8207 -99103 8287 -99075
rect 8207 -99155 8221 -99103
rect 8273 -99155 8287 -99103
rect 8207 -99179 8287 -99155
rect 8390 -98373 8404 -98293
rect 8687 -98303 8767 -98279
rect 8687 -98355 8701 -98303
rect 8753 -98355 8767 -98303
rect 8390 -99085 8470 -98373
rect 8687 -98383 8767 -98355
rect 8687 -98435 8701 -98383
rect 8753 -98435 8767 -98383
rect 8687 -98463 8767 -98435
rect 8687 -98515 8701 -98463
rect 8753 -98515 8767 -98463
rect 8498 -98807 8578 -98651
rect 8687 -98943 8767 -98515
rect 8687 -98995 8701 -98943
rect 8753 -98995 8767 -98943
rect 8687 -99023 8767 -98995
rect 8687 -99075 8701 -99023
rect 8753 -99075 8767 -99023
rect 8390 -99165 8404 -99085
rect 8687 -99103 8767 -99075
rect 8687 -99155 8701 -99103
rect 8753 -99155 8767 -99103
rect 8687 -99179 8767 -99155
rect 10615 -99299 10636 -99277
rect 10614 -99402 10635 -99380
rect 10880 -106534 10901 -106512
rect 10879 -106661 10900 -106639
rect 10610 -107819 10631 -107818
rect 10609 -107838 10631 -107819
rect 10610 -107840 10631 -107838
rect 10609 -107946 10630 -107924
rect 2840 -109396 2864 -109344
rect 2916 -109396 2944 -109344
rect 2996 -109396 3024 -109344
rect 3076 -109396 3090 -109344
rect 2840 -109410 3090 -109396
rect 10841 -112239 10862 -112217
rect 10842 -112360 10863 -112338
rect 10837 -115921 10858 -115899
rect 10840 -116043 10861 -116021
rect 1206 -141182 1286 -117880
rect 2840 -118864 3090 -118850
rect 2840 -118916 2864 -118864
rect 2916 -118916 2944 -118864
rect 2996 -118916 3024 -118864
rect 3076 -118916 3090 -118864
rect 2840 -140146 3090 -118916
rect 10607 -120336 10628 -120314
rect 10612 -120442 10633 -120420
rect 10876 -121620 10897 -121598
rect 10877 -121745 10898 -121723
rect 4461 -130670 4541 -128392
rect 10616 -128879 10637 -128857
rect 10614 -128984 10635 -128962
rect 8207 -129105 8287 -129081
rect 8207 -129157 8221 -129105
rect 8273 -129157 8287 -129105
rect 8207 -129185 8287 -129157
rect 8207 -129237 8221 -129185
rect 8273 -129237 8287 -129185
rect 8207 -129265 8287 -129237
rect 8207 -129317 8221 -129265
rect 8273 -129317 8287 -129265
rect 4577 -129611 4657 -129451
rect 8207 -129745 8287 -129317
rect 8207 -129797 8221 -129745
rect 8273 -129797 8287 -129745
rect 8207 -129825 8287 -129797
rect 8207 -129877 8221 -129825
rect 8273 -129877 8287 -129825
rect 8207 -129905 8287 -129877
rect 8207 -129957 8221 -129905
rect 8273 -129957 8287 -129905
rect 8207 -129981 8287 -129957
rect 8390 -129175 8404 -129095
rect 8687 -129105 8767 -129081
rect 8687 -129157 8701 -129105
rect 8753 -129157 8767 -129105
rect 8390 -129887 8470 -129175
rect 8687 -129185 8767 -129157
rect 8687 -129237 8701 -129185
rect 8753 -129237 8767 -129185
rect 8687 -129265 8767 -129237
rect 8687 -129317 8701 -129265
rect 8753 -129317 8767 -129265
rect 8498 -129609 8578 -129453
rect 8687 -129745 8767 -129317
rect 8687 -129797 8701 -129745
rect 8753 -129797 8767 -129745
rect 8687 -129825 8767 -129797
rect 8687 -129877 8701 -129825
rect 8753 -129877 8767 -129825
rect 8390 -129967 8404 -129887
rect 8687 -129905 8767 -129877
rect 8687 -129957 8701 -129905
rect 8753 -129957 8767 -129905
rect 8687 -129981 8767 -129957
rect 10613 -130099 10634 -130077
rect 10612 -130205 10633 -130183
rect 10880 -137336 10901 -137314
rect 10877 -137462 10898 -137440
rect 10611 -138641 10632 -138619
rect 10610 -138747 10631 -138725
rect 2840 -140198 2864 -140146
rect 2916 -140198 2944 -140146
rect 2996 -140198 3024 -140146
rect 3076 -140198 3090 -140146
rect 2840 -140212 3090 -140198
rect 10838 -143042 10859 -143020
rect 10839 -143164 10860 -143142
rect 10836 -146722 10857 -146700
rect 10837 -146844 10858 -146822
rect 1206 -171984 1286 -148682
rect 2840 -149666 3090 -149652
rect 2840 -149718 2864 -149666
rect 2916 -149718 2944 -149666
rect 2996 -149718 3024 -149666
rect 3076 -149718 3090 -149666
rect 2840 -170948 3090 -149718
rect 10608 -151139 10629 -151117
rect 10611 -151244 10632 -151222
rect 10878 -152423 10899 -152401
rect 10878 -152549 10899 -152527
rect 4461 -161472 4541 -159194
rect 10611 -159680 10632 -159658
rect 10616 -159786 10637 -159764
rect 8207 -159907 8287 -159883
rect 8207 -159959 8221 -159907
rect 8273 -159959 8287 -159907
rect 8207 -159987 8287 -159959
rect 8207 -160039 8221 -159987
rect 8273 -160039 8287 -159987
rect 8207 -160067 8287 -160039
rect 8207 -160119 8221 -160067
rect 8273 -160119 8287 -160067
rect 4577 -160413 4657 -160253
rect 8207 -160547 8287 -160119
rect 8207 -160599 8221 -160547
rect 8273 -160599 8287 -160547
rect 8207 -160627 8287 -160599
rect 8207 -160679 8221 -160627
rect 8273 -160679 8287 -160627
rect 8207 -160707 8287 -160679
rect 8207 -160759 8221 -160707
rect 8273 -160759 8287 -160707
rect 8207 -160783 8287 -160759
rect 8390 -159977 8404 -159897
rect 8687 -159907 8767 -159883
rect 8687 -159959 8701 -159907
rect 8753 -159959 8767 -159907
rect 8390 -160689 8470 -159977
rect 8687 -159987 8767 -159959
rect 8687 -160039 8701 -159987
rect 8753 -160039 8767 -159987
rect 8687 -160067 8767 -160039
rect 8687 -160119 8701 -160067
rect 8753 -160119 8767 -160067
rect 8498 -160411 8578 -160255
rect 8687 -160547 8767 -160119
rect 8687 -160599 8701 -160547
rect 8753 -160599 8767 -160547
rect 8687 -160627 8767 -160599
rect 8687 -160679 8701 -160627
rect 8753 -160679 8767 -160627
rect 8390 -160769 8404 -160689
rect 8687 -160707 8767 -160679
rect 8687 -160759 8701 -160707
rect 8753 -160759 8767 -160707
rect 8687 -160783 8767 -160759
rect 10615 -160900 10637 -160880
rect 10616 -160902 10637 -160900
rect 10614 -161007 10635 -160985
rect 10881 -168118 10902 -168117
rect 10881 -168137 10903 -168118
rect 10881 -168139 10902 -168137
rect 10878 -168265 10899 -168243
rect 10611 -169443 10632 -169421
rect 10610 -169549 10631 -169527
rect 2840 -171000 2864 -170948
rect 2916 -171000 2944 -170948
rect 2996 -171000 3024 -170948
rect 3076 -171000 3090 -170948
rect 2840 -171014 3090 -171000
rect 10839 -173824 10860 -173822
rect 10839 -173843 10861 -173824
rect 10839 -173844 10860 -173843
rect 10840 -173965 10861 -173943
rect 10840 -177526 10861 -177504
rect 10841 -177646 10862 -177624
rect 1206 -202786 1286 -179484
rect 2840 -180468 3090 -180454
rect 2840 -180520 2864 -180468
rect 2916 -180520 2944 -180468
rect 2996 -180520 3024 -180468
rect 3076 -180520 3090 -180468
rect 2840 -201750 3090 -180520
rect 10608 -181941 10629 -181919
rect 10611 -182046 10632 -182024
rect 10878 -183212 10898 -183205
rect 10878 -183225 10905 -183212
rect 10884 -183234 10905 -183225
rect 10883 -183338 10902 -183330
rect 10883 -183349 10908 -183338
rect 10887 -183360 10908 -183349
rect 4461 -192274 4541 -189996
rect 10615 -190483 10636 -190460
rect 10616 -190588 10637 -190566
rect 8207 -190709 8287 -190685
rect 8207 -190761 8221 -190709
rect 8273 -190761 8287 -190709
rect 8207 -190789 8287 -190761
rect 8207 -190841 8221 -190789
rect 8273 -190841 8287 -190789
rect 8207 -190869 8287 -190841
rect 8207 -190921 8221 -190869
rect 8273 -190921 8287 -190869
rect 4577 -191215 4657 -191055
rect 8207 -191349 8287 -190921
rect 8207 -191401 8221 -191349
rect 8273 -191401 8287 -191349
rect 8207 -191429 8287 -191401
rect 8207 -191481 8221 -191429
rect 8273 -191481 8287 -191429
rect 8207 -191509 8287 -191481
rect 8207 -191561 8221 -191509
rect 8273 -191561 8287 -191509
rect 8207 -191585 8287 -191561
rect 8390 -190779 8404 -190699
rect 8687 -190709 8767 -190685
rect 8687 -190761 8701 -190709
rect 8753 -190761 8767 -190709
rect 8390 -191491 8470 -190779
rect 8687 -190789 8767 -190761
rect 8687 -190841 8701 -190789
rect 8753 -190841 8767 -190789
rect 8687 -190869 8767 -190841
rect 8687 -190921 8701 -190869
rect 8753 -190921 8767 -190869
rect 8498 -191213 8578 -191057
rect 8687 -191349 8767 -190921
rect 8687 -191401 8701 -191349
rect 8753 -191401 8767 -191349
rect 8687 -191429 8767 -191401
rect 8687 -191481 8701 -191429
rect 8753 -191481 8767 -191429
rect 8390 -191571 8404 -191491
rect 8687 -191509 8767 -191481
rect 8687 -191561 8701 -191509
rect 8753 -191561 8767 -191509
rect 8687 -191585 8767 -191561
rect 10616 -191691 10636 -191682
rect 10616 -191702 10643 -191691
rect 10622 -191713 10643 -191702
rect 10617 -191796 10636 -191789
rect 10617 -191808 10641 -191796
rect 10620 -191818 10641 -191808
rect 10880 -198942 10901 -198920
rect 10879 -199068 10900 -199046
rect 10611 -200245 10632 -200223
rect 10611 -200351 10632 -200329
rect 2840 -201802 2864 -201750
rect 2916 -201802 2944 -201750
rect 2996 -201802 3024 -201750
rect 3076 -201802 3090 -201750
rect 2840 -201816 3090 -201802
rect 10843 -204633 10862 -204625
rect 10843 -204644 10866 -204633
rect 10845 -204655 10866 -204644
rect 10843 -204754 10863 -204746
rect 10843 -204765 10867 -204754
rect 10846 -204776 10867 -204765
rect 10841 -208307 10862 -208305
rect 10840 -208327 10862 -208307
rect 10840 -208427 10861 -208426
rect 10840 -208446 10863 -208427
rect 10840 -208448 10861 -208446
rect 1206 -233588 1286 -210286
rect 2840 -211270 3090 -211256
rect 2840 -211322 2864 -211270
rect 2916 -211322 2944 -211270
rect 2996 -211322 3024 -211270
rect 3076 -211322 3090 -211270
rect 2840 -232552 3090 -211322
rect 10611 -212743 10632 -212721
rect 10612 -212828 10633 -212827
rect 10612 -212847 10634 -212828
rect 10612 -212849 10633 -212847
rect 10879 -214027 10900 -214005
rect 10882 -214153 10903 -214131
rect 4461 -223076 4541 -220798
rect 10612 -221285 10636 -221263
rect 10615 -221390 10638 -221368
rect 8207 -221511 8287 -221487
rect 8207 -221563 8221 -221511
rect 8273 -221563 8287 -221511
rect 8207 -221591 8287 -221563
rect 8207 -221643 8221 -221591
rect 8273 -221643 8287 -221591
rect 8207 -221671 8287 -221643
rect 8207 -221723 8221 -221671
rect 8273 -221723 8287 -221671
rect 4577 -222017 4657 -221857
rect 8207 -222151 8287 -221723
rect 8207 -222203 8221 -222151
rect 8273 -222203 8287 -222151
rect 8207 -222231 8287 -222203
rect 8207 -222283 8221 -222231
rect 8273 -222283 8287 -222231
rect 8207 -222311 8287 -222283
rect 8207 -222363 8221 -222311
rect 8273 -222363 8287 -222311
rect 8207 -222387 8287 -222363
rect 8390 -221581 8404 -221501
rect 8687 -221511 8767 -221487
rect 8687 -221563 8701 -221511
rect 8753 -221563 8767 -221511
rect 8390 -222293 8470 -221581
rect 8687 -221591 8767 -221563
rect 8687 -221643 8701 -221591
rect 8753 -221643 8767 -221591
rect 8687 -221671 8767 -221643
rect 8687 -221723 8701 -221671
rect 8753 -221723 8767 -221671
rect 8498 -222015 8578 -221859
rect 8687 -222151 8767 -221723
rect 8687 -222203 8701 -222151
rect 8753 -222203 8767 -222151
rect 8687 -222231 8767 -222203
rect 8687 -222283 8701 -222231
rect 8753 -222283 8767 -222231
rect 8390 -222373 8404 -222293
rect 8687 -222311 8767 -222283
rect 8687 -222363 8701 -222311
rect 8753 -222363 8767 -222311
rect 8687 -222387 8767 -222363
rect 10617 -222506 10638 -222484
rect 10615 -222611 10636 -222589
rect 10882 -229743 10903 -229721
rect 10879 -229869 10900 -229847
rect 10612 -231047 10633 -231025
rect 10611 -231153 10632 -231131
rect 2840 -232604 2864 -232552
rect 2916 -232604 2944 -232552
rect 2996 -232604 3024 -232552
rect 3076 -232604 3090 -232552
rect 2840 -232618 3090 -232604
rect 10840 -235448 10861 -235426
rect 10841 -235569 10862 -235547
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_0
timestamp 1509269244
transform 1 0 922 0 -1 -221862
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_1
timestamp 1509269244
transform 1 0 922 0 -1 -191060
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_2
timestamp 1509269244
transform 1 0 922 0 1 -222012
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_3
timestamp 1509269244
transform 1 0 922 0 1 -191210
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_4
timestamp 1509269244
transform 1 0 922 0 -1 -160258
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_5
timestamp 1509269244
transform 1 0 922 0 1 -160408
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_6
timestamp 1509269244
transform 1 0 922 0 1 -129606
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_7
timestamp 1509269244
transform 1 0 922 0 -1 -129456
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_8
timestamp 1509269244
transform 1 0 922 0 -1 -98654
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_9
timestamp 1509269244
transform 1 0 922 0 1 -98804
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_10
timestamp 1509269244
transform 1 0 922 0 -1 -67852
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_11
timestamp 1509269244
transform 1 0 922 0 1 -68002
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_12
timestamp 1509269244
transform 1 0 922 0 -1 -6248
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_13
timestamp 1509269244
transform 1 0 922 0 1 -6398
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_14
timestamp 1509269244
transform 1 0 922 0 -1 -37050
box 0 -1 11647 15850
use EESPFAL_PRESENT_R1  EESPFAL_PRESENT_R1_15
timestamp 1509269244
transform 1 0 922 0 1 -37200
box 0 -1 11647 15850
<< labels >>
flabel metal1 s 945 7841 979 7875 2 FreeSans 2000 0 0 0 GND
port 1 nsew
rlabel locali s 927 4737 947 4756 4 k3_bar
port 2 nsew
rlabel locali s 937 4747 937 4747 4 k3_bar
port 2 nsew
rlabel locali s 928 4538 948 4557 4 x3_bar
port 3 nsew
rlabel locali s 938 4547 938 4547 4 x3_bar
port 3 nsew
rlabel locali s 929 8898 949 8917 4 x0
port 4 nsew
rlabel locali s 939 8908 939 8908 4 x0
port 4 nsew
rlabel locali s 930 8800 950 8819 4 x0_bar
port 5 nsew
rlabel locali s 940 8809 940 8809 4 x0_bar
port 5 nsew
rlabel locali s 931 8696 951 8715 4 k0
port 6 nsew
rlabel locali s 941 8706 941 8706 4 k0
port 6 nsew
rlabel locali s 928 8599 948 8618 4 k0_bar
port 7 nsew
rlabel locali s 938 8609 938 8609 4 k0_bar
port 7 nsew
rlabel locali s 933 6795 953 6815 4 x1
port 8 nsew
rlabel locali s 943 6805 943 6805 4 x1
port 8 nsew
rlabel locali s 928 7103 948 7122 4 k1_bar
port 9 nsew
rlabel locali s 938 7113 938 7113 4 k1_bar
port 9 nsew
rlabel locali s 927 7000 947 7019 4 k1
port 10 nsew
rlabel locali s 937 7010 937 7010 4 k1
port 10 nsew
rlabel locali s 932 6338 952 6357 4 k2
port 11 nsew
rlabel locali s 927 6239 947 6258 4 k2_bar
port 12 nsew
rlabel locali s 929 6538 949 6558 4 x2
port 13 nsew
rlabel locali s 928 6440 948 6459 4 x2_bar
port 14 nsew
rlabel locali s 938 6449 938 6449 4 x2_bar
port 14 nsew
rlabel locali s 939 6548 939 6548 4 x2
port 13 nsew
rlabel locali s 937 6249 937 6249 4 k2_bar
port 12 nsew
rlabel locali s 942 6348 942 6348 4 k2
port 11 nsew
rlabel locali s 928 4639 948 4658 4 k3
port 15 nsew
rlabel locali s 928 4438 948 4458 4 x3
port 16 nsew
rlabel locali s 938 4448 938 4448 4 x3
port 16 nsew
rlabel locali s 938 4649 938 4649 4 k3
port 15 nsew
rlabel locali s 950 -21362 970 -21343 4 k4
port 17 nsew
rlabel locali s 952 -19662 972 -19643 4 k5
port 18 nsew
rlabel locali s 948 -19006 968 -18987 4 k6
port 19 nsew
rlabel locali s 952 -17300 972 -17281 4 k7
port 20 nsew
rlabel locali s 949 -21266 969 -21247 4 k4_bar
port 21 nsew
rlabel locali s 943 -19763 963 -19744 4 k5_bar
port 22 nsew
rlabel locali s 932 -18903 952 -18884 4 k6_bar
port 23 nsew
rlabel locali s 954 -17404 974 -17385 4 k7_bar
port 24 nsew
rlabel locali s 953 -21564 973 -21544 4 x4
port 25 nsew
rlabel locali s 945 -19465 965 -19445 4 x5
port 26 nsew
rlabel locali s 929 -19207 949 -19187 4 x6
port 27 nsew
rlabel locali s 951 -17102 971 -17082 4 x7
port 28 nsew
rlabel locali s 949 -21464 969 -21445 4 x4_bar
port 29 nsew
rlabel locali s 948 -19564 968 -19545 4 x5_bar
port 30 nsew
rlabel locali s 952 -19104 972 -19085 4 x6_bar
port 31 nsew
rlabel locali s 954 -17203 974 -17184 4 x7_bar
port 32 nsew
rlabel locali s 964 -17194 964 -17194 4 x7_bar
port 32 nsew
rlabel locali s 962 -19095 962 -19095 4 x6_bar
port 31 nsew
rlabel locali s 958 -19555 958 -19555 4 x5_bar
port 30 nsew
rlabel locali s 959 -21455 959 -21455 4 x4_bar
port 29 nsew
rlabel locali s 961 -17092 961 -17092 4 x7
port 28 nsew
rlabel locali s 939 -19197 939 -19197 4 x6
port 27 nsew
rlabel locali s 955 -19455 955 -19455 4 x5
port 26 nsew
rlabel locali s 963 -21554 963 -21554 4 x4
port 25 nsew
rlabel locali s 964 -17394 964 -17394 4 k7_bar
port 24 nsew
rlabel locali s 942 -18893 942 -18893 4 k6_bar
port 23 nsew
rlabel locali s 953 -19753 953 -19753 4 k5_bar
port 22 nsew
rlabel locali s 959 -21256 959 -21256 4 k4_bar
port 21 nsew
rlabel locali s 962 -17290 962 -17290 4 k7
port 20 nsew
rlabel locali s 958 -18996 958 -18996 4 k6
port 19 nsew
rlabel locali s 962 -19652 962 -19652 4 k5
port 18 nsew
rlabel locali s 960 -21352 960 -21352 4 k4
port 17 nsew
rlabel locali s 947 -50007 967 -49987 4 x14
port 33 nsew
rlabel locali s 947 -48202 967 -48183 4 k15_bar
port 34 nsew
rlabel locali s 947 -49707 967 -49688 4 k14_bar
port 35 nsew
rlabel locali s 947 -50568 967 -50549 4 k13_bar
port 36 nsew
rlabel locali s 949 -52066 969 -52047 4 k12_bar
port 37 nsew
rlabel locali s 948 -50266 968 -50246 4 x13
port 38 nsew
rlabel locali s 950 -52364 970 -52344 4 x12
port 39 nsew
rlabel locali s 948 -52266 968 -52247 4 x12_bar
port 40 nsew
rlabel locali s 948 -50365 968 -50346 4 x13_bar
port 41 nsew
rlabel locali s 949 -47903 969 -47883 4 x15
port 42 nsew
rlabel locali s 953 -52164 973 -52145 4 k12
port 43 nsew
rlabel locali s 946 -48003 966 -47984 4 x15_bar
port 44 nsew
rlabel locali s 948 -49905 968 -49886 4 x14_bar
port 45 nsew
rlabel locali s 958 -49896 958 -49896 4 x14_bar
port 45 nsew
rlabel locali s 947 -48104 967 -48085 4 k15
port 46 nsew
rlabel locali s 958 -50356 958 -50356 4 x13_bar
port 41 nsew
rlabel locali s 959 -52056 959 -52056 4 k12_bar
port 37 nsew
rlabel locali s 957 -48094 957 -48094 4 k15
port 46 nsew
rlabel locali s 947 -49804 967 -49785 4 k14
port 47 nsew
rlabel locali s 947 -50465 967 -50446 4 k13
port 48 nsew
rlabel locali s 963 -52154 963 -52154 4 k12
port 43 nsew
rlabel locali s 957 -50455 957 -50455 4 k13
port 48 nsew
rlabel locali s 956 -47994 956 -47994 4 x15_bar
port 44 nsew
rlabel locali s 957 -49794 957 -49794 4 k14
port 47 nsew
rlabel locali s 959 -47893 959 -47893 4 x15
port 42 nsew
rlabel locali s 958 -52257 958 -52257 4 x12_bar
port 40 nsew
rlabel locali s 957 -50558 957 -50558 4 k13_bar
port 36 nsew
rlabel locali s 957 -49997 957 -49997 4 x14
port 33 nsew
rlabel locali s 957 -49697 957 -49697 4 k14_bar
port 35 nsew
rlabel locali s 960 -52354 960 -52354 4 x12
port 39 nsew
rlabel locali s 957 -48192 957 -48192 4 k15_bar
port 34 nsew
rlabel locali s 958 -50256 958 -50256 4 x13
port 38 nsew
rlabel locali s 950 -22004 970 -21985 4 x8_bar
port 49 nsew
rlabel locali s 960 -21995 960 -21995 4 x8_bar
port 49 nsew
rlabel locali s 950 -23899 970 -23880 4 x9_bar
port 50 nsew
rlabel locali s 953 -22101 973 -22082 4 k8
port 51 nsew
rlabel locali s 955 -24361 975 -24342 4 x10_bar
port 52 nsew
rlabel locali s 951 -23801 971 -23782 4 k9
port 53 nsew
rlabel locali s 956 -26263 976 -26244 4 x11_bar
port 54 nsew
rlabel locali s 948 -24462 968 -24443 4 k10
port 55 nsew
rlabel locali s 953 -26165 973 -26146 4 k11
port 56 nsew
rlabel locali s 951 -26365 971 -26345 4 x11
port 57 nsew
rlabel locali s 949 -24269 969 -24249 4 x10
port 58 nsew
rlabel locali s 948 -24003 968 -23983 4 x9
port 59 nsew
rlabel locali s 946 -21902 966 -21882 4 x8
port 60 nsew
rlabel locali s 950 -22200 970 -22181 4 k8_bar
port 61 nsew
rlabel locali s 956 -21892 956 -21892 4 x8
port 60 nsew
rlabel locali s 958 -23993 958 -23993 4 x9
port 59 nsew
rlabel locali s 959 -24259 959 -24259 4 x10
port 58 nsew
rlabel locali s 961 -26355 961 -26355 4 x11
port 57 nsew
rlabel locali s 949 -26063 969 -26044 4 k11_bar
port 62 nsew
rlabel locali s 951 -24565 971 -24546 4 k10_bar
port 63 nsew
rlabel locali s 949 -23704 969 -23685 4 k9_bar
port 64 nsew
rlabel locali s 960 -22190 960 -22190 4 k8_bar
port 61 nsew
rlabel locali s 959 -23694 959 -23694 4 k9_bar
port 64 nsew
rlabel locali s 961 -24555 961 -24555 4 k10_bar
port 63 nsew
rlabel locali s 959 -26053 959 -26053 4 k11_bar
port 62 nsew
rlabel locali s 963 -26155 963 -26155 4 k11
port 56 nsew
rlabel locali s 958 -24452 958 -24452 4 k10
port 55 nsew
rlabel locali s 961 -23791 961 -23791 4 k9
port 53 nsew
rlabel locali s 963 -22091 963 -22091 4 k8
port 51 nsew
rlabel locali s 966 -26254 966 -26254 4 x11_bar
port 54 nsew
rlabel locali s 965 -24352 965 -24352 4 x10_bar
port 52 nsew
rlabel locali s 960 -23890 960 -23890 4 x9_bar
port 50 nsew
rlabel locali s 949 -54806 969 -54786 4 x17
port 65 nsew
rlabel locali s 943 -52708 963 -52688 4 x16
port 66 nsew
rlabel locali s 950 -55362 970 -55343 4 k18_bar
port 67 nsew
rlabel locali s 945 -54506 965 -54487 4 k17_bar
port 68 nsew
rlabel locali s 944 -53007 964 -52988 4 k16_bar
port 69 nsew
rlabel locali s 950 -54604 970 -54585 4 k17
port 70 nsew
rlabel locali s 943 -52907 963 -52888 4 k16
port 71 nsew
rlabel locali s 949 -56968 969 -56949 4 k19
port 72 nsew
rlabel locali s 951 -55262 971 -55243 4 k18
port 73 nsew
rlabel locali s 948 -56866 968 -56847 4 k19_bar
port 74 nsew
rlabel locali s 961 -55252 961 -55252 4 k18
port 73 nsew
rlabel locali s 959 -56958 959 -56958 4 k19
port 72 nsew
rlabel locali s 947 -52807 967 -52788 4 x16_bar
port 75 nsew
rlabel locali s 948 -54702 968 -54683 4 x17_bar
port 76 nsew
rlabel locali s 954 -55162 974 -55143 4 x18_bar
port 77 nsew
rlabel locali s 946 -57064 966 -57045 4 x19_bar
port 78 nsew
rlabel locali s 953 -52897 953 -52897 4 k16
port 71 nsew
rlabel locali s 960 -54594 960 -54594 4 k17
port 70 nsew
rlabel locali s 956 -57055 956 -57055 4 x19_bar
port 78 nsew
rlabel locali s 954 -52997 954 -52997 4 k16_bar
port 69 nsew
rlabel locali s 964 -55153 964 -55153 4 x18_bar
port 77 nsew
rlabel locali s 955 -54496 955 -54496 4 k17_bar
port 68 nsew
rlabel locali s 958 -54693 958 -54693 4 x17_bar
port 76 nsew
rlabel locali s 960 -55352 960 -55352 4 k18_bar
port 67 nsew
rlabel locali s 957 -52798 957 -52798 4 x16_bar
port 75 nsew
rlabel locali s 953 -52698 953 -52698 4 x16
port 66 nsew
rlabel locali s 959 -54796 959 -54796 4 x17
port 65 nsew
rlabel locali s 952 -55066 972 -55046 4 x18
port 79 nsew
rlabel locali s 949 -57165 969 -57145 4 x19
port 80 nsew
rlabel locali s 958 -56856 958 -56856 4 k19_bar
port 74 nsew
rlabel locali s 959 -57155 959 -57155 4 x19
port 80 nsew
rlabel locali s 962 -55056 962 -55056 4 x18
port 79 nsew
rlabel locali s 948 -81166 968 -81147 4 x21_bar
port 81 nsew
rlabel locali s 947 -80706 967 -80687 4 x22_bar
port 82 nsew
rlabel locali s 957 -80697 957 -80697 4 x22_bar
port 82 nsew
rlabel locali s 950 -78807 970 -78788 4 x23_bar
port 83 nsew
rlabel locali s 958 -81157 958 -81157 4 x21_bar
port 81 nsew
rlabel locali s 952 -82867 972 -82848 4 k20_bar
port 84 nsew
rlabel locali s 953 -83068 973 -83048 4 x20_bar
port 85 nsew
rlabel locali s 948 -81369 968 -81350 4 k21_bar
port 86 nsew
rlabel locali s 945 -80509 965 -80490 4 k22_bar
port 87 nsew
rlabel locali s 945 -79009 965 -78990 4 k23_bar
port 88 nsew
rlabel locali s 949 -80606 969 -80587 4 k22
port 89 nsew
rlabel locali s 951 -81266 971 -81247 4 k21
port 90 nsew
rlabel locali s 950 -82965 970 -82946 4 k20
port 91 nsew
rlabel locali s 961 -81256 961 -81256 4 k21
port 90 nsew
rlabel locali s 959 -80596 959 -80596 4 k22
port 89 nsew
rlabel locali s 943 -78909 963 -78890 4 k23
port 92 nsew
rlabel locali s 960 -82955 960 -82955 4 k20
port 91 nsew
rlabel locali s 951 -83168 971 -83149 4 x20
port 93 nsew
rlabel locali s 949 -81067 969 -81047 4 x21
port 94 nsew
rlabel locali s 961 -83158 961 -83158 4 x20
port 93 nsew
rlabel locali s 959 -81057 959 -81057 4 x21
port 94 nsew
rlabel locali s 954 -80810 974 -80790 4 x22
port 95 nsew
rlabel locali s 950 -78707 970 -78687 4 x23
port 96 nsew
rlabel locali s 955 -78999 955 -78999 4 k23_bar
port 88 nsew
rlabel locali s 955 -80499 955 -80499 4 k22_bar
port 87 nsew
rlabel locali s 958 -81359 958 -81359 4 k21_bar
port 86 nsew
rlabel locali s 962 -82857 962 -82857 4 k20_bar
port 84 nsew
rlabel locali s 953 -78899 953 -78899 4 k23
port 92 nsew
rlabel locali s 960 -78697 960 -78697 4 x23
port 96 nsew
rlabel locali s 964 -80800 964 -80800 4 x22
port 95 nsew
rlabel locali s 960 -78798 960 -78798 4 x23_bar
port 83 nsew
rlabel locali s 963 -83058 963 -83058 4 x20_bar
port 85 nsew
rlabel locali s 946 -85606 966 -85587 4 x25
port 97 nsew
rlabel locali s 945 -83609 965 -83589 4 x24_bar
port 98 nsew
rlabel locali s 949 -83510 969 -83491 4 x24
port 99 nsew
rlabel locali s 948 -83809 968 -83790 4 k24_bar
port 100 nsew
rlabel locali s 949 -85303 969 -85284 4 k25_bar
port 101 nsew
rlabel locali s 955 -83599 955 -83599 4 x24_bar
port 98 nsew
rlabel locali s 946 -86164 966 -86145 4 k26_bar
port 102 nsew
rlabel locali s 946 -85508 966 -85488 4 x25_bar
port 103 nsew
rlabel locali s 943 -85967 963 -85947 4 x26_bar
port 104 nsew
rlabel locali s 946 -85407 966 -85388 4 k25
port 105 nsew
rlabel locali s 947 -83703 967 -83684 4 k24
port 106 nsew
rlabel locali s 957 -83694 957 -83694 4 k24
port 106 nsew
rlabel locali s 956 -85397 956 -85397 4 k25
port 105 nsew
rlabel locali s 946 -86066 966 -86047 4 k26
port 107 nsew
rlabel locali s 956 -86154 956 -86154 4 k26_bar
port 102 nsew
rlabel locali s 959 -83500 959 -83500 4 x24
port 99 nsew
rlabel locali s 959 -85293 959 -85293 4 k25_bar
port 101 nsew
rlabel locali s 956 -85596 956 -85596 4 x25
port 97 nsew
rlabel locali s 958 -83800 958 -83800 4 k24_bar
port 100 nsew
rlabel locali s 946 -85865 966 -85846 4 x26
port 108 nsew
rlabel locali s 956 -86056 956 -86056 4 k26
port 107 nsew
rlabel locali s 953 -85957 953 -85957 4 x26_bar
port 104 nsew
rlabel locali s 956 -85498 956 -85498 4 x25_bar
port 103 nsew
rlabel locali s 956 -85855 956 -85855 4 x26
port 108 nsew
rlabel locali s 948 -87968 968 -87949 4 x27
port 109 nsew
rlabel locali s 949 -87867 969 -87847 4 x27_bar
port 110 nsew
rlabel locali s 958 -87958 958 -87958 4 x27
port 109 nsew
rlabel locali s 959 -87857 959 -87857 4 x27_bar
port 110 nsew
rlabel locali s 948 -87770 968 -87751 4 k27
port 111 nsew
rlabel locali s 952 -87667 972 -87648 4 k27_bar
port 112 nsew
rlabel locali s 958 -87760 958 -87760 4 k27
port 111 nsew
rlabel locali s 962 -87657 962 -87657 4 k27_bar
port 112 nsew
rlabel locali s 949 -111410 969 -111391 4 k30
port 113 nsew
rlabel locali s 955 -111312 975 -111293 4 k30_bar
port 114 nsew
rlabel locali s 955 -111968 975 -111949 4 x29_bar
port 115 nsew
rlabel locali s 945 -112171 965 -112152 4 k29_bar
port 116 nsew
rlabel locali s 949 -113969 969 -113950 4 x28
port 117 nsew
rlabel locali s 954 -113670 974 -113651 4 k28_bar
port 118 nsew
rlabel locali s 954 -113868 974 -113848 4 x28_bar
port 119 nsew
rlabel locali s 956 -111870 976 -111850 4 x29
port 120 nsew
rlabel locali s 947 -109710 967 -109691 4 k31
port 121 nsew
rlabel locali s 964 -113660 964 -113660 4 k28_bar
port 118 nsew
rlabel locali s 959 -111401 959 -111401 4 k30
port 113 nsew
rlabel locali s 955 -112161 955 -112161 4 k29_bar
port 116 nsew
rlabel locali s 964 -113858 964 -113858 4 x28_bar
port 119 nsew
rlabel locali s 965 -111302 965 -111302 4 k30_bar
port 114 nsew
rlabel locali s 965 -111959 965 -111959 4 x29_bar
port 115 nsew
rlabel locali s 947 -109804 967 -109785 4 k31_bar
port 122 nsew
rlabel locali s 951 -111507 971 -111487 4 x30_bar
port 123 nsew
rlabel locali s 957 -109701 957 -109701 4 k31
port 121 nsew
rlabel locali s 959 -113959 959 -113959 4 x28
port 117 nsew
rlabel locali s 947 -109610 967 -109590 4 x31_bar
port 124 nsew
rlabel locali s 966 -111860 966 -111860 4 x29
port 120 nsew
rlabel locali s 948 -112070 968 -112051 4 k29
port 125 nsew
rlabel locali s 950 -111607 970 -111588 4 x30
port 126 nsew
rlabel locali s 958 -112061 958 -112061 4 k29
port 125 nsew
rlabel locali s 955 -113772 975 -113753 4 k28
port 127 nsew
rlabel locali s 965 -113762 965 -113762 4 k28
port 127 nsew
rlabel locali s 957 -109600 957 -109600 4 x31_bar
port 124 nsew
rlabel locali s 950 -109508 970 -109489 4 x31
port 128 nsew
rlabel locali s 960 -109498 960 -109498 4 x31
port 128 nsew
rlabel locali s 960 -111597 960 -111597 4 x30
port 126 nsew
rlabel locali s 961 -111497 961 -111497 4 x30_bar
port 123 nsew
rlabel locali s 957 -109794 957 -109794 4 k31_bar
port 122 nsew
rlabel locali s 926 6897 946 6916 4 x1_bar
port 129 nsew
rlabel locali s 936 6906 936 6906 4 x1_bar
port 129 nsew
rlabel locali s 953 -116867 973 -116848 4 k34
port 130 nsew
rlabel locali s 948 -118567 968 -118548 4 k35
port 131 nsew
rlabel locali s 951 -114308 971 -114288 4 x32
port 132 nsew
rlabel locali s 951 -116410 971 -116390 4 x33
port 133 nsew
rlabel locali s 946 -116670 966 -116650 4 x34
port 134 nsew
rlabel locali s 951 -118769 971 -118750 4 x35
port 135 nsew
rlabel locali s 946 -118668 966 -118648 4 x35_bar
port 136 nsew
rlabel locali s 949 -116765 969 -116746 4 x34_bar
port 137 nsew
rlabel locali s 944 -116309 964 -116290 4 x33_bar
port 138 nsew
rlabel locali s 947 -114409 967 -114390 4 x32_bar
port 139 nsew
rlabel locali s 948 -116210 968 -116191 4 k33
port 140 nsew
rlabel locali s 949 -114510 969 -114491 4 k32
port 141 nsew
rlabel locali s 959 -114501 959 -114501 4 k32
port 141 nsew
rlabel locali s 950 -114608 970 -114589 4 k32_bar
port 142 nsew
rlabel locali s 950 -118472 970 -118453 4 k35_bar
port 143 nsew
rlabel locali s 952 -116107 972 -116088 4 k33_bar
port 144 nsew
rlabel locali s 951 -116969 971 -116950 4 k34_bar
port 145 nsew
rlabel locali s 960 -118462 960 -118462 4 k35_bar
port 143 nsew
rlabel locali s 961 -118759 961 -118759 4 x35
port 135 nsew
rlabel locali s 956 -116660 956 -116660 4 x34
port 134 nsew
rlabel locali s 961 -116400 961 -116400 4 x33
port 133 nsew
rlabel locali s 961 -114298 961 -114298 4 x32
port 132 nsew
rlabel locali s 961 -116959 961 -116959 4 k34_bar
port 145 nsew
rlabel locali s 957 -114400 957 -114400 4 x32_bar
port 139 nsew
rlabel locali s 954 -116300 954 -116300 4 x33_bar
port 138 nsew
rlabel locali s 962 -116097 962 -116097 4 k33_bar
port 144 nsew
rlabel locali s 959 -116756 959 -116756 4 x34_bar
port 137 nsew
rlabel locali s 956 -118658 956 -118658 4 x35_bar
port 136 nsew
rlabel locali s 960 -114598 960 -114598 4 k32_bar
port 142 nsew
rlabel locali s 958 -116201 958 -116201 4 k33
port 140 nsew
rlabel locali s 958 -118558 958 -118558 4 k35
port 131 nsew
rlabel locali s 963 -116858 963 -116858 4 k34
port 130 nsew
rlabel locali s 943 -142412 963 -142393 4 x38
port 146 nsew
rlabel locali s 953 -142402 953 -142402 4 x38
port 146 nsew
rlabel locali s 957 -142113 977 -142094 4 k38_bar
port 147 nsew
rlabel locali s 945 -140608 965 -140589 4 k39_bar
port 148 nsew
rlabel locali s 953 -140310 973 -140291 4 x39
port 149 nsew
rlabel locali s 946 -142215 966 -142196 4 k38
port 150 nsew
rlabel locali s 950 -142673 970 -142654 4 x37
port 151 nsew
rlabel locali s 949 -144773 969 -144754 4 x36
port 152 nsew
rlabel locali s 949 -140508 969 -140489 4 k39
port 153 nsew
rlabel locali s 959 -144763 959 -144763 4 x36
port 152 nsew
rlabel locali s 960 -142663 960 -142663 4 x37
port 151 nsew
rlabel locali s 949 -144572 969 -144553 4 k36
port 154 nsew
rlabel locali s 955 -140599 955 -140599 4 k39_bar
port 148 nsew
rlabel locali s 967 -142104 967 -142104 4 k38_bar
port 147 nsew
rlabel locali s 963 -140300 963 -140300 4 x39
port 149 nsew
rlabel locali s 948 -142972 968 -142953 4 k37_bar
port 155 nsew
rlabel locali s 947 -144473 967 -144454 4 k36_bar
port 156 nsew
rlabel locali s 944 -140411 964 -140391 4 x39_bar
port 157 nsew
rlabel locali s 945 -142310 965 -142290 4 x38_bar
port 158 nsew
rlabel locali s 949 -144675 969 -144655 4 x36_bar
port 159 nsew
rlabel locali s 950 -142773 970 -142753 4 x37_bar
port 160 nsew
rlabel locali s 955 -142300 955 -142300 4 x38_bar
port 158 nsew
rlabel locali s 954 -140401 954 -140401 4 x39_bar
port 157 nsew
rlabel locali s 959 -140499 959 -140499 4 k39
port 153 nsew
rlabel locali s 956 -142206 956 -142206 4 k38
port 150 nsew
rlabel locali s 951 -142874 971 -142855 4 k37
port 161 nsew
rlabel locali s 959 -144563 959 -144563 4 k36
port 154 nsew
rlabel locali s 960 -142763 960 -142763 4 x37_bar
port 160 nsew
rlabel locali s 959 -144665 959 -144665 4 x36_bar
port 159 nsew
rlabel locali s 961 -142865 961 -142865 4 k37
port 161 nsew
rlabel locali s 957 -144463 957 -144463 4 k36_bar
port 156 nsew
rlabel locali s 958 -142963 958 -142963 4 k37_bar
port 155 nsew
rlabel locali s 948 -147110 968 -147090 4 x41_bar
port 162 nsew
rlabel locali s 951 -145210 971 -145190 4 x40_bar
port 163 nsew
rlabel locali s 947 -149571 967 -149551 4 x43
port 164 nsew
rlabel locali s 947 -147474 967 -147455 4 x42
port 165 nsew
rlabel locali s 950 -147213 970 -147194 4 x41
port 166 nsew
rlabel locali s 945 -145411 965 -145392 4 k40_bar
port 167 nsew
rlabel locali s 950 -145112 970 -145093 4 x40
port 168 nsew
rlabel locali s 949 -146910 969 -146891 4 k41_bar
port 169 nsew
rlabel locali s 946 -147770 966 -147751 4 k42_bar
port 170 nsew
rlabel locali s 945 -145311 965 -145292 4 k40
port 171 nsew
rlabel locali s 948 -149271 968 -149252 4 k43_bar
port 172 nsew
rlabel locali s 954 -147006 974 -146987 4 k41
port 173 nsew
rlabel locali s 943 -147672 963 -147653 4 k42
port 174 nsew
rlabel locali s 949 -149370 969 -149351 4 k43
port 175 nsew
rlabel locali s 958 -149262 958 -149262 4 k43_bar
port 172 nsew
rlabel locali s 956 -147761 956 -147761 4 k42_bar
port 170 nsew
rlabel locali s 959 -146901 959 -146901 4 k41_bar
port 169 nsew
rlabel locali s 955 -145402 955 -145402 4 k40_bar
port 167 nsew
rlabel locali s 961 -145200 961 -145200 4 x40_bar
port 163 nsew
rlabel locali s 958 -147100 958 -147100 4 x41_bar
port 162 nsew
rlabel locali s 946 -147571 966 -147551 4 x42_bar
port 176 nsew
rlabel locali s 946 -149474 966 -149455 4 x43_bar
port 177 nsew
rlabel locali s 959 -149361 959 -149361 4 k43
port 175 nsew
rlabel locali s 953 -147663 953 -147663 4 k42
port 174 nsew
rlabel locali s 964 -146997 964 -146997 4 k41
port 173 nsew
rlabel locali s 955 -145302 955 -145302 4 k40
port 171 nsew
rlabel locali s 956 -149465 956 -149465 4 x43_bar
port 177 nsew
rlabel locali s 960 -145102 960 -145102 4 x40
port 168 nsew
rlabel locali s 960 -147203 960 -147203 4 x41
port 166 nsew
rlabel locali s 956 -147561 956 -147561 4 x42_bar
port 176 nsew
rlabel locali s 957 -147464 957 -147464 4 x42
port 165 nsew
rlabel locali s 957 -149561 957 -149561 4 x43
port 164 nsew
rlabel locali s 944 -171413 964 -171394 4 k47_bar
port 178 nsew
rlabel locali s 946 -172913 966 -172894 4 k46_bar
port 179 nsew
rlabel locali s 946 -173773 966 -173754 4 k45_bar
port 180 nsew
rlabel locali s 949 -175272 969 -175253 4 k44_bar
port 181 nsew
rlabel locali s 947 -175576 967 -175556 4 x44
port 182 nsew
rlabel locali s 948 -171113 968 -171093 4 x47
port 183 nsew
rlabel locali s 948 -171213 968 -171194 4 x47_bar
port 184 nsew
rlabel locali s 948 -171314 968 -171295 4 k47
port 185 nsew
rlabel locali s 949 -173213 969 -173193 4 x46
port 186 nsew
rlabel locali s 948 -173013 968 -172994 4 k46
port 187 nsew
rlabel locali s 958 -173004 958 -173004 4 k46
port 187 nsew
rlabel locali s 959 -173203 959 -173203 4 x46
port 186 nsew
rlabel locali s 957 -175566 957 -175566 4 x44
port 182 nsew
rlabel locali s 946 -173676 966 -173657 4 k45
port 188 nsew
rlabel locali s 958 -171103 958 -171103 4 x47
port 183 nsew
rlabel locali s 959 -175263 959 -175263 4 k44_bar
port 181 nsew
rlabel locali s 953 -175371 973 -175352 4 k44
port 189 nsew
rlabel locali s 948 -175474 968 -175455 4 x44_bar
port 190 nsew
rlabel locali s 949 -173574 969 -173555 4 x45_bar
port 191 nsew
rlabel locali s 947 -173115 967 -173096 4 x46_bar
port 192 nsew
rlabel locali s 957 -173106 957 -173106 4 x46_bar
port 192 nsew
rlabel locali s 958 -171204 958 -171204 4 x47_bar
port 184 nsew
rlabel locali s 956 -173764 956 -173764 4 k45_bar
port 180 nsew
rlabel locali s 945 -173474 965 -173454 4 x45
port 193 nsew
rlabel locali s 956 -172904 956 -172904 4 k46_bar
port 179 nsew
rlabel locali s 958 -171305 958 -171305 4 k47
port 185 nsew
rlabel locali s 955 -173464 955 -173464 4 x45
port 193 nsew
rlabel locali s 954 -171404 954 -171404 4 k47_bar
port 178 nsew
rlabel locali s 959 -173565 959 -173565 4 x45_bar
port 191 nsew
rlabel locali s 963 -175362 963 -175362 4 k44
port 189 nsew
rlabel locali s 956 -173667 956 -173667 4 k45
port 188 nsew
rlabel locali s 958 -175465 958 -175465 4 x44_bar
port 190 nsew
rlabel locali s 950 -180276 970 -180256 4 x51_bar
port 194 nsew
rlabel locali s 946 -178372 966 -178353 4 x50_bar
port 195 nsew
rlabel locali s 944 -180073 964 -180054 4 k51_bar
port 196 nsew
rlabel locali s 949 -177814 969 -177795 4 k49
port 197 nsew
rlabel locali s 950 -176112 970 -176093 4 k48
port 198 nsew
rlabel locali s 959 -177805 959 -177805 4 k49
port 197 nsew
rlabel locali s 944 -178274 964 -178254 4 x50
port 199 nsew
rlabel locali s 943 -176210 963 -176191 4 k48_bar
port 200 nsew
rlabel locali s 951 -178013 971 -177993 4 x49
port 201 nsew
rlabel locali s 947 -176014 967 -175994 4 x48_bar
port 202 nsew
rlabel locali s 951 -175911 971 -175892 4 x48
port 203 nsew
rlabel locali s 961 -175901 961 -175901 4 x48
port 203 nsew
rlabel locali s 945 -177912 965 -177893 4 x49_bar
port 204 nsew
rlabel locali s 943 -178570 963 -178551 4 k50_bar
port 205 nsew
rlabel locali s 947 -180374 967 -180355 4 x51
port 206 nsew
rlabel locali s 957 -180365 957 -180365 4 x51
port 206 nsew
rlabel locali s 955 -177903 955 -177903 4 x49_bar
port 204 nsew
rlabel locali s 956 -178363 956 -178363 4 x50_bar
port 195 nsew
rlabel locali s 948 -178477 968 -178458 4 k50
port 207 nsew
rlabel locali s 960 -180266 960 -180266 4 x51_bar
port 194 nsew
rlabel locali s 951 -177713 971 -177694 4 k49_bar
port 208 nsew
rlabel locali s 950 -180170 970 -180151 4 k51
port 209 nsew
rlabel locali s 954 -180064 954 -180064 4 k51_bar
port 196 nsew
rlabel locali s 961 -177704 961 -177704 4 k49_bar
port 208 nsew
rlabel locali s 954 -178264 954 -178264 4 x50
port 199 nsew
rlabel locali s 953 -178561 953 -178561 4 k50_bar
port 205 nsew
rlabel locali s 960 -180161 960 -180161 4 k51
port 209 nsew
rlabel locali s 957 -176004 957 -176004 4 x48_bar
port 202 nsew
rlabel locali s 960 -176103 960 -176103 4 k48
port 198 nsew
rlabel locali s 961 -178003 961 -178003 4 x49
port 201 nsew
rlabel locali s 953 -176201 953 -176201 4 k48_bar
port 200 nsew
rlabel locali s 958 -178468 958 -178468 4 k50
port 207 nsew
rlabel locali s 947 -204015 967 -203995 4 x54
port 210 nsew
rlabel locali s 948 -202215 968 -202196 4 k55_bar
port 211 nsew
rlabel locali s 945 -201915 965 -201895 4 x55
port 212 nsew
rlabel locali s 947 -202115 967 -202096 4 k55
port 213 nsew
rlabel locali s 958 -202206 958 -202206 4 k55_bar
port 211 nsew
rlabel locali s 957 -202106 957 -202106 4 k55
port 213 nsew
rlabel locali s 946 -203916 966 -203897 4 x54_bar
port 214 nsew
rlabel locali s 949 -202015 969 -201996 4 x55_bar
port 215 nsew
rlabel locali s 947 -203716 967 -203697 4 k54_bar
port 216 nsew
rlabel locali s 956 -203907 956 -203907 4 x54_bar
port 214 nsew
rlabel locali s 959 -202006 959 -202006 4 x55_bar
port 215 nsew
rlabel locali s 955 -201905 955 -201905 4 x55
port 212 nsew
rlabel locali s 957 -203707 957 -203707 4 k54_bar
port 216 nsew
rlabel locali s 957 -204005 957 -204005 4 x54
port 210 nsew
rlabel locali s 947 -206376 967 -206357 4 x52
port 217 nsew
rlabel locali s 947 -204475 967 -204456 4 k53
port 218 nsew
rlabel locali s 947 -206178 967 -206159 4 k52
port 219 nsew
rlabel locali s 948 -204375 968 -204356 4 x53_bar
port 220 nsew
rlabel locali s 950 -204274 970 -204254 4 x53
port 221 nsew
rlabel locali s 957 -204466 957 -204466 4 k53
port 218 nsew
rlabel locali s 957 -206367 957 -206367 4 x52
port 217 nsew
rlabel locali s 952 -204576 972 -204557 4 k53_bar
port 222 nsew
rlabel locali s 962 -204567 962 -204567 4 k53_bar
port 222 nsew
rlabel locali s 949 -206074 969 -206055 4 k52_bar
port 223 nsew
rlabel locali s 960 -204264 960 -204264 4 x53
port 221 nsew
rlabel locali s 948 -203815 968 -203796 4 k54
port 224 nsew
rlabel locali s 959 -206064 959 -206064 4 k52_bar
port 223 nsew
rlabel locali s 957 -206168 957 -206168 4 k52
port 219 nsew
rlabel locali s 949 -206276 969 -206256 4 x52_bar
port 225 nsew
rlabel locali s 959 -206266 959 -206266 4 x52_bar
port 225 nsew
rlabel locali s 958 -203806 958 -203806 4 k54
port 224 nsew
rlabel locali s 958 -204366 958 -204366 4 x53_bar
port 220 nsew
rlabel locali s 948 -236979 968 -236960 4 k60
port 226 nsew
rlabel locali s 947 -234617 967 -234598 4 k62
port 227 nsew
rlabel locali s 949 -232917 969 -232898 4 k63
port 228 nsew
rlabel locali s 948 -234519 968 -234500 4 k62_bar
port 229 nsew
rlabel locali s 945 -236876 965 -236857 4 k60_bar
port 230 nsew
rlabel locali s 955 -236867 955 -236867 4 k60_bar
port 230 nsew
rlabel locali s 948 -235379 968 -235360 4 k61_bar
port 231 nsew
rlabel locali s 950 -232718 970 -232699 4 x63
port 232 nsew
rlabel locali s 957 -234608 957 -234608 4 k62
port 227 nsew
rlabel locali s 948 -233016 968 -232997 4 k63_bar
port 233 nsew
rlabel locali s 949 -237179 969 -237159 4 x60
port 234 nsew
rlabel locali s 959 -232908 959 -232908 4 k63
port 228 nsew
rlabel locali s 949 -235076 969 -235056 4 x61
port 235 nsew
rlabel locali s 950 -237079 970 -237060 4 x60_bar
port 236 nsew
rlabel locali s 960 -232708 960 -232708 4 x63
port 232 nsew
rlabel locali s 960 -237070 960 -237070 4 x60_bar
port 236 nsew
rlabel locali s 948 -232817 968 -232797 4 x63_bar
port 237 nsew
rlabel locali s 958 -233007 958 -233007 4 k63_bar
port 233 nsew
rlabel locali s 958 -235370 958 -235370 4 k61_bar
port 231 nsew
rlabel locali s 948 -235179 968 -235160 4 x61_bar
port 238 nsew
rlabel locali s 947 -235278 967 -235259 4 k61
port 239 nsew
rlabel locali s 948 -234818 968 -234798 4 x62
port 240 nsew
rlabel locali s 957 -235269 957 -235269 4 k61
port 239 nsew
rlabel locali s 948 -234718 968 -234699 4 x62_bar
port 241 nsew
rlabel locali s 958 -234510 958 -234510 4 k62_bar
port 229 nsew
rlabel locali s 959 -235066 959 -235066 4 x61
port 235 nsew
rlabel locali s 958 -236970 958 -236970 4 k60
port 226 nsew
rlabel locali s 958 -234808 958 -234808 4 x62
port 240 nsew
rlabel locali s 958 -232807 958 -232807 4 x63_bar
port 237 nsew
rlabel locali s 959 -237169 959 -237169 4 x60
port 234 nsew
rlabel locali s 958 -234709 958 -234709 4 x62_bar
port 241 nsew
rlabel locali s 958 -235170 958 -235170 4 x61_bar
port 238 nsew
rlabel locali s 947 -209273 967 -209254 4 k58
port 242 nsew
rlabel locali s 950 -206815 970 -206796 4 x56_bar
port 243 nsew
rlabel locali s 948 -211174 968 -211155 4 x59
port 244 nsew
rlabel locali s 950 -208614 970 -208595 4 k57
port 245 nsew
rlabel locali s 957 -209264 957 -209264 4 k58
port 242 nsew
rlabel locali s 948 -210875 968 -210856 4 k59_bar
port 246 nsew
rlabel locali s 946 -207015 966 -206996 4 k56_bar
port 247 nsew
rlabel locali s 946 -209373 966 -209354 4 k58_bar
port 248 nsew
rlabel locali s 958 -210865 958 -210865 4 k59_bar
port 246 nsew
rlabel locali s 946 -209173 966 -209154 4 x58_bar
port 249 nsew
rlabel locali s 960 -208605 960 -208605 4 k57
port 245 nsew
rlabel locali s 955 -206715 975 -206695 4 x56
port 250 nsew
rlabel locali s 948 -209074 968 -209054 4 x58
port 251 nsew
rlabel locali s 952 -206914 972 -206895 4 k56
port 252 nsew
rlabel locali s 949 -211076 969 -211056 4 x59_bar
port 253 nsew
rlabel locali s 965 -206705 965 -206705 4 x56
port 250 nsew
rlabel locali s 960 -206806 960 -206806 4 x56_bar
port 243 nsew
rlabel locali s 951 -208714 971 -208695 4 x57_bar
port 254 nsew
rlabel locali s 961 -208705 961 -208705 4 x57_bar
port 254 nsew
rlabel locali s 948 -208814 968 -208794 4 x57
port 255 nsew
rlabel locali s 954 -210973 974 -210954 4 k59
port 256 nsew
rlabel locali s 958 -208804 958 -208804 4 x57
port 255 nsew
rlabel locali s 956 -209164 956 -209164 4 x58_bar
port 249 nsew
rlabel locali s 964 -210963 964 -210963 4 k59
port 256 nsew
rlabel locali s 945 -208513 965 -208494 4 k57_bar
port 257 nsew
rlabel locali s 955 -208504 955 -208504 4 k57_bar
port 257 nsew
rlabel locali s 958 -211164 958 -211164 4 x59
port 244 nsew
rlabel locali s 956 -207006 956 -207006 4 k56_bar
port 247 nsew
rlabel locali s 956 -209364 956 -209364 4 k58_bar
port 248 nsew
rlabel locali s 962 -206905 962 -206905 4 k56
port 252 nsew
rlabel locali s 959 -211066 959 -211066 4 x59_bar
port 253 nsew
rlabel locali s 958 -209064 958 -209064 4 x58
port 251 nsew
flabel metal2 s 1231 9022 1261 9054 2 FreeSans 2000 0 0 0 Dis0
port 258 nsew
flabel metal2 s 4444 9020 4485 9062 2 FreeSans 2000 0 0 0 CLK1
port 259 nsew
flabel metal2 s 4566 9027 4586 9048 2 FreeSans 2000 0 0 0 Dis1
port 260 nsew
flabel metal2 s 8892 9025 8917 9053 2 FreeSans 2000 0 0 0 CLK3
port 261 nsew
flabel metal2 s 9172 9021 9203 9055 2 FreeSans 2000 0 0 0 Dis2
port 262 nsew
flabel metal2 s 9255 9021 9296 9064 2 FreeSans 2000 0 0 0 CLK2
port 263 nsew
flabel metal2 s 9355 9028 9383 9058 2 FreeSans 2000 0 0 0 Dis3
port 264 nsew
rlabel metal2 s 10842 -50758 10863 -50736 4 s12
port 265 nsew
rlabel metal2 s 10612 -46234 10633 -46212 4 s13
port 266 nsew
rlabel metal2 s 10878 -45058 10899 -45036 4 s14
port 267 nsew
rlabel metal2 s 10843 -50635 10864 -50613 4 s12_bar
port 268 nsew
rlabel metal2 s 10611 -46340 10632 -46318 4 s13_bar
port 269 nsew
rlabel metal2 s 10879 -44933 10900 -44911 4 s14_bar
port 270 nsew
rlabel metal2 s 10840 -54315 10861 -54293 4 s16
port 271 nsew
rlabel metal2 s 10613 -58839 10634 -58817 4 s17
port 272 nsew
rlabel metal2 s 10879 -60014 10900 -59992 4 s18
port 273 nsew
rlabel metal2 s 10615 -67379 10636 -67357 4 s19
port 274 nsew
rlabel metal2 s 10839 -54440 10860 -54418 4 s16_bar
port 275 nsew
rlabel metal2 s 10610 -58733 10631 -58711 4 s17_bar
port 276 nsew
rlabel metal2 s 10883 -60143 10904 -60121 4 s18_bar
port 277 nsew
rlabel metal2 s 10612 -67274 10633 -67252 4 s19_bar
port 278 nsew
rlabel metal2 s 10875 -75858 10896 -75836 4 s22
port 279 nsew
rlabel metal2 s 10614 -68497 10635 -68475 4 s23
port 280 nsew
rlabel metal2 s 10840 -81559 10861 -81537 4 s20
port 281 nsew
rlabel metal2 s 10611 -77036 10631 -77017 4 s21
port 282 nsew
rlabel metal2 s 10843 -81438 10864 -81416 4 s20_bar
port 283 nsew
rlabel metal2 s 10611 -77141 10630 -77122 4 s21_bar
port 284 nsew
rlabel metal2 s 10882 -75732 10903 -75710 4 s22_bar
port 285 nsew
rlabel metal2 s 10615 -68600 10636 -68578 4 s23_bar
port 286 nsew
rlabel metal2 s 10842 -85118 10863 -85096 4 s24
port 287 nsew
rlabel metal2 s 10611 -89640 10631 -89621 4 s25
port 288 nsew
rlabel metal2 s 10880 -90818 10901 -90796 4 s26
port 289 nsew
rlabel metal2 s 10618 -98181 10639 -98159 4 s27
port 290 nsew
rlabel metal2 s 10841 -85239 10862 -85217 4 s24_bar
port 291 nsew
rlabel metal2 s 10883 -90944 10904 -90922 4 s26_bar
port 292 nsew
rlabel metal2 s 10614 -98074 10633 -98054 4 s27_bar
port 293 nsew
rlabel metal2 s 10842 -112360 10863 -112338 4 s28
port 294 nsew
rlabel metal2 s 10609 -107838 10629 -107819 4 s29
port 295 nsew
rlabel metal2 s 10879 -106661 10900 -106639 4 s30
port 296 nsew
rlabel metal2 s 10615 -99299 10636 -99277 4 s31
port 297 nsew
rlabel metal2 s 10841 -112239 10862 -112217 4 s28_bar
port 298 nsew
rlabel metal2 s 10609 -107946 10630 -107924 4 s29_bar
port 299 nsew
rlabel metal2 s 10880 -106534 10901 -106512 4 s30_bar
port 300 nsew
rlabel metal2 s 10614 -99402 10635 -99380 4 s31_bar
port 301 nsew
rlabel metal2 s 10877 7287 10898 7309 4 s0
port 302 nsew
rlabel metal2 s 10652 2766 10673 2788 4 s1
port 303 nsew
rlabel metal2 s 10913 1586 10934 1608 4 s2
port 304 nsew
rlabel metal2 s 10653 -5776 10674 -5754 4 s3
port 305 nsew
rlabel metal2 s 10838 -19954 10859 -19932 4 s4
port 306 nsew
rlabel metal2 s 10878 -14256 10899 -14234 4 s6
port 307 nsew
rlabel metal2 s 10656 -6892 10676 -6873 4 s7
port 308 nsew
rlabel metal2 s 10838 -23515 10859 -23493 4 s8
port 309 nsew
rlabel metal2 s 10613 -28036 10634 -28014 4 s9
port 310 nsew
rlabel metal2 s 10877 -29215 10898 -29193 4 s10
port 311 nsew
rlabel metal2 s 10876 7167 10897 7189 4 s0_bar
port 312 nsew
rlabel metal2 s 10653 2870 10674 2892 4 s1_bar
port 313 nsew
rlabel metal2 s 10919 1459 10940 1481 4 s2_bar
port 314 nsew
rlabel metal2 s 10654 -5670 10674 -5650 4 s3_bar
port 315 nsew
rlabel metal2 s 10844 -19834 10865 -19812 4 s4_bar
port 316 nsew
rlabel metal2 s 10882 -14127 10903 -14105 4 s6_bar
port 317 nsew
rlabel metal2 s 10654 -6996 10674 -6976 4 s7_bar
port 318 nsew
rlabel metal2 s 10841 -23636 10862 -23614 4 s8_bar
port 319 nsew
rlabel metal2 s 10610 -27931 10631 -27909 4 s9_bar
port 320 nsew
rlabel metal2 s 10880 -29340 10901 -29318 4 s10_bar
port 321 nsew
rlabel metal2 s 10610 -15538 10631 -15516 4 s5_bar
port 322 nsew
rlabel metal2 s 10610 -15434 10631 -15412 4 s5
port 323 nsew
rlabel metal2 s 10617 -36578 10638 -36556 4 s11
port 324 nsew
rlabel metal2 s 10653 -37695 10674 -37673 4 s15
port 325 nsew
rlabel metal2 s 10616 -36470 10637 -36448 4 s11_bar
port 326 nsew
rlabel metal2 s 10651 -37799 10672 -37777 4 s15_bar
port 327 nsew
rlabel metal2 s 10606 -89535 10627 -89513 4 s25_bar
port 328 nsew
flabel metal2 s 1113 9021 1147 9055 2 FreeSans 2000 0 0 0 CLK0
port 329 nsew
rlabel metal2 s 10614 -128984 10635 -128962 4 s35
port 330 nsew
rlabel metal2 s 10616 -128879 10637 -128857 4 s35_bar
port 331 nsew
rlabel metal2 s 10843 -204765 10863 -204746 4 s52
port 332 nsew
rlabel metal2 s 10611 -200245 10632 -200223 4 s53
port 333 nsew
rlabel metal2 s 10879 -199068 10900 -199046 4 s54
port 334 nsew
rlabel metal2 s 10616 -191702 10636 -191682 4 s55
port 335 nsew
rlabel metal2 s 10840 -208327 10860 -208307 4 s56
port 336 nsew
rlabel metal2 s 10614 -212847 10634 -212828 4 s57
port 337 nsew
rlabel metal2 s 10879 -214027 10900 -214005 4 s58
port 338 nsew
rlabel metal2 s 10615 -221390 10636 -221368 4 s59
port 339 nsew
rlabel metal2 s 10841 -235569 10862 -235547 4 s60
port 340 nsew
rlabel metal2 s 10612 -231047 10633 -231025 4 s61
port 341 nsew
rlabel metal2 s 10879 -229869 10900 -229847 4 s62
port 342 nsew
rlabel metal2 s 10617 -222506 10638 -222484 4 s63
port 343 nsew
rlabel metal2 s 10837 -146844 10858 -146822 4 s40_bar
port 344 nsew
rlabel metal2 s 10608 -151139 10629 -151117 4 s41_bar
port 345 nsew
rlabel metal2 s 10878 -152549 10899 -152527 4 s42_bar
port 346 nsew
rlabel metal2 s 10611 -159680 10632 -159658 4 s43_bar
port 347 nsew
rlabel metal2 s 10842 -173843 10861 -173824 4 s44_bar
port 348 nsew
rlabel metal2 s 10610 -169549 10631 -169527 4 s45_bar
port 349 nsew
rlabel metal2 s 10884 -168137 10903 -168118 4 s46_bar
port 350 nsew
rlabel metal2 s 10614 -161007 10635 -160985 4 s47_bar
port 351 nsew
rlabel metal2 s 10841 -177646 10862 -177624 4 s48_bar
port 352 nsew
rlabel metal2 s 10608 -181941 10629 -181919 4 s49_bar
port 353 nsew
rlabel metal2 s 10883 -183349 10902 -183330 4 s50_bar
port 354 nsew
rlabel metal2 s 10615 -190482 10636 -190460 4 s51_bar
port 355 nsew
rlabel metal2 s 10843 -204644 10862 -204625 4 s52_bar
port 356 nsew
rlabel metal2 s 10611 -200351 10632 -200329 4 s53_bar
port 357 nsew
rlabel metal2 s 10880 -198942 10901 -198920 4 s54_bar
port 358 nsew
rlabel metal2 s 10617 -191808 10636 -191789 4 s55_bar
port 359 nsew
rlabel metal2 s 10844 -208446 10863 -208427 4 s56_bar
port 360 nsew
rlabel metal2 s 10611 -212743 10632 -212721 4 s57_bar
port 361 nsew
rlabel metal2 s 10882 -214153 10903 -214131 4 s58_bar
port 362 nsew
rlabel metal2 s 10612 -221285 10633 -221263 4 s59_bar
port 363 nsew
rlabel metal2 s 10840 -235448 10861 -235426 4 s60_bar
port 364 nsew
rlabel metal2 s 10611 -231153 10632 -231131 4 s61_bar
port 365 nsew
rlabel metal2 s 10882 -229743 10903 -229721 4 s62_bar
port 366 nsew
rlabel metal2 s 10615 -222611 10636 -222589 4 s63_bar
port 367 nsew
rlabel metal2 s 10612 -120442 10633 -120420 4 s33
port 368 nsew
rlabel metal2 s 10876 -121620 10897 -121598 4 s34
port 369 nsew
rlabel metal2 s 10840 -116043 10861 -116021 4 s32_bar
port 370 nsew
rlabel metal2 s 10607 -120336 10628 -120314 4 s33_bar
port 371 nsew
rlabel metal2 s 10877 -121745 10898 -121723 4 s34_bar
port 372 nsew
rlabel metal2 s 10611 -138641 10632 -138619 4 s37
port 373 nsew
rlabel metal2 s 10877 -137462 10898 -137440 4 s38
port 374 nsew
rlabel metal2 s 10613 -130099 10634 -130077 4 s39
port 375 nsew
rlabel metal2 s 10610 -138747 10631 -138725 4 s37_bar
port 376 nsew
rlabel metal2 s 10880 -137336 10901 -137314 4 s38_bar
port 377 nsew
rlabel metal2 s 10612 -130205 10633 -130183 4 s39_bar
port 378 nsew
rlabel metal2 s 10837 -115921 10858 -115899 4 s32
port 379 nsew
rlabel metal2 s 10838 -143042 10859 -143020 4 s36_bar
port 380 nsew
rlabel metal2 s 10839 -143164 10860 -143142 4 s36
port 381 nsew
rlabel metal2 s 10836 -146722 10857 -146700 4 s40
port 382 nsew
rlabel metal2 s 10611 -151244 10632 -151222 4 s41
port 383 nsew
rlabel metal2 s 10878 -152423 10899 -152401 4 s42
port 384 nsew
rlabel metal2 s 10616 -159786 10637 -159764 4 s43
port 385 nsew
rlabel metal2 s 10840 -173965 10861 -173943 4 s44
port 386 nsew
rlabel metal2 s 10611 -169443 10632 -169421 4 s45
port 387 nsew
rlabel metal2 s 10878 -168265 10899 -168243 4 s46
port 388 nsew
rlabel metal2 s 10615 -160900 10635 -160880 4 s47
port 389 nsew
rlabel metal2 s 10840 -177526 10861 -177504 4 s48
port 390 nsew
rlabel metal2 s 10611 -182046 10632 -182024 4 s49
port 391 nsew
rlabel metal2 s 10878 -183225 10898 -183205 4 s50
port 392 nsew
rlabel metal2 s 10616 -190588 10637 -190566 4 s51
port 393 nsew
<< end >>
