magic
tech sky130A
magscale 1 2
timestamp 1676579641
<< nwell >>
rect -181 1080 771 1310
rect -160 390 730 1080
<< pwell >>
rect -146 -278 716 156
rect -171 -430 761 -278
<< nmos >>
rect 0 -170 30 130
rect 150 -170 180 130
rect 540 -170 570 130
<< pmos >>
rect 0 440 30 1040
rect 150 440 180 1040
rect 540 440 570 1040
<< ndiff >>
rect -120 99 0 130
rect -120 65 -77 99
rect -43 65 0 99
rect -120 31 0 65
rect -120 -3 -77 31
rect -43 -3 0 31
rect -120 -37 0 -3
rect -120 -71 -77 -37
rect -43 -71 0 -37
rect -120 -105 0 -71
rect -120 -139 -77 -105
rect -43 -139 0 -105
rect -120 -170 0 -139
rect 30 -170 150 130
rect 180 99 300 130
rect 180 65 223 99
rect 257 65 300 99
rect 180 31 300 65
rect 180 -3 223 31
rect 257 -3 300 31
rect 180 -37 300 -3
rect 180 -71 223 -37
rect 257 -71 300 -37
rect 180 -105 300 -71
rect 180 -139 223 -105
rect 257 -139 300 -105
rect 180 -170 300 -139
rect 420 99 540 130
rect 420 65 463 99
rect 497 65 540 99
rect 420 31 540 65
rect 420 -3 463 31
rect 497 -3 540 31
rect 420 -37 540 -3
rect 420 -71 463 -37
rect 497 -71 540 -37
rect 420 -105 540 -71
rect 420 -139 463 -105
rect 497 -139 540 -105
rect 420 -170 540 -139
rect 570 99 690 130
rect 570 65 613 99
rect 647 65 690 99
rect 570 31 690 65
rect 570 -3 613 31
rect 647 -3 690 31
rect 570 -37 690 -3
rect 570 -71 613 -37
rect 647 -71 690 -37
rect 570 -105 690 -71
rect 570 -139 613 -105
rect 647 -139 690 -105
rect 570 -170 690 -139
<< pdiff >>
rect -120 995 0 1040
rect -120 961 -77 995
rect -43 961 0 995
rect -120 927 0 961
rect -120 893 -77 927
rect -43 893 0 927
rect -120 859 0 893
rect -120 825 -77 859
rect -43 825 0 859
rect -120 791 0 825
rect -120 757 -77 791
rect -43 757 0 791
rect -120 723 0 757
rect -120 689 -77 723
rect -43 689 0 723
rect -120 655 0 689
rect -120 621 -77 655
rect -43 621 0 655
rect -120 587 0 621
rect -120 553 -77 587
rect -43 553 0 587
rect -120 519 0 553
rect -120 485 -77 519
rect -43 485 0 519
rect -120 440 0 485
rect 30 995 150 1040
rect 30 961 73 995
rect 107 961 150 995
rect 30 927 150 961
rect 30 893 73 927
rect 107 893 150 927
rect 30 859 150 893
rect 30 825 73 859
rect 107 825 150 859
rect 30 791 150 825
rect 30 757 73 791
rect 107 757 150 791
rect 30 723 150 757
rect 30 689 73 723
rect 107 689 150 723
rect 30 655 150 689
rect 30 621 73 655
rect 107 621 150 655
rect 30 587 150 621
rect 30 553 73 587
rect 107 553 150 587
rect 30 519 150 553
rect 30 485 73 519
rect 107 485 150 519
rect 30 440 150 485
rect 180 995 300 1040
rect 180 961 223 995
rect 257 961 300 995
rect 180 927 300 961
rect 180 893 223 927
rect 257 893 300 927
rect 180 859 300 893
rect 180 825 223 859
rect 257 825 300 859
rect 180 791 300 825
rect 180 757 223 791
rect 257 757 300 791
rect 180 723 300 757
rect 180 689 223 723
rect 257 689 300 723
rect 180 655 300 689
rect 180 621 223 655
rect 257 621 300 655
rect 180 587 300 621
rect 180 553 223 587
rect 257 553 300 587
rect 180 519 300 553
rect 180 485 223 519
rect 257 485 300 519
rect 180 440 300 485
rect 420 995 540 1040
rect 420 961 463 995
rect 497 961 540 995
rect 420 927 540 961
rect 420 893 463 927
rect 497 893 540 927
rect 420 859 540 893
rect 420 825 463 859
rect 497 825 540 859
rect 420 791 540 825
rect 420 757 463 791
rect 497 757 540 791
rect 420 723 540 757
rect 420 689 463 723
rect 497 689 540 723
rect 420 655 540 689
rect 420 621 463 655
rect 497 621 540 655
rect 420 587 540 621
rect 420 553 463 587
rect 497 553 540 587
rect 420 519 540 553
rect 420 485 463 519
rect 497 485 540 519
rect 420 440 540 485
rect 570 995 690 1040
rect 570 961 613 995
rect 647 961 690 995
rect 570 927 690 961
rect 570 893 613 927
rect 647 893 690 927
rect 570 859 690 893
rect 570 825 613 859
rect 647 825 690 859
rect 570 791 690 825
rect 570 757 613 791
rect 647 757 690 791
rect 570 723 690 757
rect 570 689 613 723
rect 647 689 690 723
rect 570 655 690 689
rect 570 621 613 655
rect 647 621 690 655
rect 570 587 690 621
rect 570 553 613 587
rect 647 553 690 587
rect 570 519 690 553
rect 570 485 613 519
rect 647 485 690 519
rect 570 440 690 485
<< ndiffc >>
rect -77 65 -43 99
rect -77 -3 -43 31
rect -77 -71 -43 -37
rect -77 -139 -43 -105
rect 223 65 257 99
rect 223 -3 257 31
rect 223 -71 257 -37
rect 223 -139 257 -105
rect 463 65 497 99
rect 463 -3 497 31
rect 463 -71 497 -37
rect 463 -139 497 -105
rect 613 65 647 99
rect 613 -3 647 31
rect 613 -71 647 -37
rect 613 -139 647 -105
<< pdiffc >>
rect -77 961 -43 995
rect -77 893 -43 927
rect -77 825 -43 859
rect -77 757 -43 791
rect -77 689 -43 723
rect -77 621 -43 655
rect -77 553 -43 587
rect -77 485 -43 519
rect 73 961 107 995
rect 73 893 107 927
rect 73 825 107 859
rect 73 757 107 791
rect 73 689 107 723
rect 73 621 107 655
rect 73 553 107 587
rect 73 485 107 519
rect 223 961 257 995
rect 223 893 257 927
rect 223 825 257 859
rect 223 757 257 791
rect 223 689 257 723
rect 223 621 257 655
rect 223 553 257 587
rect 223 485 257 519
rect 463 961 497 995
rect 463 893 497 927
rect 463 825 497 859
rect 463 757 497 791
rect 463 689 497 723
rect 463 621 497 655
rect 463 553 497 587
rect 463 485 497 519
rect 613 961 647 995
rect 613 893 647 927
rect 613 825 647 859
rect 613 757 647 791
rect 613 689 647 723
rect 613 621 647 655
rect 613 553 647 587
rect 613 485 647 519
<< psubdiff >>
rect -145 -337 735 -304
rect -145 -371 -122 -337
rect -88 -371 -50 -337
rect -16 -371 22 -337
rect 56 -371 94 -337
rect 128 -371 166 -337
rect 200 -371 238 -337
rect 272 -371 310 -337
rect 344 -371 382 -337
rect 416 -371 454 -337
rect 488 -371 526 -337
rect 560 -371 598 -337
rect 632 -371 670 -337
rect 704 -371 735 -337
rect -145 -404 735 -371
<< nsubdiff >>
rect -145 1241 735 1274
rect -145 1207 -122 1241
rect -88 1207 -50 1241
rect -16 1207 22 1241
rect 56 1207 94 1241
rect 128 1207 166 1241
rect 200 1207 238 1241
rect 272 1207 310 1241
rect 344 1207 382 1241
rect 416 1207 454 1241
rect 488 1207 526 1241
rect 560 1207 598 1241
rect 632 1207 670 1241
rect 704 1207 735 1241
rect -145 1174 735 1207
<< psubdiffcont >>
rect -122 -371 -88 -337
rect -50 -371 -16 -337
rect 22 -371 56 -337
rect 94 -371 128 -337
rect 166 -371 200 -337
rect 238 -371 272 -337
rect 310 -371 344 -337
rect 382 -371 416 -337
rect 454 -371 488 -337
rect 526 -371 560 -337
rect 598 -371 632 -337
rect 670 -371 704 -337
<< nsubdiffcont >>
rect -122 1207 -88 1241
rect -50 1207 -16 1241
rect 22 1207 56 1241
rect 94 1207 128 1241
rect 166 1207 200 1241
rect 238 1207 272 1241
rect 310 1207 344 1241
rect 382 1207 416 1241
rect 454 1207 488 1241
rect 526 1207 560 1241
rect 598 1207 632 1241
rect 670 1207 704 1241
<< poly >>
rect 0 1040 30 1070
rect 150 1040 180 1070
rect 540 1040 570 1070
rect 0 410 30 440
rect -80 387 30 410
rect -80 353 -57 387
rect -23 353 30 387
rect -80 330 30 353
rect 0 130 30 330
rect 150 130 180 440
rect 540 410 570 440
rect 460 387 570 410
rect 460 353 483 387
rect 517 353 570 387
rect 460 330 570 353
rect 540 130 570 330
rect 0 -200 30 -170
rect 150 -200 180 -170
rect 540 -200 570 -170
rect 100 -223 180 -200
rect 100 -257 123 -223
rect 157 -257 180 -223
rect 100 -280 180 -257
<< polycont >>
rect -57 353 -23 387
rect 483 353 517 387
rect 123 -257 157 -223
<< locali >>
rect -145 1241 735 1264
rect -145 1207 -122 1241
rect -88 1207 -50 1241
rect -16 1207 22 1241
rect 56 1207 94 1241
rect 128 1207 166 1241
rect 200 1207 238 1241
rect 272 1207 310 1241
rect 344 1207 382 1241
rect 416 1207 454 1241
rect 488 1207 526 1241
rect 560 1207 598 1241
rect 632 1207 670 1241
rect 704 1207 735 1241
rect -145 1184 735 1207
rect -100 1009 -20 1020
rect -100 961 -77 1009
rect -43 961 -20 1009
rect -100 937 -20 961
rect -100 893 -77 937
rect -43 893 -20 937
rect -100 865 -20 893
rect -100 825 -77 865
rect -43 825 -20 865
rect -100 793 -20 825
rect -100 757 -77 793
rect -43 757 -20 793
rect -100 723 -20 757
rect -100 687 -77 723
rect -43 687 -20 723
rect -100 655 -20 687
rect -100 615 -77 655
rect -43 615 -20 655
rect -100 587 -20 615
rect -100 543 -77 587
rect -43 543 -20 587
rect -100 519 -20 543
rect -100 471 -77 519
rect -43 471 -20 519
rect -100 460 -20 471
rect 50 995 130 1020
rect 50 961 73 995
rect 107 961 130 995
rect 50 927 130 961
rect 50 893 73 927
rect 107 893 130 927
rect 50 859 130 893
rect 50 825 73 859
rect 107 825 130 859
rect 50 791 130 825
rect 50 757 73 791
rect 107 757 130 791
rect 50 723 130 757
rect 50 689 73 723
rect 107 689 130 723
rect 50 655 130 689
rect 50 621 73 655
rect 107 621 130 655
rect 50 587 130 621
rect 50 553 73 587
rect 107 553 130 587
rect 50 519 130 553
rect 50 485 73 519
rect 107 485 130 519
rect 50 460 130 485
rect 200 1009 280 1020
rect 200 961 223 1009
rect 257 961 280 1009
rect 200 937 280 961
rect 200 893 223 937
rect 257 893 280 937
rect 200 865 280 893
rect 200 825 223 865
rect 257 825 280 865
rect 200 793 280 825
rect 200 757 223 793
rect 257 757 280 793
rect 200 723 280 757
rect 200 687 223 723
rect 257 687 280 723
rect 200 655 280 687
rect 200 615 223 655
rect 257 615 280 655
rect 200 587 280 615
rect 200 543 223 587
rect 257 543 280 587
rect 200 519 280 543
rect 200 471 223 519
rect 257 471 280 519
rect 200 460 280 471
rect 440 1009 520 1020
rect 440 961 463 1009
rect 497 961 520 1009
rect 440 937 520 961
rect 440 893 463 937
rect 497 893 520 937
rect 440 865 520 893
rect 440 825 463 865
rect 497 825 520 865
rect 440 793 520 825
rect 440 757 463 793
rect 497 757 520 793
rect 440 723 520 757
rect 440 687 463 723
rect 497 687 520 723
rect 440 655 520 687
rect 440 615 463 655
rect 497 615 520 655
rect 440 587 520 615
rect 440 543 463 587
rect 497 543 520 587
rect 440 519 520 543
rect 440 471 463 519
rect 497 471 520 519
rect 440 460 520 471
rect 590 995 670 1020
rect 590 961 613 995
rect 647 961 670 995
rect 590 927 670 961
rect 590 893 613 927
rect 647 893 670 927
rect 590 859 670 893
rect 590 825 613 859
rect 647 825 670 859
rect 590 791 670 825
rect 590 757 613 791
rect 647 757 670 791
rect 590 723 670 757
rect 590 689 613 723
rect 647 689 670 723
rect 590 655 670 689
rect 590 621 613 655
rect 647 621 670 655
rect 590 587 670 621
rect 590 553 613 587
rect 647 553 670 587
rect 590 519 670 553
rect 590 485 613 519
rect 647 485 670 519
rect 590 460 670 485
rect -80 387 0 410
rect -80 353 -57 387
rect -23 353 0 387
rect -80 330 0 353
rect 70 390 110 460
rect 460 390 540 410
rect 70 387 540 390
rect 70 353 483 387
rect 517 353 540 387
rect 70 350 540 353
rect 220 110 260 350
rect 460 330 540 350
rect 610 110 650 460
rect -100 99 -20 110
rect -100 35 -77 99
rect -43 35 -20 99
rect -100 31 -20 35
rect -100 -71 -77 31
rect -43 -71 -20 31
rect -100 -75 -20 -71
rect -100 -139 -77 -75
rect -43 -139 -20 -75
rect -100 -150 -20 -139
rect 200 99 280 110
rect 200 65 223 99
rect 257 65 280 99
rect 200 31 280 65
rect 200 -3 223 31
rect 257 -3 280 31
rect 200 -37 280 -3
rect 200 -71 223 -37
rect 257 -71 280 -37
rect 200 -105 280 -71
rect 200 -139 223 -105
rect 257 -139 280 -105
rect 200 -150 280 -139
rect 440 99 520 110
rect 440 35 463 99
rect 497 35 520 99
rect 440 31 520 35
rect 440 -71 463 31
rect 497 -71 520 31
rect 440 -75 520 -71
rect 440 -139 463 -75
rect 497 -139 520 -75
rect 440 -150 520 -139
rect 590 99 670 110
rect 590 65 613 99
rect 647 65 670 99
rect 590 31 670 65
rect 590 -3 613 31
rect 647 -3 670 31
rect 590 -37 670 -3
rect 590 -71 613 -37
rect 647 -71 670 -37
rect 590 -105 670 -71
rect 590 -139 613 -105
rect 647 -139 670 -105
rect 590 -150 670 -139
rect 100 -223 180 -200
rect 100 -257 123 -223
rect 157 -257 180 -223
rect 100 -280 180 -257
rect -145 -337 735 -314
rect -145 -371 -122 -337
rect -88 -371 -50 -337
rect -16 -371 22 -337
rect 56 -371 94 -337
rect 128 -371 166 -337
rect 200 -371 238 -337
rect 272 -371 310 -337
rect 344 -371 382 -337
rect 416 -371 454 -337
rect 488 -371 526 -337
rect 560 -371 598 -337
rect 632 -371 670 -337
rect 704 -371 735 -337
rect -145 -394 735 -371
<< viali >>
rect -122 1207 -88 1241
rect -50 1207 -16 1241
rect 22 1207 56 1241
rect 94 1207 128 1241
rect 166 1207 200 1241
rect 238 1207 272 1241
rect 310 1207 344 1241
rect 382 1207 416 1241
rect 454 1207 488 1241
rect 526 1207 560 1241
rect 598 1207 632 1241
rect 670 1207 704 1241
rect -77 995 -43 1009
rect -77 975 -43 995
rect -77 927 -43 937
rect -77 903 -43 927
rect -77 859 -43 865
rect -77 831 -43 859
rect -77 791 -43 793
rect -77 759 -43 791
rect -77 689 -43 721
rect -77 687 -43 689
rect -77 621 -43 649
rect -77 615 -43 621
rect -77 553 -43 577
rect -77 543 -43 553
rect -77 485 -43 505
rect -77 471 -43 485
rect 223 995 257 1009
rect 223 975 257 995
rect 223 927 257 937
rect 223 903 257 927
rect 223 859 257 865
rect 223 831 257 859
rect 223 791 257 793
rect 223 759 257 791
rect 223 689 257 721
rect 223 687 257 689
rect 223 621 257 649
rect 223 615 257 621
rect 223 553 257 577
rect 223 543 257 553
rect 223 485 257 505
rect 223 471 257 485
rect 463 995 497 1009
rect 463 975 497 995
rect 463 927 497 937
rect 463 903 497 927
rect 463 859 497 865
rect 463 831 497 859
rect 463 791 497 793
rect 463 759 497 791
rect 463 689 497 721
rect 463 687 497 689
rect 463 621 497 649
rect 463 615 497 621
rect 463 553 497 577
rect 463 543 497 553
rect 463 485 497 505
rect 463 471 497 485
rect -77 65 -43 69
rect -77 35 -43 65
rect -77 -37 -43 -3
rect -77 -105 -43 -75
rect -77 -109 -43 -105
rect 463 65 497 69
rect 463 35 497 65
rect 463 -37 497 -3
rect 463 -105 497 -75
rect 463 -109 497 -105
rect -122 -371 -88 -337
rect -50 -371 -16 -337
rect 22 -371 56 -337
rect 94 -371 128 -337
rect 166 -371 200 -337
rect 238 -371 272 -337
rect 310 -371 344 -337
rect 382 -371 416 -337
rect 454 -371 488 -337
rect 526 -371 560 -337
rect 598 -371 632 -337
rect 670 -371 704 -337
<< metal1 >>
rect -145 1241 735 1274
rect -145 1207 -122 1241
rect -88 1207 -50 1241
rect -16 1207 22 1241
rect 56 1207 94 1241
rect 128 1207 166 1241
rect 200 1207 238 1241
rect 272 1207 310 1241
rect 344 1207 382 1241
rect 416 1207 454 1241
rect 488 1207 526 1241
rect 560 1207 598 1241
rect 632 1207 670 1241
rect 704 1207 735 1241
rect -145 1174 735 1207
rect -80 1020 -40 1174
rect 221 1020 261 1174
rect 460 1020 500 1174
rect -100 1009 -20 1020
rect -100 975 -77 1009
rect -43 975 -20 1009
rect -100 937 -20 975
rect -100 903 -77 937
rect -43 903 -20 937
rect -100 865 -20 903
rect -100 831 -77 865
rect -43 831 -20 865
rect -100 793 -20 831
rect -100 759 -77 793
rect -43 759 -20 793
rect -100 721 -20 759
rect -100 687 -77 721
rect -43 687 -20 721
rect -100 649 -20 687
rect -100 615 -77 649
rect -43 615 -20 649
rect -100 577 -20 615
rect -100 543 -77 577
rect -43 543 -20 577
rect -100 505 -20 543
rect -100 471 -77 505
rect -43 471 -20 505
rect -100 460 -20 471
rect 200 1009 280 1020
rect 200 975 223 1009
rect 257 975 280 1009
rect 200 937 280 975
rect 200 903 223 937
rect 257 903 280 937
rect 200 865 280 903
rect 200 831 223 865
rect 257 831 280 865
rect 200 793 280 831
rect 200 759 223 793
rect 257 759 280 793
rect 200 721 280 759
rect 200 687 223 721
rect 257 687 280 721
rect 200 649 280 687
rect 200 615 223 649
rect 257 615 280 649
rect 200 577 280 615
rect 200 543 223 577
rect 257 543 280 577
rect 200 505 280 543
rect 200 471 223 505
rect 257 471 280 505
rect 200 460 280 471
rect 440 1009 520 1020
rect 440 975 463 1009
rect 497 975 520 1009
rect 440 937 520 975
rect 440 903 463 937
rect 497 903 520 937
rect 440 865 520 903
rect 440 831 463 865
rect 497 831 520 865
rect 440 793 520 831
rect 440 759 463 793
rect 497 759 520 793
rect 440 721 520 759
rect 440 687 463 721
rect 497 687 520 721
rect 440 649 520 687
rect 440 615 463 649
rect 497 615 520 649
rect 440 577 520 615
rect 440 543 463 577
rect 497 543 520 577
rect 440 505 520 543
rect 440 471 463 505
rect 497 471 520 505
rect 440 460 520 471
rect -100 69 -20 110
rect -100 35 -77 69
rect -43 35 -20 69
rect -100 -3 -20 35
rect -100 -37 -77 -3
rect -43 -37 -20 -3
rect -100 -75 -20 -37
rect -100 -109 -77 -75
rect -43 -109 -20 -75
rect -100 -150 -20 -109
rect 440 69 520 110
rect 440 35 463 69
rect 497 35 520 69
rect 440 -3 520 35
rect 440 -37 463 -3
rect 497 -37 520 -3
rect 440 -75 520 -37
rect 440 -109 463 -75
rect 497 -109 520 -75
rect 440 -150 520 -109
rect -80 -304 -40 -150
rect 460 -304 500 -150
rect -145 -337 735 -304
rect -145 -371 -122 -337
rect -88 -371 -50 -337
rect -16 -371 22 -337
rect 56 -371 94 -337
rect 128 -371 166 -337
rect 200 -371 238 -337
rect 272 -371 310 -337
rect 344 -371 382 -337
rect 416 -371 454 -337
rect 488 -371 526 -337
rect 560 -371 598 -337
rect 632 -371 670 -337
rect 704 -371 735 -337
rect -145 -404 735 -371
<< labels >>
rlabel metal1 s 235 -374 275 -334 4 GND!
port 1 nsew
rlabel metal1 s 235 1204 275 1244 4 VDD
port 2 nsew
flabel locali s 613 353 647 387 2 FreeSans 2000 0 0 0 AND
port 3 nsew
flabel locali s 123 -257 157 -223 2 FreeSans 2000 0 0 0 A
port 4 nsew
flabel locali s -57 353 -23 387 2 FreeSans 2000 0 0 0 B
port 5 nsew
<< properties >>
string path 2.400 5.100 2.400 5.870 
<< end >>
