magic
tech sky130A
magscale 1 2
timestamp 1676906723
<< nwell >>
rect 252 1190 701 1420
rect 330 500 680 1190
<< pwell >>
rect 344 -168 666 266
rect 262 -320 702 -168
<< nmos >>
rect 490 -60 520 240
<< pmos >>
rect 490 550 520 1150
<< ndiff >>
rect 370 209 490 240
rect 370 175 413 209
rect 447 175 490 209
rect 370 141 490 175
rect 370 107 413 141
rect 447 107 490 141
rect 370 73 490 107
rect 370 39 413 73
rect 447 39 490 73
rect 370 5 490 39
rect 370 -29 413 5
rect 447 -29 490 5
rect 370 -60 490 -29
rect 520 209 640 240
rect 520 175 563 209
rect 597 175 640 209
rect 520 141 640 175
rect 520 107 563 141
rect 597 107 640 141
rect 520 73 640 107
rect 520 39 563 73
rect 597 39 640 73
rect 520 5 640 39
rect 520 -29 563 5
rect 597 -29 640 5
rect 520 -60 640 -29
<< pdiff >>
rect 370 1105 490 1150
rect 370 1071 413 1105
rect 447 1071 490 1105
rect 370 1037 490 1071
rect 370 1003 413 1037
rect 447 1003 490 1037
rect 370 969 490 1003
rect 370 935 413 969
rect 447 935 490 969
rect 370 901 490 935
rect 370 867 413 901
rect 447 867 490 901
rect 370 833 490 867
rect 370 799 413 833
rect 447 799 490 833
rect 370 765 490 799
rect 370 731 413 765
rect 447 731 490 765
rect 370 697 490 731
rect 370 663 413 697
rect 447 663 490 697
rect 370 629 490 663
rect 370 595 413 629
rect 447 595 490 629
rect 370 550 490 595
rect 520 1105 640 1150
rect 520 1071 563 1105
rect 597 1071 640 1105
rect 520 1037 640 1071
rect 520 1003 563 1037
rect 597 1003 640 1037
rect 520 969 640 1003
rect 520 935 563 969
rect 597 935 640 969
rect 520 901 640 935
rect 520 867 563 901
rect 597 867 640 901
rect 520 833 640 867
rect 520 799 563 833
rect 597 799 640 833
rect 520 765 640 799
rect 520 731 563 765
rect 597 731 640 765
rect 520 697 640 731
rect 520 663 563 697
rect 597 663 640 697
rect 520 629 640 663
rect 520 595 563 629
rect 597 595 640 629
rect 520 550 640 595
<< ndiffc >>
rect 413 175 447 209
rect 413 107 447 141
rect 413 39 447 73
rect 413 -29 447 5
rect 563 175 597 209
rect 563 107 597 141
rect 563 39 597 73
rect 563 -29 597 5
<< pdiffc >>
rect 413 1071 447 1105
rect 413 1003 447 1037
rect 413 935 447 969
rect 413 867 447 901
rect 413 799 447 833
rect 413 731 447 765
rect 413 663 447 697
rect 413 595 447 629
rect 563 1071 597 1105
rect 563 1003 597 1037
rect 563 935 597 969
rect 563 867 597 901
rect 563 799 597 833
rect 563 731 597 765
rect 563 663 597 697
rect 563 595 597 629
<< psubdiff >>
rect 288 -227 676 -194
rect 288 -261 326 -227
rect 360 -261 398 -227
rect 432 -261 470 -227
rect 504 -261 542 -227
rect 576 -261 614 -227
rect 648 -261 676 -227
rect 288 -294 676 -261
<< nsubdiff >>
rect 288 1351 665 1384
rect 288 1317 326 1351
rect 360 1317 398 1351
rect 432 1317 470 1351
rect 504 1317 542 1351
rect 576 1317 614 1351
rect 648 1317 665 1351
rect 288 1284 665 1317
<< psubdiffcont >>
rect 326 -261 360 -227
rect 398 -261 432 -227
rect 470 -261 504 -227
rect 542 -261 576 -227
rect 614 -261 648 -227
<< nsubdiffcont >>
rect 326 1317 360 1351
rect 398 1317 432 1351
rect 470 1317 504 1351
rect 542 1317 576 1351
rect 614 1317 648 1351
<< poly >>
rect 490 1150 520 1180
rect 490 520 520 550
rect 410 497 520 520
rect 410 463 433 497
rect 467 463 520 497
rect 410 440 520 463
rect 490 240 520 440
rect 490 -90 520 -60
<< polycont >>
rect 433 463 467 497
<< locali >>
rect 288 1351 665 1374
rect 288 1317 326 1351
rect 360 1317 398 1351
rect 432 1317 470 1351
rect 504 1317 542 1351
rect 576 1317 614 1351
rect 648 1317 665 1351
rect 288 1294 665 1317
rect 390 1119 470 1130
rect 390 1071 413 1119
rect 447 1071 470 1119
rect 390 1047 470 1071
rect 390 1003 413 1047
rect 447 1003 470 1047
rect 390 975 470 1003
rect 390 935 413 975
rect 447 935 470 975
rect 390 903 470 935
rect 390 867 413 903
rect 447 867 470 903
rect 390 833 470 867
rect 390 797 413 833
rect 447 797 470 833
rect 390 765 470 797
rect 390 725 413 765
rect 447 725 470 765
rect 390 697 470 725
rect 390 653 413 697
rect 447 653 470 697
rect 390 629 470 653
rect 390 581 413 629
rect 447 581 470 629
rect 390 570 470 581
rect 540 1105 620 1130
rect 540 1071 563 1105
rect 597 1071 620 1105
rect 540 1037 620 1071
rect 540 1003 563 1037
rect 597 1003 620 1037
rect 540 969 620 1003
rect 540 935 563 969
rect 597 935 620 969
rect 540 901 620 935
rect 540 867 563 901
rect 597 867 620 901
rect 540 833 620 867
rect 540 799 563 833
rect 597 799 620 833
rect 540 765 620 799
rect 540 731 563 765
rect 597 731 620 765
rect 540 697 620 731
rect 540 663 563 697
rect 597 663 620 697
rect 540 629 620 663
rect 540 595 563 629
rect 597 595 620 629
rect 540 570 620 595
rect 410 500 490 520
rect 288 497 490 500
rect 288 463 433 497
rect 467 463 490 497
rect 288 460 490 463
rect 410 440 490 460
rect 560 220 600 570
rect 390 209 470 220
rect 390 145 413 209
rect 447 145 470 209
rect 390 141 470 145
rect 390 39 413 141
rect 447 39 470 141
rect 390 35 470 39
rect 390 -29 413 35
rect 447 -29 470 35
rect 390 -40 470 -29
rect 540 209 620 220
rect 540 175 563 209
rect 597 175 620 209
rect 540 141 620 175
rect 540 107 563 141
rect 597 107 620 141
rect 540 73 620 107
rect 540 39 563 73
rect 597 39 620 73
rect 540 5 620 39
rect 540 -29 563 5
rect 597 -29 620 5
rect 540 -40 620 -29
rect 288 -227 676 -204
rect 288 -261 326 -227
rect 360 -261 398 -227
rect 432 -261 470 -227
rect 504 -261 542 -227
rect 576 -261 614 -227
rect 648 -261 676 -227
rect 288 -284 676 -261
<< viali >>
rect 326 1317 360 1351
rect 398 1317 432 1351
rect 470 1317 504 1351
rect 542 1317 576 1351
rect 614 1317 648 1351
rect 413 1105 447 1119
rect 413 1085 447 1105
rect 413 1037 447 1047
rect 413 1013 447 1037
rect 413 969 447 975
rect 413 941 447 969
rect 413 901 447 903
rect 413 869 447 901
rect 413 799 447 831
rect 413 797 447 799
rect 413 731 447 759
rect 413 725 447 731
rect 413 663 447 687
rect 413 653 447 663
rect 413 595 447 615
rect 413 581 447 595
rect 413 175 447 179
rect 413 145 447 175
rect 413 73 447 107
rect 413 5 447 35
rect 413 1 447 5
rect 326 -261 360 -227
rect 398 -261 432 -227
rect 470 -261 504 -227
rect 542 -261 576 -227
rect 614 -261 648 -227
<< metal1 >>
rect 288 1351 665 1384
rect 288 1317 326 1351
rect 360 1317 398 1351
rect 432 1317 470 1351
rect 504 1317 542 1351
rect 576 1317 614 1351
rect 648 1317 665 1351
rect 288 1284 665 1317
rect 410 1130 450 1284
rect 390 1119 470 1130
rect 390 1085 413 1119
rect 447 1085 470 1119
rect 390 1047 470 1085
rect 390 1013 413 1047
rect 447 1013 470 1047
rect 390 975 470 1013
rect 390 941 413 975
rect 447 941 470 975
rect 390 903 470 941
rect 390 869 413 903
rect 447 869 470 903
rect 390 831 470 869
rect 390 797 413 831
rect 447 797 470 831
rect 390 759 470 797
rect 390 725 413 759
rect 447 725 470 759
rect 390 687 470 725
rect 390 653 413 687
rect 447 653 470 687
rect 390 615 470 653
rect 390 581 413 615
rect 447 581 470 615
rect 390 570 470 581
rect 390 179 470 220
rect 390 145 413 179
rect 447 145 470 179
rect 390 107 470 145
rect 390 73 413 107
rect 447 73 470 107
rect 390 35 470 73
rect 390 1 413 35
rect 447 1 470 35
rect 390 -40 470 1
rect 410 -194 450 -40
rect 288 -227 676 -194
rect 288 -261 326 -227
rect 360 -261 398 -227
rect 432 -261 470 -227
rect 504 -261 542 -227
rect 576 -261 614 -227
rect 648 -261 676 -227
rect 288 -294 676 -261
<< labels >>
flabel locali s 433 463 467 497 2 FreeSans 2500 0 0 0 A
port 1 nsew
flabel locali s 563 368 597 402 2 FreeSans 3125 0 0 0 OUT
port 2 nsew
flabel metal1 s 470 1317 504 1351 2 FreeSans 2500 0 0 0 VDD
port 3 nsew
flabel metal1 s 470 -261 504 -227 2 FreeSans 2500 0 0 0 GND
port 4 nsew
<< end >>
