magic
tech sky130A
magscale 1 2
timestamp 1670883550
<< xpolycontact >>
rect -35 332 35 764
rect -35 -764 35 -332
<< xpolyres >>
rect -35 -332 35 332
<< viali >>
rect -19 349 19 746
rect -19 -746 19 -349
<< metal1 >>
rect -25 746 25 758
rect -25 349 -19 746
rect 19 349 25 746
rect -25 337 25 349
rect -25 -349 25 -337
rect -25 -746 -19 -349
rect 19 -746 25 -349
rect -25 -758 25 -746
<< res0p35 >>
rect -37 -334 37 334
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 3.32 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 20.046k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
