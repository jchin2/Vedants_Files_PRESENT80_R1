magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -10 -10 30 30
<< l67d20 >>
rect -10 -10 30 30
<< l67d44 >>
rect 2 2 19 19
<< l68d20 >>
rect -10 -10 30 30
<< l69d20 >>
rect -10 -10 30 30
<< end >>
