* NGSPICE file created from EESPFAL_4in_XOR_flat.ext - technology: sky130A

.subckt EESPFAL_4in_XOR_flat x0 x0_bar k0 k0_bar x1 x1_bar k1 k1_bar x2 x2_bar k2
+ k2_bar x3 x3_bar k3 k3_bar XOR0_bar XOR0 XOR1_bar XOR1 XOR2_bar XOR2 XOR3_bar XOR3
+ GND Dis CLK
X0 XOR1_bar.t5 XOR1.t6 CLK.t42 CLK.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 XOR2_bar.t5 XOR2.t6 CLK.t27 CLK.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_420_n1950# k2_bar.t0 XOR2.t1 GND.t35 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X3 CLK.t11 XOR0.t6 XOR0_bar.t2 CLK.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 XOR0_bar.t3 Dis.t0 GND.t21 GND.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 CLK.t31 x2.t0 a_420_n1950# GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 XOR3_bar.t3 Dis.t1 GND.t2 GND.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n840_410# x0.t0 CLK.t23 GND.t18 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n840_n2630# x3.t0 CLK.t35 GND.t31 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X9 XOR3.t2 XOR3_bar.t6 CLK.t14 CLK.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_n1140_410# k0_bar.t0 XOR0_bar.t4 GND.t27 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X11 XOR2.t2 XOR2_bar.t6 GND.t36 GND.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK.t19 x3_bar.t0 a_n1140_n2630# GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X13 a_420_410# k0_bar.t1 XOR0.t1 GND.t19 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X14 GND.t20 Dis.t2 XOR0.t2 GND.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_720_n270# x1_bar.t0 CLK.t28 GND.t4 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X16 XOR1.t3 k1.t0 a_720_n270# GND.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 XOR0.t4 XOR0_bar.t6 CLK.t34 CLK.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_n840_n270# x1.t0 CLK.t38 GND.t18 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X19 GND.t8 Dis.t3 XOR1.t2 GND.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X20 a_720_410# x0_bar.t0 CLK.t12 GND.t4 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X21 a_720_n2630# x3_bar.t1 CLK.t22 GND.t17 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X22 CLK.t3 x1_bar.t1 a_n1140_n270# GND.t3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X23 XOR3.t4 k3.t0 a_720_n2630# GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X24 CLK.t25 XOR2.t7 XOR2_bar.t4 CLK.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X25 a_n1140_n1950# k2_bar.t1 XOR2_bar.t0 GND.t34 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X26 XOR1.t5 XOR1_bar.t6 GND.t38 GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X27 CLK.t8 XOR1_bar.t7 XOR1.t1 CLK.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X28 GND.t6 XOR3.t6 XOR3_bar.t0 GND.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X29 CLK.t18 XOR3_bar.t7 XOR3.t1 CLK.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X30 GND.t13 Dis.t4 XOR2.t4 GND.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X31 XOR3_bar.t4 k3.t1 a_n840_n2630# GND.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X32 XOR0_bar.t1 XOR0.t7 CLK.t16 CLK.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X33 a_n1140_n270# k1_bar.t0 XOR1_bar.t2 GND.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X34 a_420_n2630# k3_bar.t0 XOR3.t5 GND.t35 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X35 XOR3_bar.t1 XOR3.t7 CLK.t21 CLK.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X36 GND.t39 XOR1.t7 XOR1_bar.t3 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X37 XOR1.t0 XOR1_bar.t8 CLK.t2 CLK.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X38 XOR2.t3 XOR2_bar.t7 CLK.t9 CLK.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X39 XOR2_bar.t2 Dis.t5 GND.t30 GND.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X40 CLK.t32 x3.t1 a_420_n2630# GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X41 CLK.t7 XOR0_bar.t7 XOR0.t0 CLK.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X42 CLK.t40 x2_bar.t0 a_n1140_n1950# GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X43 a_n840_n1950# x2.t1 CLK.t43 GND.t31 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X44 XOR3.t0 XOR3_bar.t8 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X45 XOR0_bar.t5 k0.t0 a_n840_410# GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X46 GND.t23 XOR0.t8 XOR0_bar.t0 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X47 CLK.t36 x0_bar.t1 a_n1140_410# GND.t3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X48 CLK.t41 XOR1.t8 XOR1_bar.t4 CLK.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X49 a_720_n1950# x2_bar.t1 CLK.t39 GND.t17 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X50 XOR2.t5 k2.t0 a_720_n1950# GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X51 XOR0.t3 XOR0_bar.t8 GND.t25 GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X52 XOR1_bar.t0 Dis.t6 GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X53 CLK.t5 XOR2_bar.t8 XOR2.t0 CLK.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X54 a_n1140_n2630# k3_bar.t1 XOR3_bar.t5 GND.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X55 CLK.t0 x0.t1 a_420_410# GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X56 CLK.t30 XOR3.t8 XOR3_bar.t2 CLK.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X57 GND.t37 XOR2.t8 XOR2_bar.t3 GND.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X58 a_420_n270# k1_bar.t1 XOR1.t4 GND.t19 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X59 XOR2_bar.t1 k2.t1 a_n840_n1950# GND.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X60 GND.t12 Dis.t7 XOR3.t3 GND.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X61 XOR0.t5 k0.t1 a_720_410# GND.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X62 XOR1_bar.t1 k1.t1 a_n840_n270# GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X63 CLK.t37 x1.t1 a_420_n270# GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
R0 XOR1.t8 XOR1.t6 819.4
R1 XOR1.n5 XOR1.t8 514.133
R2 XOR1.n5 XOR1.t7 305.266
R3 XOR1.n3 XOR1.n2 192
R4 XOR1.n4 XOR1.n1 166.734
R5 XOR1.n4 XOR1.n3 105.6
R6 XOR1.n2 XOR1.t3 97.937
R7 XOR1.n3 XOR1.t4 97.937
R8 XOR1.n6 XOR1.n5 76
R9 XOR1.n4 XOR1.n0 73.937
R10 XOR1.n6 XOR1.n4 57.6
R11 XOR1.n1 XOR1.t1 39.4
R12 XOR1.n1 XOR1.t0 39.4
R13 XOR1.n0 XOR1.t2 24
R14 XOR1.n0 XOR1.t5 24
R15 XOR1.n2 XOR1 9.92
R16 XOR1 XOR1.n6 3.2
R17 CLK.n93 CLK.t18 44.338
R18 CLK.n64 CLK.t21 44.338
R19 CLK.n209 CLK.t8 44.338
R20 CLK.n180 CLK.t42 44.338
R21 CLK.n337 CLK.t16 44.337
R22 CLK.n280 CLK.t7 44.337
R23 CLK.n209 CLK.t5 44.337
R24 CLK.n180 CLK.t27 44.337
R25 CLK.n0 CLK.t34 39.4
R26 CLK.n0 CLK.t11 39.4
R27 CLK.n25 CLK.t14 39.4
R28 CLK.n25 CLK.t30 39.4
R29 CLK.n140 CLK.t9 39.4
R30 CLK.n140 CLK.t25 39.4
R31 CLK.n139 CLK.t2 39.4
R32 CLK.n139 CLK.t41 39.4
R33 CLK.n281 CLK.t6 24.568
R34 CLK.n338 CLK.t15 24.568
R35 CLK.n89 CLK.t17 24.568
R36 CLK.n65 CLK.t20 24.568
R37 CLK.n297 CLK.t23 24
R38 CLK.n297 CLK.t36 24
R39 CLK.n4 CLK.t28 24
R40 CLK.n4 CLK.t37 24
R41 CLK.n10 CLK.t22 24
R42 CLK.n10 CLK.t32 24
R43 CLK.n26 CLK.t35 24
R44 CLK.n26 CLK.t19 24
R45 CLK.n8 CLK.t39 24
R46 CLK.n8 CLK.t31 24
R47 CLK.n142 CLK.t43 24
R48 CLK.n142 CLK.t40 24
R49 CLK.n141 CLK.t38 24
R50 CLK.n141 CLK.t3 24
R51 CLK.n2 CLK.t12 24
R52 CLK.n2 CLK.t0 24
R53 CLK.n205 CLK.t4 14.843
R54 CLK.n181 CLK.t26 14.843
R55 CLK.n79 CLK.n76 12.8
R56 CLK.n195 CLK.n192 12.8
R57 CLK.n15 CLK.n14 8.855
R58 CLK.n19 CLK.n18 8.855
R59 CLK.n18 CLK.n17 8.855
R60 CLK.n23 CLK.n22 8.855
R61 CLK.n22 CLK.n21 8.855
R62 CLK.n116 CLK.n115 8.855
R63 CLK.n115 CLK.n114 8.855
R64 CLK.n112 CLK.n111 8.855
R65 CLK.n111 CLK.n110 8.855
R66 CLK.n108 CLK.n107 8.855
R67 CLK.n107 CLK.n106 8.855
R68 CLK.n104 CLK.n103 8.855
R69 CLK.n103 CLK.n102 8.855
R70 CLK.n100 CLK.n99 8.855
R71 CLK.n99 CLK.n98 8.855
R72 CLK.n96 CLK.n95 8.855
R73 CLK.n95 CLK.n94 8.855
R74 CLK.n91 CLK.n90 8.855
R75 CLK.n90 CLK.n89 8.855
R76 CLK.n87 CLK.n86 8.855
R77 CLK.n86 CLK.n85 8.855
R78 CLK.n83 CLK.n82 8.855
R79 CLK.n82 CLK.n81 8.855
R80 CLK.n79 CLK.n78 8.855
R81 CLK.n78 CLK.n77 8.855
R82 CLK.n76 CLK.n75 8.855
R83 CLK.n75 CLK.n74 8.855
R84 CLK.n71 CLK.n70 8.855
R85 CLK.n70 CLK.n69 8.855
R86 CLK.n67 CLK.n66 8.855
R87 CLK.n66 CLK.n65 8.855
R88 CLK.n62 CLK.n61 8.855
R89 CLK.n61 CLK.n60 8.855
R90 CLK.n58 CLK.n57 8.855
R91 CLK.n57 CLK.n56 8.855
R92 CLK.n54 CLK.n53 8.855
R93 CLK.n53 CLK.n52 8.855
R94 CLK.n50 CLK.n49 8.855
R95 CLK.n49 CLK.n48 8.855
R96 CLK.n46 CLK.n45 8.855
R97 CLK.n45 CLK.n44 8.855
R98 CLK.n42 CLK.n41 8.855
R99 CLK.n41 CLK.n40 8.855
R100 CLK.n37 CLK.n36 8.855
R101 CLK.n36 CLK.n35 8.855
R102 CLK.n33 CLK.n32 8.855
R103 CLK.n32 CLK.n31 8.855
R104 CLK.n29 CLK.n28 8.855
R105 CLK.n129 CLK.n128 8.855
R106 CLK.n133 CLK.n132 8.855
R107 CLK.n132 CLK.n131 8.855
R108 CLK.n137 CLK.n136 8.855
R109 CLK.n136 CLK.n135 8.855
R110 CLK.n232 CLK.n231 8.855
R111 CLK.n231 CLK.n230 8.855
R112 CLK.n228 CLK.n227 8.855
R113 CLK.n227 CLK.n226 8.855
R114 CLK.n224 CLK.n223 8.855
R115 CLK.n223 CLK.n222 8.855
R116 CLK.n220 CLK.n219 8.855
R117 CLK.n219 CLK.n218 8.855
R118 CLK.n216 CLK.n215 8.855
R119 CLK.n215 CLK.n214 8.855
R120 CLK.n212 CLK.n211 8.855
R121 CLK.n211 CLK.n210 8.855
R122 CLK.n207 CLK.n206 8.855
R123 CLK.n206 CLK.n205 8.855
R124 CLK.n203 CLK.n202 8.855
R125 CLK.n202 CLK.n201 8.855
R126 CLK.n199 CLK.n198 8.855
R127 CLK.n198 CLK.n197 8.855
R128 CLK.n195 CLK.n194 8.855
R129 CLK.n194 CLK.n193 8.855
R130 CLK.n192 CLK.n191 8.855
R131 CLK.n191 CLK.n190 8.855
R132 CLK.n187 CLK.n186 8.855
R133 CLK.n186 CLK.n185 8.855
R134 CLK.n183 CLK.n182 8.855
R135 CLK.n182 CLK.n181 8.855
R136 CLK.n178 CLK.n177 8.855
R137 CLK.n177 CLK.n176 8.855
R138 CLK.n174 CLK.n173 8.855
R139 CLK.n173 CLK.n172 8.855
R140 CLK.n170 CLK.n169 8.855
R141 CLK.n169 CLK.n168 8.855
R142 CLK.n166 CLK.n165 8.855
R143 CLK.n165 CLK.n164 8.855
R144 CLK.n162 CLK.n161 8.855
R145 CLK.n161 CLK.n160 8.855
R146 CLK.n158 CLK.n157 8.855
R147 CLK.n157 CLK.n156 8.855
R148 CLK.n153 CLK.n152 8.855
R149 CLK.n152 CLK.n151 8.855
R150 CLK.n149 CLK.n148 8.855
R151 CLK.n148 CLK.n147 8.855
R152 CLK.n145 CLK.n144 8.855
R153 CLK.n245 CLK.n244 8.855
R154 CLK.n249 CLK.n248 8.855
R155 CLK.n248 CLK.n247 8.855
R156 CLK.n253 CLK.n252 8.855
R157 CLK.n252 CLK.n251 8.855
R158 CLK.n258 CLK.n257 8.855
R159 CLK.n257 CLK.n256 8.855
R160 CLK.n262 CLK.n261 8.855
R161 CLK.n261 CLK.n260 8.855
R162 CLK.n266 CLK.n265 8.855
R163 CLK.n265 CLK.n264 8.855
R164 CLK.n270 CLK.n269 8.855
R165 CLK.n269 CLK.n268 8.855
R166 CLK.n274 CLK.n273 8.855
R167 CLK.n273 CLK.n272 8.855
R168 CLK.n278 CLK.n277 8.855
R169 CLK.n277 CLK.n276 8.855
R170 CLK.n283 CLK.n282 8.855
R171 CLK.n282 CLK.n281 8.855
R172 CLK.n287 CLK.n286 8.855
R173 CLK.n286 CLK.n285 8.855
R174 CLK.n291 CLK.n290 8.855
R175 CLK.n290 CLK.n289 8.855
R176 CLK.n295 CLK.n294 8.855
R177 CLK.n294 CLK.n293 8.855
R178 CLK.n348 CLK.n347 8.855
R179 CLK.n347 CLK.n346 8.855
R180 CLK.n344 CLK.n343 8.855
R181 CLK.n343 CLK.n342 8.855
R182 CLK.n340 CLK.n339 8.855
R183 CLK.n339 CLK.n338 8.855
R184 CLK.n335 CLK.n334 8.855
R185 CLK.n334 CLK.n333 8.855
R186 CLK.n331 CLK.n330 8.855
R187 CLK.n330 CLK.n329 8.855
R188 CLK.n327 CLK.n326 8.855
R189 CLK.n326 CLK.n325 8.855
R190 CLK.n323 CLK.n322 8.855
R191 CLK.n322 CLK.n321 8.855
R192 CLK.n319 CLK.n318 8.855
R193 CLK.n318 CLK.n317 8.855
R194 CLK.n315 CLK.n314 8.855
R195 CLK.n314 CLK.n313 8.855
R196 CLK.n310 CLK.n309 8.855
R197 CLK.n309 CLK.n308 8.855
R198 CLK.n306 CLK.n305 8.855
R199 CLK.n305 CLK.n304 8.855
R200 CLK.n302 CLK.n301 8.855
R201 CLK.n289 CLK.t33 8.189
R202 CLK.n346 CLK.t10 8.189
R203 CLK.n81 CLK.t13 8.189
R204 CLK.n74 CLK.t29 8.189
R205 CLK.n312 CLK.n297 6.776
R206 CLK.n39 CLK.n26 6.776
R207 CLK.n155 CLK.n142 6.776
R208 CLK.n155 CLK.n141 6.776
R209 CLK.n123 CLK.n9 6.754
R210 CLK.n239 CLK.n3 6.754
R211 CLK.n197 CLK.t1 4.947
R212 CLK.n190 CLK.t24 4.947
R213 CLK.n296 CLK.n0 4.938
R214 CLK.n80 CLK.n25 4.938
R215 CLK.n196 CLK.n139 4.938
R216 CLK.n196 CLK.n140 4.938
R217 CLK.n20 CLK.n19 4.65
R218 CLK.n24 CLK.n23 4.65
R219 CLK.n117 CLK.n116 4.65
R220 CLK.n113 CLK.n112 4.65
R221 CLK.n109 CLK.n108 4.65
R222 CLK.n105 CLK.n104 4.65
R223 CLK.n101 CLK.n100 4.65
R224 CLK.n97 CLK.n96 4.65
R225 CLK.n92 CLK.n91 4.65
R226 CLK.n88 CLK.n87 4.65
R227 CLK.n84 CLK.n83 4.65
R228 CLK.n80 CLK.n79 4.65
R229 CLK.n76 CLK.n73 4.65
R230 CLK.n72 CLK.n71 4.65
R231 CLK.n68 CLK.n67 4.65
R232 CLK.n63 CLK.n62 4.65
R233 CLK.n59 CLK.n58 4.65
R234 CLK.n55 CLK.n54 4.65
R235 CLK.n51 CLK.n50 4.65
R236 CLK.n47 CLK.n46 4.65
R237 CLK.n43 CLK.n42 4.65
R238 CLK.n38 CLK.n37 4.65
R239 CLK.n34 CLK.n33 4.65
R240 CLK.n120 CLK.n12 4.65
R241 CLK.n126 CLK.n7 4.65
R242 CLK.n125 CLK.n124 4.65
R243 CLK.n134 CLK.n133 4.65
R244 CLK.n138 CLK.n137 4.65
R245 CLK.n233 CLK.n232 4.65
R246 CLK.n229 CLK.n228 4.65
R247 CLK.n225 CLK.n224 4.65
R248 CLK.n221 CLK.n220 4.65
R249 CLK.n217 CLK.n216 4.65
R250 CLK.n213 CLK.n212 4.65
R251 CLK.n208 CLK.n207 4.65
R252 CLK.n204 CLK.n203 4.65
R253 CLK.n200 CLK.n199 4.65
R254 CLK.n196 CLK.n195 4.65
R255 CLK.n192 CLK.n189 4.65
R256 CLK.n188 CLK.n187 4.65
R257 CLK.n184 CLK.n183 4.65
R258 CLK.n179 CLK.n178 4.65
R259 CLK.n175 CLK.n174 4.65
R260 CLK.n171 CLK.n170 4.65
R261 CLK.n167 CLK.n166 4.65
R262 CLK.n163 CLK.n162 4.65
R263 CLK.n159 CLK.n158 4.65
R264 CLK.n154 CLK.n153 4.65
R265 CLK.n150 CLK.n149 4.65
R266 CLK.n236 CLK.n6 4.65
R267 CLK.n242 CLK.n1 4.65
R268 CLK.n241 CLK.n240 4.65
R269 CLK.n250 CLK.n249 4.65
R270 CLK.n254 CLK.n253 4.65
R271 CLK.n259 CLK.n258 4.65
R272 CLK.n263 CLK.n262 4.65
R273 CLK.n267 CLK.n266 4.65
R274 CLK.n271 CLK.n270 4.65
R275 CLK.n275 CLK.n274 4.65
R276 CLK.n279 CLK.n278 4.65
R277 CLK.n284 CLK.n283 4.65
R278 CLK.n288 CLK.n287 4.65
R279 CLK.n292 CLK.n291 4.65
R280 CLK.n296 CLK.n295 4.65
R281 CLK.n349 CLK.n348 4.65
R282 CLK.n345 CLK.n344 4.65
R283 CLK.n341 CLK.n340 4.65
R284 CLK.n336 CLK.n335 4.65
R285 CLK.n332 CLK.n331 4.65
R286 CLK.n328 CLK.n327 4.65
R287 CLK.n324 CLK.n323 4.65
R288 CLK.n320 CLK.n319 4.65
R289 CLK.n316 CLK.n315 4.65
R290 CLK.n311 CLK.n310 4.65
R291 CLK.n307 CLK.n306 4.65
R292 CLK.n303 CLK.n302 4.65
R293 CLK.n6 CLK.n5 3.715
R294 CLK.n12 CLK.n11 3.715
R295 CLK.n122 CLK.n121 3.039
R296 CLK.n238 CLK.n237 3.039
R297 CLK.n299 CLK.n298 3.037
R298 CLK.n246 CLK.n245 2.682
R299 CLK.n16 CLK.n15 2.682
R300 CLK.n30 CLK.n29 2.682
R301 CLK.n130 CLK.n129 2.682
R302 CLK.n146 CLK.n145 2.682
R303 CLK.n5 CLK.n4 2.57
R304 CLK.n11 CLK.n10 2.57
R305 CLK.n9 CLK.n8 2.57
R306 CLK.n3 CLK.n2 2.57
R307 CLK.n123 CLK.n122 2.224
R308 CLK.n239 CLK.n238 2.224
R309 CLK.n119 CLK.n118 2.203
R310 CLK.n234 CLK.n126 2.203
R311 CLK.n235 CLK.n234 2.203
R312 CLK.n255 CLK.n242 2.203
R313 CLK.n128 CLK.n127 1.722
R314 CLK.n144 CLK.n143 1.722
R315 CLK.n244 CLK.n243 1.655
R316 CLK.n14 CLK.n13 1.655
R317 CLK.n28 CLK.n27 1.655
R318 CLK.n301 CLK.n300 1.655
R319 CLK.n250 CLK.n246 1.096
R320 CLK.n20 CLK.n16 1.095
R321 CLK.n34 CLK.n30 1.095
R322 CLK.n134 CLK.n130 1.095
R323 CLK.n150 CLK.n146 1.095
R324 CLK.n299 CLK 0.764
R325 CLK.n120 CLK.n119 0.125
R326 CLK.n126 CLK.n125 0.125
R327 CLK.n236 CLK.n235 0.125
R328 CLK.n242 CLK.n241 0.125
R329 CLK.n125 CLK.n123 0.12
R330 CLK.n241 CLK.n239 0.12
R331 CLK.n122 CLK.n120 0.119
R332 CLK.n238 CLK.n236 0.119
R333 CLK.n24 CLK.n20 0.1
R334 CLK.n117 CLK.n113 0.1
R335 CLK.n113 CLK.n109 0.1
R336 CLK.n109 CLK.n105 0.1
R337 CLK.n105 CLK.n101 0.1
R338 CLK.n101 CLK.n97 0.1
R339 CLK.n92 CLK.n88 0.1
R340 CLK.n88 CLK.n84 0.1
R341 CLK.n84 CLK.n80 0.1
R342 CLK.n73 CLK.n72 0.1
R343 CLK.n72 CLK.n68 0.1
R344 CLK.n63 CLK.n59 0.1
R345 CLK.n59 CLK.n55 0.1
R346 CLK.n55 CLK.n51 0.1
R347 CLK.n51 CLK.n47 0.1
R348 CLK.n47 CLK.n43 0.1
R349 CLK.n38 CLK.n34 0.1
R350 CLK.n138 CLK.n134 0.1
R351 CLK.n233 CLK.n229 0.1
R352 CLK.n229 CLK.n225 0.1
R353 CLK.n225 CLK.n221 0.1
R354 CLK.n221 CLK.n217 0.1
R355 CLK.n217 CLK.n213 0.1
R356 CLK.n208 CLK.n204 0.1
R357 CLK.n204 CLK.n200 0.1
R358 CLK.n200 CLK.n196 0.1
R359 CLK.n189 CLK.n188 0.1
R360 CLK.n188 CLK.n184 0.1
R361 CLK.n179 CLK.n175 0.1
R362 CLK.n175 CLK.n171 0.1
R363 CLK.n171 CLK.n167 0.1
R364 CLK.n167 CLK.n163 0.1
R365 CLK.n163 CLK.n159 0.1
R366 CLK.n154 CLK.n150 0.1
R367 CLK.n254 CLK.n250 0.1
R368 CLK.n263 CLK.n259 0.1
R369 CLK.n267 CLK.n263 0.1
R370 CLK.n271 CLK.n267 0.1
R371 CLK.n275 CLK.n271 0.1
R372 CLK.n279 CLK.n275 0.1
R373 CLK.n288 CLK.n284 0.1
R374 CLK.n292 CLK.n288 0.1
R375 CLK.n296 CLK.n292 0.1
R376 CLK.n349 CLK.n345 0.1
R377 CLK.n345 CLK.n341 0.1
R378 CLK.n336 CLK.n332 0.1
R379 CLK.n332 CLK.n328 0.1
R380 CLK.n328 CLK.n324 0.1
R381 CLK.n324 CLK.n320 0.1
R382 CLK.n320 CLK.n316 0.1
R383 CLK.n311 CLK.n307 0.1
R384 CLK.n307 CLK.n303 0.1
R385 CLK.n303 CLK.n299 0.095
R386 CLK.n118 CLK.n117 0.075
R387 CLK.n93 CLK.n92 0.075
R388 CLK.n73 EESPFAL_XOR_v3_0/CLK 0.075
R389 CLK.n68 CLK.n64 0.075
R390 CLK.n43 CLK.n39 0.075
R391 CLK.n234 CLK.n233 0.075
R392 CLK.n209 CLK.n208 0.075
R393 CLK.n189 EESPFAL_XOR_v3_2/CLK 0.075
R394 CLK.n184 CLK.n180 0.075
R395 CLK.n159 CLK.n155 0.075
R396 CLK.n259 CLK.n255 0.075
R397 CLK.n284 CLK.n280 0.075
R398 CLK CLK.n349 0.075
R399 CLK.n341 CLK.n337 0.075
R400 CLK.n316 CLK.n312 0.075
R401 CLK.n118 CLK.n24 0.025
R402 CLK.n97 CLK.n93 0.025
R403 CLK.n80 EESPFAL_XOR_v3_0/CLK 0.025
R404 CLK.n64 CLK.n63 0.025
R405 CLK.n39 CLK.n38 0.025
R406 CLK.n234 CLK.n138 0.025
R407 CLK.n213 CLK.n209 0.025
R408 CLK.n196 EESPFAL_XOR_v3_2/CLK 0.025
R409 CLK.n180 CLK.n179 0.025
R410 CLK.n155 CLK.n154 0.025
R411 CLK.n255 CLK.n254 0.025
R412 CLK.n280 CLK.n279 0.025
R413 CLK CLK.n296 0.025
R414 CLK.n337 CLK.n336 0.025
R415 CLK.n312 CLK.n311 0.025
R416 XOR1_bar.t8 XOR1_bar.t7 819.4
R417 XOR1_bar.n0 XOR1_bar.t6 506.1
R418 XOR1_bar.n0 XOR1_bar.t8 313.3
R419 XOR1_bar.n2 XOR1_bar.t2 273.936
R420 XOR1_bar.n7 XOR1_bar 220.4
R421 XOR1_bar.n5 XOR1_bar.n4 128.334
R422 XOR1_bar.n3 XOR1_bar.n2 105.6
R423 XOR1_bar.n2 XOR1_bar.t1 81.937
R424 XOR1_bar.n3 XOR1_bar.n1 57.937
R425 XOR1_bar.n6 XOR1_bar.n5 57.6
R426 XOR1_bar.n5 XOR1_bar.n3 41.6
R427 XOR1_bar.n4 XOR1_bar.t4 39.4
R428 XOR1_bar.n4 XOR1_bar.t5 39.4
R429 XOR1_bar.n1 XOR1_bar.t3 24
R430 XOR1_bar.n1 XOR1_bar.t0 24
R431 XOR1_bar.n6 XOR1_bar.n0 8.764
R432 XOR1_bar.n7 XOR1_bar.n6 4.65
R433 XOR1_bar XOR1_bar.n7 0.031
R434 XOR2.t7 XOR2.t6 819.4
R435 XOR2.n5 XOR2.t7 514.133
R436 XOR2.n5 XOR2.t8 305.266
R437 XOR2.n3 XOR2.n2 192
R438 XOR2.n4 XOR2.n0 166.734
R439 XOR2.n4 XOR2.n3 105.6
R440 XOR2.n3 XOR2.t1 97.937
R441 XOR2.n2 XOR2.t5 97.937
R442 XOR2.n6 XOR2.n5 76
R443 XOR2.n4 XOR2.n1 73.937
R444 XOR2.n6 XOR2.n4 57.6
R445 XOR2.n0 XOR2.t0 39.4
R446 XOR2.n0 XOR2.t3 39.4
R447 XOR2.n1 XOR2.t4 24
R448 XOR2.n1 XOR2.t2 24
R449 XOR2.n2 XOR2 10.56
R450 XOR2 XOR2.n6 3.2
R451 XOR2_bar.t7 XOR2_bar.t8 819.4
R452 XOR2_bar.n0 XOR2_bar.t6 506.1
R453 XOR2_bar.n0 XOR2_bar.t7 313.3
R454 XOR2_bar.n3 XOR2_bar.t0 273.936
R455 XOR2_bar.n7 XOR2_bar 221.04
R456 XOR2_bar.n5 XOR2_bar.n1 128.334
R457 XOR2_bar.n4 XOR2_bar.n3 105.6
R458 XOR2_bar.n3 XOR2_bar.t1 81.937
R459 XOR2_bar.n4 XOR2_bar.n2 57.937
R460 XOR2_bar.n6 XOR2_bar.n5 57.6
R461 XOR2_bar.n5 XOR2_bar.n4 41.6
R462 XOR2_bar.n1 XOR2_bar.t4 39.4
R463 XOR2_bar.n1 XOR2_bar.t5 39.4
R464 XOR2_bar.n2 XOR2_bar.t3 24
R465 XOR2_bar.n2 XOR2_bar.t2 24
R466 XOR2_bar.n6 XOR2_bar.n0 8.764
R467 XOR2_bar.n7 XOR2_bar.n6 4.65
R468 XOR2_bar XOR2_bar.n7 0.031
R469 k2_bar.n0 k2_bar.t0 810.772
R470 k2_bar.n0 k2_bar.t1 694.566
R471 k2_bar k2_bar.n0 25.6
R472 GND.n93 GND.n92 341.085
R473 GND.n101 GND.n85 341.085
R474 GND.n103 GND.n102 341.085
R475 GND.n112 GND.n79 341.085
R476 GND.n113 GND.n112 341.085
R477 GND.n114 GND.n113 341.085
R478 GND.n125 GND.n73 341.085
R479 GND.n128 GND.n127 341.085
R480 GND.n138 GND.n137 341.085
R481 GND.n140 GND.n138 341.085
R482 GND.n140 GND.n139 341.085
R483 GND.n149 GND.n148 341.085
R484 GND.n151 GND.n150 341.085
R485 GND.n160 GND.n159 341.085
R486 GND.t19 GND.n79 319.767
R487 GND.n126 GND.t24 319.767
R488 GND.t22 GND.n126 319.767
R489 GND.n139 GND.t32 319.767
R490 GND.n102 GND.t0 277.131
R491 GND.t7 GND.n73 277.131
R492 GND.n127 GND.t9 277.131
R493 GND.t18 GND.n149 277.131
R494 GND.t4 GND.n85 234.496
R495 GND.n150 GND.t3 234.496
R496 GND.n92 GND.t33 191.86
R497 GND.t27 GND.n160 191.86
R498 GND.t33 GND.n91 158.378
R499 GND.n161 GND.t27 158.378
R500 GND.n5 GND.t29 158.378
R501 GND.n163 GND.t34 158.378
R502 GND.n91 GND.n90 157.6
R503 GND.n94 GND.n90 157.6
R504 GND.n94 GND.n86 157.6
R505 GND.n100 GND.n86 157.6
R506 GND.n100 GND.n84 157.6
R507 GND.n104 GND.n84 157.6
R508 GND.n104 GND.n80 157.6
R509 GND.n111 GND.n80 157.6
R510 GND.n111 GND.n78 157.6
R511 GND.n115 GND.n78 157.6
R512 GND.n115 GND.n74 157.6
R513 GND.n124 GND.n74 157.6
R514 GND.n124 GND.n72 157.6
R515 GND.n129 GND.n72 157.6
R516 GND.n129 GND.n69 157.6
R517 GND.n136 GND.n69 157.6
R518 GND.n136 GND.n68 157.6
R519 GND.n141 GND.n68 157.6
R520 GND.n141 GND.n64 157.6
R521 GND.n147 GND.n64 157.6
R522 GND.n147 GND.n63 157.6
R523 GND.n152 GND.n63 157.6
R524 GND.n152 GND.n58 157.6
R525 GND.n158 GND.n58 157.6
R526 GND.n158 GND.n57 157.6
R527 GND.n161 GND.n57 157.6
R528 GND.n93 GND.t4 106.589
R529 GND.n159 GND.t3 106.589
R530 GND.n7 GND.t17 106.589
R531 GND.n169 GND.t16 106.589
R532 GND.t0 GND.n101 63.953
R533 GND.n114 GND.t7 63.953
R534 GND.n137 GND.t9 63.953
R535 GND.n151 GND.t18 63.953
R536 GND.n15 GND.t26 63.953
R537 GND.n40 GND.t11 63.953
R538 GND.n202 GND.t1 63.953
R539 GND.n177 GND.t31 63.953
R540 GND.n164 GND 35.195
R541 GND GND.n162 31.551
R542 GND.n76 GND.t20 29.103
R543 GND.n133 GND.t21 29.103
R544 GND.n39 GND.t13 29.103
R545 GND.n201 GND.t30 29.103
R546 GND.n76 GND.t8 29.102
R547 GND.n133 GND.t10 29.102
R548 GND.n39 GND.t12 29.102
R549 GND.n201 GND.t2 29.102
R550 GND.n120 GND.t38 24
R551 GND.n120 GND.t39 24
R552 GND.n119 GND.t25 24
R553 GND.n119 GND.t23 24
R554 GND.n1 GND.t15 24
R555 GND.n1 GND.t6 24
R556 GND.n0 GND.t36 24
R557 GND.n0 GND.t37 24
R558 GND.n103 GND.t19 21.317
R559 GND.t24 GND.n125 21.317
R560 GND.n128 GND.t22 21.317
R561 GND.n148 GND.t32 21.317
R562 GND.n23 GND.t35 21.317
R563 GND.n48 GND.t14 21.317
R564 GND.n210 GND.t5 21.317
R565 GND.n185 GND.t28 21.317
R566 GND.n95 GND.n89 12.8
R567 GND.n95 GND.n87 12.8
R568 GND.n99 GND.n87 12.8
R569 GND.n99 GND.n83 12.8
R570 GND.n105 GND.n83 12.8
R571 GND.n105 GND.n81 12.8
R572 GND.n110 GND.n81 12.8
R573 GND.n110 GND.n77 12.8
R574 GND.n116 GND.n77 12.8
R575 GND.n116 GND.n75 12.8
R576 GND.n123 GND.n75 12.8
R577 GND.n123 GND.n71 12.8
R578 GND.n130 GND.n71 12.8
R579 GND.n130 GND.n70 12.8
R580 GND.n135 GND.n70 12.8
R581 GND.n135 GND.n67 12.8
R582 GND.n142 GND.n67 12.8
R583 GND.n142 GND.n65 12.8
R584 GND.n146 GND.n65 12.8
R585 GND.n146 GND.n62 12.8
R586 GND.n153 GND.n62 12.8
R587 GND.n153 GND.n59 12.8
R588 GND.n157 GND.n59 12.8
R589 GND.n157 GND.n60 12.8
R590 GND.n6 GND.n5 11.894
R591 GND.n91 GND.n88 11.894
R592 GND.n90 GND.n89 9.154
R593 GND.n92 GND.n90 9.154
R594 GND.n95 GND.n94 9.154
R595 GND.n94 GND.n93 9.154
R596 GND.n87 GND.n86 9.154
R597 GND.n86 GND.n85 9.154
R598 GND.n100 GND.n99 9.154
R599 GND.n101 GND.n100 9.154
R600 GND.n84 GND.n83 9.154
R601 GND.n102 GND.n84 9.154
R602 GND.n105 GND.n104 9.154
R603 GND.n104 GND.n103 9.154
R604 GND.n81 GND.n80 9.154
R605 GND.n80 GND.n79 9.154
R606 GND.n111 GND.n110 9.154
R607 GND.n112 GND.n111 9.154
R608 GND.n78 GND.n77 9.154
R609 GND.n113 GND.n78 9.154
R610 GND.n116 GND.n115 9.154
R611 GND.n115 GND.n114 9.154
R612 GND.n75 GND.n74 9.154
R613 GND.n74 GND.n73 9.154
R614 GND.n124 GND.n123 9.154
R615 GND.n125 GND.n124 9.154
R616 GND.n72 GND.n71 9.154
R617 GND.n126 GND.n72 9.154
R618 GND.n130 GND.n129 9.154
R619 GND.n129 GND.n128 9.154
R620 GND.n70 GND.n69 9.154
R621 GND.n127 GND.n69 9.154
R622 GND.n136 GND.n135 9.154
R623 GND.n137 GND.n136 9.154
R624 GND.n68 GND.n67 9.154
R625 GND.n138 GND.n68 9.154
R626 GND.n142 GND.n141 9.154
R627 GND.n141 GND.n140 9.154
R628 GND.n65 GND.n64 9.154
R629 GND.n139 GND.n64 9.154
R630 GND.n147 GND.n146 9.154
R631 GND.n148 GND.n147 9.154
R632 GND.n63 GND.n62 9.154
R633 GND.n149 GND.n63 9.154
R634 GND.n153 GND.n152 9.154
R635 GND.n152 GND.n151 9.154
R636 GND.n59 GND.n58 9.154
R637 GND.n150 GND.n58 9.154
R638 GND.n158 GND.n157 9.154
R639 GND.n159 GND.n158 9.154
R640 GND.n60 GND.n57 9.154
R641 GND.n160 GND.n57 9.154
R642 GND.n162 GND.n161 9.154
R643 GND.n164 GND.n163 9.154
R644 GND.n4 GND.n3 9.154
R645 GND.n3 GND.n2 9.154
R646 GND.n9 GND.n8 9.154
R647 GND.n8 GND.n7 9.154
R648 GND.n13 GND.n12 9.154
R649 GND.n12 GND.n11 9.154
R650 GND.n17 GND.n16 9.154
R651 GND.n16 GND.n15 9.154
R652 GND.n21 GND.n20 9.154
R653 GND.n20 GND.n19 9.154
R654 GND.n25 GND.n24 9.154
R655 GND.n24 GND.n23 9.154
R656 GND.n29 GND.n28 9.154
R657 GND.n28 GND.n27 9.154
R658 GND.n33 GND.n32 9.154
R659 GND.n32 GND.n31 9.154
R660 GND.n37 GND.n36 9.154
R661 GND.n36 GND.n35 9.154
R662 GND.n42 GND.n41 9.154
R663 GND.n41 GND.n40 9.154
R664 GND.n46 GND.n45 9.154
R665 GND.n45 GND.n44 9.154
R666 GND.n50 GND.n49 9.154
R667 GND.n49 GND.n48 9.154
R668 GND.n54 GND.n53 9.154
R669 GND.n53 GND.n52 9.154
R670 GND.n212 GND.n211 9.154
R671 GND.n211 GND.n210 9.154
R672 GND.n208 GND.n207 9.154
R673 GND.n207 GND.n206 9.154
R674 GND.n204 GND.n203 9.154
R675 GND.n203 GND.n202 9.154
R676 GND.n199 GND.n198 9.154
R677 GND.n198 GND.n197 9.154
R678 GND.n195 GND.n194 9.154
R679 GND.n194 GND.n193 9.154
R680 GND.n191 GND.n190 9.154
R681 GND.n190 GND.n189 9.154
R682 GND.n187 GND.n186 9.154
R683 GND.n186 GND.n185 9.154
R684 GND.n183 GND.n182 9.154
R685 GND.n182 GND.n181 9.154
R686 GND.n179 GND.n178 9.154
R687 GND.n178 GND.n177 9.154
R688 GND.n175 GND.n174 9.154
R689 GND.n174 GND.n173 9.154
R690 GND.n171 GND.n170 9.154
R691 GND.n170 GND.n169 9.154
R692 GND.n167 GND.n166 9.154
R693 GND.n166 GND.n165 9.154
R694 GND.n121 GND.n120 5.103
R695 GND.n121 GND.n119 5.103
R696 GND.n55 GND.n1 5.103
R697 GND.n55 GND.n0 5.103
R698 GND.n96 GND.n95 4.65
R699 GND.n97 GND.n87 4.65
R700 GND.n99 GND.n98 4.65
R701 GND.n83 GND.n82 4.65
R702 GND.n106 GND.n105 4.65
R703 GND.n107 GND.n81 4.65
R704 GND.n110 GND.n109 4.65
R705 GND.n108 GND.n77 4.65
R706 GND.n117 GND.n116 4.65
R707 GND.n118 GND.n75 4.65
R708 GND.n123 GND.n122 4.65
R709 GND.n121 GND.n71 4.65
R710 GND.n131 GND.n130 4.65
R711 GND.n132 GND.n70 4.65
R712 GND.n135 GND.n134 4.65
R713 GND.n67 GND.n66 4.65
R714 GND.n143 GND.n142 4.65
R715 GND.n144 GND.n65 4.65
R716 GND.n146 GND.n145 4.65
R717 GND.n62 GND.n61 4.65
R718 GND.n154 GND.n153 4.65
R719 GND.n155 GND.n59 4.65
R720 GND.n157 GND.n156 4.65
R721 GND.n10 GND.n9 4.65
R722 GND.n14 GND.n13 4.65
R723 GND.n18 GND.n17 4.65
R724 GND.n22 GND.n21 4.65
R725 GND.n26 GND.n25 4.65
R726 GND.n30 GND.n29 4.65
R727 GND.n34 GND.n33 4.65
R728 GND.n38 GND.n37 4.65
R729 GND.n43 GND.n42 4.65
R730 GND.n47 GND.n46 4.65
R731 GND.n51 GND.n50 4.65
R732 GND.n55 GND.n54 4.65
R733 GND.n213 GND.n212 4.65
R734 GND.n209 GND.n208 4.65
R735 GND.n205 GND.n204 4.65
R736 GND.n200 GND.n199 4.65
R737 GND.n196 GND.n195 4.65
R738 GND.n192 GND.n191 4.65
R739 GND.n188 GND.n187 4.65
R740 GND.n184 GND.n183 4.65
R741 GND.n180 GND.n179 4.65
R742 GND.n176 GND.n175 4.65
R743 GND.n172 GND.n171 4.65
R744 GND.n162 GND.n56 2.739
R745 GND.n168 GND.n164 2.739
R746 GND.n6 GND.n4 2.682
R747 GND.n89 GND.n88 2.682
R748 GND.n60 GND.n56 2.682
R749 GND.n168 GND.n167 2.682
R750 GND.n10 GND.n6 1.096
R751 GND.n96 GND.n88 1.095
R752 GND.n156 GND.n56 1.095
R753 GND.n172 GND.n168 1.095
R754 GND.n97 GND.n96 0.1
R755 GND.n98 GND.n97 0.1
R756 GND.n98 GND.n82 0.1
R757 GND.n106 GND.n82 0.1
R758 GND.n107 GND.n106 0.1
R759 GND.n109 GND.n107 0.1
R760 GND.n109 GND.n108 0.1
R761 GND.n118 GND.n117 0.1
R762 GND.n122 GND.n118 0.1
R763 GND.n122 GND.n121 0.1
R764 GND.n132 GND.n131 0.1
R765 GND.n134 GND.n132 0.1
R766 GND.n143 GND.n66 0.1
R767 GND.n144 GND.n143 0.1
R768 GND.n145 GND.n144 0.1
R769 GND.n145 GND.n61 0.1
R770 GND.n154 GND.n61 0.1
R771 GND.n155 GND.n154 0.1
R772 GND.n156 GND.n155 0.1
R773 GND.n14 GND.n10 0.1
R774 GND.n18 GND.n14 0.1
R775 GND.n22 GND.n18 0.1
R776 GND.n26 GND.n22 0.1
R777 GND.n30 GND.n26 0.1
R778 GND.n34 GND.n30 0.1
R779 GND.n38 GND.n34 0.1
R780 GND.n47 GND.n43 0.1
R781 GND.n51 GND.n47 0.1
R782 GND.n55 GND.n51 0.1
R783 GND.n213 GND.n209 0.1
R784 GND.n209 GND.n205 0.1
R785 GND.n200 GND.n196 0.1
R786 GND.n196 GND.n192 0.1
R787 GND.n192 GND.n188 0.1
R788 GND.n188 GND.n184 0.1
R789 GND.n184 GND.n180 0.1
R790 GND.n180 GND.n176 0.1
R791 GND.n176 GND.n172 0.1
R792 GND.n117 GND.n76 0.075
R793 GND.n131 GND 0.075
R794 GND.n134 GND.n133 0.075
R795 GND.n43 GND.n39 0.075
R796 EESPFAL_XOR_v3_0/GND GND.n213 0.075
R797 GND.n205 GND.n201 0.075
R798 GND.n108 GND.n76 0.025
R799 GND.n121 GND 0.025
R800 GND.n133 GND.n66 0.025
R801 GND.n39 GND.n38 0.025
R802 EESPFAL_XOR_v3_0/GND GND.n55 0.025
R803 GND.n201 GND.n200 0.025
R804 XOR0.t6 XOR0.t7 819.4
R805 XOR0.n5 XOR0.t6 514.133
R806 XOR0.n5 XOR0.t8 305.266
R807 XOR0.n3 XOR0.n2 192
R808 XOR0.n4 XOR0.n0 166.734
R809 XOR0.n4 XOR0.n3 105.6
R810 XOR0.n3 XOR0.t1 97.937
R811 XOR0.n2 XOR0.t5 97.937
R812 XOR0.n6 XOR0.n5 76
R813 XOR0.n4 XOR0.n1 73.937
R814 XOR0.n6 XOR0.n4 57.6
R815 XOR0.n0 XOR0.t0 39.4
R816 XOR0.n0 XOR0.t4 39.4
R817 XOR0.n1 XOR0.t2 24
R818 XOR0.n1 XOR0.t3 24
R819 XOR0.n2 XOR0 9.6
R820 XOR0 XOR0.n6 3.2
R821 XOR0_bar.t6 XOR0_bar.t7 819.4
R822 XOR0_bar.n0 XOR0_bar.t8 506.1
R823 XOR0_bar.n0 XOR0_bar.t6 313.3
R824 XOR0_bar.n3 XOR0_bar.t4 273.936
R825 XOR0_bar.n7 XOR0_bar 220.08
R826 XOR0_bar.n5 XOR0_bar.n1 128.334
R827 XOR0_bar.n4 XOR0_bar.n3 105.6
R828 XOR0_bar.n3 XOR0_bar.t5 81.937
R829 XOR0_bar.n4 XOR0_bar.n2 57.937
R830 XOR0_bar.n6 XOR0_bar.n5 57.6
R831 XOR0_bar.n5 XOR0_bar.n4 41.6
R832 XOR0_bar.n1 XOR0_bar.t2 39.4
R833 XOR0_bar.n1 XOR0_bar.t1 39.4
R834 XOR0_bar.n2 XOR0_bar.t0 24
R835 XOR0_bar.n2 XOR0_bar.t3 24
R836 XOR0_bar.n6 XOR0_bar.n0 8.764
R837 XOR0_bar.n7 XOR0_bar.n6 4.65
R838 XOR0_bar XOR0_bar.n7 0.031
R839 Dis.n3 Dis.t2 504.5
R840 Dis.n2 Dis.t3 504.5
R841 Dis.n1 Dis.t4 504.5
R842 Dis.n0 Dis.t7 504.5
R843 Dis.n3 Dis.t0 389.3
R844 Dis.n2 Dis.t6 389.3
R845 Dis.n1 Dis.t5 389.3
R846 Dis.n0 Dis.t1 389.3
R847 EESPFAL_XOR_v3_0/Dis Dis.n6 220.082
R848 Dis.n4 Dis 219.457
R849 Dis.n5 EESPFAL_XOR_v3_2/Dis 219.456
R850 Dis.n6 EESPFAL_XOR_v3_1/Dis 219.456
R851 Dis.n6 Dis.n5 6.502
R852 Dis Dis.n3 3.2
R853 EESPFAL_XOR_v3_2/Dis Dis.n2 3.2
R854 EESPFAL_XOR_v3_1/Dis Dis.n1 3.2
R855 EESPFAL_XOR_v3_0/Dis Dis.n0 3.2
R856 Dis.n4 Dis 3.199
R857 Dis.n5 Dis.n4 0.625
R858 x2.n0 x2.t1 1176.57
R859 x2.n0 x2.t0 1149.49
R860 x2 x2.n0 128
R861 XOR3_bar.t6 XOR3_bar.t7 819.4
R862 XOR3_bar.n0 XOR3_bar.t8 506.1
R863 XOR3_bar.n0 XOR3_bar.t6 313.3
R864 XOR3_bar.n2 XOR3_bar.t5 273.936
R865 XOR3_bar.n7 XOR3_bar 221.36
R866 XOR3_bar.n5 XOR3_bar.n4 128.334
R867 XOR3_bar.n3 XOR3_bar.n2 105.6
R868 XOR3_bar.n2 XOR3_bar.t4 81.937
R869 XOR3_bar.n3 XOR3_bar.n1 57.937
R870 XOR3_bar.n6 XOR3_bar.n5 57.6
R871 XOR3_bar.n5 XOR3_bar.n3 41.6
R872 XOR3_bar.n4 XOR3_bar.t2 39.4
R873 XOR3_bar.n4 XOR3_bar.t1 39.4
R874 XOR3_bar.n1 XOR3_bar.t0 24
R875 XOR3_bar.n1 XOR3_bar.t3 24
R876 XOR3_bar.n6 XOR3_bar.n0 8.764
R877 XOR3_bar.n7 XOR3_bar.n6 4.65
R878 XOR3_bar XOR3_bar.n7 0.031
R879 x0.n0 x0.t0 1176.57
R880 x0.n0 x0.t1 1149.49
R881 x0 x0.n0 128
R882 x3.n0 x3.t0 1176.57
R883 x3.n0 x3.t1 1149.49
R884 x3 x3.n0 128
R885 XOR3.t8 XOR3.t7 819.4
R886 XOR3.n5 XOR3.t8 514.133
R887 XOR3.n5 XOR3.t6 305.266
R888 XOR3.n3 XOR3.n2 192
R889 XOR3.n4 XOR3.n1 166.734
R890 XOR3.n4 XOR3.n3 105.6
R891 XOR3.n2 XOR3.t4 97.937
R892 XOR3.n3 XOR3.t5 97.937
R893 XOR3.n6 XOR3.n5 76
R894 XOR3.n4 XOR3.n0 73.937
R895 XOR3.n6 XOR3.n4 57.6
R896 XOR3.n1 XOR3.t1 39.4
R897 XOR3.n1 XOR3.t2 39.4
R898 XOR3.n0 XOR3.t3 24
R899 XOR3.n0 XOR3.t0 24
R900 XOR3.n2 XOR3 10.88
R901 XOR3 XOR3.n6 3.2
R902 k0_bar.n0 k0_bar.t1 810.772
R903 k0_bar.n0 k0_bar.t0 694.566
R904 k0_bar k0_bar.n0 25.6
R905 x3_bar.n0 x3_bar.t1 1072.24
R906 x3_bar.n0 x3_bar.t0 1015.9
R907 x3_bar x3_bar.n0 86.4
R908 x1_bar.n0 x1_bar.t0 1072.24
R909 x1_bar.n0 x1_bar.t1 1015.9
R910 x1_bar x1_bar.n0 86.4
R911 k1.n0 k1.t0 800.452
R912 k1.n0 k1.t1 787.997
R913 k1 k1.n0 169.6
R914 x1.n0 x1.t0 1176.57
R915 x1.n0 x1.t1 1149.49
R916 x1 x1.n0 128
R917 x0_bar.n0 x0_bar.t0 1072.24
R918 x0_bar.n0 x0_bar.t1 1015.9
R919 x0_bar x0_bar.n0 86.4
R920 k3.n0 k3.t0 800.452
R921 k3.n0 k3.t1 787.997
R922 k3 k3.n0 169.6
R923 k1_bar.n0 k1_bar.t1 810.772
R924 k1_bar.n0 k1_bar.t0 694.566
R925 k1_bar k1_bar.n0 25.6
R926 k3_bar.n0 k3_bar.t0 810.772
R927 k3_bar.n0 k3_bar.t1 694.566
R928 k3_bar k3_bar.n0 25.6
R929 x2_bar.n0 x2_bar.t1 1072.24
R930 x2_bar.n0 x2_bar.t0 1015.9
R931 x2_bar x2_bar.n0 86.4
R932 k0.n0 k0.t1 800.452
R933 k0.n0 k0.t0 787.997
R934 k0 k0.n0 169.6
R935 k2.n0 k2.t0 800.452
R936 k2.n0 k2.t1 787.997
R937 k2 k2.n0 169.6
C0 k1 x2_bar 0.01fF
C1 k2 XOR1 0.03fF
C2 a_720_n1950# XOR3_bar 0.00fF
C3 Dis XOR3_bar 0.26fF
C4 x1 XOR3 0.00fF
C5 CLK x3 1.11fF
C6 XOR2 a_420_n2630# 0.00fF
C7 k1_bar a_n840_410# 0.00fF
C8 CLK k0 0.37fF
C9 x0 x0_bar 1.56fF
C10 CLK a_720_410# 0.02fF
C11 x2 a_n840_410# 0.00fF
C12 a_n840_n2630# x3_bar 0.00fF
C13 CLK a_n840_n1950# 0.01fF
C14 XOR2_bar x2_bar 0.06fF
C15 k3 XOR3 0.07fF
C16 x1_bar XOR3_bar 0.00fF
C17 k2 XOR3 0.01fF
C18 k1 k0 0.01fF
C19 CLK XOR1 0.73fF
C20 k1 a_720_410# 0.00fF
C21 XOR1_bar a_n840_410# 0.00fF
C22 k1 a_n840_n1950# 0.00fF
C23 k3_bar a_n840_n2630# 0.00fF
C24 k1 XOR1 0.08fF
C25 XOR2_bar x3 0.00fF
C26 CLK a_n1140_410# 0.02fF
C27 XOR0 k0_bar 0.07fF
C28 a_n1140_n1950# x2_bar 0.00fF
C29 XOR2 a_720_n270# 0.00fF
C30 k3 a_720_n2630# 0.00fF
C31 Dis a_n840_410# 0.01fF
C32 k2 a_720_n2630# 0.00fF
C33 x0_bar x2_bar 0.00fF
C34 k1 a_n1140_410# 0.00fF
C35 CLK XOR3 0.68fF
C36 a_n840_n1950# XOR2_bar 0.01fF
C37 XOR1 XOR2_bar 0.03fF
C38 a_n1140_n1950# x3 0.00fF
C39 x0 a_420_410# 0.00fF
C40 x1_bar a_n840_410# 0.00fF
C41 a_420_n2630# XOR3_bar 0.00fF
C42 x0 a_n840_n270# 0.00fF
C43 k3_bar x3_bar 0.09fF
C44 x0 a_420_n270# 0.00fF
C45 CLK a_720_n2630# 0.02fF
C46 x0_bar k0 1.55fF
C47 XOR0 XOR2 0.00fF
C48 x0_bar a_720_410# 0.00fF
C49 XOR2_bar XOR3 0.01fF
C50 x0_bar XOR1 0.00fF
C51 x2_bar a_420_410# 0.00fF
C52 x3_bar a_n1140_n2630# 0.00fF
C53 a_n840_n270# x2_bar 0.00fF
C54 x0_bar a_n1140_410# 0.00fF
C55 k2_bar x2_bar 0.10fF
C56 a_420_n270# x2_bar 0.00fF
C57 XOR2_bar a_720_n2630# 0.00fF
C58 x0 k1_bar 0.00fF
C59 k3_bar a_n1140_n2630# 0.00fF
C60 x0 x2 0.00fF
C61 k0 a_420_410# 0.00fF
C62 k2_bar x3 0.00fF
C63 k3 x1 0.00fF
C64 x1 k2 0.01fF
C65 x0 XOR1_bar 0.00fF
C66 k0 a_n840_n270# 0.00fF
C67 XOR0_bar k0_bar 0.30fF
C68 XOR1 a_420_410# 0.00fF
C69 a_420_n270# k0 0.00fF
C70 k2_bar a_n840_n1950# 0.00fF
C71 k3 k2 0.01fF
C72 a_n840_n270# XOR1 0.00fF
C73 x2_bar k1_bar 0.01fF
C74 x0 Dis 0.03fF
C75 k2_bar XOR1 0.00fF
C76 x2_bar x2 1.56fF
C77 a_420_n270# XOR1 0.01fF
C78 CLK x1 1.03fF
C79 XOR1_bar x2_bar 0.03fF
C80 x0 x1_bar 0.00fF
C81 a_420_n1950# x3_bar 0.00fF
C82 x2 x3 0.01fF
C83 x1 k1 0.15fF
C84 XOR2 x3_bar 0.00fF
C85 k2_bar XOR3 0.02fF
C86 k3 CLK 0.37fF
C87 a_720_n1950# x2_bar 0.00fF
C88 k0 k1_bar 0.00fF
C89 XOR0_bar XOR2 0.00fF
C90 CLK k2 0.54fF
C91 k0 x2 0.00fF
C92 Dis x2_bar 0.03fF
C93 a_n840_n1950# k1_bar 0.00fF
C94 XOR0 a_n840_410# 0.00fF
C95 k3_bar a_420_n1950# 0.00fF
C96 a_n840_n1950# x2 0.00fF
C97 k3_bar XOR2 0.02fF
C98 a_n840_n2630# XOR3_bar 0.01fF
C99 XOR1 k1_bar 0.07fF
C100 k1 k2 0.04fF
C101 XOR1 x2 0.01fF
C102 k0 XOR1_bar 0.01fF
C103 x1 XOR2_bar 0.02fF
C104 x1_bar x2_bar 0.04fF
C105 XOR0_bar a_n1140_n270# 0.00fF
C106 XOR1_bar a_720_410# 0.00fF
C107 a_n840_n1950# XOR1_bar 0.00fF
C108 Dis x3 0.01fF
C109 a_n1140_410# k1_bar 0.00fF
C110 XOR1_bar XOR1 0.78fF
C111 a_n1140_410# x2 0.00fF
C112 k0 Dis 0.04fF
C113 k3 XOR2_bar 0.01fF
C114 k2 XOR2_bar 0.10fF
C115 Dis a_n840_n1950# 0.01fF
C116 a_n1140_n1950# x1 0.00fF
C117 x1_bar x3 0.00fF
C118 a_720_n1950# XOR1 0.00fF
C119 a_n1140_410# XOR1_bar 0.00fF
C120 XOR3 x2 0.00fF
C121 CLK k1 0.54fF
C122 Dis XOR1 0.11fF
C123 x1 x0_bar 0.00fF
C124 x1_bar k0 0.00fF
C125 x3_bar XOR3_bar 0.05fF
C126 x1_bar a_720_410# 0.00fF
C127 x1_bar a_n840_n1950# 0.00fF
C128 k3 a_n1140_n1950# 0.00fF
C129 XOR1_bar XOR3 0.00fF
C130 Dis a_n1140_410# 0.02fF
C131 a_n1140_n1950# k2 0.00fF
C132 x1_bar XOR1 0.03fF
C133 CLK XOR2_bar 1.06fF
C134 a_420_n2630# x2_bar 0.00fF
C135 a_720_n1950# XOR3 0.00fF
C136 k3_bar XOR3_bar 0.30fF
C137 Dis XOR3 0.09fF
C138 x1_bar a_n1140_410# 0.00fF
C139 k1 XOR2_bar 0.03fF
C140 k0_bar a_n1140_n270# 0.00fF
C141 a_420_n2630# x3 0.00fF
C142 x1_bar XOR3 0.00fF
C143 CLK a_n1140_n1950# 0.01fF
C144 a_n1140_n2630# XOR3_bar 0.01fF
C145 x1 a_420_410# 0.00fF
C146 CLK x0_bar 0.49fF
C147 a_n1140_n1950# k1 0.00fF
C148 x1 a_n840_n270# 0.00fF
C149 a_720_n270# x2_bar 0.00fF
C150 a_420_n1950# XOR2 0.01fF
C151 XOR0_bar a_n840_410# 0.01fF
C152 x1 k2_bar 0.01fF
C153 a_420_n270# x1 0.00fF
C154 k1 x0_bar 0.00fF
C155 x0 XOR0 0.03fF
C156 x1_bar a_720_n2630# 0.00fF
C157 k3 k2_bar 0.00fF
C158 k2 a_n840_n270# 0.00fF
C159 k2_bar k2 1.30fF
C160 a_n1140_n1950# XOR2_bar 0.01fF
C161 a_420_n270# k2 0.00fF
C162 k0 a_720_n270# 0.00fF
C163 a_420_n2630# XOR3 0.01fF
C164 CLK a_420_410# 0.02fF
C165 XOR0 x2_bar 0.00fF
C166 XOR1 a_720_n270# 0.01fF
C167 x1 k1_bar 0.06fF
C168 x1 x2 0.29fF
C169 CLK a_n840_n270# 0.01fF
C170 CLK k2_bar 0.25fF
C171 k1 a_420_410# 0.00fF
C172 a_420_n270# CLK 0.02fF
C173 a_420_n1950# XOR3_bar 0.00fF
C174 k1 a_n840_n270# 0.00fF
C175 x1 XOR1_bar 0.05fF
C176 k2 k1_bar 0.01fF
C177 k2_bar k1 0.01fF
C178 XOR2 XOR3_bar 0.01fF
C179 k3 x2 0.00fF
C180 k0_bar a_n840_410# 0.00fF
C181 a_420_n270# k1 0.00fF
C182 k2 x2 0.15fF
C183 XOR0 k0 0.07fF
C184 XOR0 a_720_410# 0.01fF
C185 x1 Dis 0.04fF
C186 k2 XOR1_bar 0.03fF
C187 XOR0 XOR1 0.02fF
C188 a_n840_n270# XOR2_bar 0.00fF
C189 k2_bar XOR2_bar 0.30fF
C190 a_n840_n2630# x2_bar 0.00fF
C191 k3 a_720_n1950# 0.00fF
C192 a_420_n270# XOR2_bar 0.00fF
C193 a_720_n1950# k2 0.00fF
C194 CLK k1_bar 0.25fF
C195 k3 Dis 0.02fF
C196 x1_bar x1 1.56fF
C197 XOR0 a_n1140_410# 0.00fF
C198 Dis k2 0.05fF
C199 CLK x2 1.03fF
C200 x0 XOR0_bar 0.05fF
C201 k1 k1_bar 1.30fF
C202 x0_bar a_420_410# 0.00fF
C203 a_n840_n2630# x3 0.00fF
C204 k1 x2 0.01fF
C205 CLK XOR1_bar 1.06fF
C206 k3 x1_bar 0.00fF
C207 a_n1140_n1950# k2_bar 0.00fF
C208 x1_bar k2 0.01fF
C209 x0_bar a_n840_n270# 0.00fF
C210 a_420_n270# x0_bar 0.00fF
C211 k1 XOR1_bar 0.10fF
C212 CLK a_720_n1950# 0.02fF
C213 CLK Dis 1.17fF
C214 XOR2_bar k1_bar 0.01fF
C215 x2_bar x3_bar 0.01fF
C216 XOR2_bar x2 0.05fF
C217 a_720_n1950# k1 0.00fF
C218 XOR0_bar x2_bar 0.00fF
C219 k1 Dis 0.05fF
C220 x1 a_420_n2630# 0.00fF
C221 CLK x1_bar 0.57fF
C222 XOR1_bar XOR2_bar 0.05fF
C223 k3_bar x2_bar 0.00fF
C224 x3_bar x3 1.56fF
C225 a_n1140_n1950# k1_bar 0.00fF
C226 a_n1140_n1950# x2 0.00fF
C227 x1_bar k1 1.55fF
C228 a_720_n1950# XOR2_bar 0.00fF
C229 a_n840_n2630# XOR3 0.00fF
C230 k3 a_420_n2630# 0.00fF
C231 x0_bar k1_bar 0.00fF
C232 k2 a_420_n2630# 0.00fF
C233 Dis XOR2_bar 0.32fF
C234 x0_bar x2 0.00fF
C235 a_n840_n1950# x3_bar 0.00fF
C236 XOR0_bar k0 0.09fF
C237 k3_bar x3 0.06fF
C238 x0 k0_bar 0.06fF
C239 x2_bar a_n1140_n2630# 0.00fF
C240 a_n1140_n1950# XOR1_bar 0.00fF
C241 XOR0_bar a_720_410# 0.00fF
C242 k2_bar a_n840_n270# 0.00fF
C243 x0_bar XOR1_bar 0.00fF
C244 a_420_n270# k2_bar 0.00fF
C245 x1_bar XOR2_bar 0.03fF
C246 XOR0_bar XOR1 0.01fF
C247 k3_bar a_n840_n1950# 0.00fF
C248 a_n1140_n1950# Dis 0.02fF
C249 x3 a_n1140_n2630# 0.00fF
C250 CLK a_420_n2630# 0.02fF
C251 XOR0_bar a_n1140_410# 0.01fF
C252 x0_bar Dis 0.03fF
C253 k2 a_720_n270# 0.00fF
C254 XOR3 x3_bar 0.03fF
C255 k0_bar x2_bar 0.00fF
C256 a_n1140_n1950# x1_bar 0.00fF
C257 k1_bar a_420_410# 0.00fF
C258 x2 a_420_410# 0.00fF
C259 x1_bar x0_bar 0.01fF
C260 a_n840_n270# k1_bar 0.00fF
C261 k2_bar k1_bar 0.01fF
C262 k3_bar XOR3 0.07fF
C263 XOR0 x1 0.00fF
C264 a_n840_n270# x2 0.00fF
C265 a_420_n270# k1_bar 0.00fF
C266 k2_bar x2 0.06fF
C267 XOR1_bar a_420_410# 0.00fF
C268 a_420_n270# x2 0.00fF
C269 a_720_n2630# x3_bar 0.00fF
C270 a_420_n2630# XOR2_bar 0.00fF
C271 CLK a_720_n270# 0.02fF
C272 x0 a_n1140_n270# 0.00fF
C273 k0 k0_bar 1.30fF
C274 XOR1_bar a_n840_n270# 0.01fF
C275 k2_bar XOR1_bar 0.01fF
C276 a_420_n270# XOR1_bar 0.00fF
C277 k1 a_720_n270# 0.00fF
C278 Dis a_420_410# 0.00fF
C279 XOR3 a_n1140_n2630# 0.00fF
C280 a_420_n1950# x2_bar 0.00fF
C281 XOR2 x2_bar 0.03fF
C282 k0_bar XOR1 0.02fF
C283 Dis a_n840_n270# 0.01fF
C284 k2_bar Dis 0.06fF
C285 a_420_n270# Dis 0.00fF
C286 x1_bar a_420_410# 0.00fF
C287 a_n1140_410# k0_bar 0.00fF
C288 a_420_n1950# x3 0.00fF
C289 x2 k1_bar 0.01fF
C290 XOR2 x3 0.00fF
C291 a_n1140_n270# x2_bar 0.00fF
C292 a_720_n270# XOR2_bar 0.00fF
C293 x1 a_n840_n2630# 0.00fF
C294 x1_bar a_n840_n270# 0.00fF
C295 x1_bar k2_bar 0.01fF
C296 CLK XOR0 0.68fF
C297 a_420_n270# x1_bar 0.00fF
C298 XOR1_bar k1_bar 0.30fF
C299 XOR0 k1 0.01fF
C300 a_n840_n1950# XOR2 0.00fF
C301 XOR1_bar x2 0.02fF
C302 k3 a_n840_n2630# 0.00fF
C303 a_420_n1950# XOR1 0.00fF
C304 k2 a_n840_n2630# 0.00fF
C305 XOR2 XOR1 0.03fF
C306 Dis k1_bar 0.06fF
C307 k0 a_n1140_n270# 0.00fF
C308 x0_bar a_720_n270# 0.00fF
C309 Dis x2 0.04fF
C310 x2_bar XOR3_bar 0.00fF
C311 XOR0 XOR2_bar 0.00fF
C312 a_720_n1950# XOR1_bar 0.00fF
C313 XOR1 a_n1140_n270# 0.00fF
C314 x1 x3_bar 0.00fF
C315 x1_bar k1_bar 0.09fF
C316 Dis XOR1_bar 0.33fF
C317 a_420_n1950# XOR3 0.00fF
C318 XOR2 XOR3 0.02fF
C319 x1_bar x2 0.01fF
C320 x1 XOR0_bar 0.00fF
C321 x0 a_n840_410# 0.00fF
C322 k2_bar a_420_n2630# 0.00fF
C323 CLK a_n840_n2630# 0.01fF
C324 x3 XOR3_bar 0.05fF
C325 k3 x3_bar 1.55fF
C326 k3_bar x1 0.00fF
C327 x1_bar XOR1_bar 0.06fF
C328 k2 x3_bar 0.00fF
C329 XOR0 x0_bar 0.03fF
C330 a_n840_n1950# XOR3_bar 0.00fF
C331 XOR2 a_720_n2630# 0.00fF
C332 x1_bar a_720_n1950# 0.00fF
C333 k3 k3_bar 1.30fF
C334 x1_bar Dis 0.03fF
C335 k3_bar k2 0.00fF
C336 XOR1 XOR3_bar 0.00fF
C337 x2_bar a_n840_410# 0.00fF
C338 x1 a_n1140_n2630# 0.00fF
C339 a_n840_n2630# XOR2_bar 0.00fF
C340 CLK x3_bar 0.48fF
C341 a_420_n2630# x2 0.00fF
C342 CLK XOR0_bar 1.01fF
C343 k3 a_n1140_n2630# 0.00fF
C344 k2 a_n1140_n2630# 0.00fF
C345 XOR3 XOR3_bar 0.78fF
C346 CLK k3_bar 0.25fF
C347 k1 XOR0_bar 0.01fF
C348 k0 a_n840_410# 0.00fF
C349 x1 k0_bar 0.00fF
C350 XOR0 a_420_410# 0.01fF
C351 XOR2_bar x3_bar 0.00fF
C352 a_420_n270# XOR0 0.00fF
C353 a_720_n2630# XOR3_bar 0.00fF
C354 CLK a_n1140_n2630# 0.02fF
C355 XOR0_bar XOR2_bar 0.00fF
C356 x1_bar a_420_n2630# 0.00fF
C357 k3_bar XOR2_bar 0.02fF
C358 XOR1_bar a_720_n270# 0.00fF
C359 a_n1140_n1950# x3_bar 0.00fF
C360 x1 a_420_n1950# 0.00fF
C361 x1 XOR2 0.01fF
C362 CLK k0_bar 0.25fF
C363 XOR0_bar x0_bar 0.05fF
C364 XOR2_bar a_n1140_n2630# 0.00fF
C365 XOR0 k1_bar 0.02fF
C366 a_n1140_n1950# k3_bar 0.00fF
C367 k3 a_420_n1950# 0.00fF
C368 k3 XOR2 0.01fF
C369 XOR0 x2 0.00fF
C370 a_420_n1950# k2 0.00fF
C371 k2_bar a_n840_n2630# 0.00fF
C372 x1 a_n1140_n270# 0.00fF
C373 k2 XOR2 0.08fF
C374 k1 k0_bar 0.00fF
C375 x1_bar a_720_n270# 0.00fF
C376 x0 x2_bar 0.00fF
C377 XOR0 XOR1_bar 0.01fF
C378 k2 a_n1140_n270# 0.00fF
C379 XOR0 Dis 0.11fF
C380 CLK a_420_n1950# 0.02fF
C381 CLK XOR2 0.73fF
C382 XOR0_bar a_420_410# 0.00fF
C383 k1 a_420_n1950# 0.00fF
C384 x1 XOR3_bar 0.00fF
C385 x0 k0 0.15fF
C386 k2_bar x3_bar 0.00fF
C387 k1 XOR2 0.03fF
C388 XOR0 x1_bar 0.00fF
C389 XOR0_bar a_n840_n270# 0.00fF
C390 a_n840_n2630# x2 0.00fF
C391 CLK a_n1140_n270# 0.01fF
C392 a_420_n270# XOR0_bar 0.00fF
C393 x0 XOR1 0.00fF
C394 x0_bar k0_bar 0.10fF
C395 k3 XOR3_bar 0.09fF
C396 k3_bar k2_bar 0.05fF
C397 k2 XOR3_bar 0.01fF
C398 k1 a_n1140_n270# 0.00fF
C399 x2_bar x3 0.00fF
C400 a_420_n1950# XOR2_bar 0.00fF
C401 x0 a_n1140_410# 0.00fF
C402 XOR2 XOR2_bar 0.78fF
C403 k0 x2_bar 0.00fF
C404 Dis a_n840_n2630# 0.00fF
C405 x2_bar a_720_410# 0.00fF
C406 a_n840_n1950# x2_bar 0.00fF
C407 k2_bar a_n1140_n2630# 0.00fF
C408 x1 a_n840_410# 0.00fF
C409 a_n1140_n270# XOR2_bar 0.00fF
C410 XOR1 x2_bar 0.02fF
C411 x3_bar x2 0.00fF
C412 CLK XOR3_bar 1.00fF
C413 XOR0_bar k1_bar 0.02fF
C414 a_n1140_n1950# XOR2 0.00fF
C415 x1_bar a_n840_n2630# 0.00fF
C416 XOR0_bar x2 0.00fF
C417 a_n840_n1950# x3 0.00fF
C418 a_n1140_410# x2_bar 0.00fF
C419 k0_bar a_420_410# 0.00fF
C420 k3_bar x2 0.00fF
C421 XOR0_bar XOR1_bar 0.02fF
C422 k0 a_720_410# 0.00fF
C423 k0_bar a_n840_n270# 0.00fF
C424 a_720_n1950# x3_bar 0.00fF
C425 x2_bar XOR3 0.00fF
C426 a_420_n270# k0_bar 0.00fF
C427 x0_bar a_n1140_n270# 0.00fF
C428 k0 XOR1 0.01fF
C429 Dis x3_bar 0.01fF
C430 XOR1 a_720_410# 0.00fF
C431 XOR0_bar Dis 0.32fF
C432 XOR2_bar XOR3_bar 0.02fF
C433 x2 a_n1140_n2630# 0.00fF
C434 XOR0 a_720_n270# 0.00fF
C435 k0 a_n1140_410# 0.00fF
C436 XOR3 x3 0.03fF
C437 x1_bar x3_bar 0.00fF
C438 k3_bar Dis 0.03fF
C439 CLK a_n840_410# 0.01fF
C440 x2_bar a_720_n2630# 0.00fF
C441 x1_bar XOR0_bar 0.00fF
C442 k1 a_n840_410# 0.00fF
C443 a_n1140_n1950# XOR3_bar 0.00fF
C444 x1_bar k3_bar 0.00fF
C445 k2_bar a_420_n1950# 0.00fF
C446 k0_bar k1_bar 0.05fF
C447 k2_bar XOR2 0.07fF
C448 XOR1 XOR3 0.00fF
C449 Dis a_n1140_n2630# 0.01fF
C450 a_420_n270# XOR2 0.00fF
C451 k0_bar x2 0.00fF
C452 k0_bar XOR1_bar 0.02fF
C453 k2_bar a_n1140_n270# 0.00fF
C454 x1_bar a_n1140_n2630# 0.00fF
C455 a_420_n2630# x3_bar 0.00fF
C456 x0 x1 0.01fF
C457 Dis k0_bar 0.06fF
C458 a_420_n1950# k1_bar 0.00fF
C459 XOR2 k1_bar 0.00fF
C460 a_420_n1950# x2 0.00fF
C461 k3_bar a_420_n2630# 0.00fF
C462 XOR2 x2 0.03fF
C463 x0_bar a_n840_410# 0.00fF
C464 x1_bar k0_bar 0.00fF
C465 XOR3 a_720_n2630# 0.01fF
C466 a_420_n1950# XOR1_bar 0.00fF
C467 XOR1_bar XOR2 0.03fF
C468 k2_bar XOR3_bar 0.02fF
C469 a_n1140_n270# k1_bar 0.00fF
C470 a_n1140_n270# x2 0.00fF
C471 x1 x2_bar 0.01fF
C472 XOR0_bar a_720_n270# 0.00fF
C473 a_720_n1950# XOR2 0.01fF
C474 Dis a_420_n1950# 0.00fF
C475 Dis XOR2 0.11fF
C476 XOR1_bar a_n1140_n270# 0.01fF
C477 k3 x2_bar 0.00fF
C478 x0 CLK 1.11fF
C479 k2 x2_bar 1.55fF
C480 x1 x3 0.00fF
C481 x1_bar a_420_n1950# 0.00fF
C482 x1_bar XOR2 0.02fF
C483 x0 k1 0.00fF
C484 Dis a_n1140_n270# 0.02fF
C485 x1 k0 0.00fF
C486 x1 a_n840_n1950# 0.00fF
C487 k3 x3 0.15fF
C488 x2 XOR3_bar 0.00fF
C489 k2 x3 0.00fF
C490 x1 XOR1 0.03fF
C491 XOR0 XOR0_bar 0.78fF
C492 x1_bar a_n1140_n270# 0.00fF
C493 CLK x2_bar 0.58fF
C494 XOR1_bar XOR3_bar 0.00fF
C495 k3 a_n840_n1950# 0.00fF
C496 a_n840_n1950# k2 0.00fF
C497 x1 a_n1140_410# 0.00fF
C498 a_720_n2630# GND 0.01fF
C499 a_420_n2630# GND 0.02fF
C500 a_n840_n2630# GND 0.02fF
C501 a_n1140_n2630# GND 0.01fF
C502 XOR3_bar GND 1.14fF
C503 XOR3 GND 1.03fF
C504 k3 GND 0.65fF
C505 x3 GND 0.69fF
C506 x3_bar GND 0.55fF
C507 k3_bar GND 0.66fF
C508 a_720_n1950# GND 0.01fF
C509 a_420_n1950# GND 0.02fF
C510 a_n840_n1950# GND 0.02fF
C511 a_n1140_n1950# GND 0.02fF
C512 k2 GND 0.60fF
C513 k2_bar GND 0.66fF
C514 x2_bar GND 0.53fF
C515 XOR2_bar GND 1.09fF
C516 XOR2 GND 0.99fF
C517 x2 GND 0.56fF
C518 a_720_n270# GND 0.01fF
C519 a_420_n270# GND 0.02fF
C520 a_n840_n270# GND 0.02fF
C521 a_n1140_n270# GND 0.02fF
C522 XOR1_bar GND 1.09fF
C523 XOR1 GND 0.99fF
C524 k1 GND 0.60fF
C525 x1 GND 0.56fF
C526 x1_bar GND 0.53fF
C527 k1_bar GND 0.66fF
C528 a_720_410# GND 0.01fF
C529 a_420_410# GND 0.02fF
C530 a_n840_410# GND 0.02fF
C531 a_n1140_410# GND 0.01fF
C532 Dis GND 7.23fF
C533 k0 GND 0.65fF
C534 k0_bar GND 0.65fF
C535 x0_bar GND 0.55fF
C536 XOR0_bar GND 1.14fF
C537 XOR0 GND 1.03fF
C538 x0 GND 0.68fF
C539 CLK GND 14.90fF
C540 Dis.t7 GND 0.17fF
C541 Dis.t1 GND 0.11fF
C542 Dis.n0 GND 0.43fF $ **FLOATING
C543 Dis.t4 GND 0.17fF
C544 Dis.t5 GND 0.11fF
C545 Dis.n1 GND 0.43fF $ **FLOATING
C546 EESPFAL_XOR_v3_1/Dis GND 0.21fF $ **FLOATING
C547 Dis.t3 GND 0.17fF
C548 Dis.t6 GND 0.11fF
C549 Dis.n2 GND 0.43fF $ **FLOATING
C550 EESPFAL_XOR_v3_2/Dis GND 0.21fF $ **FLOATING
C551 Dis.t2 GND 0.17fF
C552 Dis.t0 GND 0.11fF
C553 Dis.n3 GND 0.43fF $ **FLOATING
C554 Dis.n4 GND 0.62fF $ **FLOATING
C555 Dis.n5 GND 0.90fF $ **FLOATING
C556 Dis.n6 GND 1.26fF $ **FLOATING
C557 EESPFAL_XOR_v3_0/Dis GND 0.21fF $ **FLOATING
C558 CLK.t34 GND 0.02fF
C559 CLK.t11 GND 0.02fF
C560 CLK.n0 GND 0.06fF $ **FLOATING
C561 CLK.t7 GND 0.03fF
C562 CLK.n1 GND 0.02fF $ **FLOATING
C563 CLK.t12 GND 0.02fF
C564 CLK.t0 GND 0.02fF
C565 CLK.n2 GND 0.04fF $ **FLOATING
C566 CLK.n3 GND 0.01fF $ **FLOATING
C567 CLK.t28 GND 0.02fF
C568 CLK.t37 GND 0.02fF
C569 CLK.n4 GND 0.04fF $ **FLOATING
C570 CLK.n5 GND 0.01fF $ **FLOATING
C571 CLK.n6 GND 0.01fF $ **FLOATING
C572 CLK.n7 GND 0.02fF $ **FLOATING
C573 CLK.t39 GND 0.02fF
C574 CLK.t31 GND 0.02fF
C575 CLK.n8 GND 0.04fF $ **FLOATING
C576 CLK.n9 GND 0.01fF $ **FLOATING
C577 CLK.t22 GND 0.02fF
C578 CLK.t32 GND 0.02fF
C579 CLK.n10 GND 0.04fF $ **FLOATING
C580 CLK.n11 GND 0.01fF $ **FLOATING
C581 CLK.n12 GND 0.01fF $ **FLOATING
C582 CLK.n13 GND 0.05fF $ **FLOATING
C583 CLK.n14 GND 0.02fF $ **FLOATING
C584 CLK.n15 GND 0.01fF $ **FLOATING
C585 CLK.n16 GND 0.12fF $ **FLOATING
C586 CLK.n17 GND 0.04fF $ **FLOATING
C587 CLK.n18 GND 0.02fF $ **FLOATING
C588 CLK.n19 GND 0.01fF $ **FLOATING
C589 CLK.n20 GND 0.06fF $ **FLOATING
C590 CLK.n21 GND 0.03fF $ **FLOATING
C591 CLK.n22 GND 0.02fF $ **FLOATING
C592 CLK.n23 GND 0.01fF $ **FLOATING
C593 CLK.n24 GND 0.01fF $ **FLOATING
C594 CLK.t18 GND 0.03fF
C595 CLK.t14 GND 0.02fF
C596 CLK.t30 GND 0.02fF
C597 CLK.n25 GND 0.06fF $ **FLOATING
C598 EESPFAL_XOR_v3_0/CLK GND 0.01fF $ **FLOATING
C599 CLK.t21 GND 0.03fF
C600 CLK.t35 GND 0.02fF
C601 CLK.t19 GND 0.02fF
C602 CLK.n26 GND 0.09fF $ **FLOATING
C603 CLK.n27 GND 0.05fF $ **FLOATING
C604 CLK.n28 GND 0.02fF $ **FLOATING
C605 CLK.n29 GND 0.01fF $ **FLOATING
C606 CLK.n30 GND 0.12fF $ **FLOATING
C607 CLK.n31 GND 0.04fF $ **FLOATING
C608 CLK.n32 GND 0.02fF $ **FLOATING
C609 CLK.n33 GND 0.01fF $ **FLOATING
C610 CLK.n34 GND 0.06fF $ **FLOATING
C611 CLK.n35 GND 0.03fF $ **FLOATING
C612 CLK.n36 GND 0.02fF $ **FLOATING
C613 CLK.n37 GND 0.01fF $ **FLOATING
C614 CLK.n38 GND 0.01fF $ **FLOATING
C615 CLK.n39 GND 0.11fF $ **FLOATING
C616 CLK.n40 GND 0.03fF $ **FLOATING
C617 CLK.n41 GND 0.02fF $ **FLOATING
C618 CLK.n42 GND 0.01fF $ **FLOATING
C619 CLK.n43 GND 0.02fF $ **FLOATING
C620 CLK.n44 GND 0.03fF $ **FLOATING
C621 CLK.n45 GND 0.02fF $ **FLOATING
C622 CLK.n46 GND 0.01fF $ **FLOATING
C623 CLK.n47 GND 0.02fF $ **FLOATING
C624 CLK.n48 GND 0.03fF $ **FLOATING
C625 CLK.n49 GND 0.02fF $ **FLOATING
C626 CLK.n50 GND 0.01fF $ **FLOATING
C627 CLK.n51 GND 0.02fF $ **FLOATING
C628 CLK.n52 GND 0.03fF $ **FLOATING
C629 CLK.n53 GND 0.02fF $ **FLOATING
C630 CLK.n54 GND 0.01fF $ **FLOATING
C631 CLK.n55 GND 0.02fF $ **FLOATING
C632 CLK.n56 GND 0.08fF $ **FLOATING
C633 CLK.n57 GND 0.02fF $ **FLOATING
C634 CLK.n58 GND 0.01fF $ **FLOATING
C635 CLK.n59 GND 0.02fF $ **FLOATING
C636 CLK.n60 GND 0.11fF $ **FLOATING
C637 CLK.n61 GND 0.02fF $ **FLOATING
C638 CLK.n62 GND 0.01fF $ **FLOATING
C639 CLK.n63 GND 0.01fF $ **FLOATING
C640 CLK.n64 GND 0.18fF $ **FLOATING
C641 CLK.t20 GND 0.05fF
C642 CLK.n65 GND 0.06fF $ **FLOATING
C643 CLK.n66 GND 0.02fF $ **FLOATING
C644 CLK.n67 GND 0.01fF $ **FLOATING
C645 CLK.n68 GND 0.02fF $ **FLOATING
C646 CLK.n69 GND 0.10fF $ **FLOATING
C647 CLK.n70 GND 0.02fF $ **FLOATING
C648 CLK.n71 GND 0.01fF $ **FLOATING
C649 CLK.n72 GND 0.02fF $ **FLOATING
C650 CLK.n73 GND 0.02fF $ **FLOATING
C651 CLK.t29 GND 0.05fF
C652 CLK.n74 GND 0.06fF $ **FLOATING
C653 CLK.n75 GND 0.02fF $ **FLOATING
C654 CLK.n76 GND 0.01fF $ **FLOATING
C655 CLK.n77 GND 0.10fF $ **FLOATING
C656 CLK.n78 GND 0.02fF $ **FLOATING
C657 CLK.n79 GND 0.01fF $ **FLOATING
C658 CLK.n80 GND 0.10fF $ **FLOATING
C659 CLK.t13 GND 0.05fF
C660 CLK.n81 GND 0.06fF $ **FLOATING
C661 CLK.n82 GND 0.02fF $ **FLOATING
C662 CLK.n83 GND 0.01fF $ **FLOATING
C663 CLK.n84 GND 0.02fF $ **FLOATING
C664 CLK.n85 GND 0.10fF $ **FLOATING
C665 CLK.n86 GND 0.02fF $ **FLOATING
C666 CLK.n87 GND 0.01fF $ **FLOATING
C667 CLK.n88 GND 0.02fF $ **FLOATING
C668 CLK.t17 GND 0.05fF
C669 CLK.n89 GND 0.06fF $ **FLOATING
C670 CLK.n90 GND 0.02fF $ **FLOATING
C671 CLK.n91 GND 0.01fF $ **FLOATING
C672 CLK.n92 GND 0.02fF $ **FLOATING
C673 CLK.n93 GND 0.18fF $ **FLOATING
C674 CLK.n94 GND 0.11fF $ **FLOATING
C675 CLK.n95 GND 0.02fF $ **FLOATING
C676 CLK.n96 GND 0.01fF $ **FLOATING
C677 CLK.n97 GND 0.01fF $ **FLOATING
C678 CLK.n98 GND 0.08fF $ **FLOATING
C679 CLK.n99 GND 0.02fF $ **FLOATING
C680 CLK.n100 GND 0.01fF $ **FLOATING
C681 CLK.n101 GND 0.02fF $ **FLOATING
C682 CLK.n102 GND 0.03fF $ **FLOATING
C683 CLK.n103 GND 0.02fF $ **FLOATING
C684 CLK.n104 GND 0.01fF $ **FLOATING
C685 CLK.n105 GND 0.02fF $ **FLOATING
C686 CLK.n106 GND 0.03fF $ **FLOATING
C687 CLK.n107 GND 0.02fF $ **FLOATING
C688 CLK.n108 GND 0.01fF $ **FLOATING
C689 CLK.n109 GND 0.02fF $ **FLOATING
C690 CLK.n110 GND 0.03fF $ **FLOATING
C691 CLK.n111 GND 0.02fF $ **FLOATING
C692 CLK.n112 GND 0.01fF $ **FLOATING
C693 CLK.n113 GND 0.02fF $ **FLOATING
C694 CLK.n114 GND 0.03fF $ **FLOATING
C695 CLK.n115 GND 0.02fF $ **FLOATING
C696 CLK.n116 GND 0.01fF $ **FLOATING
C697 CLK.n117 GND 0.02fF $ **FLOATING
C698 CLK.n118 GND 0.04fF $ **FLOATING
C699 CLK.n119 GND 0.05fF $ **FLOATING
C700 CLK.n120 GND 0.01fF $ **FLOATING
C701 CLK.n121 GND 0.01fF $ **FLOATING
C702 CLK.n122 GND 0.07fF $ **FLOATING
C703 CLK.n123 GND 0.07fF $ **FLOATING
C704 CLK.n124 GND 0.01fF $ **FLOATING
C705 CLK.n125 GND 0.01fF $ **FLOATING
C706 CLK.n126 GND 0.05fF $ **FLOATING
C707 CLK.n127 GND 0.05fF $ **FLOATING
C708 CLK.n128 GND 0.02fF $ **FLOATING
C709 CLK.n129 GND 0.01fF $ **FLOATING
C710 CLK.n130 GND 0.13fF $ **FLOATING
C711 CLK.n131 GND 0.04fF $ **FLOATING
C712 CLK.n132 GND 0.02fF $ **FLOATING
C713 CLK.n133 GND 0.01fF $ **FLOATING
C714 CLK.n134 GND 0.06fF $ **FLOATING
C715 CLK.n135 GND 0.04fF $ **FLOATING
C716 CLK.n136 GND 0.02fF $ **FLOATING
C717 CLK.n137 GND 0.01fF $ **FLOATING
C718 CLK.n138 GND 0.01fF $ **FLOATING
C719 CLK.t8 GND 0.03fF
C720 CLK.t5 GND 0.03fF
C721 CLK.t2 GND 0.02fF
C722 CLK.t41 GND 0.02fF
C723 CLK.n139 GND 0.06fF $ **FLOATING
C724 CLK.t9 GND 0.02fF
C725 CLK.t25 GND 0.02fF
C726 CLK.n140 GND 0.06fF $ **FLOATING
C727 EESPFAL_XOR_v3_2/CLK GND 0.01fF $ **FLOATING
C728 CLK.t42 GND 0.03fF
C729 CLK.t27 GND 0.03fF
C730 CLK.t38 GND 0.02fF
C731 CLK.t3 GND 0.02fF
C732 CLK.n141 GND 0.09fF $ **FLOATING
C733 CLK.t43 GND 0.02fF
C734 CLK.t40 GND 0.02fF
C735 CLK.n142 GND 0.09fF $ **FLOATING
C736 CLK.n143 GND 0.05fF $ **FLOATING
C737 CLK.n144 GND 0.02fF $ **FLOATING
C738 CLK.n145 GND 0.01fF $ **FLOATING
C739 CLK.n146 GND 0.13fF $ **FLOATING
C740 CLK.n147 GND 0.04fF $ **FLOATING
C741 CLK.n148 GND 0.02fF $ **FLOATING
C742 CLK.n149 GND 0.01fF $ **FLOATING
C743 CLK.n150 GND 0.06fF $ **FLOATING
C744 CLK.n151 GND 0.04fF $ **FLOATING
C745 CLK.n152 GND 0.02fF $ **FLOATING
C746 CLK.n153 GND 0.01fF $ **FLOATING
C747 CLK.n154 GND 0.01fF $ **FLOATING
C748 CLK.n155 GND 0.22fF $ **FLOATING
C749 CLK.n156 GND 0.04fF $ **FLOATING
C750 CLK.n157 GND 0.02fF $ **FLOATING
C751 CLK.n158 GND 0.01fF $ **FLOATING
C752 CLK.n159 GND 0.02fF $ **FLOATING
C753 CLK.n160 GND 0.04fF $ **FLOATING
C754 CLK.n161 GND 0.02fF $ **FLOATING
C755 CLK.n162 GND 0.01fF $ **FLOATING
C756 CLK.n163 GND 0.02fF $ **FLOATING
C757 CLK.n164 GND 0.04fF $ **FLOATING
C758 CLK.n165 GND 0.02fF $ **FLOATING
C759 CLK.n166 GND 0.01fF $ **FLOATING
C760 CLK.n167 GND 0.02fF $ **FLOATING
C761 CLK.n168 GND 0.04fF $ **FLOATING
C762 CLK.n169 GND 0.02fF $ **FLOATING
C763 CLK.n170 GND 0.01fF $ **FLOATING
C764 CLK.n171 GND 0.02fF $ **FLOATING
C765 CLK.n172 GND 0.13fF $ **FLOATING
C766 CLK.n173 GND 0.02fF $ **FLOATING
C767 CLK.n174 GND 0.01fF $ **FLOATING
C768 CLK.n175 GND 0.02fF $ **FLOATING
C769 CLK.n176 GND 0.18fF $ **FLOATING
C770 CLK.n177 GND 0.02fF $ **FLOATING
C771 CLK.n178 GND 0.01fF $ **FLOATING
C772 CLK.n179 GND 0.01fF $ **FLOATING
C773 CLK.n180 GND 0.34fF $ **FLOATING
C774 CLK.t26 GND 0.09fF
C775 CLK.n181 GND 0.10fF $ **FLOATING
C776 CLK.n182 GND 0.02fF $ **FLOATING
C777 CLK.n183 GND 0.01fF $ **FLOATING
C778 CLK.n184 GND 0.02fF $ **FLOATING
C779 CLK.n185 GND 0.16fF $ **FLOATING
C780 CLK.n186 GND 0.02fF $ **FLOATING
C781 CLK.n187 GND 0.01fF $ **FLOATING
C782 CLK.n188 GND 0.02fF $ **FLOATING
C783 CLK.n189 GND 0.02fF $ **FLOATING
C784 CLK.t24 GND 0.09fF
C785 CLK.n190 GND 0.09fF $ **FLOATING
C786 CLK.n191 GND 0.02fF $ **FLOATING
C787 CLK.n192 GND 0.01fF $ **FLOATING
C788 CLK.n193 GND 0.16fF $ **FLOATING
C789 CLK.n194 GND 0.02fF $ **FLOATING
C790 CLK.n195 GND 0.01fF $ **FLOATING
C791 CLK.n196 GND 0.20fF $ **FLOATING
C792 CLK.t1 GND 0.09fF
C793 CLK.n197 GND 0.09fF $ **FLOATING
C794 CLK.n198 GND 0.02fF $ **FLOATING
C795 CLK.n199 GND 0.01fF $ **FLOATING
C796 CLK.n200 GND 0.02fF $ **FLOATING
C797 CLK.n201 GND 0.16fF $ **FLOATING
C798 CLK.n202 GND 0.02fF $ **FLOATING
C799 CLK.n203 GND 0.01fF $ **FLOATING
C800 CLK.n204 GND 0.02fF $ **FLOATING
C801 CLK.t4 GND 0.09fF
C802 CLK.n205 GND 0.10fF $ **FLOATING
C803 CLK.n206 GND 0.02fF $ **FLOATING
C804 CLK.n207 GND 0.01fF $ **FLOATING
C805 CLK.n208 GND 0.02fF $ **FLOATING
C806 CLK.n209 GND 0.34fF $ **FLOATING
C807 CLK.n210 GND 0.18fF $ **FLOATING
C808 CLK.n211 GND 0.02fF $ **FLOATING
C809 CLK.n212 GND 0.01fF $ **FLOATING
C810 CLK.n213 GND 0.01fF $ **FLOATING
C811 CLK.n214 GND 0.13fF $ **FLOATING
C812 CLK.n215 GND 0.02fF $ **FLOATING
C813 CLK.n216 GND 0.01fF $ **FLOATING
C814 CLK.n217 GND 0.02fF $ **FLOATING
C815 CLK.n218 GND 0.04fF $ **FLOATING
C816 CLK.n219 GND 0.02fF $ **FLOATING
C817 CLK.n220 GND 0.01fF $ **FLOATING
C818 CLK.n221 GND 0.02fF $ **FLOATING
C819 CLK.n222 GND 0.04fF $ **FLOATING
C820 CLK.n223 GND 0.02fF $ **FLOATING
C821 CLK.n224 GND 0.01fF $ **FLOATING
C822 CLK.n225 GND 0.02fF $ **FLOATING
C823 CLK.n226 GND 0.04fF $ **FLOATING
C824 CLK.n227 GND 0.02fF $ **FLOATING
C825 CLK.n228 GND 0.01fF $ **FLOATING
C826 CLK.n229 GND 0.02fF $ **FLOATING
C827 CLK.n230 GND 0.04fF $ **FLOATING
C828 CLK.n231 GND 0.02fF $ **FLOATING
C829 CLK.n232 GND 0.01fF $ **FLOATING
C830 CLK.n233 GND 0.02fF $ **FLOATING
C831 CLK.n234 GND 0.07fF $ **FLOATING
C832 CLK.n235 GND 0.05fF $ **FLOATING
C833 CLK.n236 GND 0.01fF $ **FLOATING
C834 CLK.n237 GND 0.01fF $ **FLOATING
C835 CLK.n238 GND 0.07fF $ **FLOATING
C836 CLK.n239 GND 0.07fF $ **FLOATING
C837 CLK.n240 GND 0.01fF $ **FLOATING
C838 CLK.n241 GND 0.01fF $ **FLOATING
C839 CLK.n242 GND 0.05fF $ **FLOATING
C840 CLK.n243 GND 0.05fF $ **FLOATING
C841 CLK.n244 GND 0.02fF $ **FLOATING
C842 CLK.n245 GND 0.01fF $ **FLOATING
C843 CLK.n246 GND 0.12fF $ **FLOATING
C844 CLK.n247 GND 0.04fF $ **FLOATING
C845 CLK.n248 GND 0.02fF $ **FLOATING
C846 CLK.n249 GND 0.01fF $ **FLOATING
C847 CLK.n250 GND 0.06fF $ **FLOATING
C848 CLK.n251 GND 0.03fF $ **FLOATING
C849 CLK.n252 GND 0.02fF $ **FLOATING
C850 CLK.n253 GND 0.01fF $ **FLOATING
C851 CLK.n254 GND 0.01fF $ **FLOATING
C852 CLK.n255 GND 0.04fF $ **FLOATING
C853 CLK.n256 GND 0.03fF $ **FLOATING
C854 CLK.n257 GND 0.02fF $ **FLOATING
C855 CLK.n258 GND 0.01fF $ **FLOATING
C856 CLK.n259 GND 0.02fF $ **FLOATING
C857 CLK.n260 GND 0.03fF $ **FLOATING
C858 CLK.n261 GND 0.02fF $ **FLOATING
C859 CLK.n262 GND 0.01fF $ **FLOATING
C860 CLK.n263 GND 0.02fF $ **FLOATING
C861 CLK.n264 GND 0.03fF $ **FLOATING
C862 CLK.n265 GND 0.02fF $ **FLOATING
C863 CLK.n266 GND 0.01fF $ **FLOATING
C864 CLK.n267 GND 0.02fF $ **FLOATING
C865 CLK.n268 GND 0.03fF $ **FLOATING
C866 CLK.n269 GND 0.02fF $ **FLOATING
C867 CLK.n270 GND 0.01fF $ **FLOATING
C868 CLK.n271 GND 0.02fF $ **FLOATING
C869 CLK.n272 GND 0.08fF $ **FLOATING
C870 CLK.n273 GND 0.02fF $ **FLOATING
C871 CLK.n274 GND 0.01fF $ **FLOATING
C872 CLK.n275 GND 0.02fF $ **FLOATING
C873 CLK.n276 GND 0.11fF $ **FLOATING
C874 CLK.n277 GND 0.02fF $ **FLOATING
C875 CLK.n278 GND 0.01fF $ **FLOATING
C876 CLK.n279 GND 0.01fF $ **FLOATING
C877 CLK.n280 GND 0.18fF $ **FLOATING
C878 CLK.t6 GND 0.05fF
C879 CLK.n281 GND 0.06fF $ **FLOATING
C880 CLK.n282 GND 0.02fF $ **FLOATING
C881 CLK.n283 GND 0.01fF $ **FLOATING
C882 CLK.n284 GND 0.02fF $ **FLOATING
C883 CLK.n285 GND 0.10fF $ **FLOATING
C884 CLK.n286 GND 0.02fF $ **FLOATING
C885 CLK.n287 GND 0.01fF $ **FLOATING
C886 CLK.n288 GND 0.02fF $ **FLOATING
C887 CLK.t33 GND 0.05fF
C888 CLK.n289 GND 0.06fF $ **FLOATING
C889 CLK.n290 GND 0.02fF $ **FLOATING
C890 CLK.n291 GND 0.01fF $ **FLOATING
C891 CLK.n292 GND 0.02fF $ **FLOATING
C892 CLK.n293 GND 0.10fF $ **FLOATING
C893 CLK.n294 GND 0.02fF $ **FLOATING
C894 CLK.n295 GND 0.01fF $ **FLOATING
C895 CLK.n296 GND 0.10fF $ **FLOATING
C896 CLK.t16 GND 0.03fF
C897 CLK.t23 GND 0.02fF
C898 CLK.t36 GND 0.02fF
C899 CLK.n297 GND 0.09fF $ **FLOATING
C900 CLK.n298 GND 0.12fF $ **FLOATING
C901 CLK.n299 GND 0.03fF $ **FLOATING
C902 CLK.n300 GND 0.05fF $ **FLOATING
C903 CLK.n301 GND 0.02fF $ **FLOATING
C904 CLK.n302 GND 0.01fF $ **FLOATING
C905 CLK.n303 GND 0.02fF $ **FLOATING
C906 CLK.n304 GND 0.04fF $ **FLOATING
C907 CLK.n305 GND 0.02fF $ **FLOATING
C908 CLK.n306 GND 0.01fF $ **FLOATING
C909 CLK.n307 GND 0.02fF $ **FLOATING
C910 CLK.n308 GND 0.03fF $ **FLOATING
C911 CLK.n309 GND 0.02fF $ **FLOATING
C912 CLK.n310 GND 0.01fF $ **FLOATING
C913 CLK.n311 GND 0.01fF $ **FLOATING
C914 CLK.n312 GND 0.11fF $ **FLOATING
C915 CLK.n313 GND 0.03fF $ **FLOATING
C916 CLK.n314 GND 0.02fF $ **FLOATING
C917 CLK.n315 GND 0.01fF $ **FLOATING
C918 CLK.n316 GND 0.02fF $ **FLOATING
C919 CLK.n317 GND 0.03fF $ **FLOATING
C920 CLK.n318 GND 0.02fF $ **FLOATING
C921 CLK.n319 GND 0.01fF $ **FLOATING
C922 CLK.n320 GND 0.02fF $ **FLOATING
C923 CLK.n321 GND 0.03fF $ **FLOATING
C924 CLK.n322 GND 0.02fF $ **FLOATING
C925 CLK.n323 GND 0.01fF $ **FLOATING
C926 CLK.n324 GND 0.02fF $ **FLOATING
C927 CLK.n325 GND 0.03fF $ **FLOATING
C928 CLK.n326 GND 0.02fF $ **FLOATING
C929 CLK.n327 GND 0.01fF $ **FLOATING
C930 CLK.n328 GND 0.02fF $ **FLOATING
C931 CLK.n329 GND 0.08fF $ **FLOATING
C932 CLK.n330 GND 0.02fF $ **FLOATING
C933 CLK.n331 GND 0.01fF $ **FLOATING
C934 CLK.n332 GND 0.02fF $ **FLOATING
C935 CLK.n333 GND 0.11fF $ **FLOATING
C936 CLK.n334 GND 0.02fF $ **FLOATING
C937 CLK.n335 GND 0.01fF $ **FLOATING
C938 CLK.n336 GND 0.01fF $ **FLOATING
C939 CLK.n337 GND 0.18fF $ **FLOATING
C940 CLK.t15 GND 0.05fF
C941 CLK.n338 GND 0.06fF $ **FLOATING
C942 CLK.n339 GND 0.02fF $ **FLOATING
C943 CLK.n340 GND 0.01fF $ **FLOATING
C944 CLK.n341 GND 0.02fF $ **FLOATING
C945 CLK.n342 GND 0.10fF $ **FLOATING
C946 CLK.n343 GND 0.02fF $ **FLOATING
C947 CLK.n344 GND 0.01fF $ **FLOATING
C948 CLK.n345 GND 0.02fF $ **FLOATING
C949 CLK.t10 GND 0.05fF
C950 CLK.n346 GND 0.06fF $ **FLOATING
C951 CLK.n347 GND 0.02fF $ **FLOATING
C952 CLK.n348 GND 0.01fF $ **FLOATING
C953 CLK.n349 GND 0.02fF $ **FLOATING
.ends

