magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -805 0 -115 50
<< l67d20 >>
rect -805 5 -115 45
<< l66d44 >>
rect -775 17 -758 34
rect -741 17 -724 34
rect -707 17 -690 34
rect -673 17 -656 34
rect -639 17 -622 34
rect -605 17 -588 34
rect -571 17 -554 34
rect -537 17 -520 34
rect -503 17 -486 34
rect -469 17 -452 34
rect -435 17 -418 34
rect -401 17 -384 34
rect -367 17 -350 34
rect -333 17 -316 34
rect -299 17 -282 34
rect -265 17 -248 34
rect -231 17 -214 34
rect -197 17 -180 34
rect -163 17 -146 34
<< l67d44 >>
rect -775 17 -758 34
rect -739 17 -722 34
rect -703 17 -686 34
rect -667 17 -650 34
rect -631 17 -614 34
rect -595 17 -578 34
rect -559 17 -542 34
rect -523 17 -506 34
rect -487 17 -470 34
rect -451 17 -434 34
rect -415 17 -398 34
rect -379 17 -362 34
rect -343 17 -326 34
rect -307 17 -290 34
rect -271 17 -254 34
rect -235 17 -218 34
rect -199 17 -182 34
rect -163 17 -146 34
<< l68d20 >>
rect -805 0 -115 50
<< end >>
