magic
tech sky130A
magscale 1 2
timestamp 1671080676
<< pwell >>
rect -1796 34 -624 926
<< nmoslvt >>
rect -1530 60 -1430 900
rect -1310 60 -1210 900
rect -1090 60 -990 900
rect -870 60 -770 900
<< ndiff >>
rect -1650 876 -1530 900
rect -1650 842 -1607 876
rect -1573 842 -1530 876
rect -1650 808 -1530 842
rect -1650 774 -1607 808
rect -1573 774 -1530 808
rect -1650 740 -1530 774
rect -1650 706 -1607 740
rect -1573 706 -1530 740
rect -1650 672 -1530 706
rect -1650 638 -1607 672
rect -1573 638 -1530 672
rect -1650 604 -1530 638
rect -1650 570 -1607 604
rect -1573 570 -1530 604
rect -1650 536 -1530 570
rect -1650 502 -1607 536
rect -1573 502 -1530 536
rect -1650 468 -1530 502
rect -1650 434 -1607 468
rect -1573 434 -1530 468
rect -1650 400 -1530 434
rect -1650 366 -1607 400
rect -1573 366 -1530 400
rect -1650 332 -1530 366
rect -1650 298 -1607 332
rect -1573 298 -1530 332
rect -1650 264 -1530 298
rect -1650 230 -1607 264
rect -1573 230 -1530 264
rect -1650 196 -1530 230
rect -1650 162 -1607 196
rect -1573 162 -1530 196
rect -1650 128 -1530 162
rect -1650 94 -1607 128
rect -1573 94 -1530 128
rect -1650 60 -1530 94
rect -1430 876 -1310 900
rect -1430 842 -1387 876
rect -1353 842 -1310 876
rect -1430 808 -1310 842
rect -1430 774 -1387 808
rect -1353 774 -1310 808
rect -1430 740 -1310 774
rect -1430 706 -1387 740
rect -1353 706 -1310 740
rect -1430 672 -1310 706
rect -1430 638 -1387 672
rect -1353 638 -1310 672
rect -1430 604 -1310 638
rect -1430 570 -1387 604
rect -1353 570 -1310 604
rect -1430 536 -1310 570
rect -1430 502 -1387 536
rect -1353 502 -1310 536
rect -1430 468 -1310 502
rect -1430 434 -1387 468
rect -1353 434 -1310 468
rect -1430 400 -1310 434
rect -1430 366 -1387 400
rect -1353 366 -1310 400
rect -1430 332 -1310 366
rect -1430 298 -1387 332
rect -1353 298 -1310 332
rect -1430 264 -1310 298
rect -1430 230 -1387 264
rect -1353 230 -1310 264
rect -1430 196 -1310 230
rect -1430 162 -1387 196
rect -1353 162 -1310 196
rect -1430 128 -1310 162
rect -1430 94 -1387 128
rect -1353 94 -1310 128
rect -1430 60 -1310 94
rect -1210 876 -1090 900
rect -1210 842 -1167 876
rect -1133 842 -1090 876
rect -1210 808 -1090 842
rect -1210 774 -1167 808
rect -1133 774 -1090 808
rect -1210 740 -1090 774
rect -1210 706 -1167 740
rect -1133 706 -1090 740
rect -1210 672 -1090 706
rect -1210 638 -1167 672
rect -1133 638 -1090 672
rect -1210 604 -1090 638
rect -1210 570 -1167 604
rect -1133 570 -1090 604
rect -1210 536 -1090 570
rect -1210 502 -1167 536
rect -1133 502 -1090 536
rect -1210 468 -1090 502
rect -1210 434 -1167 468
rect -1133 434 -1090 468
rect -1210 400 -1090 434
rect -1210 366 -1167 400
rect -1133 366 -1090 400
rect -1210 332 -1090 366
rect -1210 298 -1167 332
rect -1133 298 -1090 332
rect -1210 264 -1090 298
rect -1210 230 -1167 264
rect -1133 230 -1090 264
rect -1210 196 -1090 230
rect -1210 162 -1167 196
rect -1133 162 -1090 196
rect -1210 128 -1090 162
rect -1210 94 -1167 128
rect -1133 94 -1090 128
rect -1210 60 -1090 94
rect -990 876 -870 900
rect -990 842 -947 876
rect -913 842 -870 876
rect -990 808 -870 842
rect -990 774 -947 808
rect -913 774 -870 808
rect -990 740 -870 774
rect -990 706 -947 740
rect -913 706 -870 740
rect -990 672 -870 706
rect -990 638 -947 672
rect -913 638 -870 672
rect -990 604 -870 638
rect -990 570 -947 604
rect -913 570 -870 604
rect -990 536 -870 570
rect -990 502 -947 536
rect -913 502 -870 536
rect -990 468 -870 502
rect -990 434 -947 468
rect -913 434 -870 468
rect -990 400 -870 434
rect -990 366 -947 400
rect -913 366 -870 400
rect -990 332 -870 366
rect -990 298 -947 332
rect -913 298 -870 332
rect -990 264 -870 298
rect -990 230 -947 264
rect -913 230 -870 264
rect -990 196 -870 230
rect -990 162 -947 196
rect -913 162 -870 196
rect -990 128 -870 162
rect -990 94 -947 128
rect -913 94 -870 128
rect -990 60 -870 94
rect -770 876 -650 900
rect -770 842 -727 876
rect -693 842 -650 876
rect -770 808 -650 842
rect -770 774 -727 808
rect -693 774 -650 808
rect -770 740 -650 774
rect -770 706 -727 740
rect -693 706 -650 740
rect -770 672 -650 706
rect -770 638 -727 672
rect -693 638 -650 672
rect -770 604 -650 638
rect -770 570 -727 604
rect -693 570 -650 604
rect -770 536 -650 570
rect -770 502 -727 536
rect -693 502 -650 536
rect -770 468 -650 502
rect -770 434 -727 468
rect -693 434 -650 468
rect -770 400 -650 434
rect -770 366 -727 400
rect -693 366 -650 400
rect -770 332 -650 366
rect -770 298 -727 332
rect -693 298 -650 332
rect -770 264 -650 298
rect -770 230 -727 264
rect -693 230 -650 264
rect -770 196 -650 230
rect -770 162 -727 196
rect -693 162 -650 196
rect -770 128 -650 162
rect -770 94 -727 128
rect -693 94 -650 128
rect -770 60 -650 94
<< ndiffc >>
rect -1607 842 -1573 876
rect -1607 774 -1573 808
rect -1607 706 -1573 740
rect -1607 638 -1573 672
rect -1607 570 -1573 604
rect -1607 502 -1573 536
rect -1607 434 -1573 468
rect -1607 366 -1573 400
rect -1607 298 -1573 332
rect -1607 230 -1573 264
rect -1607 162 -1573 196
rect -1607 94 -1573 128
rect -1387 842 -1353 876
rect -1387 774 -1353 808
rect -1387 706 -1353 740
rect -1387 638 -1353 672
rect -1387 570 -1353 604
rect -1387 502 -1353 536
rect -1387 434 -1353 468
rect -1387 366 -1353 400
rect -1387 298 -1353 332
rect -1387 230 -1353 264
rect -1387 162 -1353 196
rect -1387 94 -1353 128
rect -1167 842 -1133 876
rect -1167 774 -1133 808
rect -1167 706 -1133 740
rect -1167 638 -1133 672
rect -1167 570 -1133 604
rect -1167 502 -1133 536
rect -1167 434 -1133 468
rect -1167 366 -1133 400
rect -1167 298 -1133 332
rect -1167 230 -1133 264
rect -1167 162 -1133 196
rect -1167 94 -1133 128
rect -947 842 -913 876
rect -947 774 -913 808
rect -947 706 -913 740
rect -947 638 -913 672
rect -947 570 -913 604
rect -947 502 -913 536
rect -947 434 -913 468
rect -947 366 -913 400
rect -947 298 -913 332
rect -947 230 -913 264
rect -947 162 -913 196
rect -947 94 -913 128
rect -727 842 -693 876
rect -727 774 -693 808
rect -727 706 -693 740
rect -727 638 -693 672
rect -727 570 -693 604
rect -727 502 -693 536
rect -727 434 -693 468
rect -727 366 -693 400
rect -727 298 -693 332
rect -727 230 -693 264
rect -727 162 -693 196
rect -727 94 -693 128
<< psubdiff >>
rect -1770 876 -1650 900
rect -1770 842 -1727 876
rect -1693 842 -1650 876
rect -1770 808 -1650 842
rect -1770 774 -1727 808
rect -1693 774 -1650 808
rect -1770 740 -1650 774
rect -1770 706 -1727 740
rect -1693 706 -1650 740
rect -1770 672 -1650 706
rect -1770 638 -1727 672
rect -1693 638 -1650 672
rect -1770 604 -1650 638
rect -1770 570 -1727 604
rect -1693 570 -1650 604
rect -1770 536 -1650 570
rect -1770 502 -1727 536
rect -1693 502 -1650 536
rect -1770 468 -1650 502
rect -1770 434 -1727 468
rect -1693 434 -1650 468
rect -1770 400 -1650 434
rect -1770 366 -1727 400
rect -1693 366 -1650 400
rect -1770 332 -1650 366
rect -1770 298 -1727 332
rect -1693 298 -1650 332
rect -1770 264 -1650 298
rect -1770 230 -1727 264
rect -1693 230 -1650 264
rect -1770 196 -1650 230
rect -1770 162 -1727 196
rect -1693 162 -1650 196
rect -1770 128 -1650 162
rect -1770 94 -1727 128
rect -1693 94 -1650 128
rect -1770 60 -1650 94
<< psubdiffcont >>
rect -1727 842 -1693 876
rect -1727 774 -1693 808
rect -1727 706 -1693 740
rect -1727 638 -1693 672
rect -1727 570 -1693 604
rect -1727 502 -1693 536
rect -1727 434 -1693 468
rect -1727 366 -1693 400
rect -1727 298 -1693 332
rect -1727 230 -1693 264
rect -1727 162 -1693 196
rect -1727 94 -1693 128
<< poly >>
rect -1530 950 -770 980
rect -1530 900 -1430 950
rect -1310 900 -1210 950
rect -1090 900 -990 950
rect -870 900 -770 950
rect -1530 30 -1430 60
rect -1310 30 -1210 60
rect -1090 30 -990 60
rect -870 30 -770 60
<< locali >>
rect -1390 920 -910 960
rect -1390 880 -1350 920
rect -950 880 -910 920
rect -1750 876 -1670 880
rect -1750 842 -1727 876
rect -1693 842 -1670 876
rect -1750 808 -1670 842
rect -1750 774 -1727 808
rect -1693 774 -1670 808
rect -1750 740 -1670 774
rect -1750 706 -1727 740
rect -1693 706 -1670 740
rect -1750 672 -1670 706
rect -1750 638 -1727 672
rect -1693 638 -1670 672
rect -1750 604 -1670 638
rect -1750 570 -1727 604
rect -1693 570 -1670 604
rect -1750 536 -1670 570
rect -1750 502 -1727 536
rect -1693 502 -1670 536
rect -1750 468 -1670 502
rect -1750 434 -1727 468
rect -1693 434 -1670 468
rect -1750 400 -1670 434
rect -1750 366 -1727 400
rect -1693 366 -1670 400
rect -1750 332 -1670 366
rect -1750 298 -1727 332
rect -1693 298 -1670 332
rect -1750 264 -1670 298
rect -1750 230 -1727 264
rect -1693 230 -1670 264
rect -1750 196 -1670 230
rect -1750 162 -1727 196
rect -1693 162 -1670 196
rect -1750 128 -1670 162
rect -1750 94 -1727 128
rect -1693 94 -1670 128
rect -1750 80 -1670 94
rect -1630 876 -1550 880
rect -1630 842 -1607 876
rect -1573 842 -1550 876
rect -1630 808 -1550 842
rect -1630 774 -1607 808
rect -1573 774 -1550 808
rect -1630 740 -1550 774
rect -1630 706 -1607 740
rect -1573 706 -1550 740
rect -1630 672 -1550 706
rect -1630 638 -1607 672
rect -1573 638 -1550 672
rect -1630 604 -1550 638
rect -1630 570 -1607 604
rect -1573 570 -1550 604
rect -1630 536 -1550 570
rect -1630 502 -1607 536
rect -1573 502 -1550 536
rect -1630 468 -1550 502
rect -1630 434 -1607 468
rect -1573 434 -1550 468
rect -1630 400 -1550 434
rect -1630 366 -1607 400
rect -1573 366 -1550 400
rect -1630 332 -1550 366
rect -1630 298 -1607 332
rect -1573 298 -1550 332
rect -1630 264 -1550 298
rect -1630 230 -1607 264
rect -1573 230 -1550 264
rect -1630 196 -1550 230
rect -1630 162 -1607 196
rect -1573 162 -1550 196
rect -1630 128 -1550 162
rect -1630 94 -1607 128
rect -1573 94 -1550 128
rect -1630 80 -1550 94
rect -1410 876 -1330 880
rect -1410 842 -1387 876
rect -1353 842 -1330 876
rect -1410 808 -1330 842
rect -1410 774 -1387 808
rect -1353 774 -1330 808
rect -1410 740 -1330 774
rect -1410 706 -1387 740
rect -1353 706 -1330 740
rect -1410 672 -1330 706
rect -1410 638 -1387 672
rect -1353 638 -1330 672
rect -1410 604 -1330 638
rect -1410 570 -1387 604
rect -1353 570 -1330 604
rect -1410 536 -1330 570
rect -1410 502 -1387 536
rect -1353 502 -1330 536
rect -1410 468 -1330 502
rect -1410 434 -1387 468
rect -1353 434 -1330 468
rect -1410 400 -1330 434
rect -1410 366 -1387 400
rect -1353 366 -1330 400
rect -1410 332 -1330 366
rect -1410 298 -1387 332
rect -1353 298 -1330 332
rect -1410 264 -1330 298
rect -1410 230 -1387 264
rect -1353 230 -1330 264
rect -1410 196 -1330 230
rect -1410 162 -1387 196
rect -1353 162 -1330 196
rect -1410 128 -1330 162
rect -1410 94 -1387 128
rect -1353 94 -1330 128
rect -1410 80 -1330 94
rect -1190 876 -1110 880
rect -1190 842 -1167 876
rect -1133 842 -1110 876
rect -1190 808 -1110 842
rect -1190 774 -1167 808
rect -1133 774 -1110 808
rect -1190 740 -1110 774
rect -1190 706 -1167 740
rect -1133 706 -1110 740
rect -1190 672 -1110 706
rect -1190 638 -1167 672
rect -1133 638 -1110 672
rect -1190 604 -1110 638
rect -1190 570 -1167 604
rect -1133 570 -1110 604
rect -1190 536 -1110 570
rect -1190 502 -1167 536
rect -1133 502 -1110 536
rect -1190 468 -1110 502
rect -1190 434 -1167 468
rect -1133 434 -1110 468
rect -1190 400 -1110 434
rect -1190 366 -1167 400
rect -1133 366 -1110 400
rect -1190 332 -1110 366
rect -1190 298 -1167 332
rect -1133 298 -1110 332
rect -1190 264 -1110 298
rect -1190 230 -1167 264
rect -1133 230 -1110 264
rect -1190 196 -1110 230
rect -1190 162 -1167 196
rect -1133 162 -1110 196
rect -1190 128 -1110 162
rect -1190 94 -1167 128
rect -1133 94 -1110 128
rect -1190 80 -1110 94
rect -970 876 -890 880
rect -970 842 -947 876
rect -913 842 -890 876
rect -970 808 -890 842
rect -970 774 -947 808
rect -913 774 -890 808
rect -970 740 -890 774
rect -970 706 -947 740
rect -913 706 -890 740
rect -970 672 -890 706
rect -970 638 -947 672
rect -913 638 -890 672
rect -970 604 -890 638
rect -970 570 -947 604
rect -913 570 -890 604
rect -970 536 -890 570
rect -970 502 -947 536
rect -913 502 -890 536
rect -970 468 -890 502
rect -970 434 -947 468
rect -913 434 -890 468
rect -970 400 -890 434
rect -970 366 -947 400
rect -913 366 -890 400
rect -970 332 -890 366
rect -970 298 -947 332
rect -913 298 -890 332
rect -970 264 -890 298
rect -970 230 -947 264
rect -913 230 -890 264
rect -970 196 -890 230
rect -970 162 -947 196
rect -913 162 -890 196
rect -970 128 -890 162
rect -970 94 -947 128
rect -913 94 -890 128
rect -970 80 -890 94
rect -750 876 -670 880
rect -750 842 -727 876
rect -693 842 -670 876
rect -750 808 -670 842
rect -750 774 -727 808
rect -693 774 -670 808
rect -750 740 -670 774
rect -750 706 -727 740
rect -693 706 -670 740
rect -750 672 -670 706
rect -750 638 -727 672
rect -693 638 -670 672
rect -750 604 -670 638
rect -750 570 -727 604
rect -693 570 -670 604
rect -750 536 -670 570
rect -750 502 -727 536
rect -693 502 -670 536
rect -750 468 -670 502
rect -750 434 -727 468
rect -693 434 -670 468
rect -750 400 -670 434
rect -750 366 -727 400
rect -693 366 -670 400
rect -750 332 -670 366
rect -750 298 -727 332
rect -693 298 -670 332
rect -750 264 -670 298
rect -750 230 -727 264
rect -693 230 -670 264
rect -750 196 -670 230
rect -750 162 -727 196
rect -693 162 -670 196
rect -750 128 -670 162
rect -750 94 -727 128
rect -693 94 -670 128
rect -750 80 -670 94
rect -1610 40 -1570 80
rect -1170 40 -1130 80
rect -730 40 -690 80
rect -1610 0 -690 40
<< end >>
