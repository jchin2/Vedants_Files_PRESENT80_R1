magic
tech sky130a
timestamp 1670961910
<< checkpaint >>
rect -9 -152 9 152
<< l67d20 >>
rect -9 -152 9 152
<< l67d13 >>
rect -9 -123 9 123
<< end >>
