* NGSPICE file created from EESPFAL_XOR_v3.ext - technology: sky130A

.subckt EESPFAL_XOR_v3 A A_bar B B_bar OUT OUT_bar Dis GND CLK
X0 CLK OUT OUT_bar CLK sky130_fd_pr__pfet_01v8 ad=2.7e+12p pd=1.26e+07u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u M=2
X1 OUT_bar Dis GND GND sky130_fd_pr__nfet_01v8 ad=2.7e+12p pd=1.26e+07u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X2 a_n840_410# A CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=7.5e+12p ps=3.22e+07u w=1.5e+06u l=150000u
X3 a_n1140_410# B_bar OUT_bar GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_420_410# B_bar OUT GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X5 GND Dis OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 OUT OUT_bar CLK CLK sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u M=2
X7 a_720_410# A_bar CLK GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 OUT_bar B a_n840_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 GND OUT OUT_bar GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 CLK A_bar a_n1140_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 OUT OUT_bar GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 CLK A a_420_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 OUT B a_720_410# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

