magic
tech sky130A
magscale 1 2
timestamp 1672691392
<< nwell >>
rect -2670 1540 -590 1730
rect -2040 1150 -1220 1540
<< pwell >>
rect -2646 526 -614 966
rect -2656 374 -604 526
<< nmos >>
rect -2500 640 -2470 940
rect -2350 640 -2320 940
rect -2200 640 -2170 940
rect -1870 640 -1840 940
rect -1720 640 -1690 940
rect -1570 640 -1540 940
rect -1420 640 -1390 940
rect -1090 640 -1060 940
rect -940 640 -910 940
rect -790 640 -760 940
<< pmos >>
rect -1870 1200 -1840 1500
rect -1720 1200 -1690 1500
rect -1570 1200 -1540 1500
rect -1420 1200 -1390 1500
<< ndiff >>
rect -2620 867 -2500 940
rect -2620 833 -2577 867
rect -2543 833 -2500 867
rect -2620 787 -2500 833
rect -2620 753 -2577 787
rect -2543 753 -2500 787
rect -2620 707 -2500 753
rect -2620 673 -2577 707
rect -2543 673 -2500 707
rect -2620 640 -2500 673
rect -2470 867 -2350 940
rect -2470 833 -2427 867
rect -2393 833 -2350 867
rect -2470 787 -2350 833
rect -2470 753 -2427 787
rect -2393 753 -2350 787
rect -2470 707 -2350 753
rect -2470 673 -2427 707
rect -2393 673 -2350 707
rect -2470 640 -2350 673
rect -2320 867 -2200 940
rect -2320 833 -2277 867
rect -2243 833 -2200 867
rect -2320 787 -2200 833
rect -2320 753 -2277 787
rect -2243 753 -2200 787
rect -2320 707 -2200 753
rect -2320 673 -2277 707
rect -2243 673 -2200 707
rect -2320 640 -2200 673
rect -2170 867 -2050 940
rect -2170 833 -2127 867
rect -2093 833 -2050 867
rect -2170 787 -2050 833
rect -2170 753 -2127 787
rect -2093 753 -2050 787
rect -2170 707 -2050 753
rect -2170 673 -2127 707
rect -2093 673 -2050 707
rect -2170 640 -2050 673
rect -1990 867 -1870 940
rect -1990 833 -1947 867
rect -1913 833 -1870 867
rect -1990 787 -1870 833
rect -1990 753 -1947 787
rect -1913 753 -1870 787
rect -1990 707 -1870 753
rect -1990 673 -1947 707
rect -1913 673 -1870 707
rect -1990 640 -1870 673
rect -1840 867 -1720 940
rect -1840 833 -1797 867
rect -1763 833 -1720 867
rect -1840 787 -1720 833
rect -1840 753 -1797 787
rect -1763 753 -1720 787
rect -1840 707 -1720 753
rect -1840 673 -1797 707
rect -1763 673 -1720 707
rect -1840 640 -1720 673
rect -1690 867 -1570 940
rect -1690 833 -1647 867
rect -1613 833 -1570 867
rect -1690 787 -1570 833
rect -1690 753 -1647 787
rect -1613 753 -1570 787
rect -1690 707 -1570 753
rect -1690 673 -1647 707
rect -1613 673 -1570 707
rect -1690 640 -1570 673
rect -1540 867 -1420 940
rect -1540 833 -1497 867
rect -1463 833 -1420 867
rect -1540 787 -1420 833
rect -1540 753 -1497 787
rect -1463 753 -1420 787
rect -1540 707 -1420 753
rect -1540 673 -1497 707
rect -1463 673 -1420 707
rect -1540 640 -1420 673
rect -1390 867 -1270 940
rect -1390 833 -1347 867
rect -1313 833 -1270 867
rect -1390 787 -1270 833
rect -1390 753 -1347 787
rect -1313 753 -1270 787
rect -1390 707 -1270 753
rect -1390 673 -1347 707
rect -1313 673 -1270 707
rect -1390 640 -1270 673
rect -1210 867 -1090 940
rect -1210 833 -1167 867
rect -1133 833 -1090 867
rect -1210 787 -1090 833
rect -1210 753 -1167 787
rect -1133 753 -1090 787
rect -1210 707 -1090 753
rect -1210 673 -1167 707
rect -1133 673 -1090 707
rect -1210 640 -1090 673
rect -1060 640 -940 940
rect -910 640 -790 940
rect -760 867 -640 940
rect -760 833 -717 867
rect -683 833 -640 867
rect -760 787 -640 833
rect -760 753 -717 787
rect -683 753 -640 787
rect -760 707 -640 753
rect -760 673 -717 707
rect -683 673 -640 707
rect -760 640 -640 673
<< pdiff >>
rect -1990 1427 -1870 1500
rect -1990 1393 -1947 1427
rect -1913 1393 -1870 1427
rect -1990 1347 -1870 1393
rect -1990 1313 -1947 1347
rect -1913 1313 -1870 1347
rect -1990 1267 -1870 1313
rect -1990 1233 -1947 1267
rect -1913 1233 -1870 1267
rect -1990 1200 -1870 1233
rect -1840 1427 -1720 1500
rect -1840 1393 -1797 1427
rect -1763 1393 -1720 1427
rect -1840 1347 -1720 1393
rect -1840 1313 -1797 1347
rect -1763 1313 -1720 1347
rect -1840 1267 -1720 1313
rect -1840 1233 -1797 1267
rect -1763 1233 -1720 1267
rect -1840 1200 -1720 1233
rect -1690 1427 -1570 1500
rect -1690 1393 -1647 1427
rect -1613 1393 -1570 1427
rect -1690 1347 -1570 1393
rect -1690 1313 -1647 1347
rect -1613 1313 -1570 1347
rect -1690 1267 -1570 1313
rect -1690 1233 -1647 1267
rect -1613 1233 -1570 1267
rect -1690 1200 -1570 1233
rect -1540 1427 -1420 1500
rect -1540 1393 -1497 1427
rect -1463 1393 -1420 1427
rect -1540 1347 -1420 1393
rect -1540 1313 -1497 1347
rect -1463 1313 -1420 1347
rect -1540 1267 -1420 1313
rect -1540 1233 -1497 1267
rect -1463 1233 -1420 1267
rect -1540 1200 -1420 1233
rect -1390 1427 -1270 1500
rect -1390 1393 -1347 1427
rect -1313 1393 -1270 1427
rect -1390 1347 -1270 1393
rect -1390 1313 -1347 1347
rect -1313 1313 -1270 1347
rect -1390 1267 -1270 1313
rect -1390 1233 -1347 1267
rect -1313 1233 -1270 1267
rect -1390 1200 -1270 1233
<< ndiffc >>
rect -2577 833 -2543 867
rect -2577 753 -2543 787
rect -2577 673 -2543 707
rect -2427 833 -2393 867
rect -2427 753 -2393 787
rect -2427 673 -2393 707
rect -2277 833 -2243 867
rect -2277 753 -2243 787
rect -2277 673 -2243 707
rect -2127 833 -2093 867
rect -2127 753 -2093 787
rect -2127 673 -2093 707
rect -1947 833 -1913 867
rect -1947 753 -1913 787
rect -1947 673 -1913 707
rect -1797 833 -1763 867
rect -1797 753 -1763 787
rect -1797 673 -1763 707
rect -1647 833 -1613 867
rect -1647 753 -1613 787
rect -1647 673 -1613 707
rect -1497 833 -1463 867
rect -1497 753 -1463 787
rect -1497 673 -1463 707
rect -1347 833 -1313 867
rect -1347 753 -1313 787
rect -1347 673 -1313 707
rect -1167 833 -1133 867
rect -1167 753 -1133 787
rect -1167 673 -1133 707
rect -717 833 -683 867
rect -717 753 -683 787
rect -717 673 -683 707
<< pdiffc >>
rect -1947 1393 -1913 1427
rect -1947 1313 -1913 1347
rect -1947 1233 -1913 1267
rect -1797 1393 -1763 1427
rect -1797 1313 -1763 1347
rect -1797 1233 -1763 1267
rect -1647 1393 -1613 1427
rect -1647 1313 -1613 1347
rect -1647 1233 -1613 1267
rect -1497 1393 -1463 1427
rect -1497 1313 -1463 1347
rect -1497 1233 -1463 1267
rect -1347 1393 -1313 1427
rect -1347 1313 -1313 1347
rect -1347 1233 -1313 1267
<< psubdiff >>
rect -2630 467 -630 500
rect -2630 433 -2607 467
rect -2573 433 -2527 467
rect -2493 433 -2447 467
rect -2413 433 -2367 467
rect -2333 433 -2287 467
rect -2253 433 -2207 467
rect -2173 433 -2127 467
rect -2093 433 -2047 467
rect -2013 433 -1967 467
rect -1933 433 -1887 467
rect -1853 433 -1807 467
rect -1773 433 -1727 467
rect -1693 433 -1647 467
rect -1613 433 -1567 467
rect -1533 433 -1487 467
rect -1453 433 -1407 467
rect -1373 433 -1327 467
rect -1293 433 -1247 467
rect -1213 433 -1167 467
rect -1133 433 -1087 467
rect -1053 433 -1007 467
rect -973 433 -927 467
rect -893 433 -847 467
rect -813 433 -767 467
rect -733 433 -687 467
rect -653 433 -630 467
rect -2630 400 -630 433
<< nsubdiff >>
rect -2630 1647 -630 1680
rect -2630 1613 -2607 1647
rect -2573 1613 -2527 1647
rect -2493 1613 -2447 1647
rect -2413 1613 -2367 1647
rect -2333 1613 -2287 1647
rect -2253 1613 -2207 1647
rect -2173 1613 -2127 1647
rect -2093 1613 -2047 1647
rect -2013 1613 -1967 1647
rect -1933 1613 -1887 1647
rect -1853 1613 -1807 1647
rect -1773 1613 -1727 1647
rect -1693 1613 -1647 1647
rect -1613 1613 -1567 1647
rect -1533 1613 -1487 1647
rect -1453 1613 -1407 1647
rect -1373 1613 -1327 1647
rect -1293 1613 -1247 1647
rect -1213 1613 -1167 1647
rect -1133 1613 -1087 1647
rect -1053 1613 -1007 1647
rect -973 1613 -927 1647
rect -893 1613 -847 1647
rect -813 1613 -767 1647
rect -733 1613 -687 1647
rect -653 1613 -630 1647
rect -2630 1580 -630 1613
<< psubdiffcont >>
rect -2607 433 -2573 467
rect -2527 433 -2493 467
rect -2447 433 -2413 467
rect -2367 433 -2333 467
rect -2287 433 -2253 467
rect -2207 433 -2173 467
rect -2127 433 -2093 467
rect -2047 433 -2013 467
rect -1967 433 -1933 467
rect -1887 433 -1853 467
rect -1807 433 -1773 467
rect -1727 433 -1693 467
rect -1647 433 -1613 467
rect -1567 433 -1533 467
rect -1487 433 -1453 467
rect -1407 433 -1373 467
rect -1327 433 -1293 467
rect -1247 433 -1213 467
rect -1167 433 -1133 467
rect -1087 433 -1053 467
rect -1007 433 -973 467
rect -927 433 -893 467
rect -847 433 -813 467
rect -767 433 -733 467
rect -687 433 -653 467
<< nsubdiffcont >>
rect -2607 1613 -2573 1647
rect -2527 1613 -2493 1647
rect -2447 1613 -2413 1647
rect -2367 1613 -2333 1647
rect -2287 1613 -2253 1647
rect -2207 1613 -2173 1647
rect -2127 1613 -2093 1647
rect -2047 1613 -2013 1647
rect -1967 1613 -1933 1647
rect -1887 1613 -1853 1647
rect -1807 1613 -1773 1647
rect -1727 1613 -1693 1647
rect -1647 1613 -1613 1647
rect -1567 1613 -1533 1647
rect -1487 1613 -1453 1647
rect -1407 1613 -1373 1647
rect -1327 1613 -1293 1647
rect -1247 1613 -1213 1647
rect -1167 1613 -1133 1647
rect -1087 1613 -1053 1647
rect -1007 1613 -973 1647
rect -927 1613 -893 1647
rect -847 1613 -813 1647
rect -767 1613 -733 1647
rect -687 1613 -653 1647
<< poly >>
rect -1870 1530 -1690 1560
rect -1870 1500 -1840 1530
rect -1720 1500 -1690 1530
rect -1570 1530 -1390 1560
rect -1570 1500 -1540 1530
rect -1420 1500 -1390 1530
rect -840 1527 -760 1550
rect -840 1493 -817 1527
rect -783 1493 -760 1527
rect -840 1470 -760 1493
rect -990 1407 -910 1430
rect -990 1373 -967 1407
rect -933 1373 -910 1407
rect -990 1350 -910 1373
rect -1120 1287 -1040 1310
rect -1120 1253 -1097 1287
rect -1063 1253 -1040 1287
rect -1120 1230 -1040 1253
rect -1870 1170 -1840 1200
rect -2420 1117 -2320 1140
rect -2420 1083 -2397 1117
rect -2363 1083 -2320 1117
rect -2420 1060 -2320 1083
rect -2250 1137 -2170 1160
rect -2250 1103 -2227 1137
rect -2193 1103 -2170 1137
rect -2250 1080 -2170 1103
rect -2550 1037 -2470 1060
rect -2550 1003 -2527 1037
rect -2493 1003 -2470 1037
rect -2550 980 -2470 1003
rect -2500 940 -2470 980
rect -2350 940 -2320 1060
rect -2200 940 -2170 1080
rect -1720 1045 -1690 1200
rect -1570 1170 -1540 1200
rect -1420 1170 -1390 1200
rect -1620 1147 -1540 1170
rect -1620 1113 -1597 1147
rect -1563 1113 -1540 1147
rect -1620 1090 -1540 1113
rect -1720 1022 -1640 1045
rect -1720 988 -1697 1022
rect -1663 988 -1640 1022
rect -1870 940 -1840 970
rect -1720 965 -1640 988
rect -1720 940 -1690 965
rect -1570 940 -1540 1090
rect -1420 940 -1390 970
rect -1090 940 -1060 1230
rect -940 940 -910 1350
rect -790 940 -760 1470
rect -2500 610 -2470 640
rect -2350 610 -2320 640
rect -2200 610 -2170 640
rect -1870 610 -1840 640
rect -1720 610 -1690 640
rect -1570 610 -1540 640
rect -1420 610 -1390 640
rect -1090 610 -1060 640
rect -940 610 -910 640
rect -790 610 -760 640
rect -1870 587 -1790 610
rect -1870 553 -1847 587
rect -1813 553 -1790 587
rect -1870 530 -1790 553
rect -1470 587 -1390 610
rect -1470 553 -1447 587
rect -1413 553 -1390 587
rect -1470 530 -1390 553
<< polycont >>
rect -817 1493 -783 1527
rect -967 1373 -933 1407
rect -1097 1253 -1063 1287
rect -2397 1083 -2363 1117
rect -2227 1103 -2193 1137
rect -2527 1003 -2493 1037
rect -1597 1113 -1563 1147
rect -1697 988 -1663 1022
rect -1847 553 -1813 587
rect -1447 553 -1413 587
<< locali >>
rect -2630 1647 -630 1670
rect -2630 1613 -2607 1647
rect -2573 1613 -2527 1647
rect -2493 1613 -2447 1647
rect -2413 1613 -2367 1647
rect -2333 1613 -2287 1647
rect -2253 1613 -2207 1647
rect -2173 1613 -2127 1647
rect -2093 1613 -2047 1647
rect -2013 1613 -1967 1647
rect -1933 1613 -1887 1647
rect -1853 1613 -1807 1647
rect -1773 1613 -1727 1647
rect -1693 1613 -1647 1647
rect -1613 1613 -1567 1647
rect -1533 1613 -1487 1647
rect -1453 1613 -1407 1647
rect -1373 1613 -1327 1647
rect -1293 1613 -1247 1647
rect -1213 1613 -1167 1647
rect -1133 1613 -1087 1647
rect -1053 1613 -1007 1647
rect -973 1613 -927 1647
rect -893 1613 -847 1647
rect -813 1613 -767 1647
rect -733 1613 -687 1647
rect -653 1613 -630 1647
rect -2630 1590 -630 1613
rect -2210 1530 -2130 1550
rect -2620 1527 -2130 1530
rect -2620 1493 -2187 1527
rect -2153 1493 -2130 1527
rect -2620 1490 -2130 1493
rect -2210 1470 -2130 1490
rect -840 1527 -760 1550
rect -840 1493 -817 1527
rect -783 1493 -760 1527
rect -840 1470 -760 1493
rect -2120 1410 -2040 1430
rect -2620 1407 -2040 1410
rect -2620 1373 -2097 1407
rect -2063 1373 -2040 1407
rect -2620 1370 -2040 1373
rect -2120 1350 -2040 1370
rect -1970 1427 -1890 1460
rect -1970 1393 -1947 1427
rect -1913 1393 -1890 1427
rect -1970 1347 -1890 1393
rect -1970 1313 -1947 1347
rect -1913 1313 -1890 1347
rect -2150 1300 -2070 1310
rect -2620 1287 -2070 1300
rect -2620 1260 -2127 1287
rect -2150 1253 -2127 1260
rect -2093 1253 -2070 1287
rect -2150 1230 -2070 1253
rect -1970 1267 -1890 1313
rect -1970 1233 -1947 1267
rect -1913 1233 -1890 1267
rect -2620 1180 -2190 1220
rect -1970 1210 -1890 1233
rect -1820 1427 -1740 1460
rect -1820 1393 -1797 1427
rect -1763 1393 -1740 1427
rect -1820 1347 -1740 1393
rect -1820 1313 -1797 1347
rect -1763 1313 -1740 1347
rect -1820 1267 -1740 1313
rect -1820 1233 -1797 1267
rect -1763 1233 -1740 1267
rect -1820 1200 -1740 1233
rect -1670 1427 -1590 1460
rect -1670 1393 -1647 1427
rect -1613 1393 -1590 1427
rect -1670 1347 -1590 1393
rect -1670 1313 -1647 1347
rect -1613 1313 -1590 1347
rect -1670 1267 -1590 1313
rect -1670 1233 -1647 1267
rect -1613 1233 -1590 1267
rect -1670 1210 -1590 1233
rect -1520 1427 -1440 1460
rect -1520 1393 -1497 1427
rect -1463 1393 -1440 1427
rect -1520 1347 -1440 1393
rect -1520 1313 -1497 1347
rect -1463 1313 -1440 1347
rect -1520 1267 -1440 1313
rect -1520 1233 -1497 1267
rect -1463 1233 -1440 1267
rect -1520 1200 -1440 1233
rect -1370 1427 -1290 1460
rect -1370 1393 -1347 1427
rect -1313 1393 -1290 1427
rect -1370 1347 -1290 1393
rect -990 1407 -910 1430
rect -990 1373 -967 1407
rect -933 1373 -910 1407
rect -990 1350 -910 1373
rect -1370 1313 -1347 1347
rect -1313 1313 -1290 1347
rect -1370 1267 -1290 1313
rect -1370 1233 -1347 1267
rect -1313 1233 -1290 1267
rect -1370 1210 -1290 1233
rect -1120 1287 -1040 1310
rect -1120 1253 -1097 1287
rect -1063 1253 -1040 1287
rect -1120 1230 -1040 1253
rect -2250 1160 -2190 1180
rect -2620 1117 -2340 1140
rect -2620 1100 -2397 1117
rect -2420 1083 -2397 1100
rect -2363 1083 -2340 1117
rect -2420 1060 -2340 1083
rect -2250 1137 -2170 1160
rect -2250 1103 -2227 1137
rect -2193 1103 -2170 1137
rect -2250 1080 -2170 1103
rect -1800 1150 -1760 1200
rect -1620 1150 -1540 1170
rect -1800 1147 -1540 1150
rect -1800 1113 -1597 1147
rect -1563 1113 -1540 1147
rect -1800 1110 -1540 1113
rect -2550 1040 -2470 1060
rect -2620 1037 -2470 1040
rect -2620 1003 -2527 1037
rect -2493 1003 -2470 1037
rect -2620 1000 -2470 1003
rect -2550 980 -2470 1000
rect -1800 980 -1760 1110
rect -1620 1090 -1540 1110
rect -2430 940 -1760 980
rect -1720 1030 -1640 1045
rect -1500 1030 -1460 1200
rect -1220 1150 -1140 1170
rect -1220 1147 -640 1150
rect -1220 1113 -1197 1147
rect -1163 1113 -640 1147
rect -1220 1110 -640 1113
rect -1220 1090 -1140 1110
rect -1720 1022 -640 1030
rect -1720 988 -1697 1022
rect -1663 990 -640 1022
rect -1663 988 -1640 990
rect -1720 965 -1640 988
rect -2430 900 -2390 940
rect -2130 900 -2090 940
rect -1800 900 -1760 940
rect -1500 900 -1460 990
rect -1170 900 -1130 990
rect -2600 867 -2520 900
rect -2600 833 -2577 867
rect -2543 833 -2520 867
rect -2600 787 -2520 833
rect -2600 753 -2577 787
rect -2543 753 -2520 787
rect -2600 707 -2520 753
rect -2600 673 -2577 707
rect -2543 673 -2520 707
rect -2600 650 -2520 673
rect -2450 867 -2370 900
rect -2450 833 -2427 867
rect -2393 833 -2370 867
rect -2450 787 -2370 833
rect -2450 753 -2427 787
rect -2393 753 -2370 787
rect -2450 707 -2370 753
rect -2450 673 -2427 707
rect -2393 673 -2370 707
rect -2450 650 -2370 673
rect -2300 867 -2220 900
rect -2300 833 -2277 867
rect -2243 833 -2220 867
rect -2300 787 -2220 833
rect -2300 753 -2277 787
rect -2243 753 -2220 787
rect -2300 707 -2220 753
rect -2300 673 -2277 707
rect -2243 673 -2220 707
rect -2300 650 -2220 673
rect -2150 867 -2070 900
rect -2150 833 -2127 867
rect -2093 833 -2070 867
rect -2150 787 -2070 833
rect -2150 753 -2127 787
rect -2093 753 -2070 787
rect -2150 707 -2070 753
rect -2150 673 -2127 707
rect -2093 673 -2070 707
rect -2150 650 -2070 673
rect -1970 867 -1890 900
rect -1970 833 -1947 867
rect -1913 833 -1890 867
rect -1970 787 -1890 833
rect -1970 753 -1947 787
rect -1913 753 -1890 787
rect -1970 707 -1890 753
rect -1970 673 -1947 707
rect -1913 673 -1890 707
rect -1970 650 -1890 673
rect -1820 867 -1740 900
rect -1820 833 -1797 867
rect -1763 833 -1740 867
rect -1820 787 -1740 833
rect -1820 753 -1797 787
rect -1763 753 -1740 787
rect -1820 707 -1740 753
rect -1820 673 -1797 707
rect -1763 673 -1740 707
rect -1820 650 -1740 673
rect -1670 867 -1590 900
rect -1670 833 -1647 867
rect -1613 833 -1590 867
rect -1670 787 -1590 833
rect -1670 753 -1647 787
rect -1613 753 -1590 787
rect -1670 707 -1590 753
rect -1670 673 -1647 707
rect -1613 673 -1590 707
rect -1670 650 -1590 673
rect -1520 867 -1440 900
rect -1520 833 -1497 867
rect -1463 833 -1440 867
rect -1520 787 -1440 833
rect -1520 753 -1497 787
rect -1463 753 -1440 787
rect -1520 707 -1440 753
rect -1520 673 -1497 707
rect -1463 673 -1440 707
rect -1520 650 -1440 673
rect -1370 867 -1290 900
rect -1370 833 -1347 867
rect -1313 833 -1290 867
rect -1370 787 -1290 833
rect -1370 753 -1347 787
rect -1313 753 -1290 787
rect -1370 707 -1290 753
rect -1370 673 -1347 707
rect -1313 673 -1290 707
rect -1370 650 -1290 673
rect -1190 867 -1110 900
rect -1190 833 -1167 867
rect -1133 833 -1110 867
rect -1190 787 -1110 833
rect -1190 753 -1167 787
rect -1133 753 -1110 787
rect -1190 707 -1110 753
rect -1190 673 -1167 707
rect -1133 673 -1110 707
rect -1190 650 -1110 673
rect -740 867 -660 900
rect -740 833 -717 867
rect -683 833 -660 867
rect -740 787 -660 833
rect -740 753 -717 787
rect -683 753 -660 787
rect -740 707 -660 753
rect -740 673 -717 707
rect -683 673 -660 707
rect -740 650 -660 673
rect -1870 590 -1790 610
rect -1470 590 -1390 610
rect -2620 587 -1390 590
rect -2620 553 -1847 587
rect -1813 553 -1447 587
rect -1413 553 -1390 587
rect -2620 550 -1390 553
rect -1870 530 -1790 550
rect -1470 530 -1390 550
rect -2630 467 -630 490
rect -2630 433 -2607 467
rect -2573 433 -2527 467
rect -2493 433 -2447 467
rect -2413 433 -2367 467
rect -2333 433 -2287 467
rect -2253 433 -2207 467
rect -2173 433 -2127 467
rect -2093 433 -2047 467
rect -2013 433 -1967 467
rect -1933 433 -1887 467
rect -1853 433 -1807 467
rect -1773 433 -1727 467
rect -1693 433 -1647 467
rect -1613 433 -1567 467
rect -1533 433 -1487 467
rect -1453 433 -1407 467
rect -1373 433 -1327 467
rect -1293 433 -1247 467
rect -1213 433 -1167 467
rect -1133 433 -1087 467
rect -1053 433 -1007 467
rect -973 433 -927 467
rect -893 433 -847 467
rect -813 433 -767 467
rect -733 433 -687 467
rect -653 433 -630 467
rect -2630 410 -630 433
<< viali >>
rect -2607 1613 -2573 1647
rect -2527 1613 -2493 1647
rect -2447 1613 -2413 1647
rect -2367 1613 -2333 1647
rect -2287 1613 -2253 1647
rect -2207 1613 -2173 1647
rect -2127 1613 -2093 1647
rect -2047 1613 -2013 1647
rect -1967 1613 -1933 1647
rect -1887 1613 -1853 1647
rect -1807 1613 -1773 1647
rect -1727 1613 -1693 1647
rect -1647 1613 -1613 1647
rect -1567 1613 -1533 1647
rect -1487 1613 -1453 1647
rect -1407 1613 -1373 1647
rect -1327 1613 -1293 1647
rect -1247 1613 -1213 1647
rect -1167 1613 -1133 1647
rect -1087 1613 -1053 1647
rect -1007 1613 -973 1647
rect -927 1613 -893 1647
rect -847 1613 -813 1647
rect -767 1613 -733 1647
rect -687 1613 -653 1647
rect -2187 1493 -2153 1527
rect -817 1493 -783 1527
rect -2097 1373 -2063 1407
rect -1947 1393 -1913 1427
rect -1947 1313 -1913 1347
rect -2127 1253 -2093 1287
rect -1947 1233 -1913 1267
rect -1647 1393 -1613 1427
rect -1647 1313 -1613 1347
rect -1647 1233 -1613 1267
rect -1347 1393 -1313 1427
rect -967 1373 -933 1407
rect -1347 1313 -1313 1347
rect -1347 1233 -1313 1267
rect -1097 1253 -1063 1287
rect -1597 1113 -1563 1147
rect -1197 1113 -1163 1147
rect -2577 833 -2543 867
rect -2577 753 -2543 787
rect -2577 673 -2543 707
rect -2277 833 -2243 867
rect -2277 753 -2243 787
rect -2277 673 -2243 707
rect -1947 833 -1913 867
rect -1947 753 -1913 787
rect -1947 673 -1913 707
rect -1647 833 -1613 867
rect -1647 753 -1613 787
rect -1647 673 -1613 707
rect -1347 833 -1313 867
rect -1347 753 -1313 787
rect -1347 673 -1313 707
rect -717 833 -683 867
rect -717 753 -683 787
rect -717 673 -683 707
rect -2607 433 -2573 467
rect -2527 433 -2493 467
rect -2447 433 -2413 467
rect -2367 433 -2333 467
rect -2287 433 -2253 467
rect -2207 433 -2173 467
rect -2127 433 -2093 467
rect -2047 433 -2013 467
rect -1967 433 -1933 467
rect -1887 433 -1853 467
rect -1807 433 -1773 467
rect -1727 433 -1693 467
rect -1647 433 -1613 467
rect -1567 433 -1533 467
rect -1487 433 -1453 467
rect -1407 433 -1373 467
rect -1327 433 -1293 467
rect -1247 433 -1213 467
rect -1167 433 -1133 467
rect -1087 433 -1053 467
rect -1007 433 -973 467
rect -927 433 -893 467
rect -847 433 -813 467
rect -767 433 -733 467
rect -687 433 -653 467
<< metal1 >>
rect -2630 1647 -630 1680
rect -2630 1613 -2607 1647
rect -2573 1613 -2527 1647
rect -2493 1613 -2447 1647
rect -2413 1613 -2367 1647
rect -2333 1613 -2287 1647
rect -2253 1613 -2207 1647
rect -2173 1613 -2127 1647
rect -2093 1613 -2047 1647
rect -2013 1613 -1967 1647
rect -1933 1613 -1887 1647
rect -1853 1613 -1807 1647
rect -1773 1613 -1727 1647
rect -1693 1613 -1647 1647
rect -1613 1613 -1567 1647
rect -1533 1613 -1487 1647
rect -1453 1613 -1407 1647
rect -1373 1613 -1327 1647
rect -1293 1613 -1247 1647
rect -1213 1613 -1167 1647
rect -1133 1613 -1087 1647
rect -1053 1613 -1007 1647
rect -973 1613 -927 1647
rect -893 1613 -847 1647
rect -813 1613 -767 1647
rect -733 1613 -687 1647
rect -653 1613 -630 1647
rect -2630 1580 -630 1613
rect -2580 900 -2540 1580
rect -2280 900 -2240 1580
rect -2210 1536 -2130 1550
rect -2210 1484 -2196 1536
rect -2144 1484 -2130 1536
rect -2210 1470 -2130 1484
rect -2120 1416 -2040 1430
rect -2120 1364 -2106 1416
rect -2054 1364 -2040 1416
rect -2120 1350 -2040 1364
rect -1970 1427 -1890 1580
rect -1970 1393 -1947 1427
rect -1913 1393 -1890 1427
rect -1970 1347 -1890 1393
rect -1970 1313 -1947 1347
rect -1913 1313 -1890 1347
rect -2150 1296 -2070 1310
rect -2150 1244 -2136 1296
rect -2084 1244 -2070 1296
rect -2150 1230 -2070 1244
rect -1970 1267 -1890 1313
rect -1970 1233 -1947 1267
rect -1913 1233 -1890 1267
rect -1970 1210 -1890 1233
rect -1670 1427 -1590 1580
rect -1670 1393 -1647 1427
rect -1613 1393 -1590 1427
rect -1670 1347 -1590 1393
rect -1670 1313 -1647 1347
rect -1613 1313 -1590 1347
rect -1670 1267 -1590 1313
rect -1670 1233 -1647 1267
rect -1613 1233 -1590 1267
rect -1670 1210 -1590 1233
rect -1370 1427 -1290 1580
rect -840 1536 -760 1550
rect -840 1484 -826 1536
rect -774 1484 -760 1536
rect -840 1470 -760 1484
rect -1370 1393 -1347 1427
rect -1313 1393 -1290 1427
rect -1370 1347 -1290 1393
rect -990 1416 -910 1430
rect -990 1364 -976 1416
rect -924 1364 -910 1416
rect -990 1350 -910 1364
rect -1370 1313 -1347 1347
rect -1313 1313 -1290 1347
rect -1370 1267 -1290 1313
rect -1370 1233 -1347 1267
rect -1313 1233 -1290 1267
rect -1370 1210 -1290 1233
rect -1120 1296 -1040 1310
rect -1120 1244 -1106 1296
rect -1054 1244 -1040 1296
rect -1120 1230 -1040 1244
rect -1620 1150 -1540 1170
rect -1220 1150 -1140 1170
rect -1620 1147 -1140 1150
rect -1620 1113 -1597 1147
rect -1563 1113 -1197 1147
rect -1163 1113 -1140 1147
rect -1620 1110 -1140 1113
rect -1620 1090 -1540 1110
rect -1220 1090 -1140 1110
rect -720 900 -680 1580
rect -2600 867 -2520 900
rect -2600 833 -2577 867
rect -2543 833 -2520 867
rect -2600 787 -2520 833
rect -2600 753 -2577 787
rect -2543 753 -2520 787
rect -2600 707 -2520 753
rect -2600 673 -2577 707
rect -2543 673 -2520 707
rect -2600 650 -2520 673
rect -2300 867 -2220 900
rect -2300 833 -2277 867
rect -2243 833 -2220 867
rect -2300 787 -2220 833
rect -2300 753 -2277 787
rect -2243 753 -2220 787
rect -2300 707 -2220 753
rect -2300 673 -2277 707
rect -2243 673 -2220 707
rect -2300 650 -2220 673
rect -1970 867 -1890 900
rect -1970 833 -1947 867
rect -1913 833 -1890 867
rect -1970 787 -1890 833
rect -1970 753 -1947 787
rect -1913 753 -1890 787
rect -1970 707 -1890 753
rect -1970 673 -1947 707
rect -1913 673 -1890 707
rect -1970 650 -1890 673
rect -1670 867 -1590 900
rect -1670 833 -1647 867
rect -1613 833 -1590 867
rect -1670 787 -1590 833
rect -1670 753 -1647 787
rect -1613 753 -1590 787
rect -1670 707 -1590 753
rect -1670 673 -1647 707
rect -1613 673 -1590 707
rect -1670 650 -1590 673
rect -1370 867 -1290 900
rect -1370 833 -1347 867
rect -1313 833 -1290 867
rect -1370 787 -1290 833
rect -1370 753 -1347 787
rect -1313 753 -1290 787
rect -1370 707 -1290 753
rect -1370 673 -1347 707
rect -1313 673 -1290 707
rect -1370 650 -1290 673
rect -740 867 -660 900
rect -740 833 -717 867
rect -683 833 -660 867
rect -740 787 -660 833
rect -740 753 -717 787
rect -683 753 -660 787
rect -740 707 -660 753
rect -740 673 -717 707
rect -683 673 -660 707
rect -740 650 -660 673
rect -1950 500 -1910 650
rect -1650 500 -1610 650
rect -1350 500 -1310 650
rect -2630 467 -630 500
rect -2630 433 -2607 467
rect -2573 433 -2527 467
rect -2493 433 -2447 467
rect -2413 433 -2367 467
rect -2333 433 -2287 467
rect -2253 433 -2207 467
rect -2173 433 -2127 467
rect -2093 433 -2047 467
rect -2013 433 -1967 467
rect -1933 433 -1887 467
rect -1853 433 -1807 467
rect -1773 433 -1727 467
rect -1693 433 -1647 467
rect -1613 433 -1567 467
rect -1533 433 -1487 467
rect -1453 433 -1407 467
rect -1373 433 -1327 467
rect -1293 433 -1247 467
rect -1213 433 -1167 467
rect -1133 433 -1087 467
rect -1053 433 -1007 467
rect -973 433 -927 467
rect -893 433 -847 467
rect -813 433 -767 467
rect -733 433 -687 467
rect -653 433 -630 467
rect -2630 400 -630 433
<< via1 >>
rect -2196 1527 -2144 1536
rect -2196 1493 -2187 1527
rect -2187 1493 -2153 1527
rect -2153 1493 -2144 1527
rect -2196 1484 -2144 1493
rect -2106 1407 -2054 1416
rect -2106 1373 -2097 1407
rect -2097 1373 -2063 1407
rect -2063 1373 -2054 1407
rect -2106 1364 -2054 1373
rect -2136 1287 -2084 1296
rect -2136 1253 -2127 1287
rect -2127 1253 -2093 1287
rect -2093 1253 -2084 1287
rect -2136 1244 -2084 1253
rect -826 1527 -774 1536
rect -826 1493 -817 1527
rect -817 1493 -783 1527
rect -783 1493 -774 1527
rect -826 1484 -774 1493
rect -976 1407 -924 1416
rect -976 1373 -967 1407
rect -967 1373 -933 1407
rect -933 1373 -924 1407
rect -976 1364 -924 1373
rect -1106 1287 -1054 1296
rect -1106 1253 -1097 1287
rect -1097 1253 -1063 1287
rect -1063 1253 -1054 1287
rect -1106 1244 -1054 1253
<< metal2 >>
rect -2210 1536 -2130 1550
rect -2210 1484 -2196 1536
rect -2144 1530 -2130 1536
rect -840 1536 -760 1550
rect -840 1530 -826 1536
rect -2144 1490 -826 1530
rect -2144 1484 -2130 1490
rect -2210 1470 -2130 1484
rect -840 1484 -826 1490
rect -774 1484 -760 1536
rect -840 1470 -760 1484
rect -2120 1416 -2040 1430
rect -2120 1364 -2106 1416
rect -2054 1410 -2040 1416
rect -990 1416 -910 1430
rect -990 1410 -976 1416
rect -2054 1370 -976 1410
rect -2054 1364 -2040 1370
rect -2120 1350 -2040 1364
rect -990 1364 -976 1370
rect -924 1364 -910 1416
rect -990 1350 -910 1364
rect -2150 1296 -2070 1310
rect -2150 1244 -2136 1296
rect -2084 1290 -2070 1296
rect -1120 1296 -1040 1310
rect -1120 1290 -1106 1296
rect -2084 1250 -1106 1290
rect -2084 1244 -2070 1250
rect -2150 1230 -2070 1244
rect -1120 1244 -1106 1250
rect -1054 1244 -1040 1296
rect -1120 1230 -1040 1244
<< labels >>
rlabel locali s -1700 985 -1660 1025 4 OUT
port 1 nsew
rlabel locali s -2610 1500 -2590 1520 4 A
port 2 nsew
rlabel locali s -2610 1190 -2590 1210 4 A_bar
port 3 nsew
rlabel locali s -2610 1380 -2590 1400 4 B
port 4 nsew
rlabel locali s -2610 1110 -2590 1130 4 B_bar
port 5 nsew
rlabel locali s -2610 1270 -2590 1290 4 C
port 6 nsew
rlabel locali s -2610 1010 -2590 1030 4 C_bar
port 7 nsew
rlabel locali s -1850 550 -1810 590 4 Dis
port 8 nsew
rlabel metal1 s -1600 1110 -1560 1150 4 OUT_bar
port 9 nsew
rlabel metal1 s -1650 430 -1610 470 4 GND!
port 10 nsew
rlabel metal1 s -1650 1610 -1610 1650 4 CLK
port 11 nsew
<< properties >>
string path -7.400 4.500 -7.400 4.700 
<< end >>
