magic
tech sky130A
magscale 1 2
timestamp 1671041739
<< nwell >>
rect -240 170 1180 1430
<< pmoslvt >>
rect 90 380 190 1220
rect 310 380 410 1220
rect 530 380 630 1220
rect 750 380 850 1220
<< pdiff >>
rect -30 1186 90 1220
rect -30 1152 13 1186
rect 47 1152 90 1186
rect -30 1118 90 1152
rect -30 1084 13 1118
rect 47 1084 90 1118
rect -30 1050 90 1084
rect -30 1016 13 1050
rect 47 1016 90 1050
rect -30 982 90 1016
rect -30 948 13 982
rect 47 948 90 982
rect -30 914 90 948
rect -30 880 13 914
rect 47 880 90 914
rect -30 846 90 880
rect -30 812 13 846
rect 47 812 90 846
rect -30 778 90 812
rect -30 744 13 778
rect 47 744 90 778
rect -30 710 90 744
rect -30 676 13 710
rect 47 676 90 710
rect -30 642 90 676
rect -30 608 13 642
rect 47 608 90 642
rect -30 574 90 608
rect -30 540 13 574
rect 47 540 90 574
rect -30 506 90 540
rect -30 472 13 506
rect 47 472 90 506
rect -30 438 90 472
rect -30 404 13 438
rect 47 404 90 438
rect -30 380 90 404
rect 190 1186 310 1220
rect 190 1152 233 1186
rect 267 1152 310 1186
rect 190 1118 310 1152
rect 190 1084 233 1118
rect 267 1084 310 1118
rect 190 1050 310 1084
rect 190 1016 233 1050
rect 267 1016 310 1050
rect 190 982 310 1016
rect 190 948 233 982
rect 267 948 310 982
rect 190 914 310 948
rect 190 880 233 914
rect 267 880 310 914
rect 190 846 310 880
rect 190 812 233 846
rect 267 812 310 846
rect 190 778 310 812
rect 190 744 233 778
rect 267 744 310 778
rect 190 710 310 744
rect 190 676 233 710
rect 267 676 310 710
rect 190 642 310 676
rect 190 608 233 642
rect 267 608 310 642
rect 190 574 310 608
rect 190 540 233 574
rect 267 540 310 574
rect 190 506 310 540
rect 190 472 233 506
rect 267 472 310 506
rect 190 438 310 472
rect 190 404 233 438
rect 267 404 310 438
rect 190 380 310 404
rect 410 1186 530 1220
rect 410 1152 453 1186
rect 487 1152 530 1186
rect 410 1118 530 1152
rect 410 1084 453 1118
rect 487 1084 530 1118
rect 410 1050 530 1084
rect 410 1016 453 1050
rect 487 1016 530 1050
rect 410 982 530 1016
rect 410 948 453 982
rect 487 948 530 982
rect 410 914 530 948
rect 410 880 453 914
rect 487 880 530 914
rect 410 846 530 880
rect 410 812 453 846
rect 487 812 530 846
rect 410 778 530 812
rect 410 744 453 778
rect 487 744 530 778
rect 410 710 530 744
rect 410 676 453 710
rect 487 676 530 710
rect 410 642 530 676
rect 410 608 453 642
rect 487 608 530 642
rect 410 574 530 608
rect 410 540 453 574
rect 487 540 530 574
rect 410 506 530 540
rect 410 472 453 506
rect 487 472 530 506
rect 410 438 530 472
rect 410 404 453 438
rect 487 404 530 438
rect 410 380 530 404
rect 630 1186 750 1220
rect 630 1152 673 1186
rect 707 1152 750 1186
rect 630 1118 750 1152
rect 630 1084 673 1118
rect 707 1084 750 1118
rect 630 1050 750 1084
rect 630 1016 673 1050
rect 707 1016 750 1050
rect 630 982 750 1016
rect 630 948 673 982
rect 707 948 750 982
rect 630 914 750 948
rect 630 880 673 914
rect 707 880 750 914
rect 630 846 750 880
rect 630 812 673 846
rect 707 812 750 846
rect 630 778 750 812
rect 630 744 673 778
rect 707 744 750 778
rect 630 710 750 744
rect 630 676 673 710
rect 707 676 750 710
rect 630 642 750 676
rect 630 608 673 642
rect 707 608 750 642
rect 630 574 750 608
rect 630 540 673 574
rect 707 540 750 574
rect 630 506 750 540
rect 630 472 673 506
rect 707 472 750 506
rect 630 438 750 472
rect 630 404 673 438
rect 707 404 750 438
rect 630 380 750 404
rect 850 1186 970 1220
rect 850 1152 893 1186
rect 927 1152 970 1186
rect 850 1118 970 1152
rect 850 1084 893 1118
rect 927 1084 970 1118
rect 850 1050 970 1084
rect 850 1016 893 1050
rect 927 1016 970 1050
rect 850 982 970 1016
rect 850 948 893 982
rect 927 948 970 982
rect 850 914 970 948
rect 850 880 893 914
rect 927 880 970 914
rect 850 846 970 880
rect 850 812 893 846
rect 927 812 970 846
rect 850 778 970 812
rect 850 744 893 778
rect 927 744 970 778
rect 850 710 970 744
rect 850 676 893 710
rect 927 676 970 710
rect 850 642 970 676
rect 850 608 893 642
rect 927 608 970 642
rect 850 574 970 608
rect 850 540 893 574
rect 927 540 970 574
rect 850 506 970 540
rect 850 472 893 506
rect 927 472 970 506
rect 850 438 970 472
rect 850 404 893 438
rect 927 404 970 438
rect 850 380 970 404
<< pdiffc >>
rect 13 1152 47 1186
rect 13 1084 47 1118
rect 13 1016 47 1050
rect 13 948 47 982
rect 13 880 47 914
rect 13 812 47 846
rect 13 744 47 778
rect 13 676 47 710
rect 13 608 47 642
rect 13 540 47 574
rect 13 472 47 506
rect 13 404 47 438
rect 233 1152 267 1186
rect 233 1084 267 1118
rect 233 1016 267 1050
rect 233 948 267 982
rect 233 880 267 914
rect 233 812 267 846
rect 233 744 267 778
rect 233 676 267 710
rect 233 608 267 642
rect 233 540 267 574
rect 233 472 267 506
rect 233 404 267 438
rect 453 1152 487 1186
rect 453 1084 487 1118
rect 453 1016 487 1050
rect 453 948 487 982
rect 453 880 487 914
rect 453 812 487 846
rect 453 744 487 778
rect 453 676 487 710
rect 453 608 487 642
rect 453 540 487 574
rect 453 472 487 506
rect 453 404 487 438
rect 673 1152 707 1186
rect 673 1084 707 1118
rect 673 1016 707 1050
rect 673 948 707 982
rect 673 880 707 914
rect 673 812 707 846
rect 673 744 707 778
rect 673 676 707 710
rect 673 608 707 642
rect 673 540 707 574
rect 673 472 707 506
rect 673 404 707 438
rect 893 1152 927 1186
rect 893 1084 927 1118
rect 893 1016 927 1050
rect 893 948 927 982
rect 893 880 927 914
rect 893 812 927 846
rect 893 744 927 778
rect 893 676 927 710
rect 893 608 927 642
rect 893 540 927 574
rect 893 472 927 506
rect 893 404 927 438
<< nsubdiff >>
rect -150 1186 -30 1220
rect -150 1152 -107 1186
rect -73 1152 -30 1186
rect -150 1118 -30 1152
rect -150 1084 -107 1118
rect -73 1084 -30 1118
rect -150 1050 -30 1084
rect -150 1016 -107 1050
rect -73 1016 -30 1050
rect -150 982 -30 1016
rect -150 948 -107 982
rect -73 948 -30 982
rect -150 914 -30 948
rect -150 880 -107 914
rect -73 880 -30 914
rect -150 846 -30 880
rect -150 812 -107 846
rect -73 812 -30 846
rect -150 778 -30 812
rect -150 744 -107 778
rect -73 744 -30 778
rect -150 710 -30 744
rect -150 676 -107 710
rect -73 676 -30 710
rect -150 642 -30 676
rect -150 608 -107 642
rect -73 608 -30 642
rect -150 574 -30 608
rect -150 540 -107 574
rect -73 540 -30 574
rect -150 506 -30 540
rect -150 472 -107 506
rect -73 472 -30 506
rect -150 438 -30 472
rect -150 404 -107 438
rect -73 404 -30 438
rect -150 380 -30 404
<< nsubdiffcont >>
rect -107 1152 -73 1186
rect -107 1084 -73 1118
rect -107 1016 -73 1050
rect -107 948 -73 982
rect -107 880 -73 914
rect -107 812 -73 846
rect -107 744 -73 778
rect -107 676 -73 710
rect -107 608 -73 642
rect -107 540 -73 574
rect -107 472 -73 506
rect -107 404 -73 438
<< poly >>
rect 90 1250 850 1280
rect 90 1220 190 1250
rect 310 1220 410 1250
rect 530 1220 630 1250
rect 750 1220 850 1250
rect 90 330 190 380
rect 310 330 410 380
rect 530 330 630 380
rect 750 330 850 380
<< locali >>
rect 10 1240 930 1280
rect 10 1200 50 1240
rect 450 1200 490 1240
rect 890 1200 930 1240
rect -130 1186 -50 1200
rect -130 1152 -107 1186
rect -73 1152 -50 1186
rect -130 1118 -50 1152
rect -130 1084 -107 1118
rect -73 1084 -50 1118
rect -130 1050 -50 1084
rect -130 1016 -107 1050
rect -73 1016 -50 1050
rect -130 982 -50 1016
rect -130 948 -107 982
rect -73 948 -50 982
rect -130 914 -50 948
rect -130 880 -107 914
rect -73 880 -50 914
rect -130 846 -50 880
rect -130 812 -107 846
rect -73 812 -50 846
rect -130 778 -50 812
rect -130 744 -107 778
rect -73 744 -50 778
rect -130 710 -50 744
rect -130 676 -107 710
rect -73 676 -50 710
rect -130 642 -50 676
rect -130 608 -107 642
rect -73 608 -50 642
rect -130 574 -50 608
rect -130 540 -107 574
rect -73 540 -50 574
rect -130 506 -50 540
rect -130 472 -107 506
rect -73 472 -50 506
rect -130 438 -50 472
rect -130 404 -107 438
rect -73 404 -50 438
rect -130 400 -50 404
rect -10 1186 70 1200
rect -10 1152 13 1186
rect 47 1152 70 1186
rect -10 1118 70 1152
rect -10 1084 13 1118
rect 47 1084 70 1118
rect -10 1050 70 1084
rect -10 1016 13 1050
rect 47 1016 70 1050
rect -10 982 70 1016
rect -10 948 13 982
rect 47 948 70 982
rect -10 914 70 948
rect -10 880 13 914
rect 47 880 70 914
rect -10 846 70 880
rect -10 812 13 846
rect 47 812 70 846
rect -10 778 70 812
rect -10 744 13 778
rect 47 744 70 778
rect -10 710 70 744
rect -10 676 13 710
rect 47 676 70 710
rect -10 642 70 676
rect -10 608 13 642
rect 47 608 70 642
rect -10 574 70 608
rect -10 540 13 574
rect 47 540 70 574
rect -10 506 70 540
rect -10 472 13 506
rect 47 472 70 506
rect -10 438 70 472
rect -10 404 13 438
rect 47 404 70 438
rect -10 400 70 404
rect 210 1186 290 1200
rect 210 1152 233 1186
rect 267 1152 290 1186
rect 210 1118 290 1152
rect 210 1084 233 1118
rect 267 1084 290 1118
rect 210 1050 290 1084
rect 210 1016 233 1050
rect 267 1016 290 1050
rect 210 982 290 1016
rect 210 948 233 982
rect 267 948 290 982
rect 210 914 290 948
rect 210 880 233 914
rect 267 880 290 914
rect 210 846 290 880
rect 210 812 233 846
rect 267 812 290 846
rect 210 778 290 812
rect 210 744 233 778
rect 267 744 290 778
rect 210 710 290 744
rect 210 676 233 710
rect 267 676 290 710
rect 210 642 290 676
rect 210 608 233 642
rect 267 608 290 642
rect 210 574 290 608
rect 210 540 233 574
rect 267 540 290 574
rect 210 506 290 540
rect 210 472 233 506
rect 267 472 290 506
rect 210 438 290 472
rect 210 404 233 438
rect 267 404 290 438
rect 210 400 290 404
rect 430 1186 510 1200
rect 430 1152 453 1186
rect 487 1152 510 1186
rect 430 1118 510 1152
rect 430 1084 453 1118
rect 487 1084 510 1118
rect 430 1050 510 1084
rect 430 1016 453 1050
rect 487 1016 510 1050
rect 430 982 510 1016
rect 430 948 453 982
rect 487 948 510 982
rect 430 914 510 948
rect 430 880 453 914
rect 487 880 510 914
rect 430 846 510 880
rect 430 812 453 846
rect 487 812 510 846
rect 430 778 510 812
rect 430 744 453 778
rect 487 744 510 778
rect 430 710 510 744
rect 430 676 453 710
rect 487 676 510 710
rect 430 642 510 676
rect 430 608 453 642
rect 487 608 510 642
rect 430 574 510 608
rect 430 540 453 574
rect 487 540 510 574
rect 430 506 510 540
rect 430 472 453 506
rect 487 472 510 506
rect 430 438 510 472
rect 430 404 453 438
rect 487 404 510 438
rect 430 400 510 404
rect 650 1186 730 1200
rect 650 1152 673 1186
rect 707 1152 730 1186
rect 650 1118 730 1152
rect 650 1084 673 1118
rect 707 1084 730 1118
rect 650 1050 730 1084
rect 650 1016 673 1050
rect 707 1016 730 1050
rect 650 982 730 1016
rect 650 948 673 982
rect 707 948 730 982
rect 650 914 730 948
rect 650 880 673 914
rect 707 880 730 914
rect 650 846 730 880
rect 650 812 673 846
rect 707 812 730 846
rect 650 778 730 812
rect 650 744 673 778
rect 707 744 730 778
rect 650 710 730 744
rect 650 676 673 710
rect 707 676 730 710
rect 650 642 730 676
rect 650 608 673 642
rect 707 608 730 642
rect 650 574 730 608
rect 650 540 673 574
rect 707 540 730 574
rect 650 506 730 540
rect 650 472 673 506
rect 707 472 730 506
rect 650 438 730 472
rect 650 404 673 438
rect 707 404 730 438
rect 650 400 730 404
rect 870 1186 950 1200
rect 870 1152 893 1186
rect 927 1152 950 1186
rect 870 1118 950 1152
rect 870 1084 893 1118
rect 927 1084 950 1118
rect 870 1050 950 1084
rect 870 1016 893 1050
rect 927 1016 950 1050
rect 870 982 950 1016
rect 870 948 893 982
rect 927 948 950 982
rect 870 914 950 948
rect 870 880 893 914
rect 927 880 950 914
rect 870 846 950 880
rect 870 812 893 846
rect 927 812 950 846
rect 870 778 950 812
rect 870 744 893 778
rect 927 744 950 778
rect 870 710 950 744
rect 870 676 893 710
rect 927 676 950 710
rect 870 642 950 676
rect 870 608 893 642
rect 927 608 950 642
rect 870 574 950 608
rect 870 540 893 574
rect 927 540 950 574
rect 870 506 950 540
rect 870 472 893 506
rect 927 472 950 506
rect 870 438 950 472
rect 870 404 893 438
rect 927 404 950 438
rect 870 400 950 404
rect 230 360 270 400
rect 670 360 710 400
rect 230 320 710 360
<< end >>
