* SPICE3 file created from CMOS_NOR.ext - technology: sky130A

.subckt CMOS_NOR A B NOR VP VN
X0 VN B NOR VN sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X1 NOR A VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_30_430# A VP VP sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X3 NOR B a_30_430# VP sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
.ends

