magic
tech sky130A
magscale 1 2
timestamp 1675786016
<< nwell >>
rect -949 486 811 676
rect -479 96 341 486
<< pwell >>
rect -935 -680 797 -88
<< nmos >>
rect -789 -414 -759 -114
rect -639 -414 -609 -114
rect -309 -414 -279 -114
rect -159 -414 -129 -114
rect -9 -414 21 -114
rect 141 -414 171 -114
rect 471 -414 501 -114
rect 621 -414 651 -114
<< pmos >>
rect -309 146 -279 446
rect -159 146 -129 446
rect -9 146 21 446
rect 141 146 171 446
<< ndiff >>
rect -909 -187 -789 -114
rect -909 -221 -866 -187
rect -832 -221 -789 -187
rect -909 -267 -789 -221
rect -909 -301 -866 -267
rect -832 -301 -789 -267
rect -909 -347 -789 -301
rect -909 -381 -866 -347
rect -832 -381 -789 -347
rect -909 -414 -789 -381
rect -759 -187 -639 -114
rect -759 -221 -716 -187
rect -682 -221 -639 -187
rect -759 -267 -639 -221
rect -759 -301 -716 -267
rect -682 -301 -639 -267
rect -759 -347 -639 -301
rect -759 -381 -716 -347
rect -682 -381 -639 -347
rect -759 -414 -639 -381
rect -609 -187 -489 -114
rect -609 -221 -566 -187
rect -532 -221 -489 -187
rect -609 -267 -489 -221
rect -609 -301 -566 -267
rect -532 -301 -489 -267
rect -609 -347 -489 -301
rect -609 -381 -566 -347
rect -532 -381 -489 -347
rect -609 -414 -489 -381
rect -429 -187 -309 -114
rect -429 -221 -386 -187
rect -352 -221 -309 -187
rect -429 -267 -309 -221
rect -429 -301 -386 -267
rect -352 -301 -309 -267
rect -429 -347 -309 -301
rect -429 -381 -386 -347
rect -352 -381 -309 -347
rect -429 -414 -309 -381
rect -279 -187 -159 -114
rect -279 -221 -236 -187
rect -202 -221 -159 -187
rect -279 -267 -159 -221
rect -279 -301 -236 -267
rect -202 -301 -159 -267
rect -279 -347 -159 -301
rect -279 -381 -236 -347
rect -202 -381 -159 -347
rect -279 -414 -159 -381
rect -129 -187 -9 -114
rect -129 -221 -86 -187
rect -52 -221 -9 -187
rect -129 -267 -9 -221
rect -129 -301 -86 -267
rect -52 -301 -9 -267
rect -129 -347 -9 -301
rect -129 -381 -86 -347
rect -52 -381 -9 -347
rect -129 -414 -9 -381
rect 21 -187 141 -114
rect 21 -221 64 -187
rect 98 -221 141 -187
rect 21 -267 141 -221
rect 21 -301 64 -267
rect 98 -301 141 -267
rect 21 -347 141 -301
rect 21 -381 64 -347
rect 98 -381 141 -347
rect 21 -414 141 -381
rect 171 -187 291 -114
rect 171 -221 214 -187
rect 248 -221 291 -187
rect 171 -267 291 -221
rect 171 -301 214 -267
rect 248 -301 291 -267
rect 171 -347 291 -301
rect 171 -381 214 -347
rect 248 -381 291 -347
rect 171 -414 291 -381
rect 351 -187 471 -114
rect 351 -221 394 -187
rect 428 -221 471 -187
rect 351 -267 471 -221
rect 351 -301 394 -267
rect 428 -301 471 -267
rect 351 -347 471 -301
rect 351 -381 394 -347
rect 428 -381 471 -347
rect 351 -414 471 -381
rect 501 -414 621 -114
rect 651 -187 771 -114
rect 651 -221 694 -187
rect 728 -221 771 -187
rect 651 -267 771 -221
rect 651 -301 694 -267
rect 728 -301 771 -267
rect 651 -347 771 -301
rect 651 -381 694 -347
rect 728 -381 771 -347
rect 651 -414 771 -381
<< pdiff >>
rect -429 373 -309 446
rect -429 339 -386 373
rect -352 339 -309 373
rect -429 293 -309 339
rect -429 259 -386 293
rect -352 259 -309 293
rect -429 213 -309 259
rect -429 179 -386 213
rect -352 179 -309 213
rect -429 146 -309 179
rect -279 373 -159 446
rect -279 339 -236 373
rect -202 339 -159 373
rect -279 293 -159 339
rect -279 259 -236 293
rect -202 259 -159 293
rect -279 213 -159 259
rect -279 179 -236 213
rect -202 179 -159 213
rect -279 146 -159 179
rect -129 373 -9 446
rect -129 339 -86 373
rect -52 339 -9 373
rect -129 293 -9 339
rect -129 259 -86 293
rect -52 259 -9 293
rect -129 213 -9 259
rect -129 179 -86 213
rect -52 179 -9 213
rect -129 146 -9 179
rect 21 373 141 446
rect 21 339 64 373
rect 98 339 141 373
rect 21 293 141 339
rect 21 259 64 293
rect 98 259 141 293
rect 21 213 141 259
rect 21 179 64 213
rect 98 179 141 213
rect 21 146 141 179
rect 171 373 291 446
rect 171 339 214 373
rect 248 339 291 373
rect 171 293 291 339
rect 171 259 214 293
rect 248 259 291 293
rect 171 213 291 259
rect 171 179 214 213
rect 248 179 291 213
rect 171 146 291 179
<< ndiffc >>
rect -866 -221 -832 -187
rect -866 -301 -832 -267
rect -866 -381 -832 -347
rect -716 -221 -682 -187
rect -716 -301 -682 -267
rect -716 -381 -682 -347
rect -566 -221 -532 -187
rect -566 -301 -532 -267
rect -566 -381 -532 -347
rect -386 -221 -352 -187
rect -386 -301 -352 -267
rect -386 -381 -352 -347
rect -236 -221 -202 -187
rect -236 -301 -202 -267
rect -236 -381 -202 -347
rect -86 -221 -52 -187
rect -86 -301 -52 -267
rect -86 -381 -52 -347
rect 64 -221 98 -187
rect 64 -301 98 -267
rect 64 -381 98 -347
rect 214 -221 248 -187
rect 214 -301 248 -267
rect 214 -381 248 -347
rect 394 -221 428 -187
rect 394 -301 428 -267
rect 394 -381 428 -347
rect 694 -221 728 -187
rect 694 -301 728 -267
rect 694 -381 728 -347
<< pdiffc >>
rect -386 339 -352 373
rect -386 259 -352 293
rect -386 179 -352 213
rect -236 339 -202 373
rect -236 259 -202 293
rect -236 179 -202 213
rect -86 339 -52 373
rect -86 259 -52 293
rect -86 179 -52 213
rect 64 339 98 373
rect 64 259 98 293
rect 64 179 98 213
rect 214 339 248 373
rect 214 259 248 293
rect 214 179 248 213
<< psubdiff >>
rect -909 -587 771 -554
rect -909 -621 -886 -587
rect -852 -621 -806 -587
rect -772 -621 -726 -587
rect -692 -621 -646 -587
rect -612 -621 -566 -587
rect -532 -621 -486 -587
rect -452 -621 -406 -587
rect -372 -621 -326 -587
rect -292 -621 -246 -587
rect -212 -621 -166 -587
rect -132 -621 -86 -587
rect -52 -621 -6 -587
rect 28 -621 74 -587
rect 108 -621 154 -587
rect 188 -621 234 -587
rect 268 -621 314 -587
rect 348 -621 394 -587
rect 428 -621 474 -587
rect 508 -621 554 -587
rect 588 -621 634 -587
rect 668 -621 714 -587
rect 748 -621 771 -587
rect -909 -654 771 -621
<< nsubdiff >>
rect -909 593 771 626
rect -909 559 -886 593
rect -852 559 -806 593
rect -772 559 -726 593
rect -692 559 -646 593
rect -612 559 -566 593
rect -532 559 -486 593
rect -452 559 -406 593
rect -372 559 -326 593
rect -292 559 -246 593
rect -212 559 -166 593
rect -132 559 -86 593
rect -52 559 -6 593
rect 28 559 74 593
rect 108 559 154 593
rect 188 559 234 593
rect 268 559 314 593
rect 348 559 394 593
rect 428 559 474 593
rect 508 559 554 593
rect 588 559 634 593
rect 668 559 714 593
rect 748 559 771 593
rect -909 526 771 559
<< psubdiffcont >>
rect -886 -621 -852 -587
rect -806 -621 -772 -587
rect -726 -621 -692 -587
rect -646 -621 -612 -587
rect -566 -621 -532 -587
rect -486 -621 -452 -587
rect -406 -621 -372 -587
rect -326 -621 -292 -587
rect -246 -621 -212 -587
rect -166 -621 -132 -587
rect -86 -621 -52 -587
rect -6 -621 28 -587
rect 74 -621 108 -587
rect 154 -621 188 -587
rect 234 -621 268 -587
rect 314 -621 348 -587
rect 394 -621 428 -587
rect 474 -621 508 -587
rect 554 -621 588 -587
rect 634 -621 668 -587
rect 714 -621 748 -587
<< nsubdiffcont >>
rect -886 559 -852 593
rect -806 559 -772 593
rect -726 559 -692 593
rect -646 559 -612 593
rect -566 559 -532 593
rect -486 559 -452 593
rect -406 559 -372 593
rect -326 559 -292 593
rect -246 559 -212 593
rect -166 559 -132 593
rect -86 559 -52 593
rect -6 559 28 593
rect 74 559 108 593
rect 154 559 188 593
rect 234 559 268 593
rect 314 559 348 593
rect 394 559 428 593
rect 474 559 508 593
rect 554 559 588 593
rect 634 559 668 593
rect 714 559 748 593
<< poly >>
rect -309 476 -129 506
rect -309 446 -279 476
rect -159 446 -129 476
rect -9 476 171 506
rect -9 446 21 476
rect 141 446 171 476
rect -689 143 -609 166
rect 571 363 651 386
rect 571 329 594 363
rect 628 329 651 363
rect 571 306 651 329
rect 421 243 501 266
rect 421 209 444 243
rect 478 209 501 243
rect 421 186 501 209
rect -689 109 -666 143
rect -632 109 -609 143
rect -309 116 -279 146
rect -689 86 -609 109
rect -839 43 -759 66
rect -839 9 -816 43
rect -782 9 -759 43
rect -839 -14 -759 9
rect -789 -114 -759 -14
rect -639 -114 -609 86
rect -159 -9 -129 146
rect -9 116 21 146
rect 141 116 171 146
rect -59 93 21 116
rect -59 59 -36 93
rect -2 59 21 93
rect -59 36 21 59
rect -159 -32 -79 -9
rect -159 -66 -136 -32
rect -102 -66 -79 -32
rect -309 -114 -279 -84
rect -159 -89 -79 -66
rect -159 -114 -129 -89
rect -9 -114 21 36
rect 141 -114 171 -84
rect 471 -114 501 186
rect 621 -114 651 306
rect -789 -444 -759 -414
rect -639 -444 -609 -414
rect -309 -444 -279 -414
rect -159 -444 -129 -414
rect -9 -444 21 -414
rect 141 -444 171 -414
rect 471 -444 501 -414
rect 621 -444 651 -414
rect -309 -467 -229 -444
rect -309 -501 -286 -467
rect -252 -501 -229 -467
rect -309 -524 -229 -501
rect 91 -467 171 -444
rect 91 -501 114 -467
rect 148 -501 171 -467
rect 91 -524 171 -501
<< polycont >>
rect 594 329 628 363
rect 444 209 478 243
rect -666 109 -632 143
rect -816 9 -782 43
rect -36 59 -2 93
rect -136 -66 -102 -32
rect -286 -501 -252 -467
rect 114 -501 148 -467
<< locali >>
rect -909 593 771 616
rect -909 559 -886 593
rect -852 559 -806 593
rect -772 559 -726 593
rect -692 559 -646 593
rect -612 559 -566 593
rect -532 559 -486 593
rect -452 559 -406 593
rect -372 559 -326 593
rect -292 559 -246 593
rect -212 559 -166 593
rect -132 559 -86 593
rect -52 559 -6 593
rect 28 559 74 593
rect 108 559 154 593
rect 188 559 234 593
rect 268 559 314 593
rect 348 559 394 593
rect 428 559 474 593
rect 508 559 554 593
rect 588 559 634 593
rect 668 559 714 593
rect 748 559 771 593
rect -909 536 771 559
rect -559 366 -479 386
rect -909 363 -479 366
rect -909 329 -536 363
rect -502 329 -479 363
rect -909 326 -479 329
rect -559 306 -479 326
rect -409 373 -329 406
rect -409 339 -386 373
rect -352 339 -329 373
rect -409 293 -329 339
rect -559 246 -479 266
rect -909 243 -479 246
rect -909 209 -536 243
rect -502 209 -479 243
rect -909 206 -479 209
rect -559 186 -479 206
rect -409 259 -386 293
rect -352 259 -329 293
rect -409 213 -329 259
rect -409 179 -386 213
rect -352 179 -329 213
rect -689 146 -609 166
rect -409 156 -329 179
rect -259 373 -179 406
rect -259 339 -236 373
rect -202 339 -179 373
rect -259 293 -179 339
rect -259 259 -236 293
rect -202 259 -179 293
rect -259 213 -179 259
rect -259 179 -236 213
rect -202 179 -179 213
rect -259 146 -179 179
rect -109 373 -29 406
rect -109 339 -86 373
rect -52 339 -29 373
rect -109 293 -29 339
rect -109 259 -86 293
rect -52 259 -29 293
rect -109 213 -29 259
rect -109 179 -86 213
rect -52 179 -29 213
rect -109 156 -29 179
rect 41 373 121 406
rect 41 339 64 373
rect 98 339 121 373
rect 41 293 121 339
rect 41 259 64 293
rect 98 259 121 293
rect 41 213 121 259
rect 41 179 64 213
rect 98 179 121 213
rect 41 146 121 179
rect 191 373 271 406
rect 191 339 214 373
rect 248 339 271 373
rect 191 293 271 339
rect 571 363 651 386
rect 571 329 594 363
rect 628 329 651 363
rect 571 306 651 329
rect 191 259 214 293
rect 248 259 271 293
rect 191 213 271 259
rect 191 179 214 213
rect 248 179 271 213
rect 421 243 501 266
rect 421 209 444 243
rect 478 209 501 243
rect 421 186 501 209
rect 191 156 271 179
rect -909 143 -609 146
rect -909 109 -666 143
rect -632 109 -609 143
rect -909 106 -609 109
rect -689 86 -609 106
rect -239 96 -199 146
rect -59 96 21 116
rect -239 93 21 96
rect -839 46 -759 66
rect -909 43 -759 46
rect -909 9 -816 43
rect -782 9 -759 43
rect -909 6 -759 9
rect -839 -14 -759 6
rect -239 59 -36 93
rect -2 59 21 93
rect -239 56 21 59
rect -239 -74 -199 56
rect -59 36 21 56
rect -869 -114 -199 -74
rect -159 -24 -79 -9
rect 61 -24 101 146
rect 341 96 421 116
rect 341 93 771 96
rect 341 59 364 93
rect 398 59 771 93
rect 341 56 771 59
rect 341 36 421 56
rect -159 -32 771 -24
rect -159 -66 -136 -32
rect -102 -64 771 -32
rect -102 -66 -79 -64
rect -159 -89 -79 -66
rect -869 -154 -829 -114
rect -569 -154 -529 -114
rect -238 -154 -199 -114
rect 61 -154 101 -64
rect 391 -154 431 -64
rect -889 -187 -809 -154
rect -889 -221 -866 -187
rect -832 -221 -809 -187
rect -889 -267 -809 -221
rect -889 -301 -866 -267
rect -832 -301 -809 -267
rect -889 -347 -809 -301
rect -889 -381 -866 -347
rect -832 -381 -809 -347
rect -889 -404 -809 -381
rect -739 -187 -659 -154
rect -739 -221 -716 -187
rect -682 -221 -659 -187
rect -739 -267 -659 -221
rect -739 -301 -716 -267
rect -682 -301 -659 -267
rect -739 -347 -659 -301
rect -739 -381 -716 -347
rect -682 -381 -659 -347
rect -739 -404 -659 -381
rect -589 -187 -509 -154
rect -589 -221 -566 -187
rect -532 -221 -509 -187
rect -589 -267 -509 -221
rect -589 -301 -566 -267
rect -532 -301 -509 -267
rect -589 -347 -509 -301
rect -589 -381 -566 -347
rect -532 -381 -509 -347
rect -589 -404 -509 -381
rect -409 -187 -329 -154
rect -409 -221 -386 -187
rect -352 -221 -329 -187
rect -409 -267 -329 -221
rect -409 -301 -386 -267
rect -352 -301 -329 -267
rect -409 -347 -329 -301
rect -409 -381 -386 -347
rect -352 -381 -329 -347
rect -409 -404 -329 -381
rect -259 -187 -179 -154
rect -259 -221 -236 -187
rect -202 -221 -179 -187
rect -259 -267 -179 -221
rect -259 -301 -236 -267
rect -202 -301 -179 -267
rect -259 -347 -179 -301
rect -259 -381 -236 -347
rect -202 -381 -179 -347
rect -259 -404 -179 -381
rect -109 -187 -29 -154
rect -109 -221 -86 -187
rect -52 -221 -29 -187
rect -109 -267 -29 -221
rect -109 -301 -86 -267
rect -52 -301 -29 -267
rect -109 -347 -29 -301
rect -109 -381 -86 -347
rect -52 -381 -29 -347
rect -109 -404 -29 -381
rect 41 -187 121 -154
rect 41 -221 64 -187
rect 98 -221 121 -187
rect 41 -267 121 -221
rect 41 -301 64 -267
rect 98 -301 121 -267
rect 41 -347 121 -301
rect 41 -381 64 -347
rect 98 -381 121 -347
rect 41 -404 121 -381
rect 191 -187 271 -154
rect 191 -221 214 -187
rect 248 -221 271 -187
rect 191 -267 271 -221
rect 191 -301 214 -267
rect 248 -301 271 -267
rect 191 -347 271 -301
rect 191 -381 214 -347
rect 248 -381 271 -347
rect 191 -404 271 -381
rect 371 -187 451 -154
rect 371 -221 394 -187
rect 428 -221 451 -187
rect 371 -267 451 -221
rect 371 -301 394 -267
rect 428 -301 451 -267
rect 371 -347 451 -301
rect 371 -381 394 -347
rect 428 -381 451 -347
rect 371 -404 451 -381
rect 671 -187 751 -154
rect 671 -221 694 -187
rect 728 -221 751 -187
rect 671 -267 751 -221
rect 671 -301 694 -267
rect 728 -301 751 -267
rect 671 -347 751 -301
rect 671 -381 694 -347
rect 728 -381 751 -347
rect 671 -404 751 -381
rect -309 -464 -229 -444
rect 91 -464 171 -444
rect -909 -467 171 -464
rect -909 -501 -286 -467
rect -252 -501 114 -467
rect 148 -501 171 -467
rect -909 -504 171 -501
rect -309 -524 -229 -504
rect 91 -524 171 -504
rect -909 -587 771 -564
rect -909 -621 -886 -587
rect -852 -621 -806 -587
rect -772 -621 -726 -587
rect -692 -621 -646 -587
rect -612 -621 -566 -587
rect -532 -621 -486 -587
rect -452 -621 -406 -587
rect -372 -621 -326 -587
rect -292 -621 -246 -587
rect -212 -621 -166 -587
rect -132 -621 -86 -587
rect -52 -621 -6 -587
rect 28 -621 74 -587
rect 108 -621 154 -587
rect 188 -621 234 -587
rect 268 -621 314 -587
rect 348 -621 394 -587
rect 428 -621 474 -587
rect 508 -621 554 -587
rect 588 -621 634 -587
rect 668 -621 714 -587
rect 748 -621 771 -587
rect -909 -644 771 -621
<< viali >>
rect -886 559 -852 593
rect -806 559 -772 593
rect -726 559 -692 593
rect -646 559 -612 593
rect -566 559 -532 593
rect -486 559 -452 593
rect -406 559 -372 593
rect -326 559 -292 593
rect -246 559 -212 593
rect -166 559 -132 593
rect -86 559 -52 593
rect -6 559 28 593
rect 74 559 108 593
rect 154 559 188 593
rect 234 559 268 593
rect 314 559 348 593
rect 394 559 428 593
rect 474 559 508 593
rect 554 559 588 593
rect 634 559 668 593
rect 714 559 748 593
rect -536 329 -502 363
rect -386 339 -352 373
rect -536 209 -502 243
rect -386 259 -352 293
rect -386 179 -352 213
rect -86 339 -52 373
rect -86 259 -52 293
rect -86 179 -52 213
rect 214 339 248 373
rect 594 329 628 363
rect 214 259 248 293
rect 214 179 248 213
rect 444 209 478 243
rect -36 59 -2 93
rect 364 59 398 93
rect -716 -221 -682 -187
rect -716 -301 -682 -267
rect -716 -381 -682 -347
rect -386 -221 -352 -187
rect -386 -301 -352 -267
rect -386 -381 -352 -347
rect -86 -221 -52 -187
rect -86 -301 -52 -267
rect -86 -381 -52 -347
rect 214 -221 248 -187
rect 214 -301 248 -267
rect 214 -381 248 -347
rect 694 -221 728 -187
rect 694 -301 728 -267
rect 694 -381 728 -347
rect -886 -621 -852 -587
rect -806 -621 -772 -587
rect -726 -621 -692 -587
rect -646 -621 -612 -587
rect -566 -621 -532 -587
rect -486 -621 -452 -587
rect -406 -621 -372 -587
rect -326 -621 -292 -587
rect -246 -621 -212 -587
rect -166 -621 -132 -587
rect -86 -621 -52 -587
rect -6 -621 28 -587
rect 74 -621 108 -587
rect 154 -621 188 -587
rect 234 -621 268 -587
rect 314 -621 348 -587
rect 394 -621 428 -587
rect 474 -621 508 -587
rect 554 -621 588 -587
rect 634 -621 668 -587
rect 714 -621 748 -587
<< metal1 >>
rect -909 593 771 626
rect -909 559 -886 593
rect -852 559 -806 593
rect -772 559 -726 593
rect -692 559 -646 593
rect -612 559 -566 593
rect -532 559 -486 593
rect -452 559 -406 593
rect -372 559 -326 593
rect -292 559 -246 593
rect -212 559 -166 593
rect -132 559 -86 593
rect -52 559 -6 593
rect 28 559 74 593
rect 108 559 154 593
rect 188 559 234 593
rect 268 559 314 593
rect 348 559 394 593
rect 428 559 474 593
rect 508 559 554 593
rect 588 559 634 593
rect 668 559 714 593
rect 748 559 771 593
rect -909 526 771 559
rect -719 -154 -679 526
rect -559 372 -479 386
rect -559 320 -545 372
rect -493 320 -479 372
rect -559 306 -479 320
rect -409 373 -329 526
rect -409 339 -386 373
rect -352 339 -329 373
rect -409 293 -329 339
rect -559 252 -479 266
rect -559 200 -545 252
rect -493 200 -479 252
rect -559 186 -479 200
rect -409 259 -386 293
rect -352 259 -329 293
rect -409 213 -329 259
rect -409 179 -386 213
rect -352 179 -329 213
rect -409 156 -329 179
rect -109 373 -29 526
rect -109 339 -86 373
rect -52 339 -29 373
rect -109 293 -29 339
rect -109 259 -86 293
rect -52 259 -29 293
rect -109 213 -29 259
rect -109 179 -86 213
rect -52 179 -29 213
rect -109 156 -29 179
rect 191 373 271 526
rect 191 339 214 373
rect 248 339 271 373
rect 191 293 271 339
rect 571 372 651 386
rect 571 320 585 372
rect 637 320 651 372
rect 571 306 651 320
rect 191 259 214 293
rect 248 259 271 293
rect 191 213 271 259
rect 191 179 214 213
rect 248 179 271 213
rect 421 252 501 266
rect 421 200 435 252
rect 487 200 501 252
rect 421 186 501 200
rect 191 156 271 179
rect -59 96 21 116
rect 341 96 421 116
rect -59 93 421 96
rect -59 59 -36 93
rect -2 59 364 93
rect 398 59 421 93
rect -59 56 421 59
rect -59 36 21 56
rect 341 36 421 56
rect 691 -154 731 526
rect -739 -187 -659 -154
rect -739 -221 -716 -187
rect -682 -221 -659 -187
rect -739 -267 -659 -221
rect -739 -301 -716 -267
rect -682 -301 -659 -267
rect -739 -347 -659 -301
rect -739 -381 -716 -347
rect -682 -381 -659 -347
rect -739 -404 -659 -381
rect -409 -187 -329 -154
rect -409 -221 -386 -187
rect -352 -221 -329 -187
rect -409 -267 -329 -221
rect -409 -301 -386 -267
rect -352 -301 -329 -267
rect -409 -347 -329 -301
rect -409 -381 -386 -347
rect -352 -381 -329 -347
rect -409 -404 -329 -381
rect -109 -187 -29 -154
rect -109 -221 -86 -187
rect -52 -221 -29 -187
rect -109 -267 -29 -221
rect -109 -301 -86 -267
rect -52 -301 -29 -267
rect -109 -347 -29 -301
rect -109 -381 -86 -347
rect -52 -381 -29 -347
rect -109 -404 -29 -381
rect 191 -187 271 -154
rect 191 -221 214 -187
rect 248 -221 271 -187
rect 191 -267 271 -221
rect 191 -301 214 -267
rect 248 -301 271 -267
rect 191 -347 271 -301
rect 191 -381 214 -347
rect 248 -381 271 -347
rect 191 -404 271 -381
rect 671 -187 751 -154
rect 671 -221 694 -187
rect 728 -221 751 -187
rect 671 -267 751 -221
rect 671 -301 694 -267
rect 728 -301 751 -267
rect 671 -347 751 -301
rect 671 -381 694 -347
rect 728 -381 751 -347
rect 671 -404 751 -381
rect -389 -554 -349 -404
rect -89 -554 -49 -404
rect 211 -554 251 -404
rect -909 -587 771 -554
rect -909 -621 -886 -587
rect -852 -621 -806 -587
rect -772 -621 -726 -587
rect -692 -621 -646 -587
rect -612 -621 -566 -587
rect -532 -621 -486 -587
rect -452 -621 -406 -587
rect -372 -621 -326 -587
rect -292 -621 -246 -587
rect -212 -621 -166 -587
rect -132 -621 -86 -587
rect -52 -621 -6 -587
rect 28 -621 74 -587
rect 108 -621 154 -587
rect 188 -621 234 -587
rect 268 -621 314 -587
rect 348 -621 394 -587
rect 428 -621 474 -587
rect 508 -621 554 -587
rect 588 -621 634 -587
rect 668 -621 714 -587
rect 748 -621 771 -587
rect -909 -654 771 -621
<< via1 >>
rect -545 363 -493 372
rect -545 329 -536 363
rect -536 329 -502 363
rect -502 329 -493 363
rect -545 320 -493 329
rect -545 243 -493 252
rect -545 209 -536 243
rect -536 209 -502 243
rect -502 209 -493 243
rect -545 200 -493 209
rect 585 363 637 372
rect 585 329 594 363
rect 594 329 628 363
rect 628 329 637 363
rect 585 320 637 329
rect 435 243 487 252
rect 435 209 444 243
rect 444 209 478 243
rect 478 209 487 243
rect 435 200 487 209
<< metal2 >>
rect -559 372 -479 386
rect -559 320 -545 372
rect -493 366 -479 372
rect 571 372 651 386
rect 571 366 585 372
rect -493 326 585 366
rect -493 320 -479 326
rect -559 306 -479 320
rect 571 320 585 326
rect 637 320 651 372
rect 571 306 651 320
rect -559 252 -479 266
rect -559 200 -545 252
rect -493 246 -479 252
rect 421 252 501 266
rect 421 246 435 252
rect -493 206 435 246
rect -493 200 -479 206
rect -559 186 -479 200
rect 421 200 435 206
rect 487 200 501 252
rect 421 186 501 200
<< labels >>
rlabel metal1 s -39 56 1 96 4 OUT_bar
port 1 nsew
rlabel metal1 s -89 -624 -49 -584 4 GND!
port 2 nsew
rlabel metal1 s -89 556 -49 596 4 CLK
port 3 nsew
rlabel locali s -139 -69 -99 -29 4 OUT
port 4 nsew
rlabel locali s -899 336 -879 356 4 A
port 5 nsew
rlabel locali s -899 116 -879 136 4 A_bar
port 6 nsew
rlabel locali s -899 216 -879 236 4 B
port 7 nsew
rlabel locali s -899 16 -879 36 4 B_bar
port 8 nsew
rlabel locali s -289 -504 -249 -464 4 Dis
port 9 nsew
<< end >>
