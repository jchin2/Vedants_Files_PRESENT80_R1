magic
tech sky130A
magscale 1 2
timestamp 1670882924
<< xpolycontact >>
rect -194 156 -124 588
rect -194 -588 -124 -156
rect 124 156 194 588
rect 124 -588 194 -156
<< xpolyres >>
rect -194 -156 -124 156
rect 124 -156 194 156
<< viali >>
rect -178 173 -140 570
rect 140 173 178 570
rect -178 -570 -140 -173
rect 140 -570 178 -173
<< metal1 >>
rect -184 570 -134 582
rect -184 173 -178 570
rect -140 173 -134 570
rect -184 161 -134 173
rect 134 570 184 582
rect 134 173 140 570
rect 178 173 184 570
rect 134 161 184 173
rect -184 -173 -134 -161
rect -184 -570 -178 -173
rect -140 -570 -134 -173
rect -184 -582 -134 -570
rect 134 -173 184 -161
rect 134 -570 140 -173
rect 178 -570 184 -173
rect 134 -582 184 -570
<< res0p35 >>
rect -196 -158 -122 158
rect 122 -158 196 158
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.56 m 1 nx 2 wmin 0.350 lmin 0.50 rho 2000 val 9.989k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
