magic
tech sky130A
timestamp 1671306811
<< end >>
