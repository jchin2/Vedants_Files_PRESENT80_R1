magic
tech sky130A
timestamp 1666721195
<< nwell >>
rect -545 520 215 610
rect -295 185 -25 520
<< nmos >>
rect -440 -70 -425 80
rect -275 -70 -260 80
rect -200 -70 -185 80
rect -125 -70 -110 80
rect -50 -70 -35 80
rect 115 -70 130 80
<< pmos >>
rect -200 210 -185 510
rect -125 210 -110 510
<< ndiff >>
rect -500 45 -440 80
rect -500 25 -480 45
rect -460 25 -440 45
rect -500 5 -440 25
rect -500 -15 -480 5
rect -460 -15 -440 5
rect -500 -35 -440 -15
rect -500 -55 -480 -35
rect -460 -55 -440 -35
rect -500 -70 -440 -55
rect -425 45 -365 80
rect -425 25 -405 45
rect -385 25 -365 45
rect -425 5 -365 25
rect -425 -15 -405 5
rect -385 -15 -365 5
rect -425 -35 -365 -15
rect -425 -55 -405 -35
rect -385 -55 -365 -35
rect -425 -70 -365 -55
rect -335 45 -275 80
rect -335 25 -315 45
rect -295 25 -275 45
rect -335 5 -275 25
rect -335 -15 -315 5
rect -295 -15 -275 5
rect -335 -35 -275 -15
rect -335 -55 -315 -35
rect -295 -55 -275 -35
rect -335 -70 -275 -55
rect -260 45 -200 80
rect -260 25 -240 45
rect -220 25 -200 45
rect -260 5 -200 25
rect -260 -15 -240 5
rect -220 -15 -200 5
rect -260 -35 -200 -15
rect -260 -55 -240 -35
rect -220 -55 -200 -35
rect -260 -70 -200 -55
rect -185 45 -125 80
rect -185 25 -165 45
rect -145 25 -125 45
rect -185 5 -125 25
rect -185 -15 -165 5
rect -145 -15 -125 5
rect -185 -35 -125 -15
rect -185 -55 -165 -35
rect -145 -55 -125 -35
rect -185 -70 -125 -55
rect -110 45 -50 80
rect -110 25 -90 45
rect -70 25 -50 45
rect -110 5 -50 25
rect -110 -15 -90 5
rect -70 -15 -50 5
rect -110 -35 -50 -15
rect -110 -55 -90 -35
rect -70 -55 -50 -35
rect -110 -70 -50 -55
rect -35 45 25 80
rect -35 25 -15 45
rect 5 25 25 45
rect -35 5 25 25
rect -35 -15 -15 5
rect 5 -15 25 5
rect -35 -35 25 -15
rect -35 -55 -15 -35
rect 5 -55 25 -35
rect -35 -70 25 -55
rect 55 45 115 80
rect 55 25 75 45
rect 95 25 115 45
rect 55 5 115 25
rect 55 -15 75 5
rect 95 -15 115 5
rect 55 -35 115 -15
rect 55 -55 75 -35
rect 95 -55 115 -35
rect 55 -70 115 -55
rect 130 45 190 80
rect 130 25 150 45
rect 170 25 190 45
rect 130 5 190 25
rect 130 -15 150 5
rect 170 -15 190 5
rect 130 -35 190 -15
rect 130 -55 150 -35
rect 170 -55 190 -35
rect 130 -70 190 -55
<< pdiff >>
rect -260 485 -200 510
rect -260 465 -240 485
rect -220 465 -200 485
rect -260 445 -200 465
rect -260 425 -240 445
rect -220 425 -200 445
rect -260 405 -200 425
rect -260 385 -240 405
rect -220 385 -200 405
rect -260 365 -200 385
rect -260 345 -240 365
rect -220 345 -200 365
rect -260 325 -200 345
rect -260 305 -240 325
rect -220 305 -200 325
rect -260 285 -200 305
rect -260 265 -240 285
rect -220 265 -200 285
rect -260 245 -200 265
rect -260 225 -240 245
rect -220 225 -200 245
rect -260 210 -200 225
rect -185 485 -125 510
rect -185 465 -165 485
rect -145 465 -125 485
rect -185 445 -125 465
rect -185 425 -165 445
rect -145 425 -125 445
rect -185 405 -125 425
rect -185 385 -165 405
rect -145 385 -125 405
rect -185 365 -125 385
rect -185 345 -165 365
rect -145 345 -125 365
rect -185 325 -125 345
rect -185 305 -165 325
rect -145 305 -125 325
rect -185 285 -125 305
rect -185 265 -165 285
rect -145 265 -125 285
rect -185 245 -125 265
rect -185 225 -165 245
rect -145 225 -125 245
rect -185 210 -125 225
rect -110 485 -50 510
rect -110 465 -90 485
rect -70 465 -50 485
rect -110 445 -50 465
rect -110 425 -90 445
rect -70 425 -50 445
rect -110 405 -50 425
rect -110 385 -90 405
rect -70 385 -50 405
rect -110 365 -50 385
rect -110 345 -90 365
rect -70 345 -50 365
rect -110 325 -50 345
rect -110 305 -90 325
rect -70 305 -50 325
rect -110 285 -50 305
rect -110 265 -90 285
rect -70 265 -50 285
rect -110 245 -50 265
rect -110 225 -90 245
rect -70 225 -50 245
rect -110 210 -50 225
<< ndiffc >>
rect -480 25 -460 45
rect -480 -15 -460 5
rect -480 -55 -460 -35
rect -405 25 -385 45
rect -405 -15 -385 5
rect -405 -55 -385 -35
rect -315 25 -295 45
rect -315 -15 -295 5
rect -315 -55 -295 -35
rect -240 25 -220 45
rect -240 -15 -220 5
rect -240 -55 -220 -35
rect -165 25 -145 45
rect -165 -15 -145 5
rect -165 -55 -145 -35
rect -90 25 -70 45
rect -90 -15 -70 5
rect -90 -55 -70 -35
rect -15 25 5 45
rect -15 -15 5 5
rect -15 -55 5 -35
rect 75 25 95 45
rect 75 -15 95 5
rect 75 -55 95 -35
rect 150 25 170 45
rect 150 -15 170 5
rect 150 -55 170 -35
<< pdiffc >>
rect -240 465 -220 485
rect -240 425 -220 445
rect -240 385 -220 405
rect -240 345 -220 365
rect -240 305 -220 325
rect -240 265 -220 285
rect -240 225 -220 245
rect -165 465 -145 485
rect -165 425 -145 445
rect -165 385 -145 405
rect -165 345 -145 365
rect -165 305 -145 325
rect -165 265 -145 285
rect -165 225 -145 245
rect -90 465 -70 485
rect -90 425 -70 445
rect -90 385 -70 405
rect -90 345 -70 365
rect -90 305 -70 325
rect -90 265 -70 285
rect -90 225 -70 245
<< psubdiff >>
rect -505 -205 195 -190
rect -505 -225 -485 -205
rect -465 -225 -445 -205
rect -425 -225 -405 -205
rect -385 -225 -365 -205
rect -345 -225 -325 -205
rect -305 -225 -285 -205
rect -265 -225 -245 -205
rect -225 -225 -205 -205
rect -185 -225 -165 -205
rect -145 -225 -125 -205
rect -105 -225 -85 -205
rect -65 -225 -45 -205
rect -25 -225 -5 -205
rect 15 -225 35 -205
rect 55 -225 75 -205
rect 95 -225 115 -205
rect 135 -225 155 -205
rect 175 -225 195 -205
rect -505 -240 195 -225
<< nsubdiff >>
rect -525 575 195 590
rect -525 555 -485 575
rect -465 555 -445 575
rect -425 555 -405 575
rect -385 555 -365 575
rect -345 555 -325 575
rect -305 555 -285 575
rect -265 555 -245 575
rect -225 555 -205 575
rect -185 555 -165 575
rect -145 555 -125 575
rect -105 555 -85 575
rect -65 555 -45 575
rect -25 555 -5 575
rect 15 555 35 575
rect 55 555 75 575
rect 95 555 115 575
rect 135 555 155 575
rect 175 555 195 575
rect -525 540 195 555
<< psubdiffcont >>
rect -485 -225 -465 -205
rect -445 -225 -425 -205
rect -405 -225 -385 -205
rect -365 -225 -345 -205
rect -325 -225 -305 -205
rect -285 -225 -265 -205
rect -245 -225 -225 -205
rect -205 -225 -185 -205
rect -165 -225 -145 -205
rect -125 -225 -105 -205
rect -85 -225 -65 -205
rect -45 -225 -25 -205
rect -5 -225 15 -205
rect 35 -225 55 -205
rect 75 -225 95 -205
rect 115 -225 135 -205
rect 155 -225 175 -205
<< nsubdiffcont >>
rect -485 555 -465 575
rect -445 555 -425 575
rect -405 555 -385 575
rect -365 555 -345 575
rect -325 555 -305 575
rect -285 555 -265 575
rect -245 555 -225 575
rect -205 555 -185 575
rect -165 555 -145 575
rect -125 555 -105 575
rect -85 555 -65 575
rect -45 555 -25 575
rect -5 555 15 575
rect 35 555 55 575
rect 75 555 95 575
rect 115 555 135 575
rect 155 555 175 575
<< poly >>
rect -200 510 -185 525
rect -125 510 -110 525
rect -200 135 -185 210
rect -125 195 -110 210
rect -150 185 -110 195
rect -150 165 -140 185
rect -120 165 -110 185
rect -150 155 -110 165
rect -465 125 -425 135
rect -465 105 -455 125
rect -435 105 -425 125
rect -465 95 -425 105
rect -200 125 -160 135
rect -200 105 -190 125
rect -170 105 -160 125
rect -200 95 -160 105
rect -440 80 -425 95
rect -275 80 -260 95
rect -200 80 -185 95
rect -125 80 -110 155
rect -50 80 -35 95
rect 115 80 130 95
rect -440 -85 -425 -70
rect -275 -85 -260 -70
rect -200 -85 -185 -70
rect -125 -85 -110 -70
rect -50 -85 -35 -70
rect -275 -95 -235 -85
rect -275 -115 -265 -95
rect -245 -115 -235 -95
rect -275 -125 -235 -115
rect -75 -95 -35 -85
rect -75 -115 -65 -95
rect -45 -115 -35 -95
rect -75 -125 -35 -115
rect 115 -135 130 -70
rect 105 -145 145 -135
rect 105 -165 115 -145
rect 135 -165 145 -145
rect 105 -175 145 -165
<< polycont >>
rect -140 165 -120 185
rect -455 105 -435 125
rect -190 105 -170 125
rect -265 -115 -245 -95
rect -65 -115 -45 -95
rect 115 -165 135 -145
<< locali >>
rect -525 575 195 585
rect -525 555 -485 575
rect -465 555 -445 575
rect -425 555 -405 575
rect -385 555 -365 575
rect -345 555 -325 575
rect -305 555 -285 575
rect -265 555 -245 575
rect -225 555 -205 575
rect -185 555 -165 575
rect -145 555 -125 575
rect -105 555 -85 575
rect -65 555 -45 575
rect -25 555 -5 575
rect 15 555 35 575
rect 55 555 75 575
rect 95 555 115 575
rect 135 555 155 575
rect 175 555 195 575
rect -525 545 195 555
rect -250 485 -210 495
rect -250 465 -240 485
rect -220 465 -210 485
rect -250 445 -210 465
rect -250 425 -240 445
rect -220 425 -210 445
rect -250 405 -210 425
rect -250 385 -240 405
rect -220 385 -210 405
rect -250 365 -210 385
rect -250 345 -240 365
rect -220 345 -210 365
rect -250 325 -210 345
rect -250 305 -240 325
rect -220 305 -210 325
rect -250 285 -210 305
rect -250 265 -240 285
rect -220 265 -210 285
rect -250 245 -210 265
rect -250 225 -240 245
rect -220 225 -210 245
rect -250 210 -210 225
rect -175 485 -135 495
rect -175 465 -165 485
rect -145 465 -135 485
rect -175 445 -135 465
rect -175 425 -165 445
rect -145 425 -135 445
rect -175 405 -135 425
rect -175 385 -165 405
rect -145 385 -135 405
rect -175 365 -135 385
rect -175 345 -165 365
rect -145 345 -135 365
rect -175 325 -135 345
rect -175 305 -165 325
rect -145 305 -135 325
rect -175 285 -135 305
rect -175 265 -165 285
rect -145 265 -135 285
rect -175 245 -135 265
rect -175 225 -165 245
rect -145 225 -135 245
rect -175 215 -135 225
rect -100 485 -60 495
rect -100 465 -90 485
rect -70 465 -60 485
rect -100 445 -60 465
rect -100 425 -90 445
rect -70 425 -60 445
rect -100 405 -60 425
rect -100 385 -90 405
rect -70 385 -60 405
rect -100 365 -60 385
rect -100 345 -90 365
rect -70 345 -60 365
rect -100 325 -60 345
rect -100 305 -90 325
rect -70 305 -60 325
rect -100 285 -60 305
rect -100 265 -90 285
rect -70 265 -60 285
rect -100 245 -60 265
rect -100 225 -90 245
rect -70 225 -60 245
rect -100 210 -60 225
rect -375 185 -335 195
rect -520 165 -365 185
rect -345 165 -335 185
rect -375 155 -335 165
rect -240 185 -220 210
rect -150 185 -110 195
rect -240 165 -140 185
rect -120 165 -110 185
rect -465 125 -425 135
rect -520 105 -455 125
rect -435 105 -425 125
rect -240 120 -220 165
rect -150 155 -110 165
rect -465 95 -425 105
rect -405 100 -220 120
rect -405 60 -385 100
rect -240 80 -220 100
rect -200 125 -160 135
rect -90 125 -70 210
rect -25 185 15 195
rect -25 165 -15 185
rect 5 165 210 185
rect -25 155 15 165
rect -200 105 -190 125
rect -170 105 210 125
rect -200 95 -160 105
rect -90 80 -70 105
rect -490 45 -450 60
rect -490 25 -480 45
rect -460 25 -450 45
rect -490 5 -450 25
rect -490 -15 -480 5
rect -460 -15 -450 5
rect -490 -35 -450 -15
rect -490 -55 -480 -35
rect -460 -55 -450 -35
rect -490 -65 -450 -55
rect -415 45 -375 60
rect -415 25 -405 45
rect -385 25 -375 45
rect -415 5 -375 25
rect -415 -15 -405 5
rect -385 -15 -375 5
rect -415 -35 -375 -15
rect -415 -55 -405 -35
rect -385 -55 -375 -35
rect -415 -65 -375 -55
rect -325 45 -285 60
rect -325 25 -315 45
rect -295 25 -285 45
rect -325 5 -285 25
rect -325 -15 -315 5
rect -295 -15 -285 5
rect -325 -35 -285 -15
rect -325 -55 -315 -35
rect -295 -55 -285 -35
rect -325 -65 -285 -55
rect -250 45 -210 80
rect -250 25 -240 45
rect -220 25 -210 45
rect -250 5 -210 25
rect -250 -15 -240 5
rect -220 -15 -210 5
rect -250 -35 -210 -15
rect -250 -55 -240 -35
rect -220 -55 -210 -35
rect -250 -65 -210 -55
rect -175 45 -135 60
rect -175 25 -165 45
rect -145 25 -135 45
rect -175 5 -135 25
rect -175 -15 -165 5
rect -145 -15 -135 5
rect -175 -35 -135 -15
rect -175 -55 -165 -35
rect -145 -55 -135 -35
rect -175 -65 -135 -55
rect -100 45 -60 80
rect 150 60 170 105
rect -100 25 -90 45
rect -70 25 -60 45
rect -100 5 -60 25
rect -100 -15 -90 5
rect -70 -15 -60 5
rect -100 -35 -60 -15
rect -100 -55 -90 -35
rect -70 -55 -60 -35
rect -100 -65 -60 -55
rect -25 45 15 60
rect -25 25 -15 45
rect 5 25 15 45
rect -25 5 15 25
rect -25 -15 -15 5
rect 5 -15 15 5
rect -25 -35 15 -15
rect -25 -55 -15 -35
rect 5 -55 15 -35
rect -25 -65 15 -55
rect 65 45 105 60
rect 65 25 75 45
rect 95 25 105 45
rect 65 5 105 25
rect 65 -15 75 5
rect 95 -15 105 5
rect 65 -35 105 -15
rect 65 -55 75 -35
rect 95 -55 105 -35
rect 65 -65 105 -55
rect 140 45 180 60
rect 140 25 150 45
rect 170 25 180 45
rect 140 5 180 25
rect 140 -15 150 5
rect 170 -15 180 5
rect 140 -35 180 -15
rect 140 -55 150 -35
rect 170 -55 180 -35
rect 140 -65 180 -55
rect -275 -95 -235 -85
rect -75 -95 -35 -85
rect -520 -115 -265 -95
rect -245 -115 -65 -95
rect -45 -115 -35 -95
rect -275 -125 -235 -115
rect -75 -125 -35 -115
rect -375 -145 -335 -135
rect 105 -145 145 -135
rect -375 -165 -365 -145
rect -345 -165 115 -145
rect 135 -165 145 -145
rect -375 -175 -335 -165
rect 105 -175 145 -165
rect -505 -205 195 -195
rect -505 -225 -485 -205
rect -465 -225 -445 -205
rect -425 -225 -405 -205
rect -385 -225 -365 -205
rect -345 -225 -325 -205
rect -305 -225 -285 -205
rect -265 -225 -245 -205
rect -225 -225 -205 -205
rect -185 -225 -165 -205
rect -145 -225 -125 -205
rect -105 -225 -85 -205
rect -65 -225 -45 -205
rect -25 -225 -5 -205
rect 15 -225 35 -205
rect 55 -225 75 -205
rect 95 -225 115 -205
rect 135 -225 155 -205
rect 175 -225 195 -205
rect -505 -235 195 -225
<< viali >>
rect -485 555 -465 575
rect -445 555 -425 575
rect -405 555 -385 575
rect -365 555 -345 575
rect -325 555 -305 575
rect -285 555 -265 575
rect -245 555 -225 575
rect -205 555 -185 575
rect -165 555 -145 575
rect -125 555 -105 575
rect -85 555 -65 575
rect -45 555 -25 575
rect -5 555 15 575
rect 35 555 55 575
rect 75 555 95 575
rect 115 555 135 575
rect 155 555 175 575
rect -165 465 -145 485
rect -165 425 -145 445
rect -165 385 -145 405
rect -165 345 -145 365
rect -165 305 -145 325
rect -165 265 -145 285
rect -165 225 -145 245
rect -365 165 -345 185
rect -140 165 -120 185
rect -15 165 5 185
rect -480 25 -460 45
rect -480 -15 -460 5
rect -480 -55 -460 -35
rect -315 25 -295 45
rect -315 -15 -295 5
rect -315 -55 -295 -35
rect -165 25 -145 45
rect -165 -15 -145 5
rect -165 -55 -145 -35
rect -15 25 5 45
rect -15 -15 5 5
rect -15 -55 5 -35
rect 75 25 95 45
rect 75 -15 95 5
rect 75 -55 95 -35
rect -365 -165 -345 -145
rect -485 -225 -465 -205
rect -445 -225 -425 -205
rect -405 -225 -385 -205
rect -365 -225 -345 -205
rect -325 -225 -305 -205
rect -285 -225 -265 -205
rect -245 -225 -225 -205
rect -205 -225 -185 -205
rect -165 -225 -145 -205
rect -125 -225 -105 -205
rect -85 -225 -65 -205
rect -45 -225 -25 -205
rect -5 -225 15 -205
rect 35 -225 55 -205
rect 75 -225 95 -205
rect 115 -225 135 -205
rect 155 -225 175 -205
<< metal1 >>
rect -525 575 195 590
rect -525 555 -485 575
rect -465 555 -445 575
rect -425 555 -405 575
rect -385 555 -365 575
rect -345 555 -325 575
rect -305 555 -285 575
rect -265 555 -245 575
rect -225 555 -205 575
rect -185 555 -165 575
rect -145 555 -125 575
rect -105 555 -85 575
rect -65 555 -45 575
rect -25 555 -5 575
rect 15 555 35 575
rect 55 555 75 575
rect 95 555 115 575
rect 135 555 155 575
rect 175 555 195 575
rect -525 540 195 555
rect -480 60 -460 540
rect -165 495 -145 540
rect -175 485 -135 495
rect -175 465 -165 485
rect -145 465 -135 485
rect -175 445 -135 465
rect -175 425 -165 445
rect -145 425 -135 445
rect -175 405 -135 425
rect -175 385 -165 405
rect -145 385 -135 405
rect -175 365 -135 385
rect -175 345 -165 365
rect -145 345 -135 365
rect -175 325 -135 345
rect -175 305 -165 325
rect -145 305 -135 325
rect -175 285 -135 305
rect -175 265 -165 285
rect -145 265 -135 285
rect -175 245 -135 265
rect -175 225 -165 245
rect -145 225 -135 245
rect -175 215 -135 225
rect -375 185 -335 195
rect -375 165 -365 185
rect -345 165 -335 185
rect -375 155 -335 165
rect -150 185 -110 195
rect -25 185 15 195
rect -150 165 -140 185
rect -120 165 -15 185
rect 5 165 15 185
rect -150 155 -110 165
rect -25 155 15 165
rect -490 45 -450 60
rect -490 25 -480 45
rect -460 25 -450 45
rect -490 5 -450 25
rect -490 -15 -480 5
rect -460 -15 -450 5
rect -490 -35 -450 -15
rect -490 -55 -480 -35
rect -460 -55 -450 -35
rect -490 -65 -450 -55
rect -365 -135 -345 155
rect 80 60 100 540
rect -325 45 -285 60
rect -325 25 -315 45
rect -295 25 -285 45
rect -325 5 -285 25
rect -325 -15 -315 5
rect -295 -15 -285 5
rect -325 -35 -285 -15
rect -325 -55 -315 -35
rect -295 -55 -285 -35
rect -325 -65 -285 -55
rect -175 45 -135 60
rect -175 25 -165 45
rect -145 25 -135 45
rect -175 5 -135 25
rect -175 -15 -165 5
rect -145 -15 -135 5
rect -175 -35 -135 -15
rect -175 -55 -165 -35
rect -145 -55 -135 -35
rect -175 -65 -135 -55
rect -25 45 15 60
rect -25 25 -15 45
rect 5 25 15 45
rect -25 5 15 25
rect -25 -15 -15 5
rect 5 -15 15 5
rect -25 -35 15 -15
rect -25 -55 -15 -35
rect 5 -55 15 -35
rect -25 -65 15 -55
rect 65 45 105 60
rect 65 25 75 45
rect 95 25 105 45
rect 65 5 105 25
rect 65 -15 75 5
rect 95 -15 105 5
rect 65 -35 105 -15
rect 65 -55 75 -35
rect 95 -55 105 -35
rect 65 -65 105 -55
rect -375 -145 -335 -135
rect -375 -165 -365 -145
rect -345 -165 -335 -145
rect -375 -175 -335 -165
rect -315 -190 -295 -65
rect -165 -190 -145 -65
rect -15 -190 5 -65
rect -520 -205 210 -190
rect -520 -225 -485 -205
rect -465 -225 -445 -205
rect -425 -225 -405 -205
rect -385 -225 -365 -205
rect -345 -225 -325 -205
rect -305 -225 -285 -205
rect -265 -225 -245 -205
rect -225 -225 -205 -205
rect -185 -225 -165 -205
rect -145 -225 -125 -205
rect -105 -225 -85 -205
rect -65 -225 -45 -205
rect -25 -225 -5 -205
rect 15 -225 35 -205
rect 55 -225 75 -205
rect 95 -225 115 -205
rect 135 -225 155 -205
rect 175 -225 210 -205
rect -520 -240 210 -225
<< labels >>
rlabel locali 195 110 205 120 3 OUT_bar
port 3 e
rlabel locali -515 -110 -505 -100 7 Dis
port 5 w
rlabel locali 195 170 205 180 3 OUT
port 2 e
rlabel metal1 -515 -220 -505 -210 1 GND!
port 6 n
rlabel metal1 -520 560 -510 570 7 CLK
port 4 w
rlabel locali -515 170 -505 180 7 A
port 0 w
rlabel locali -515 110 -505 120 7 A_bar
port 1 w
<< end >>
