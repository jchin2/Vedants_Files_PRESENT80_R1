magic
tech sky130A
magscale 1 2
timestamp 1677167040
<< locali >>
rect -2970 1399 -2890 1422
rect -2970 1365 -2947 1399
rect -2913 1365 -2890 1399
rect -2970 1330 -2890 1365
rect -2970 1327 -1920 1330
rect -2970 1293 -2947 1327
rect -2913 1293 -1920 1327
rect -2970 1290 -1920 1293
rect -1706 1326 -1554 1346
rect -1706 1323 -1480 1326
rect -2970 1255 -2890 1290
rect -1706 1289 -1683 1323
rect -1649 1289 -1611 1323
rect -1577 1289 -1480 1323
rect -1706 1286 -1480 1289
rect -1706 1266 -1554 1286
rect -2970 1221 -2947 1255
rect -2913 1221 -2890 1255
rect -2970 1198 -2890 1221
rect -2856 665 -2776 688
rect -2856 631 -2833 665
rect -2799 631 -2776 665
rect -2856 596 -2776 631
rect -2856 593 -2400 596
rect -2856 559 -2833 593
rect -2799 559 -2400 593
rect -2856 556 -2400 559
rect -1520 590 -1480 1286
rect -2856 521 -2776 556
rect -1520 550 -897 590
rect -167 556 315 596
rect 1045 550 1527 590
rect 2197 525 2277 548
rect -3654 474 -3574 497
rect -3654 440 -3631 474
rect -3597 440 -3574 474
rect -2856 487 -2833 521
rect -2799 487 -2776 521
rect -2856 464 -2776 487
rect -81 499 -1 522
rect -81 465 -58 499
rect -24 465 -1 499
rect -81 442 -1 465
rect 2197 491 2220 525
rect 2254 491 2277 525
rect 2197 453 2277 491
rect -3654 405 -3574 440
rect -3654 402 -2370 405
rect -3654 368 -3631 402
rect -3597 368 -2370 402
rect -3654 365 -2370 368
rect -3654 330 -3574 365
rect -3654 296 -3631 330
rect -3597 296 -3574 330
rect -3654 273 -3574 296
rect -3540 49 -3460 72
rect -3540 15 -3517 49
rect -3483 15 -3460 49
rect -3540 -20 -3460 15
rect -2816 -8 -2588 32
rect -2816 -20 -2776 -8
rect -3540 -23 -2776 -20
rect -3540 -57 -3517 -23
rect -3483 -57 -2776 -23
rect -2628 -20 -2588 -8
rect -1706 -19 -1554 4
rect -3540 -60 -2776 -57
rect -3540 -95 -3460 -60
rect -3540 -129 -3517 -95
rect -3483 -129 -3460 -95
rect -3540 -152 -3460 -129
rect -2742 -65 -2662 -42
rect -2628 -60 -1920 -20
rect -1706 -53 -1683 -19
rect -1649 -53 -1611 -19
rect -1577 -20 -1554 -19
rect -61 -20 -21 442
rect 2197 419 2220 453
rect 2254 419 2277 453
rect 2197 396 2277 419
rect -1577 -53 -717 -20
rect -1706 -60 -717 -53
rect -61 -60 495 -20
rect 1164 -60 1707 -20
rect -2742 -99 -2719 -65
rect -2685 -99 -2662 -65
rect -1706 -76 -1554 -60
rect -2742 -114 -2662 -99
rect -2742 -137 -2520 -114
rect -2856 -179 -2776 -156
rect -2856 -213 -2833 -179
rect -2799 -213 -2776 -179
rect -2856 -251 -2776 -213
rect -2856 -285 -2833 -251
rect -2799 -285 -2776 -251
rect -2742 -171 -2719 -137
rect -2685 -171 -2520 -137
rect -2742 -194 -2520 -171
rect -2742 -209 -2662 -194
rect -2742 -243 -2719 -209
rect -2685 -243 -2662 -209
rect -2742 -266 -2662 -243
rect -1481 -248 -1329 -232
rect -2856 -300 -2776 -285
rect -2628 -288 -1920 -248
rect -1481 -255 -717 -248
rect -2628 -300 -2588 -288
rect -2856 -323 -2588 -300
rect -1481 -289 -1458 -255
rect -1424 -289 -1386 -255
rect -1352 -288 -717 -255
rect -60 -288 495 -248
rect -1352 -289 -1329 -288
rect -1481 -312 -1329 -289
rect -2856 -357 -2833 -323
rect -2799 -340 -2588 -323
rect -2799 -357 -2776 -340
rect -2856 -380 -2776 -357
rect -60 -358 -20 -288
rect 1164 -358 1204 -60
rect -167 -398 -20 -358
rect 1065 -398 1204 -358
rect -2970 -604 -2890 -581
rect -2970 -638 -2947 -604
rect -2913 -638 -2890 -604
rect -2970 -673 -2890 -638
rect -2970 -676 -2370 -673
rect -2970 -710 -2947 -676
rect -2913 -710 -2370 -676
rect -2970 -713 -2370 -710
rect -1419 -701 -1339 -678
rect -2970 -748 -2890 -713
rect -3540 -795 -3460 -772
rect -3540 -829 -3517 -795
rect -3483 -829 -3460 -795
rect -2970 -782 -2947 -748
rect -2913 -782 -2890 -748
rect -2970 -805 -2890 -782
rect -1419 -735 -1396 -701
rect -1362 -735 -1339 -701
rect -1419 -773 -1339 -735
rect -3540 -864 -3460 -829
rect -1691 -827 -1611 -804
rect -1691 -861 -1668 -827
rect -1634 -861 -1611 -827
rect -1419 -807 -1396 -773
rect -1362 -807 -1339 -773
rect -1419 -830 -1339 -807
rect -81 -701 -1 -678
rect -81 -735 -58 -701
rect -24 -735 -1 -701
rect -81 -773 -1 -735
rect -81 -807 -58 -773
rect -24 -807 -1 -773
rect -81 -830 -1 -807
rect -3540 -867 -2400 -864
rect -3540 -901 -3517 -867
rect -3483 -901 -2400 -867
rect -1691 -884 -1611 -861
rect -1691 -898 -1671 -884
rect -1295 -898 -897 -858
rect -61 -864 -21 -830
rect -3540 -904 -2400 -901
rect -3540 -939 -3460 -904
rect -3540 -973 -3517 -939
rect -3483 -973 -3460 -939
rect -3540 -996 -3460 -973
rect -3654 -1529 -3574 -1506
rect -3654 -1563 -3631 -1529
rect -3597 -1563 -3574 -1529
rect -3654 -1598 -3574 -1563
rect -1481 -1594 -1329 -1574
rect -1295 -1594 -1255 -898
rect -61 -904 324 -864
rect -1481 -1597 -1255 -1594
rect -3654 -1601 -1920 -1598
rect -3654 -1635 -3631 -1601
rect -3597 -1635 -1920 -1601
rect -3654 -1638 -1920 -1635
rect -1481 -1631 -1458 -1597
rect -1424 -1631 -1386 -1597
rect -1352 -1631 -1255 -1597
rect -1481 -1634 -1255 -1631
rect -3654 -1673 -3574 -1638
rect -1481 -1654 -1329 -1634
rect -3654 -1707 -3631 -1673
rect -3597 -1707 -3574 -1673
rect -3654 -1730 -3574 -1707
<< viali >>
rect -2947 1365 -2913 1399
rect -2947 1293 -2913 1327
rect -1683 1289 -1649 1323
rect -1611 1289 -1577 1323
rect -2947 1221 -2913 1255
rect -2833 631 -2799 665
rect -2833 559 -2799 593
rect -3631 440 -3597 474
rect -2833 487 -2799 521
rect -58 465 -24 499
rect 2220 491 2254 525
rect -3631 368 -3597 402
rect -3631 296 -3597 330
rect -3517 15 -3483 49
rect -3517 -57 -3483 -23
rect -3517 -129 -3483 -95
rect -1683 -53 -1649 -19
rect -1611 -53 -1577 -19
rect 2220 419 2254 453
rect -2719 -99 -2685 -65
rect -2833 -213 -2799 -179
rect -2833 -285 -2799 -251
rect -2719 -171 -2685 -137
rect -2719 -243 -2685 -209
rect -1458 -289 -1424 -255
rect -1386 -289 -1352 -255
rect -2833 -357 -2799 -323
rect -2947 -638 -2913 -604
rect -2947 -710 -2913 -676
rect -3517 -829 -3483 -795
rect -2947 -782 -2913 -748
rect -1396 -735 -1362 -701
rect -1668 -861 -1634 -827
rect -1396 -807 -1362 -773
rect -58 -735 -24 -701
rect -58 -807 -24 -773
rect -3517 -901 -3483 -867
rect -3517 -973 -3483 -939
rect -3631 -1563 -3597 -1529
rect -3631 -1635 -3597 -1601
rect -1458 -1631 -1424 -1597
rect -1386 -1631 -1352 -1597
rect -3631 -1707 -3597 -1673
<< metal1 >>
rect -3654 474 -3574 1474
rect -3654 440 -3631 474
rect -3597 440 -3574 474
rect -3654 402 -3574 440
rect -3654 368 -3631 402
rect -3597 368 -3574 402
rect -3654 330 -3574 368
rect -3654 296 -3631 330
rect -3597 296 -3574 330
rect -3654 -1529 -3574 296
rect -3654 -1563 -3631 -1529
rect -3597 -1563 -3574 -1529
rect -3654 -1601 -3574 -1563
rect -3654 -1635 -3631 -1601
rect -3597 -1635 -3574 -1601
rect -3654 -1673 -3574 -1635
rect -3654 -1707 -3631 -1673
rect -3597 -1707 -3574 -1673
rect -3654 -1783 -3574 -1707
rect -3540 49 -3460 1474
rect -3540 15 -3517 49
rect -3483 15 -3460 49
rect -3540 -23 -3460 15
rect -3540 -57 -3517 -23
rect -3483 -57 -3460 -23
rect -3540 -95 -3460 -57
rect -3540 -129 -3517 -95
rect -3483 -129 -3460 -95
rect -3540 -795 -3460 -129
rect -3540 -829 -3517 -795
rect -3483 -829 -3460 -795
rect -3540 -867 -3460 -829
rect -3540 -901 -3517 -867
rect -3483 -901 -3460 -867
rect -3540 -939 -3460 -901
rect -3540 -973 -3517 -939
rect -3483 -973 -3460 -939
rect -3540 -1783 -3460 -973
rect -3426 1400 -3346 1474
rect -3426 1348 -3412 1400
rect -3360 1348 -3346 1400
rect -3426 1332 -3346 1348
rect -3426 1280 -3412 1332
rect -3360 1280 -3346 1332
rect -3426 1264 -3346 1280
rect -3426 1212 -3412 1264
rect -3360 1212 -3346 1264
rect -3426 -1783 -3346 1212
rect -3312 -1524 -3232 1474
rect -3312 -1576 -3298 -1524
rect -3246 -1576 -3232 -1524
rect -3312 -1592 -3232 -1576
rect -3312 -1644 -3298 -1592
rect -3246 -1644 -3232 -1592
rect -3312 -1660 -3232 -1644
rect -3312 -1712 -3298 -1660
rect -3246 -1712 -3232 -1660
rect -3312 -1783 -3232 -1712
rect -3198 -178 -3118 1474
rect -3198 -230 -3184 -178
rect -3132 -230 -3118 -178
rect -3198 -246 -3118 -230
rect -3198 -298 -3184 -246
rect -3132 -298 -3118 -246
rect -3198 -314 -3118 -298
rect -3198 -366 -3184 -314
rect -3132 -366 -3118 -314
rect -3198 -1782 -3118 -366
rect -3084 58 -3004 1474
rect -3084 6 -3070 58
rect -3018 6 -3004 58
rect -3084 -10 -3004 6
rect -3084 -62 -3070 -10
rect -3018 -62 -3004 -10
rect -3084 -78 -3004 -62
rect -3084 -130 -3070 -78
rect -3018 -130 -3004 -78
rect -3084 -1783 -3004 -130
rect -2970 1399 -2890 1474
rect -2970 1365 -2947 1399
rect -2913 1365 -2890 1399
rect -2970 1327 -2890 1365
rect -2970 1293 -2947 1327
rect -2913 1293 -2890 1327
rect -2970 1255 -2890 1293
rect -2970 1221 -2947 1255
rect -2913 1221 -2890 1255
rect -2970 -604 -2890 1221
rect -2970 -638 -2947 -604
rect -2913 -638 -2890 -604
rect -2970 -676 -2890 -638
rect -2970 -710 -2947 -676
rect -2913 -710 -2890 -676
rect -2970 -748 -2890 -710
rect -2970 -782 -2947 -748
rect -2913 -782 -2890 -748
rect -2970 -1782 -2890 -782
rect -2856 665 -2776 1474
rect -2856 631 -2833 665
rect -2799 631 -2776 665
rect -2856 593 -2776 631
rect -2856 559 -2833 593
rect -2799 559 -2776 593
rect -2856 521 -2776 559
rect -2856 487 -2833 521
rect -2799 487 -2776 521
rect -2856 -179 -2776 487
rect -2856 -213 -2833 -179
rect -2799 -213 -2776 -179
rect -2856 -251 -2776 -213
rect -2856 -285 -2833 -251
rect -2799 -285 -2776 -251
rect -2856 -323 -2776 -285
rect -2856 -357 -2833 -323
rect -2799 -357 -2776 -323
rect -2856 -1782 -2776 -357
rect -2742 -65 -2662 1474
rect -2742 -99 -2719 -65
rect -2685 -99 -2662 -65
rect -2742 -137 -2662 -99
rect -2742 -171 -2719 -137
rect -2685 -171 -2662 -137
rect -2742 -209 -2662 -171
rect -2742 -243 -2719 -209
rect -2685 -243 -2662 -209
rect -2742 -1782 -2662 -243
rect -2628 1374 -2520 1474
rect -1640 1374 -962 1474
rect -428 1374 250 1474
rect 1130 1374 1462 1474
rect -2628 -1682 -2548 1374
rect -1706 1332 -1554 1346
rect -1706 1280 -1692 1332
rect -1640 1280 -1620 1332
rect -1568 1280 -1554 1332
rect -1706 1266 -1554 1280
rect 2197 534 2277 548
rect -1676 508 -1528 522
rect -1676 456 -1662 508
rect -1610 456 -1594 508
rect -1542 502 -1528 508
rect -81 502 -1 522
rect -1542 499 -1 502
rect -1542 465 -58 499
rect -24 465 -1 499
rect -1542 462 -1 465
rect -1542 456 -1528 462
rect -1676 442 -1528 456
rect -81 442 -1 462
rect 2197 482 2211 534
rect 2263 482 2277 534
rect 2197 462 2277 482
rect 2197 410 2211 462
rect 2263 410 2277 462
rect 2197 396 2277 410
rect -1706 -10 -1554 4
rect -1706 -62 -1692 -10
rect -1640 -62 -1620 -10
rect -1568 -62 -1554 -10
rect -1706 -76 -1554 -62
rect -1283 -204 -951 -104
rect -82 -204 250 -104
rect 1130 -204 1462 -104
rect -1481 -246 -1329 -232
rect -1481 -298 -1467 -246
rect -1415 -298 -1395 -246
rect -1343 -298 -1329 -246
rect -1481 -312 -1329 -298
rect -1419 -701 -1339 -678
rect -1419 -735 -1396 -701
rect -1362 -735 -1339 -701
rect -1419 -770 -1339 -735
rect -81 -701 -1 -678
rect -81 -735 -58 -701
rect -24 -735 -1 -701
rect -81 -770 -1 -735
rect -1419 -773 -1 -770
rect -1691 -818 -1611 -804
rect -1691 -870 -1677 -818
rect -1625 -870 -1611 -818
rect -1419 -807 -1396 -773
rect -1362 -807 -58 -773
rect -24 -807 -1 -773
rect -1419 -810 -1 -807
rect -1419 -830 -1339 -810
rect -81 -830 -1 -810
rect -1691 -884 -1611 -870
rect -1481 -1588 -1329 -1574
rect -1481 -1640 -1467 -1588
rect -1415 -1640 -1395 -1588
rect -1343 -1640 -1329 -1588
rect -1481 -1654 -1329 -1640
rect -2628 -1782 -2520 -1682
rect -1294 -1782 -962 -1682
rect -82 -1782 250 -1682
<< via1 >>
rect -3412 1348 -3360 1400
rect -3412 1280 -3360 1332
rect -3412 1212 -3360 1264
rect -3298 -1576 -3246 -1524
rect -3298 -1644 -3246 -1592
rect -3298 -1712 -3246 -1660
rect -3184 -230 -3132 -178
rect -3184 -298 -3132 -246
rect -3184 -366 -3132 -314
rect -3070 6 -3018 58
rect -3070 -62 -3018 -10
rect -3070 -130 -3018 -78
rect -1692 1323 -1640 1332
rect -1692 1289 -1683 1323
rect -1683 1289 -1649 1323
rect -1649 1289 -1640 1323
rect -1692 1280 -1640 1289
rect -1620 1323 -1568 1332
rect -1620 1289 -1611 1323
rect -1611 1289 -1577 1323
rect -1577 1289 -1568 1323
rect -1620 1280 -1568 1289
rect -1662 456 -1610 508
rect -1594 456 -1542 508
rect 2211 525 2263 534
rect 2211 491 2220 525
rect 2220 491 2254 525
rect 2254 491 2263 525
rect 2211 482 2263 491
rect 2211 453 2263 462
rect 2211 419 2220 453
rect 2220 419 2254 453
rect 2254 419 2263 453
rect 2211 410 2263 419
rect -1692 -19 -1640 -10
rect -1692 -53 -1683 -19
rect -1683 -53 -1649 -19
rect -1649 -53 -1640 -19
rect -1692 -62 -1640 -53
rect -1620 -19 -1568 -10
rect -1620 -53 -1611 -19
rect -1611 -53 -1577 -19
rect -1577 -53 -1568 -19
rect -1620 -62 -1568 -53
rect -1467 -255 -1415 -246
rect -1467 -289 -1458 -255
rect -1458 -289 -1424 -255
rect -1424 -289 -1415 -255
rect -1467 -298 -1415 -289
rect -1395 -255 -1343 -246
rect -1395 -289 -1386 -255
rect -1386 -289 -1352 -255
rect -1352 -289 -1343 -255
rect -1395 -298 -1343 -289
rect -1677 -827 -1625 -818
rect -1677 -861 -1668 -827
rect -1668 -861 -1634 -827
rect -1634 -861 -1625 -827
rect -1677 -870 -1625 -861
rect -1467 -1597 -1415 -1588
rect -1467 -1631 -1458 -1597
rect -1458 -1631 -1424 -1597
rect -1424 -1631 -1415 -1597
rect -1467 -1640 -1415 -1631
rect -1395 -1597 -1343 -1588
rect -1395 -1631 -1386 -1597
rect -1386 -1631 -1352 -1597
rect -1352 -1631 -1343 -1597
rect -1395 -1640 -1343 -1631
<< metal2 >>
rect -3426 1400 -3346 1414
rect -3426 1348 -3412 1400
rect -3360 1348 -3346 1400
rect -3426 1332 -3346 1348
rect -3426 1280 -3412 1332
rect -3360 1326 -3346 1332
rect -1706 1332 -1554 1346
rect -1706 1326 -1692 1332
rect -3360 1286 -1692 1326
rect -3360 1280 -3346 1286
rect -3426 1264 -3346 1280
rect -1706 1280 -1692 1286
rect -1640 1280 -1620 1332
rect -1568 1280 -1554 1332
rect -1706 1266 -1554 1280
rect -3426 1212 -3412 1264
rect -3360 1212 -3346 1264
rect -3426 1198 -3346 1212
rect 2197 534 2277 548
rect -1676 508 -1528 522
rect -1676 456 -1662 508
rect -1610 456 -1594 508
rect -1542 456 -1528 508
rect -1676 442 -1528 456
rect 2197 482 2211 534
rect 2263 492 2277 534
rect 2263 482 2322 492
rect 2197 462 2322 482
rect 2197 410 2211 462
rect 2263 452 2322 462
rect 2263 410 2277 452
rect 2197 396 2277 410
rect -3084 58 -3004 72
rect -3084 6 -3070 58
rect -3018 6 -3004 58
rect -3084 -10 -3004 6
rect -3084 -62 -3070 -10
rect -3018 -16 -3004 -10
rect -1706 -10 -1554 4
rect -1706 -16 -1692 -10
rect -3018 -56 -1692 -16
rect -3018 -62 -3004 -56
rect -3084 -78 -3004 -62
rect -1706 -62 -1692 -56
rect -1640 -62 -1620 -10
rect -1568 -62 -1554 -10
rect -1706 -76 -1554 -62
rect -3084 -130 -3070 -78
rect -3018 -130 -3004 -78
rect -3084 -144 -3004 -130
rect -3198 -178 -3118 -164
rect -3198 -230 -3184 -178
rect -3132 -230 -3118 -178
rect -3198 -246 -3118 -230
rect -3198 -298 -3184 -246
rect -3132 -252 -3118 -246
rect -1481 -246 -1329 -232
rect -1481 -252 -1467 -246
rect -3132 -292 -1467 -252
rect -3132 -298 -3118 -292
rect -3198 -314 -3118 -298
rect -1481 -298 -1467 -292
rect -1415 -298 -1395 -246
rect -1343 -298 -1329 -246
rect -1481 -312 -1329 -298
rect -3198 -366 -3184 -314
rect -3132 -366 -3118 -314
rect -3198 -380 -3118 -366
rect -1691 -818 -1611 -804
rect -1691 -870 -1677 -818
rect -1625 -870 -1611 -818
rect -1691 -884 -1611 -870
rect -3312 -1524 -3232 -1510
rect -3312 -1576 -3298 -1524
rect -3246 -1576 -3232 -1524
rect -3312 -1592 -3232 -1576
rect -3312 -1644 -3298 -1592
rect -3246 -1598 -3232 -1592
rect -1481 -1588 -1329 -1574
rect -1481 -1598 -1467 -1588
rect -3246 -1638 -1467 -1598
rect -3246 -1644 -3232 -1638
rect -3312 -1660 -3232 -1644
rect -1481 -1640 -1467 -1638
rect -1415 -1640 -1395 -1588
rect -1343 -1640 -1329 -1588
rect -1481 -1654 -1329 -1640
rect -3312 -1712 -3298 -1660
rect -3246 -1712 -3232 -1660
rect -3312 -1726 -3232 -1712
use CMOS_AND  CMOS_AND_0
timestamp 1505768678
transform 1 0 690 0 1 640
box -476 -870 476 870
use CMOS_AND  CMOS_AND_1
timestamp 1505768678
transform 1 0 690 0 -1 -948
box -476 -870 476 870
use CMOS_AND  CMOS_AND_2
timestamp 1505768678
transform 1 0 -522 0 -1 -948
box -476 -870 476 870
use CMOS_OR  CMOS_OR_0
timestamp 1505768678
transform 1 0 1902 0 1 640
box -476 -870 476 870
use CMOS_OR  CMOS_OR_1
timestamp 1505768678
transform 1 0 -522 0 1 640
box -476 -870 476 870
use CMOS_XNOR  CMOS_XNOR_0
timestamp 1505768678
transform 1 0 -1907 0 -1 -948
box -649 -870 650 870
use CMOS_XOR  CMOS_XOR_0
timestamp 1505768678
transform 1 0 -2080 0 1 640
box -476 -870 476 870
<< labels >>
flabel metal1 s -2719 -171 -2685 -137 2 FreeSans 2500 0 0 0 GND
port 1 nsew
flabel metal1 s -3644 1408 -3583 1468 2 FreeSans 3126 0 0 0 x0
port 2 nsew
flabel metal1 s -3531 1347 -3470 1407 2 FreeSans 3126 0 0 0 x0_bar
port 3 nsew
flabel metal1 s -3416 1408 -3355 1468 2 FreeSans 3126 0 0 0 x1
port 4 nsew
flabel metal1 s -3302 1347 -3241 1407 2 FreeSans 3126 0 0 0 x1_bar
port 5 nsew
flabel metal1 s -3188 1409 -3127 1469 2 FreeSans 3126 0 0 0 x2
port 6 nsew
flabel metal1 s -3075 1348 -3014 1408 2 FreeSans 3126 0 0 0 x2_bar
port 7 nsew
flabel metal1 s -2960 1409 -2899 1469 2 FreeSans 3126 0 0 0 x3
port 8 nsew
flabel metal1 s -2846 1348 -2785 1408 2 FreeSans 3126 0 0 0 x3_bar
port 9 nsew
flabel metal1 s -2610 1408 -2576 1442 2 FreeSans 2500 0 0 0 VDD
port 10 nsew
flabel metal2 s 2220 491 2254 525 2 FreeSans 2500 0 0 0 s0
port 11 nsew
<< end >>
