**.subckt Diff_LNA_one_part
XM1 net1 net2 net3 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
L1 VDD net4 30n m=1
Vdd VDD GND 1.2
XM2 Vout VDD net1 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
VGS1 net5 GND AC 1 sin(0 0.01 2400MEG 0 0 0)
C1 VDD Vout 65f m=1
L2 net3 GND 1n m=1
R1 VDD Vout 6.9k m=1
R2 net4 Vout 17 m=1
R3 net5 net7 50 m=1
C2 net2 GND 2p m=1
I0 VDD net6 .4m
XM3 net6 net6 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
L3 net8 net2 1n m=1
C4 Vout GND 50f m=1
R4 VDD Vout 20k m=1
R5 net2 net6 10k m=1
C3 net6 GND 1pf m=1
C5 net7 net8 10p m=1
**** begin user architecture code

.lib /research/pdk/open_pdks/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.control
**tran 1ps 100n
ac lin 1k 1E9 5E9
plot db(v(Vout))
**plot v(Vout)
write Diff_LNA_one_part.raw
save all
.endc


**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
