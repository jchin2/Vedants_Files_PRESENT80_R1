* NGSPICE file created from CMOS_s1_flat.ext - technology: sky130A

.subckt CMOS_s1_flat GND x0 x0_bar x1 x1_bar x2 x2_bar x3 x3_bar s1 VDD
X0 s1.t0 a_2442_n779# GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_2592_n1689# CMOS_3in_OR_0/A VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X2 VDD.t3 x3.t0 a_1735_499# VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X3 a_2592_n111# x2_bar.t0 GND.t8 GND.t7 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_2592_499# CMOS_XOR_0/XOR a_2592_n111# GND.t22 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 CMOS_3in_OR_0/A a_1380_n1689# GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_1380_n1689# x3.t1 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X7 a_2742_n1689# CMOS_3in_OR_0/B a_2592_n1689# VDD.t35 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X8 VDD.t39 x2.t0 a_177_499# VDD.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X9 CMOS_XNOR_0/XNOR a_27_n111# VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X10 GND.t9 CMOS_3in_OR_0/A a_2442_n779# GND.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X11 a_2442_n779# CMOS_3in_OR_0/B GND.t30 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 VDD.t37 CMOS_XNOR_0/XNOR a_1380_n1689# VDD.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X13 GND.t11 x0_bar.t0 a_177_n111# GND.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X14 a_27_n111# x2.t1 a_n123_n111# GND.t35 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X15 VDD.t21 x3_bar.t0 a_n328_n1689# VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X16 a_27_n111# x0.t0 a_n123_499# VDD.t28 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X17 CMOS_3in_AND_0/OUT.t0 a_n328_n1689# GND.t29 GND.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 GND.t27 CMOS_3in_AND_0/OUT.t2 a_2442_n779# GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 VDD.t12 x0_bar.t1 a_n328_n1689# VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X20 CMOS_3in_OR_0/B a_2592_499# VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X21 a_1435_n111# x1.t0 GND.t4 GND.t3 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X22 a_1380_n779# x3.t2 GND.t32 GND.t31 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X23 a_1380_n1689# CMOS_XNOR_0/XNOR a_1380_n779# GND.t34 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X24 s1.t1 a_2442_n779# VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X25 a_1435_499# x3_bar.t1 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X26 a_n123_499# x2_bar.t1 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X27 a_n28_n779# x1.t1 a_n178_n779# GND.t25 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X28 a_n328_n1689# x3_bar.t2 a_n28_n779# GND.t20 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X29 VDD.t30 CMOS_XOR_0/XOR a_2592_499# VDD.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X30 a_n328_n1689# x1.t2 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X31 CMOS_3in_OR_0/A a_1380_n1689# VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X32 a_1735_499# x1_bar.t0 CMOS_XOR_0/XOR VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X33 a_177_499# x0_bar.t2 a_27_n111# VDD.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X34 CMOS_XOR_0/XOR x3.t3 a_1435_n111# GND.t2 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X35 a_1735_n111# x3_bar.t3 CMOS_XOR_0/XOR GND.t33 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X36 CMOS_3in_OR_0/B a_2592_499# GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X37 CMOS_3in_AND_0/OUT.t1 a_n328_n1689# VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X38 a_2442_n779# CMOS_3in_AND_0/OUT.t3 a_2742_n1689# VDD.t1 sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X39 a_n123_n111# x0.t1 GND.t24 GND.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X40 a_n178_n779# x0_bar.t3 GND.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X41 a_177_n111# x2_bar.t2 a_27_n111# GND.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X42 a_2592_499# x2_bar.t3 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X43 CMOS_XNOR_0/XNOR a_27_n111# GND.t19 GND.t18 sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X44 GND.t6 x1_bar.t1 a_1735_n111# GND.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X45 CMOS_XOR_0/XOR x1.t3 a_1435_499# VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
R0 GND.n91 GND.t18 2383.33
R1 GND.n92 GND.n91 150.98
R2 GND.n57 GND.t35 150.98
R3 GND.n126 GND.t2 150.98
R4 GND.n45 GND.t23 133.725
R5 GND.n114 GND.t3 133.725
R6 GND.n65 GND.t21 125.098
R7 GND.n134 GND.t33 125.098
R8 GND.n45 GND.t12 103.529
R9 GND.n160 GND.t7 103.529
R10 GND.n114 GND.t31 103.529
R11 GND.n73 GND.t10 99.215
R12 GND.n143 GND.t5 99.215
R13 GND.n83 GND.t28 77.647
R14 GND.n54 GND.t25 77.647
R15 GND.n4 GND.t16 77.647
R16 GND.n169 GND.t22 77.647
R17 GND.n123 GND.t34 77.647
R18 GND.n61 GND.t20 51.764
R19 GND.n13 GND.t14 51.764
R20 GND.n27 GND.t26 51.764
R21 GND.n143 GND.t0 51.764
R22 GND.n38 GND 37.93
R23 GND.n44 GND.t24 30.21
R24 GND.n39 GND.t13 30.21
R25 GND.n82 GND.t29 30.21
R26 GND.n108 GND.t32 30.21
R27 GND.n142 GND.t1 30.21
R28 GND.n26 GND.t27 30.21
R29 GND.n8 GND.t17 30.21
R30 GND.n17 GND.t15 30.21
R31 GND.n155 GND.t8 30.21
R32 GND.n147 GND.t6 30.21
R33 GND.n113 GND.t4 30.21
R34 GND.n96 GND.t19 30.21
R35 GND.n77 GND.t11 30.21
R36 GND.n35 GND.t30 24
R37 GND.n35 GND.t9 24
R38 GND.n105 GND.n104 17.263
R39 GND.n128 GND.n125 11.52
R40 GND.n59 GND.n56 11.52
R41 GND.n2 GND.n1 9.154
R42 GND.n150 GND.n149 9.154
R43 GND.n145 GND.n144 9.154
R44 GND.n144 GND.n143 9.154
R45 GND.n140 GND.n139 9.154
R46 GND.n139 GND.n138 9.154
R47 GND.n136 GND.n135 9.154
R48 GND.n135 GND.n134 9.154
R49 GND.n132 GND.n131 9.154
R50 GND.n131 GND.n130 9.154
R51 GND.n128 GND.n127 9.154
R52 GND.n127 GND.n126 9.154
R53 GND.n125 GND.n124 9.154
R54 GND.n124 GND.n123 9.154
R55 GND.n120 GND.n119 9.154
R56 GND.n119 GND.n118 9.154
R57 GND.n116 GND.n115 9.154
R58 GND.n115 GND.n114 9.154
R59 GND.n111 GND.n110 9.154
R60 GND.n6 GND.n5 9.154
R61 GND.n5 GND.n4 9.154
R62 GND.n11 GND.n10 9.154
R63 GND.n10 GND.n9 9.154
R64 GND.n15 GND.n14 9.154
R65 GND.n14 GND.n13 9.154
R66 GND.n20 GND.n19 9.154
R67 GND.n19 GND.n18 9.154
R68 GND.n24 GND.n23 9.154
R69 GND.n23 GND.n22 9.154
R70 GND.n29 GND.n28 9.154
R71 GND.n28 GND.n27 9.154
R72 GND.n33 GND.n32 9.154
R73 GND.n32 GND.n31 9.154
R74 GND.n171 GND.n170 9.154
R75 GND.n170 GND.n169 9.154
R76 GND.n167 GND.n166 9.154
R77 GND.n166 GND.n165 9.154
R78 GND.n162 GND.n161 9.154
R79 GND.n161 GND.n160 9.154
R80 GND.n158 GND.n157 9.154
R81 GND.n101 GND.n100 9.154
R82 GND.n98 GND.n97 9.154
R83 GND.n94 GND.n93 9.154
R84 GND.n93 GND.n92 9.154
R85 GND.n89 GND.n88 9.154
R86 GND.n88 GND.n87 9.154
R87 GND.n85 GND.n84 9.154
R88 GND.n84 GND.n83 9.154
R89 GND.n80 GND.n79 9.154
R90 GND.n79 GND.n78 9.154
R91 GND.n75 GND.n74 9.154
R92 GND.n74 GND.n73 9.154
R93 GND.n71 GND.n70 9.154
R94 GND.n70 GND.n69 9.154
R95 GND.n67 GND.n66 9.154
R96 GND.n66 GND.n65 9.154
R97 GND.n63 GND.n62 9.154
R98 GND.n62 GND.n61 9.154
R99 GND.n59 GND.n58 9.154
R100 GND.n58 GND.n57 9.154
R101 GND.n56 GND.n55 9.154
R102 GND.n55 GND.n54 9.154
R103 GND.n51 GND.n50 9.154
R104 GND.n50 GND.n49 9.154
R105 GND.n47 GND.n46 9.154
R106 GND.n46 GND.n45 9.154
R107 GND.n42 GND.n41 9.154
R108 GND.n1 GND.n0 8.108
R109 GND.n164 GND.n35 6.21
R110 GND.n39 GND.n38 4.706
R111 GND.n107 GND.n37 4.65
R112 GND.n151 GND.n150 4.65
R113 GND.n146 GND.n145 4.65
R114 GND.n141 GND.n140 4.65
R115 GND.n137 GND.n136 4.65
R116 GND.n133 GND.n132 4.65
R117 GND.n129 GND.n128 4.65
R118 GND.n125 GND.n122 4.65
R119 GND.n121 GND.n120 4.65
R120 GND.n117 GND.n116 4.65
R121 GND.n112 GND.n111 4.65
R122 GND.n153 GND.n152 4.65
R123 GND.n154 GND.n36 4.65
R124 GND.n7 GND.n6 4.65
R125 GND.n12 GND.n11 4.65
R126 GND.n16 GND.n15 4.65
R127 GND.n21 GND.n20 4.65
R128 GND.n25 GND.n24 4.65
R129 GND.n30 GND.n29 4.65
R130 GND.n34 GND.n33 4.65
R131 GND.n172 GND.n171 4.65
R132 GND.n168 GND.n167 4.65
R133 GND.n163 GND.n162 4.65
R134 GND.n159 GND.n158 4.65
R135 GND.n102 GND.n101 4.65
R136 GND.n99 GND.n98 4.65
R137 GND.n95 GND.n94 4.65
R138 GND.n90 GND.n89 4.65
R139 GND.n86 GND.n85 4.65
R140 GND.n81 GND.n80 4.65
R141 GND.n76 GND.n75 4.65
R142 GND.n72 GND.n71 4.65
R143 GND.n68 GND.n67 4.65
R144 GND.n64 GND.n63 4.65
R145 GND.n60 GND.n59 4.65
R146 GND.n56 GND.n53 4.65
R147 GND.n52 GND.n51 4.65
R148 GND.n48 GND.n47 4.65
R149 GND.n43 GND.n42 4.65
R150 GND.n106 GND.n105 4.65
R151 GND.n157 GND.n156 2.759
R152 GND.n3 GND.n2 2.562
R153 GND.n7 GND.n3 1.145
R154 GND.n154 GND.n153 0.525
R155 GND.n104 GND.n103 0.524
R156 GND.n107 GND.n106 0.507
R157 GND.n16 GND.n12 0.09
R158 GND.n25 GND.n21 0.09
R159 GND.n34 GND.n30 0.09
R160 GND.n172 GND.n168 0.09
R161 GND.n163 GND.n159 0.09
R162 GND.n153 GND.n151 0.09
R163 GND.n141 GND.n137 0.09
R164 GND.n137 GND.n133 0.09
R165 GND.n133 GND.n129 0.09
R166 GND.n122 GND.n121 0.09
R167 GND.n121 GND.n117 0.09
R168 GND.n106 GND.n102 0.09
R169 GND.n102 GND.n99 0.09
R170 GND.n95 GND.n90 0.09
R171 GND.n90 GND.n86 0.09
R172 GND.n76 GND.n72 0.09
R173 GND.n72 GND.n68 0.09
R174 GND.n68 GND.n64 0.09
R175 GND.n64 GND.n60 0.09
R176 GND.n53 GND.n52 0.09
R177 GND.n52 GND.n48 0.09
R178 GND.n17 GND.n16 0.078
R179 GND.n30 GND.n26 0.078
R180 GND.n146 GND.n142 0.078
R181 GND.n110 GND.n109 0.074
R182 GND.n41 GND.n40 0.074
R183 GND.n8 GND.n7 0.072
R184 GND.n99 GND.n96 0.071
R185 GND.n86 GND.n82 0.071
R186 CMOS_3in_OR_0/GND GND.n172 0.065
R187 GND.n147 GND.n146 0.065
R188 GND.n122 CMOS_XOR_0/GND 0.065
R189 GND.n77 GND.n76 0.065
R190 GND.n53 GND 0.065
R191 GND.n164 GND.n163 0.063
R192 GND.n155 GND.n154 0.056
R193 GND.n108 GND.n107 0.056
R194 GND.n117 GND.n113 0.055
R195 GND.n48 GND.n44 0.055
R196 GND.n149 GND.n148 0.047
R197 GND.n113 GND.n112 0.035
R198 GND.n44 GND.n43 0.035
R199 GND.n159 GND.n155 0.033
R200 GND.n112 GND.n108 0.033
R201 GND.n43 GND.n39 0.033
R202 GND.n168 GND.n164 0.026
R203 CMOS_3in_OR_0/GND GND.n34 0.025
R204 GND.n151 GND.n147 0.025
R205 GND.n129 CMOS_XOR_0/GND 0.025
R206 GND.n81 GND.n77 0.025
R207 GND.n60 GND 0.025
R208 GND.n96 GND.n95 0.018
R209 GND.n82 GND.n81 0.018
R210 GND.n12 GND.n8 0.017
R211 GND.n21 GND.n17 0.011
R212 GND.n26 GND.n25 0.011
R213 GND.n142 GND.n141 0.011
R214 s1.n2 s1.t1 120.552
R215 s1.n1 s1.t0 98.438
R216 s1 s1.n2 7.84
R217 s1 s1.n1 3.68
R218 s1.n1 s1.n0 3.084
R219 s1.n0 s1 0.374
R220 VDD.n30 VDD.t28 36.141
R221 VDD.n269 VDD.t0 36.141
R222 VDD.n195 VDD.t9 32.01
R223 VDD.n259 VDD.t22 32.01
R224 VDD.n213 VDD.t19 29.945
R225 VDD.n277 VDD.t4 29.945
R226 VDD.n302 VDD.t26 24.782
R227 VDD.n74 VDD.t7 24.782
R228 VDD.n121 VDD.t24 24.782
R229 VDD.n177 VDD.t11 24.782
R230 VDD.n221 VDD.t38 23.75
R231 VDD.n285 VDD.t2 23.75
R232 VDD.n194 VDD.t10 22.029
R233 VDD.n225 VDD.t39 22.029
R234 VDD.n242 VDD.t18 22.029
R235 VDD.n258 VDD.t23 22.029
R236 VDD.n289 VDD.t3 22.029
R237 VDD.n297 VDD.t27 22.029
R238 VDD.n25 VDD.t30 22.029
R239 VDD.n8 VDD.t14 22.029
R240 VDD.n41 VDD.t16 22.029
R241 VDD.n82 VDD.t8 22.029
R242 VDD.n95 VDD.t6 22.029
R243 VDD.n108 VDD.t37 22.029
R244 VDD.n129 VDD.t25 22.029
R245 VDD.n142 VDD.t34 22.029
R246 VDD.n159 VDD.t21 22.029
R247 VDD.n32 VDD.t32 19.7
R248 VDD.n32 VDD.t12 19.7
R249 VDD.n243 VDD.t17 18.586
R250 VDD.n310 VDD.t29 18.586
R251 VDD.n37 VDD.t15 18.586
R252 VDD.n66 VDD.t35 18.586
R253 VDD.n113 VDD.t36 18.586
R254 VDD.n138 VDD.t33 18.586
R255 VDD.n168 VDD.t31 18.586
R256 VDD.n4 VDD.t13 12.391
R257 VDD.n58 VDD.t1 12.391
R258 VDD.n91 VDD.t5 12.391
R259 VDD.n160 VDD.t20 12.391
R260 VDD.n207 VDD.n206 11.52
R261 VDD.n271 VDD.n268 11.52
R262 VDD.n68 VDD.n65 11.52
R263 VDD.n115 VDD.n112 11.52
R264 VDD.n170 VDD.n167 11.52
R265 VDD.n35 VDD.n34 8.855
R266 VDD.n89 VDD.n88 8.855
R267 VDD.n136 VDD.n135 8.855
R268 VDD.n140 VDD.n139 8.855
R269 VDD.n139 VDD.n138 8.855
R270 VDD.n145 VDD.n144 8.855
R271 VDD.n144 VDD.n143 8.855
R272 VDD.n149 VDD.n148 8.855
R273 VDD.n148 VDD.n147 8.855
R274 VDD.n153 VDD.n152 8.855
R275 VDD.n152 VDD.n151 8.855
R276 VDD.n157 VDD.n156 8.855
R277 VDD.n156 VDD.n155 8.855
R278 VDD.n162 VDD.n161 8.855
R279 VDD.n161 VDD.n160 8.855
R280 VDD.n167 VDD.n166 8.855
R281 VDD.n166 VDD.n165 8.855
R282 VDD.n170 VDD.n169 8.855
R283 VDD.n169 VDD.n168 8.855
R284 VDD.n174 VDD.n173 8.855
R285 VDD.n173 VDD.n172 8.855
R286 VDD.n179 VDD.n178 8.855
R287 VDD.n178 VDD.n177 8.855
R288 VDD.n183 VDD.n182 8.855
R289 VDD.n93 VDD.n92 8.855
R290 VDD.n92 VDD.n91 8.855
R291 VDD.n98 VDD.n97 8.855
R292 VDD.n97 VDD.n96 8.855
R293 VDD.n102 VDD.n101 8.855
R294 VDD.n101 VDD.n100 8.855
R295 VDD.n106 VDD.n105 8.855
R296 VDD.n105 VDD.n104 8.855
R297 VDD.n112 VDD.n111 8.855
R298 VDD.n111 VDD.n110 8.855
R299 VDD.n115 VDD.n114 8.855
R300 VDD.n114 VDD.n113 8.855
R301 VDD.n119 VDD.n118 8.855
R302 VDD.n118 VDD.n117 8.855
R303 VDD.n123 VDD.n122 8.855
R304 VDD.n122 VDD.n121 8.855
R305 VDD.n127 VDD.n126 8.855
R306 VDD.n39 VDD.n38 8.855
R307 VDD.n38 VDD.n37 8.855
R308 VDD.n44 VDD.n43 8.855
R309 VDD.n43 VDD.n42 8.855
R310 VDD.n48 VDD.n47 8.855
R311 VDD.n47 VDD.n46 8.855
R312 VDD.n52 VDD.n51 8.855
R313 VDD.n51 VDD.n50 8.855
R314 VDD.n56 VDD.n55 8.855
R315 VDD.n55 VDD.n54 8.855
R316 VDD.n60 VDD.n59 8.855
R317 VDD.n59 VDD.n58 8.855
R318 VDD.n65 VDD.n64 8.855
R319 VDD.n64 VDD.n63 8.855
R320 VDD.n68 VDD.n67 8.855
R321 VDD.n67 VDD.n66 8.855
R322 VDD.n72 VDD.n71 8.855
R323 VDD.n71 VDD.n70 8.855
R324 VDD.n76 VDD.n75 8.855
R325 VDD.n75 VDD.n74 8.855
R326 VDD.n80 VDD.n79 8.855
R327 VDD.n2 VDD.n1 8.855
R328 VDD.n6 VDD.n5 8.855
R329 VDD.n5 VDD.n4 8.855
R330 VDD.n11 VDD.n10 8.855
R331 VDD.n10 VDD.n9 8.855
R332 VDD.n15 VDD.n14 8.855
R333 VDD.n14 VDD.n13 8.855
R334 VDD.n19 VDD.n18 8.855
R335 VDD.n18 VDD.n17 8.855
R336 VDD.n23 VDD.n22 8.855
R337 VDD.n22 VDD.n21 8.855
R338 VDD.n312 VDD.n311 8.855
R339 VDD.n311 VDD.n310 8.855
R340 VDD.n308 VDD.n307 8.855
R341 VDD.n307 VDD.n306 8.855
R342 VDD.n304 VDD.n303 8.855
R343 VDD.n303 VDD.n302 8.855
R344 VDD.n300 VDD.n299 8.855
R345 VDD.n292 VDD.n291 8.855
R346 VDD.n287 VDD.n286 8.855
R347 VDD.n286 VDD.n285 8.855
R348 VDD.n283 VDD.n282 8.855
R349 VDD.n282 VDD.n281 8.855
R350 VDD.n279 VDD.n278 8.855
R351 VDD.n278 VDD.n277 8.855
R352 VDD.n275 VDD.n274 8.855
R353 VDD.n274 VDD.n273 8.855
R354 VDD.n271 VDD.n270 8.855
R355 VDD.n270 VDD.n269 8.855
R356 VDD.n268 VDD.n28 8.855
R357 VDD.n28 VDD.n27 8.855
R358 VDD.n265 VDD.n264 8.855
R359 VDD.n264 VDD.n263 8.855
R360 VDD.n261 VDD.n260 8.855
R361 VDD.n260 VDD.n259 8.855
R362 VDD.n256 VDD.n255 8.855
R363 VDD.n249 VDD.n248 8.855
R364 VDD.n245 VDD.n244 8.855
R365 VDD.n244 VDD.n243 8.855
R366 VDD.n240 VDD.n239 8.855
R367 VDD.n239 VDD.n238 8.855
R368 VDD.n236 VDD.n235 8.855
R369 VDD.n235 VDD.n234 8.855
R370 VDD.n232 VDD.n231 8.855
R371 VDD.n231 VDD.n230 8.855
R372 VDD.n228 VDD.n227 8.855
R373 VDD.n227 VDD.n226 8.855
R374 VDD.n223 VDD.n222 8.855
R375 VDD.n222 VDD.n221 8.855
R376 VDD.n219 VDD.n218 8.855
R377 VDD.n218 VDD.n217 8.855
R378 VDD.n215 VDD.n214 8.855
R379 VDD.n214 VDD.n213 8.855
R380 VDD.n211 VDD.n210 8.855
R381 VDD.n210 VDD.n209 8.855
R382 VDD.n207 VDD.n31 8.855
R383 VDD.n31 VDD.n30 8.855
R384 VDD.n206 VDD.n205 8.855
R385 VDD.n205 VDD.n204 8.855
R386 VDD.n201 VDD.n200 8.855
R387 VDD.n200 VDD.n199 8.855
R388 VDD.n197 VDD.n196 8.855
R389 VDD.n196 VDD.n195 8.855
R390 VDD.n192 VDD.n191 8.855
R391 VDD.n187 VDD.n186 4.91
R392 VDD.n186 VDD.n185 4.65
R393 VDD.n137 VDD.n136 4.65
R394 VDD.n141 VDD.n140 4.65
R395 VDD.n146 VDD.n145 4.65
R396 VDD.n150 VDD.n149 4.65
R397 VDD.n154 VDD.n153 4.65
R398 VDD.n158 VDD.n157 4.65
R399 VDD.n163 VDD.n162 4.65
R400 VDD.n167 VDD.n164 4.65
R401 VDD.n171 VDD.n170 4.65
R402 VDD.n175 VDD.n174 4.65
R403 VDD.n180 VDD.n179 4.65
R404 VDD.n184 VDD.n183 4.65
R405 VDD.n133 VDD.n132 4.65
R406 VDD.n131 VDD.n130 4.65
R407 VDD.n90 VDD.n89 4.65
R408 VDD.n94 VDD.n93 4.65
R409 VDD.n99 VDD.n98 4.65
R410 VDD.n103 VDD.n102 4.65
R411 VDD.n107 VDD.n106 4.65
R412 VDD.n112 VDD.n109 4.65
R413 VDD.n116 VDD.n115 4.65
R414 VDD.n120 VDD.n119 4.65
R415 VDD.n124 VDD.n123 4.65
R416 VDD.n128 VDD.n127 4.65
R417 VDD.n86 VDD.n85 4.65
R418 VDD.n84 VDD.n83 4.65
R419 VDD.n40 VDD.n39 4.65
R420 VDD.n45 VDD.n44 4.65
R421 VDD.n49 VDD.n48 4.65
R422 VDD.n53 VDD.n52 4.65
R423 VDD.n57 VDD.n56 4.65
R424 VDD.n61 VDD.n60 4.65
R425 VDD.n65 VDD.n62 4.65
R426 VDD.n69 VDD.n68 4.65
R427 VDD.n73 VDD.n72 4.65
R428 VDD.n77 VDD.n76 4.65
R429 VDD.n81 VDD.n80 4.65
R430 VDD.n7 VDD.n6 4.65
R431 VDD.n12 VDD.n11 4.65
R432 VDD.n16 VDD.n15 4.65
R433 VDD.n20 VDD.n19 4.65
R434 VDD.n24 VDD.n23 4.65
R435 VDD.n313 VDD.n312 4.65
R436 VDD.n309 VDD.n308 4.65
R437 VDD.n305 VDD.n304 4.65
R438 VDD.n301 VDD.n300 4.65
R439 VDD.n296 VDD.n295 4.65
R440 VDD.n294 VDD.n26 4.65
R441 VDD.n293 VDD.n292 4.65
R442 VDD.n288 VDD.n287 4.65
R443 VDD.n284 VDD.n283 4.65
R444 VDD.n280 VDD.n279 4.65
R445 VDD.n276 VDD.n275 4.65
R446 VDD.n272 VDD.n271 4.65
R447 VDD.n268 VDD.n267 4.65
R448 VDD.n266 VDD.n265 4.65
R449 VDD.n262 VDD.n261 4.65
R450 VDD.n257 VDD.n256 4.65
R451 VDD.n253 VDD.n252 4.65
R452 VDD.n251 VDD.n29 4.65
R453 VDD.n250 VDD.n249 4.65
R454 VDD.n246 VDD.n245 4.65
R455 VDD.n241 VDD.n240 4.65
R456 VDD.n237 VDD.n236 4.65
R457 VDD.n233 VDD.n232 4.65
R458 VDD.n229 VDD.n228 4.65
R459 VDD.n224 VDD.n223 4.65
R460 VDD.n220 VDD.n219 4.65
R461 VDD.n216 VDD.n215 4.65
R462 VDD.n212 VDD.n211 4.65
R463 VDD.n208 VDD.n207 4.65
R464 VDD.n206 VDD.n203 4.65
R465 VDD.n202 VDD.n201 4.65
R466 VDD.n198 VDD.n197 4.65
R467 VDD.n193 VDD.n192 4.65
R468 VDD.n189 VDD.n188 4.65
R469 VDD.n1 VDD.n0 4.288
R470 VDD.n291 VDD.n290 4.288
R471 VDD.n248 VDD.n247 4.288
R472 VDD.n34 VDD.n33 4.288
R473 VDD.n88 VDD.n87 4.288
R474 VDD.n135 VDD.n134 4.288
R475 VDD.n182 VDD.n181 4.288
R476 VDD.n126 VDD.n125 4.288
R477 VDD.n79 VDD.n78 4.288
R478 VDD.n299 VDD.n298 4.288
R479 VDD.n255 VDD.n254 4.288
R480 VDD.n191 VDD.n190 4.288
R481 VDD.n3 VDD.n2 2.562
R482 VDD.n36 VDD.n35 2.562
R483 VDD.n176 VDD.n32 2.329
R484 VDD.n7 VDD.n3 1.145
R485 VDD.n40 VDD.n36 1.145
R486 VDD.n133 VDD.n131 0.777
R487 VDD.n86 VDD.n84 0.525
R488 VDD.n296 VDD.n294 0.525
R489 VDD.n253 VDD.n251 0.507
R490 VDD.n189 VDD.n187 0.135
R491 VDD.n49 VDD.n45 0.09
R492 VDD.n53 VDD.n49 0.09
R493 VDD.n57 VDD.n53 0.09
R494 VDD.n61 VDD.n57 0.09
R495 VDD.n62 VDD.n61 0.09
R496 VDD.n73 VDD.n69 0.09
R497 VDD.n77 VDD.n73 0.09
R498 VDD.n81 VDD.n77 0.09
R499 VDD.n90 VDD.n86 0.09
R500 VDD.n94 VDD.n90 0.09
R501 VDD.n103 VDD.n99 0.09
R502 VDD.n107 VDD.n103 0.09
R503 VDD.n109 VDD.n107 0.09
R504 VDD.n120 VDD.n116 0.09
R505 VDD.n124 VDD.n120 0.09
R506 VDD.n128 VDD.n124 0.09
R507 VDD.n137 VDD.n133 0.09
R508 VDD.n141 VDD.n137 0.09
R509 VDD.n150 VDD.n146 0.09
R510 VDD.n154 VDD.n150 0.09
R511 VDD.n158 VDD.n154 0.09
R512 VDD.n164 VDD.n163 0.09
R513 VDD.n175 VDD.n171 0.09
R514 VDD.n184 VDD.n180 0.09
R515 VDD.n186 VDD.n184 0.09
R516 VDD.n16 VDD.n12 0.09
R517 VDD.n20 VDD.n16 0.09
R518 VDD.n24 VDD.n20 0.09
R519 VDD.n313 VDD.n309 0.09
R520 VDD.n309 VDD.n305 0.09
R521 VDD.n305 VDD.n301 0.09
R522 VDD.n294 VDD.n293 0.09
R523 VDD.n288 VDD.n284 0.09
R524 VDD.n284 VDD.n280 0.09
R525 VDD.n280 VDD.n276 0.09
R526 VDD.n276 VDD.n272 0.09
R527 VDD.n267 VDD.n266 0.09
R528 VDD.n266 VDD.n262 0.09
R529 VDD.n257 VDD.n253 0.09
R530 VDD.n251 VDD.n250 0.09
R531 VDD.n250 VDD.n246 0.09
R532 VDD.n241 VDD.n237 0.09
R533 VDD.n237 VDD.n233 0.09
R534 VDD.n233 VDD.n229 0.09
R535 VDD.n224 VDD.n220 0.09
R536 VDD.n220 VDD.n216 0.09
R537 VDD.n216 VDD.n212 0.09
R538 VDD.n212 VDD.n208 0.09
R539 VDD.n203 VDD.n202 0.09
R540 VDD.n202 VDD.n198 0.09
R541 VDD.n193 VDD.n189 0.09
R542 VDD.n95 VDD.n94 0.078
R543 VDD.n163 VDD.n159 0.078
R544 VDD.n8 VDD.n7 0.078
R545 VDD.n142 VDD.n141 0.071
R546 VDD.n246 VDD.n242 0.071
R547 VDD.n41 VDD.n40 0.07
R548 VDD.n69 CMOS_3in_OR_0/VDD 0.065
R549 VDD.n116 CMOS_AND_1/VDD 0.065
R550 VDD.n171 CMOS_3in_AND_0/VDD 0.065
R551 CMOS_AND_0/VDD VDD.n313 0.065
R552 VDD.n289 VDD.n288 0.065
R553 VDD.n267 CMOS_XOR_0/VDD 0.065
R554 VDD.n225 VDD.n224 0.065
R555 VDD.n203 VDD 0.065
R556 VDD.n180 VDD.n176 0.063
R557 VDD.n84 VDD.n82 0.056
R558 VDD.n131 VDD.n129 0.056
R559 VDD.n297 VDD.n296 0.056
R560 VDD.n262 VDD.n258 0.055
R561 VDD.n198 VDD.n194 0.055
R562 VDD.n258 VDD.n257 0.035
R563 VDD.n194 VDD.n193 0.035
R564 VDD.n82 VDD.n81 0.033
R565 VDD.n129 VDD.n128 0.033
R566 VDD.n301 VDD.n297 0.033
R567 VDD.n187 VDD 0.027
R568 VDD.n176 VDD.n175 0.026
R569 VDD.n62 CMOS_3in_OR_0/VDD 0.025
R570 VDD.n164 CMOS_3in_AND_0/VDD 0.025
R571 VDD.n293 VDD.n289 0.025
R572 VDD.n272 CMOS_XOR_0/VDD 0.025
R573 VDD.n229 VDD.n225 0.025
R574 VDD.n208 VDD 0.025
R575 VDD.n45 VDD.n41 0.02
R576 VDD.n146 VDD.n142 0.018
R577 VDD.n242 VDD.n241 0.018
R578 VDD.n109 VDD.n108 0.017
R579 VDD.n25 VDD.n24 0.017
R580 VDD.n99 VDD.n95 0.011
R581 VDD.n159 VDD.n158 0.011
R582 VDD.n12 VDD.n8 0.011
R583 VDD.n108 CMOS_AND_1/VDD 0.007
R584 CMOS_AND_0/VDD VDD.n25 0.007
R585 x3.t0 x3.t3 924.95
R586 x3 x3.t0 633.02
R587 x3.n0 x3.t2 579.86
R588 x3.n0 x3.t1 547.727
R589 x3 x3.n2 42.894
R590 x3.n2 x3.n1 14.2
R591 x3.n1 x3.n0 8.764
R592 x3.n1 CMOS_AND_1/B 2.72
R593 x3.n2 x3 0.157
R594 x2_bar.n0 x2_bar.t1 683.32
R595 x2_bar.n1 x2_bar.t0 579.86
R596 x2_bar.n1 x2_bar.t3 547.727
R597 x2_bar.n0 x2_bar.t2 528.72
R598 x2_bar x2_bar.n3 198.92
R599 x2_bar.n3 x2_bar.n2 19.691
R600 x2_bar.n2 x2_bar.n1 8.764
R601 x2_bar x2_bar.n0 3.68
R602 x2_bar.n2 CMOS_AND_0/B 2.72
R603 x2_bar.n3 x2_bar 1.205
R604 x2.t0 x2.t1 924.95
R605 x2 x2.t0 633.02
R606 x0_bar.t0 x0_bar.t2 1345.61
R607 x0_bar.n0 x0_bar.t3 570.366
R608 x0_bar.n0 x0_bar.t1 570.366
R609 x0_bar x0_bar.n1 507.08
R610 x0_bar x0_bar.t0 392.02
R611 x0_bar.n1 CMOS_3in_AND_0/C 339.092
R612 CMOS_3in_AND_0/C x0_bar.n0 78.72
R613 x0_bar.n1 x0_bar 2.166
R614 x3_bar.t0 x3_bar.t2 1221.07
R615 x3_bar.n0 x3_bar.t0 630.3
R616 x3_bar.n2 x3_bar.t1 616.084
R617 x3_bar.n2 x3_bar.t3 528.72
R618 x3_bar.n1 x3_bar.n0 41.005
R619 x3_bar.n2 x3_bar.n1 12.411
R620 x3_bar x3_bar.n2 3.68
R621 x3_bar.n0 CMOS_3in_AND_0/A 2.72
R622 x3_bar.n1 x3_bar 2.167
R623 x0.n0 x0.t0 993.097
R624 x0.n0 x0.t1 356.59
R625 x0 x0.n0 78.72
R626 CMOS_3in_AND_0/OUT.t3 CMOS_3in_AND_0/OUT.t2 1221.07
R627 CMOS_3in_OR_0/C CMOS_3in_AND_0/OUT.n0 787.238
R628 CMOS_3in_OR_0/C CMOS_3in_AND_0/OUT.t3 633.02
R629 CMOS_3in_AND_0/OUT CMOS_3in_AND_0/OUT.t0 117.958
R630 CMOS_3in_AND_0/OUT.n0 CMOS_3in_AND_0/OUT 91.717
R631 CMOS_3in_AND_0/OUT.n0 CMOS_3in_AND_0/OUT.t1 45.156
R632 x1.t1 x1.t2 1221.07
R633 x1.n0 x1.t3 993.097
R634 x1.n2 x1.t1 389.3
R635 x1.n0 x1.t0 356.59
R636 CMOS_3in_AND_0/B x1 355.219
R637 x1.n2 x1.n1 211.591
R638 x1.n1 x1.n0 8.764
R639 x1.n1 x1 2.72
R640 CMOS_3in_AND_0/B x1.n2 2.72
R641 x1_bar.t1 x1_bar.t0 1345.61
R642 x1_bar x1_bar.t1 392.02
C0 a_1435_n111# x1_bar 0.00fF
C1 s1 CMOS_3in_OR_0/A 0.01fF
C2 a_1735_499# CMOS_3in_OR_0/B 0.00fF
C3 a_n178_n779# x2 0.00fF
C4 VDD x3_bar 1.54fF
C5 a_n178_n779# CMOS_3in_AND_0/OUT 0.00fF
C6 a_n28_n779# x0_bar 0.00fF
C7 CMOS_XNOR_0/XNOR x0 0.00fF
C8 a_n123_n111# VDD 0.01fF
C9 s1 x1_bar 0.00fF
C10 a_1735_n111# x2_bar 0.01fF
C11 CMOS_XOR_0/XOR x3 0.35fF
C12 CMOS_XNOR_0/XNOR a_n123_499# 0.00fF
C13 a_177_n111# x0_bar 0.01fF
C14 a_1380_n1689# x2_bar 0.03fF
C15 a_n28_n779# a_n328_n1689# 0.01fF
C16 CMOS_XOR_0/XOR a_27_n111# 0.04fF
C17 a_1735_n111# VDD 0.01fF
C18 a_177_499# x0 0.00fF
C19 CMOS_XNOR_0/XNOR x3 0.09fF
C20 CMOS_XNOR_0/XNOR a_1380_n779# 0.01fF
C21 CMOS_3in_OR_0/B x1 0.00fF
C22 a_2592_499# x2_bar 0.05fF
C23 a_n28_n779# x3_bar 0.00fF
C24 a_2442_n779# CMOS_3in_AND_0/OUT 0.05fF
C25 x0 x2_bar 0.27fF
C26 a_1380_n1689# VDD 0.75fF
C27 a_177_n111# a_n328_n1689# 0.00fF
C28 CMOS_XNOR_0/XNOR a_27_n111# 0.08fF
C29 a_1735_499# x3_bar 0.00fF
C30 CMOS_XOR_0/XOR CMOS_3in_OR_0/A 0.02fF
C31 x1 x0_bar 2.62fF
C32 s1 a_2442_n779# 0.06fF
C33 a_2592_499# VDD 0.78fF
C34 a_177_499# x3 0.01fF
C35 a_n123_499# x2_bar 0.01fF
C36 VDD x0 0.09fF
C37 a_177_n111# x3_bar 0.01fF
C38 CMOS_XOR_0/XOR a_1435_499# 0.02fF
C39 CMOS_XOR_0/XOR x1_bar 0.14fF
C40 a_2592_n111# a_2442_n779# 0.00fF
C41 CMOS_3in_AND_0/OUT x2 0.00fF
C42 CMOS_XNOR_0/XNOR CMOS_3in_OR_0/A 0.00fF
C43 a_177_499# a_27_n111# 0.03fF
C44 x2_bar x3 2.91fF
C45 a_1380_n1689# a_2592_n1689# 0.00fF
C46 a_n123_499# VDD 0.05fF
C47 x1 a_n328_n1689# 0.13fF
C48 a_1380_n779# x2_bar 0.01fF
C49 a_n28_n779# a_1380_n1689# 0.00fF
C50 CMOS_XNOR_0/XNOR x1_bar 0.04fF
C51 a_1435_499# CMOS_XNOR_0/XNOR 0.01fF
C52 a_27_n111# x2_bar 0.18fF
C53 s1 CMOS_3in_AND_0/OUT 0.00fF
C54 a_2592_499# a_2592_n1689# 0.00fF
C55 VDD x3 1.93fF
C56 x1 x3_bar 0.38fF
C57 a_1735_499# a_1380_n1689# 0.00fF
C58 a_1380_n779# VDD 0.00fF
C59 a_n123_n111# x1 0.00fF
C60 a_n28_n779# x0 0.00fF
C61 a_27_n111# VDD 1.04fF
C62 a_1735_499# a_2592_499# 0.00fF
C63 a_177_499# x1_bar 0.00fF
C64 CMOS_3in_OR_0/A x2_bar 0.03fF
C65 CMOS_XOR_0/XOR a_2442_n779# 0.01fF
C66 a_1735_n111# x1 0.00fF
C67 a_177_n111# x0 0.00fF
C68 a_1435_499# x2_bar 0.00fF
C69 x1_bar x2_bar 3.79fF
C70 a_2742_n1689# VDD 0.06fF
C71 CMOS_3in_OR_0/A VDD 0.52fF
C72 a_n328_n1689# x0_bar 0.08fF
C73 CMOS_3in_OR_0/B x3_bar 0.00fF
C74 a_n178_n779# x2_bar 0.01fF
C75 a_n28_n779# x3 0.00fF
C76 CMOS_XNOR_0/XNOR a_2442_n779# 0.00fF
C77 x1 a_1380_n1689# 0.00fF
C78 CMOS_XOR_0/XOR x2 0.00fF
C79 a_1735_499# x3 0.03fF
C80 x1_bar VDD 0.20fF
C81 a_1435_499# VDD 0.06fF
C82 CMOS_XOR_0/XOR CMOS_3in_AND_0/OUT 0.00fF
C83 x0_bar x3_bar 0.13fF
C84 CMOS_XOR_0/XOR a_1435_n111# 0.01fF
C85 a_n28_n779# a_27_n111# 0.00fF
C86 a_n123_n111# x0_bar 0.01fF
C87 a_n178_n779# VDD 0.01fF
C88 a_2592_499# x1 0.00fF
C89 a_177_n111# x3 0.00fF
C90 x1 x0 0.03fF
C91 CMOS_3in_OR_0/B a_1735_n111# 0.00fF
C92 a_2592_n1689# CMOS_3in_OR_0/A 0.01fF
C93 CMOS_XNOR_0/XNOR x2 0.01fF
C94 CMOS_XNOR_0/XNOR CMOS_3in_AND_0/OUT 0.02fF
C95 a_177_n111# a_27_n111# 0.01fF
C96 a_1435_n111# CMOS_XNOR_0/XNOR 0.00fF
C97 CMOS_XOR_0/XOR a_2592_n111# 0.01fF
C98 a_n328_n1689# x3_bar 0.14fF
C99 a_n123_499# x1 0.00fF
C100 a_n123_n111# a_n328_n1689# 0.00fF
C101 a_2442_n779# x2_bar 0.02fF
C102 CMOS_3in_OR_0/B a_1380_n1689# 0.00fF
C103 a_n28_n779# x1_bar 0.00fF
C104 x1 x3 0.21fF
C105 a_177_499# x2 0.03fF
C106 a_n123_n111# x3_bar 0.01fF
C107 a_1380_n1689# x0_bar 0.00fF
C108 a_1380_n779# x1 0.00fF
C109 a_2592_499# CMOS_3in_OR_0/B 0.08fF
C110 a_2442_n779# VDD 0.54fF
C111 a_1735_499# x1_bar 0.01fF
C112 x1 a_27_n111# 0.04fF
C113 x2 x2_bar 3.61fF
C114 a_177_n111# x1_bar 0.00fF
C115 CMOS_3in_AND_0/OUT x2_bar 0.03fF
C116 x0_bar x0 3.07fF
C117 a_1435_n111# x2_bar 0.01fF
C118 a_1735_n111# x3_bar 0.00fF
C119 a_1380_n1689# a_n328_n1689# 0.00fF
C120 x2 VDD 1.01fF
C121 s1 x2_bar 0.00fF
C122 a_n123_499# x0_bar 0.01fF
C123 CMOS_3in_OR_0/B x3 0.00fF
C124 CMOS_3in_AND_0/OUT VDD 2.10fF
C125 a_2442_n779# a_2592_n1689# 0.02fF
C126 a_1435_n111# VDD 0.01fF
C127 a_1380_n1689# x3_bar 0.00fF
C128 a_2592_n111# x2_bar 0.01fF
C129 a_n328_n1689# x0 0.01fF
C130 x1_bar x1 3.48fF
C131 CMOS_XOR_0/XOR CMOS_XNOR_0/XNOR 0.05fF
C132 x0_bar x3 0.10fF
C133 s1 VDD 0.37fF
C134 a_2592_499# x3_bar 0.00fF
C135 x1 a_n178_n779# 0.01fF
C136 x0 x3_bar 0.05fF
C137 a_2592_n111# VDD 0.01fF
C138 a_n123_n111# x0 0.00fF
C139 a_27_n111# x0_bar 0.11fF
C140 CMOS_3in_AND_0/OUT a_2592_n1689# 0.01fF
C141 a_1735_n111# a_1380_n1689# 0.00fF
C142 CMOS_3in_OR_0/B a_2742_n1689# 0.00fF
C143 CMOS_3in_OR_0/B CMOS_3in_OR_0/A 0.04fF
C144 a_n28_n779# x2 0.00fF
C145 a_n328_n1689# x3 0.10fF
C146 CMOS_XOR_0/XOR a_177_499# 0.00fF
C147 a_n123_499# x3_bar 0.01fF
C148 a_n28_n779# CMOS_3in_AND_0/OUT 0.00fF
C149 a_1380_n779# a_n328_n1689# 0.00fF
C150 s1 a_2592_n1689# 0.00fF
C151 a_2592_499# a_1735_n111# 0.00fF
C152 a_1435_499# CMOS_3in_OR_0/B 0.00fF
C153 CMOS_3in_OR_0/B x1_bar 0.00fF
C154 a_n328_n1689# a_27_n111# 0.01fF
C155 CMOS_XOR_0/XOR x2_bar 0.24fF
C156 x3 x3_bar 3.31fF
C157 a_n123_n111# x3 0.00fF
C158 a_177_n111# x2 0.01fF
C159 a_1380_n779# x3_bar 0.00fF
C160 CMOS_XNOR_0/XNOR a_177_499# 0.00fF
C161 x1_bar x0_bar 0.08fF
C162 a_27_n111# x3_bar 0.25fF
C163 CMOS_XOR_0/XOR VDD 1.03fF
C164 a_n123_n111# a_27_n111# 0.01fF
C165 a_n178_n779# x0_bar 0.00fF
C166 CMOS_XNOR_0/XNOR x2_bar 0.04fF
C167 CMOS_3in_OR_0/A a_n328_n1689# 0.00fF
C168 a_1735_n111# x3 0.01fF
C169 x1 x2 0.04fF
C170 x1_bar a_n328_n1689# 0.02fF
C171 CMOS_XNOR_0/XNOR VDD 0.51fF
C172 x1 CMOS_3in_AND_0/OUT 0.09fF
C173 a_1435_n111# x1 0.00fF
C174 a_n178_n779# a_n328_n1689# 0.01fF
C175 a_1380_n1689# x3 0.06fF
C176 a_177_499# x2_bar 0.01fF
C177 CMOS_3in_OR_0/B a_2442_n779# 0.12fF
C178 a_n123_499# x0 0.00fF
C179 a_1380_n779# a_1380_n1689# 0.01fF
C180 CMOS_XOR_0/XOR a_2592_n1689# 0.00fF
C181 x1_bar x3_bar 0.34fF
C182 a_1435_499# x3_bar 0.01fF
C183 a_n123_n111# x1_bar 0.00fF
C184 a_2592_499# x3 0.01fF
C185 a_n178_n779# x3_bar 0.00fF
C186 x0 x3 0.04fF
C187 x1 a_2592_n111# 0.00fF
C188 a_177_499# VDD 0.05fF
C189 a_1735_499# CMOS_XOR_0/XOR 0.03fF
C190 a_27_n111# x0 0.02fF
C191 a_n123_499# x3 0.01fF
C192 CMOS_3in_OR_0/B CMOS_3in_AND_0/OUT 0.06fF
C193 a_177_n111# CMOS_XOR_0/XOR 0.00fF
C194 VDD x2_bar 0.80fF
C195 a_2742_n1689# a_1380_n1689# 0.00fF
C196 a_1435_n111# CMOS_3in_OR_0/B 0.00fF
C197 a_1735_n111# x1_bar 0.01fF
C198 a_1380_n1689# CMOS_3in_OR_0/A 0.07fF
C199 a_1735_499# CMOS_XNOR_0/XNOR 0.00fF
C200 x2 x0_bar 0.12fF
C201 a_n123_499# a_27_n111# 0.02fF
C202 CMOS_3in_AND_0/OUT x0_bar 0.00fF
C203 s1 CMOS_3in_OR_0/B 0.04fF
C204 a_2592_499# a_2742_n1689# 0.00fF
C205 x1_bar a_1380_n1689# 0.01fF
C206 a_1435_499# a_1380_n1689# 0.00fF
C207 a_177_n111# CMOS_XNOR_0/XNOR 0.00fF
C208 CMOS_3in_OR_0/B a_2592_n111# 0.01fF
C209 a_27_n111# x3 0.17fF
C210 a_2592_499# x1_bar 0.00fF
C211 a_2592_499# a_1435_499# 0.00fF
C212 CMOS_XOR_0/XOR x1 0.09fF
C213 x1_bar x0 0.04fF
C214 x2 a_n328_n1689# 0.02fF
C215 CMOS_3in_AND_0/OUT a_n328_n1689# 0.05fF
C216 a_n28_n779# x2_bar 0.01fF
C217 a_n178_n779# x0 0.00fF
C218 x2 x3_bar 0.09fF
C219 a_1735_499# x2_bar 0.00fF
C220 a_2592_n1689# VDD 0.06fF
C221 a_n123_499# x1_bar 0.00fF
C222 CMOS_3in_OR_0/A x3 0.02fF
C223 CMOS_XNOR_0/XNOR x1 0.08fF
C224 a_n123_n111# x2 0.01fF
C225 CMOS_3in_AND_0/OUT x3_bar 0.02fF
C226 a_1435_n111# x3_bar 0.01fF
C227 a_1380_n779# CMOS_3in_OR_0/A 0.00fF
C228 a_n28_n779# VDD 0.01fF
C229 a_177_n111# x2_bar 0.01fF
C230 x1_bar x3 0.12fF
C231 a_1435_499# x3 0.01fF
C232 a_2442_n779# a_1380_n1689# 0.01fF
C233 a_1735_499# VDD 0.06fF
C234 a_1380_n779# x1_bar 0.00fF
C235 CMOS_XOR_0/XOR CMOS_3in_OR_0/B 0.04fF
C236 a_n178_n779# x3 0.00fF
C237 a_2592_n111# x3_bar 0.00fF
C238 a_177_499# x1 0.00fF
C239 a_177_n111# VDD 0.01fF
C240 x1_bar a_27_n111# 0.04fF
C241 a_1435_499# a_27_n111# 0.00fF
C242 a_2592_499# a_2442_n779# 0.01fF
C243 CMOS_XOR_0/XOR x0_bar 0.00fF
C244 a_2742_n1689# CMOS_3in_OR_0/A 0.00fF
C245 CMOS_XNOR_0/XNOR CMOS_3in_OR_0/B 0.01fF
C246 x1 x2_bar 0.08fF
C247 CMOS_3in_AND_0/OUT a_1380_n1689# 0.10fF
C248 a_1435_n111# a_1380_n1689# 0.00fF
C249 x1_bar CMOS_3in_OR_0/A 0.00fF
C250 CMOS_XNOR_0/XNOR x0_bar 0.01fF
C251 x2 x0 0.15fF
C252 x1 VDD 0.35fF
C253 a_2592_499# CMOS_3in_AND_0/OUT 0.00fF
C254 s1 a_1380_n1689# 0.00fF
C255 a_2592_499# a_1435_n111# 0.00fF
C256 a_2442_n779# x3 0.00fF
C257 a_1435_499# x1_bar 0.00fF
C258 a_1380_n779# a_2442_n779# 0.00fF
C259 CMOS_XOR_0/XOR x3_bar 0.15fF
C260 x1_bar a_n178_n779# 0.00fF
C261 a_n123_499# x2 0.02fF
C262 CMOS_XNOR_0/XNOR a_n328_n1689# 0.00fF
C263 CMOS_3in_OR_0/B x2_bar 0.06fF
C264 a_177_499# x0_bar 0.01fF
C265 a_2592_499# a_2592_n111# 0.01fF
C266 x2 x3 0.11fF
C267 CMOS_XNOR_0/XNOR x3_bar 0.07fF
C268 CMOS_3in_AND_0/OUT x3 0.05fF
C269 x0_bar x2_bar 0.18fF
C270 a_1435_n111# x3 0.01fF
C271 CMOS_XNOR_0/XNOR a_n123_n111# 0.00fF
C272 CMOS_3in_OR_0/B VDD 0.49fF
C273 a_1380_n779# CMOS_3in_AND_0/OUT 0.01fF
C274 a_2742_n1689# a_2442_n779# 0.02fF
C275 CMOS_XOR_0/XOR a_1735_n111# 0.01fF
C276 a_n28_n779# x1 0.01fF
C277 a_2442_n779# CMOS_3in_OR_0/A 0.10fF
C278 a_177_499# a_n328_n1689# 0.00fF
C279 x2 a_27_n111# 0.34fF
C280 CMOS_3in_AND_0/OUT a_27_n111# 0.01fF
C281 a_1435_n111# a_27_n111# 0.00fF
C282 x0_bar VDD 0.28fF
C283 x1_bar a_2442_n779# 0.00fF
C284 CMOS_XOR_0/XOR a_1380_n1689# 0.01fF
C285 a_n328_n1689# x2_bar 0.06fF
C286 a_177_499# x3_bar 0.01fF
C287 a_177_n111# x1 0.00fF
C288 CMOS_XNOR_0/XNOR a_1735_n111# 0.00fF
C289 CMOS_3in_OR_0/B a_2592_n1689# 0.00fF
C290 a_2742_n1689# CMOS_3in_AND_0/OUT 0.01fF
C291 CMOS_XOR_0/XOR a_2592_499# 0.09fF
C292 CMOS_3in_AND_0/OUT CMOS_3in_OR_0/A 0.10fF
C293 CMOS_XOR_0/XOR x0 0.00fF
C294 x2_bar x3_bar 0.14fF
C295 a_n328_n1689# VDD 1.40fF
C296 CMOS_XNOR_0/XNOR a_1380_n1689# 0.05fF
C297 a_n123_n111# x2_bar 0.01fF
C298 x1_bar x2 2.67fF
C299 x1_bar CMOS_3in_AND_0/OUT 0.01fF
C300 s1 a_2742_n1689# 0.00fF
C301 a_2742_n1689# GND 0.02fF
C302 a_2592_n1689# GND 0.02fF
C303 s1 GND 0.55fF
C304 a_1380_n779# GND 0.03fF
C305 a_n28_n779# GND 0.03fF
C306 a_n178_n779# GND 0.03fF
C307 a_2442_n779# GND 0.94fF
C308 CMOS_3in_AND_0/OUT GND 0.86fF $ **FLOATING
C309 CMOS_3in_OR_0/A GND 0.58fF
C310 a_1380_n1689# GND 0.50fF
C311 a_n328_n1689# GND 0.67fF
C312 a_2592_n111# GND 0.02fF
C313 a_1735_n111# GND 0.03fF
C314 a_1435_n111# GND 0.02fF
C315 a_177_n111# GND 0.02fF
C316 a_n123_n111# GND 0.02fF
C317 CMOS_3in_OR_0/B GND 1.97fF
C318 a_1735_499# GND 0.01fF
C319 a_1435_499# GND 0.01fF
C320 CMOS_XNOR_0/XNOR GND 1.09fF
C321 a_177_499# GND 0.01fF
C322 a_n123_499# GND 0.01fF
C323 a_2592_499# GND 0.54fF
C324 CMOS_XOR_0/XOR GND 1.15fF
C325 x1_bar GND 10.39fF
C326 x1 GND 7.19fF
C327 x3_bar GND 3.75fF
C328 a_27_n111# GND 0.63fF
C329 x0_bar GND 3.88fF
C330 x0 GND 4.16fF
C331 x2_bar GND 2.58fF
C332 x3 GND 1.76fF
C333 x2 GND 5.84fF
C334 VDD GND 24.56fF
C335 x1_bar.t0 GND 0.45fF
C336 x1_bar.t1 GND 0.40fF
C337 x1.t3 GND 0.28fF
C338 x1.t0 GND 0.11fF
C339 x1.n0 GND 0.31fF $ **FLOATING
C340 x1.n1 GND 1.58fF $ **FLOATING
C341 x1.t2 GND 0.31fF
C342 x1.t1 GND 0.26fF
C343 x1.n2 GND 0.41fF $ **FLOATING
C344 CMOS_3in_AND_0/B GND 0.43fF $ **FLOATING
C345 CMOS_3in_AND_0/OUT.t2 GND 0.10fF
C346 CMOS_3in_AND_0/OUT.t3 GND 0.11fF
C347 CMOS_3in_AND_0/OUT.t1 GND 0.31fF
C348 CMOS_3in_AND_0/OUT.t0 GND 0.28fF
C349 CMOS_3in_AND_0/OUT.n0 GND 0.69fF $ **FLOATING
C350 CMOS_3in_OR_0/C GND 0.42fF $ **FLOATING
C351 x0.t0 GND 0.14fF
C352 x0.t1 GND 0.06fF
C353 x0.n0 GND 0.16fF $ **FLOATING
C354 x3_bar.t3 GND 0.17fF
C355 x3_bar.t1 GND 0.15fF
C356 x3_bar.t2 GND 0.16fF
C357 x3_bar.t0 GND 0.19fF
C358 CMOS_3in_AND_0/A GND 0.03fF $ **FLOATING
C359 x3_bar.n0 GND 0.30fF $ **FLOATING
C360 x3_bar.n1 GND 3.62fF $ **FLOATING
C361 x3_bar.n2 GND 0.98fF $ **FLOATING
C362 x0_bar.t2 GND 0.33fF
C363 x0_bar.t0 GND 0.29fF
C364 x0_bar.t3 GND 0.14fF
C365 x0_bar.t1 GND 0.21fF
C366 x0_bar.n0 GND 0.25fF $ **FLOATING
C367 CMOS_3in_AND_0/C GND 0.43fF $ **FLOATING
C368 x0_bar.n1 GND 4.42fF $ **FLOATING
C369 x2.t1 GND 0.75fF
C370 x2.t0 GND 0.50fF
C371 x2_bar.t2 GND 0.25fF
C372 x2_bar.t1 GND 0.25fF
C373 x2_bar.n0 GND 0.67fF $ **FLOATING
C374 x2_bar.t3 GND 0.22fF
C375 x2_bar.t0 GND 0.15fF
C376 x2_bar.n1 GND 0.31fF $ **FLOATING
C377 CMOS_AND_0/B GND 0.04fF $ **FLOATING
C378 x2_bar.n2 GND 1.81fF $ **FLOATING
C379 x2_bar.n3 GND 5.69fF $ **FLOATING
C380 x3.t3 GND 0.48fF
C381 x3.t0 GND 0.33fF
C382 x3.t2 GND 0.09fF
C383 x3.t1 GND 0.13fF
C384 x3.n0 GND 0.18fF $ **FLOATING
C385 CMOS_AND_1/B GND 0.02fF $ **FLOATING
C386 x3.n1 GND 0.93fF $ **FLOATING
C387 x3.n2 GND 3.66fF $ **FLOATING
C388 VDD.t30 GND 0.07fF
C389 VDD.t14 GND 0.07fF
C390 VDD.n0 GND 0.21fF $ **FLOATING
C391 VDD.n1 GND 0.02fF $ **FLOATING
C392 VDD.n2 GND 0.02fF $ **FLOATING
C393 VDD.n3 GND 0.15fF $ **FLOATING
C394 VDD.t13 GND 0.10fF
C395 VDD.n4 GND 0.10fF $ **FLOATING
C396 VDD.n5 GND 0.02fF $ **FLOATING
C397 VDD.n6 GND 0.02fF $ **FLOATING
C398 VDD.n7 GND 0.06fF $ **FLOATING
C399 VDD.n8 GND 0.38fF $ **FLOATING
C400 VDD.n9 GND 0.17fF $ **FLOATING
C401 VDD.n10 GND 0.02fF $ **FLOATING
C402 VDD.n11 GND 0.02fF $ **FLOATING
C403 VDD.n12 GND 0.01fF $ **FLOATING
C404 VDD.n13 GND 0.17fF $ **FLOATING
C405 VDD.n14 GND 0.02fF $ **FLOATING
C406 VDD.n15 GND 0.02fF $ **FLOATING
C407 VDD.n16 GND 0.02fF $ **FLOATING
C408 VDD.n17 GND 0.17fF $ **FLOATING
C409 VDD.n18 GND 0.02fF $ **FLOATING
C410 VDD.n19 GND 0.02fF $ **FLOATING
C411 VDD.n20 GND 0.02fF $ **FLOATING
C412 VDD.n21 GND 0.17fF $ **FLOATING
C413 VDD.n22 GND 0.02fF $ **FLOATING
C414 VDD.n23 GND 0.02fF $ **FLOATING
C415 VDD.n24 GND 0.01fF $ **FLOATING
C416 VDD.n25 GND 0.37fF $ **FLOATING
C417 VDD.t27 GND 0.07fF
C418 VDD.n26 GND 0.15fF $ **FLOATING
C419 VDD.t3 GND 0.07fF
C420 CMOS_XOR_0/VDD GND 0.01fF $ **FLOATING
C421 VDD.n27 GND 0.13fF $ **FLOATING
C422 VDD.n28 GND 0.02fF $ **FLOATING
C423 VDD.t23 GND 0.07fF
C424 VDD.n29 GND 0.17fF $ **FLOATING
C425 VDD.t18 GND 0.07fF
C426 VDD.t39 GND 0.07fF
C427 VDD.t28 GND 0.09fF
C428 VDD.n30 GND 0.13fF $ **FLOATING
C429 VDD.n31 GND 0.02fF $ **FLOATING
C430 VDD.t10 GND 0.07fF
C431 VDD.t32 GND 0.05fF
C432 VDD.t12 GND 0.05fF
C433 VDD.n32 GND 0.19fF $ **FLOATING
C434 CMOS_3in_AND_0/VDD GND 0.01fF $ **FLOATING
C435 VDD.t21 GND 0.07fF
C436 VDD.t34 GND 0.07fF
C437 VDD.t25 GND 0.07fF
C438 CMOS_AND_1/VDD GND 0.01fF $ **FLOATING
C439 VDD.t6 GND 0.07fF
C440 VDD.t8 GND 0.07fF
C441 CMOS_3in_OR_0/VDD GND 0.01fF $ **FLOATING
C442 VDD.t16 GND 0.07fF
C443 VDD.n33 GND 0.20fF $ **FLOATING
C444 VDD.n34 GND 0.02fF $ **FLOATING
C445 VDD.n35 GND 0.02fF $ **FLOATING
C446 VDD.n36 GND 0.17fF $ **FLOATING
C447 VDD.t15 GND 0.10fF
C448 VDD.n37 GND 0.11fF $ **FLOATING
C449 VDD.n38 GND 0.02fF $ **FLOATING
C450 VDD.n39 GND 0.02fF $ **FLOATING
C451 VDD.n40 GND 0.05fF $ **FLOATING
C452 VDD.n41 GND 0.38fF $ **FLOATING
C453 VDD.n42 GND 0.17fF $ **FLOATING
C454 VDD.n43 GND 0.02fF $ **FLOATING
C455 VDD.n44 GND 0.02fF $ **FLOATING
C456 VDD.n45 GND 0.01fF $ **FLOATING
C457 VDD.n46 GND 0.17fF $ **FLOATING
C458 VDD.n47 GND 0.02fF $ **FLOATING
C459 VDD.n48 GND 0.02fF $ **FLOATING
C460 VDD.n49 GND 0.02fF $ **FLOATING
C461 VDD.n50 GND 0.17fF $ **FLOATING
C462 VDD.n51 GND 0.02fF $ **FLOATING
C463 VDD.n52 GND 0.02fF $ **FLOATING
C464 VDD.n53 GND 0.02fF $ **FLOATING
C465 VDD.n54 GND 0.17fF $ **FLOATING
C466 VDD.n55 GND 0.02fF $ **FLOATING
C467 VDD.n56 GND 0.02fF $ **FLOATING
C468 VDD.n57 GND 0.02fF $ **FLOATING
C469 VDD.t1 GND 0.09fF
C470 VDD.n58 GND 0.10fF $ **FLOATING
C471 VDD.n59 GND 0.02fF $ **FLOATING
C472 VDD.n60 GND 0.02fF $ **FLOATING
C473 VDD.n61 GND 0.02fF $ **FLOATING
C474 VDD.n62 GND 0.01fF $ **FLOATING
C475 VDD.n63 GND 0.16fF $ **FLOATING
C476 VDD.n64 GND 0.02fF $ **FLOATING
C477 VDD.n65 GND 0.02fF $ **FLOATING
C478 VDD.t35 GND 0.09fF
C479 VDD.n66 GND 0.11fF $ **FLOATING
C480 VDD.n67 GND 0.02fF $ **FLOATING
C481 VDD.n68 GND 0.02fF $ **FLOATING
C482 VDD.n69 GND 0.02fF $ **FLOATING
C483 VDD.n70 GND 0.15fF $ **FLOATING
C484 VDD.n71 GND 0.02fF $ **FLOATING
C485 VDD.n72 GND 0.02fF $ **FLOATING
C486 VDD.n73 GND 0.02fF $ **FLOATING
C487 VDD.t7 GND 0.10fF
C488 VDD.n74 GND 0.12fF $ **FLOATING
C489 VDD.n75 GND 0.02fF $ **FLOATING
C490 VDD.n76 GND 0.02fF $ **FLOATING
C491 VDD.n77 GND 0.02fF $ **FLOATING
C492 VDD.n78 GND 0.19fF $ **FLOATING
C493 VDD.n79 GND 0.02fF $ **FLOATING
C494 VDD.n80 GND 0.02fF $ **FLOATING
C495 VDD.n81 GND 0.01fF $ **FLOATING
C496 VDD.n82 GND 0.38fF $ **FLOATING
C497 VDD.n83 GND 0.18fF $ **FLOATING
C498 VDD.n84 GND 0.06fF $ **FLOATING
C499 VDD.n85 GND 0.16fF $ **FLOATING
C500 VDD.n86 GND 0.06fF $ **FLOATING
C501 VDD.n87 GND 0.20fF $ **FLOATING
C502 VDD.n88 GND 0.02fF $ **FLOATING
C503 VDD.n89 GND 0.02fF $ **FLOATING
C504 VDD.n90 GND 0.02fF $ **FLOATING
C505 VDD.t5 GND 0.10fF
C506 VDD.n91 GND 0.10fF $ **FLOATING
C507 VDD.n92 GND 0.02fF $ **FLOATING
C508 VDD.n93 GND 0.02fF $ **FLOATING
C509 VDD.n94 GND 0.02fF $ **FLOATING
C510 VDD.n95 GND 0.38fF $ **FLOATING
C511 VDD.n96 GND 0.17fF $ **FLOATING
C512 VDD.n97 GND 0.02fF $ **FLOATING
C513 VDD.n98 GND 0.02fF $ **FLOATING
C514 VDD.n99 GND 0.01fF $ **FLOATING
C515 VDD.n100 GND 0.17fF $ **FLOATING
C516 VDD.n101 GND 0.02fF $ **FLOATING
C517 VDD.n102 GND 0.02fF $ **FLOATING
C518 VDD.n103 GND 0.02fF $ **FLOATING
C519 VDD.n104 GND 0.17fF $ **FLOATING
C520 VDD.n105 GND 0.02fF $ **FLOATING
C521 VDD.n106 GND 0.02fF $ **FLOATING
C522 VDD.n107 GND 0.02fF $ **FLOATING
C523 VDD.t37 GND 0.07fF
C524 VDD.n108 GND 0.37fF $ **FLOATING
C525 VDD.n109 GND 0.01fF $ **FLOATING
C526 VDD.n110 GND 0.17fF $ **FLOATING
C527 VDD.n111 GND 0.02fF $ **FLOATING
C528 VDD.n112 GND 0.02fF $ **FLOATING
C529 VDD.t36 GND 0.09fF
C530 VDD.n113 GND 0.11fF $ **FLOATING
C531 VDD.n114 GND 0.02fF $ **FLOATING
C532 VDD.n115 GND 0.02fF $ **FLOATING
C533 VDD.n116 GND 0.02fF $ **FLOATING
C534 VDD.n117 GND 0.15fF $ **FLOATING
C535 VDD.n118 GND 0.02fF $ **FLOATING
C536 VDD.n119 GND 0.02fF $ **FLOATING
C537 VDD.n120 GND 0.02fF $ **FLOATING
C538 VDD.t24 GND 0.10fF
C539 VDD.n121 GND 0.12fF $ **FLOATING
C540 VDD.n122 GND 0.02fF $ **FLOATING
C541 VDD.n123 GND 0.02fF $ **FLOATING
C542 VDD.n124 GND 0.02fF $ **FLOATING
C543 VDD.n125 GND 0.19fF $ **FLOATING
C544 VDD.n126 GND 0.02fF $ **FLOATING
C545 VDD.n127 GND 0.02fF $ **FLOATING
C546 VDD.n128 GND 0.01fF $ **FLOATING
C547 VDD.n129 GND 0.38fF $ **FLOATING
C548 VDD.n130 GND 0.18fF $ **FLOATING
C549 VDD.n131 GND 0.09fF $ **FLOATING
C550 VDD.n132 GND 0.17fF $ **FLOATING
C551 VDD.n133 GND 0.09fF $ **FLOATING
C552 VDD.n134 GND 0.20fF $ **FLOATING
C553 VDD.n135 GND 0.02fF $ **FLOATING
C554 VDD.n136 GND 0.02fF $ **FLOATING
C555 VDD.n137 GND 0.02fF $ **FLOATING
C556 VDD.t33 GND 0.10fF
C557 VDD.n138 GND 0.11fF $ **FLOATING
C558 VDD.n139 GND 0.02fF $ **FLOATING
C559 VDD.n140 GND 0.02fF $ **FLOATING
C560 VDD.n141 GND 0.02fF $ **FLOATING
C561 VDD.n142 GND 0.38fF $ **FLOATING
C562 VDD.n143 GND 0.17fF $ **FLOATING
C563 VDD.n144 GND 0.02fF $ **FLOATING
C564 VDD.n145 GND 0.02fF $ **FLOATING
C565 VDD.n146 GND 0.01fF $ **FLOATING
C566 VDD.n147 GND 0.17fF $ **FLOATING
C567 VDD.n148 GND 0.02fF $ **FLOATING
C568 VDD.n149 GND 0.02fF $ **FLOATING
C569 VDD.n150 GND 0.02fF $ **FLOATING
C570 VDD.n151 GND 0.17fF $ **FLOATING
C571 VDD.n152 GND 0.02fF $ **FLOATING
C572 VDD.n153 GND 0.02fF $ **FLOATING
C573 VDD.n154 GND 0.02fF $ **FLOATING
C574 VDD.n155 GND 0.17fF $ **FLOATING
C575 VDD.n156 GND 0.02fF $ **FLOATING
C576 VDD.n157 GND 0.02fF $ **FLOATING
C577 VDD.n158 GND 0.01fF $ **FLOATING
C578 VDD.n159 GND 0.38fF $ **FLOATING
C579 VDD.t20 GND 0.09fF
C580 VDD.n160 GND 0.10fF $ **FLOATING
C581 VDD.n161 GND 0.02fF $ **FLOATING
C582 VDD.n162 GND 0.02fF $ **FLOATING
C583 VDD.n163 GND 0.02fF $ **FLOATING
C584 VDD.n164 GND 0.01fF $ **FLOATING
C585 VDD.n165 GND 0.16fF $ **FLOATING
C586 VDD.n166 GND 0.02fF $ **FLOATING
C587 VDD.n167 GND 0.02fF $ **FLOATING
C588 VDD.t31 GND 0.09fF
C589 VDD.n168 GND 0.11fF $ **FLOATING
C590 VDD.n169 GND 0.02fF $ **FLOATING
C591 VDD.n170 GND 0.02fF $ **FLOATING
C592 VDD.n171 GND 0.02fF $ **FLOATING
C593 VDD.n172 GND 0.15fF $ **FLOATING
C594 VDD.n173 GND 0.02fF $ **FLOATING
C595 VDD.n174 GND 0.02fF $ **FLOATING
C596 VDD.n175 GND 0.01fF $ **FLOATING
C597 VDD.n176 GND 0.16fF $ **FLOATING
C598 VDD.t11 GND 0.10fF
C599 VDD.n177 GND 0.12fF $ **FLOATING
C600 VDD.n178 GND 0.02fF $ **FLOATING
C601 VDD.n179 GND 0.02fF $ **FLOATING
C602 VDD.n180 GND 0.02fF $ **FLOATING
C603 VDD.n181 GND 0.19fF $ **FLOATING
C604 VDD.n182 GND 0.02fF $ **FLOATING
C605 VDD.n183 GND 0.02fF $ **FLOATING
C606 VDD.n184 GND 0.02fF $ **FLOATING
C607 VDD.n185 GND 0.18fF $ **FLOATING
C608 VDD.n186 GND 0.36fF $ **FLOATING
C609 VDD.n187 GND 0.35fF $ **FLOATING
C610 VDD.n188 GND 0.11fF $ **FLOATING
C611 VDD.n189 GND 0.02fF $ **FLOATING
C612 VDD.n190 GND 0.20fF $ **FLOATING
C613 VDD.n191 GND 0.02fF $ **FLOATING
C614 VDD.n192 GND 0.02fF $ **FLOATING
C615 VDD.n193 GND 0.01fF $ **FLOATING
C616 VDD.n194 GND 0.38fF $ **FLOATING
C617 VDD.t9 GND 0.09fF
C618 VDD.n195 GND 0.13fF $ **FLOATING
C619 VDD.n196 GND 0.02fF $ **FLOATING
C620 VDD.n197 GND 0.02fF $ **FLOATING
C621 VDD.n198 GND 0.02fF $ **FLOATING
C622 VDD.n199 GND 0.14fF $ **FLOATING
C623 VDD.n200 GND 0.02fF $ **FLOATING
C624 VDD.n201 GND 0.02fF $ **FLOATING
C625 VDD.n202 GND 0.02fF $ **FLOATING
C626 VDD.n203 GND 0.02fF $ **FLOATING
C627 VDD.n204 GND 0.13fF $ **FLOATING
C628 VDD.n205 GND 0.02fF $ **FLOATING
C629 VDD.n206 GND 0.02fF $ **FLOATING
C630 VDD.n207 GND 0.02fF $ **FLOATING
C631 VDD.n208 GND 0.01fF $ **FLOATING
C632 VDD.n209 GND 0.14fF $ **FLOATING
C633 VDD.n210 GND 0.02fF $ **FLOATING
C634 VDD.n211 GND 0.02fF $ **FLOATING
C635 VDD.n212 GND 0.02fF $ **FLOATING
C636 VDD.t19 GND 0.09fF
C637 VDD.n213 GND 0.12fF $ **FLOATING
C638 VDD.n214 GND 0.02fF $ **FLOATING
C639 VDD.n215 GND 0.02fF $ **FLOATING
C640 VDD.n216 GND 0.02fF $ **FLOATING
C641 VDD.n217 GND 0.15fF $ **FLOATING
C642 VDD.n218 GND 0.02fF $ **FLOATING
C643 VDD.n219 GND 0.02fF $ **FLOATING
C644 VDD.n220 GND 0.02fF $ **FLOATING
C645 VDD.t38 GND 0.09fF
C646 VDD.n221 GND 0.12fF $ **FLOATING
C647 VDD.n222 GND 0.02fF $ **FLOATING
C648 VDD.n223 GND 0.02fF $ **FLOATING
C649 VDD.n224 GND 0.02fF $ **FLOATING
C650 VDD.n225 GND 0.38fF $ **FLOATING
C651 VDD.n226 GND 0.17fF $ **FLOATING
C652 VDD.n227 GND 0.02fF $ **FLOATING
C653 VDD.n228 GND 0.02fF $ **FLOATING
C654 VDD.n229 GND 0.01fF $ **FLOATING
C655 VDD.n230 GND 0.17fF $ **FLOATING
C656 VDD.n231 GND 0.02fF $ **FLOATING
C657 VDD.n232 GND 0.02fF $ **FLOATING
C658 VDD.n233 GND 0.02fF $ **FLOATING
C659 VDD.n234 GND 0.17fF $ **FLOATING
C660 VDD.n235 GND 0.02fF $ **FLOATING
C661 VDD.n236 GND 0.02fF $ **FLOATING
C662 VDD.n237 GND 0.02fF $ **FLOATING
C663 VDD.n238 GND 0.17fF $ **FLOATING
C664 VDD.n239 GND 0.02fF $ **FLOATING
C665 VDD.n240 GND 0.02fF $ **FLOATING
C666 VDD.n241 GND 0.01fF $ **FLOATING
C667 VDD.n242 GND 0.38fF $ **FLOATING
C668 VDD.t17 GND 0.10fF
C669 VDD.n243 GND 0.11fF $ **FLOATING
C670 VDD.n244 GND 0.02fF $ **FLOATING
C671 VDD.n245 GND 0.02fF $ **FLOATING
C672 VDD.n246 GND 0.02fF $ **FLOATING
C673 VDD.n247 GND 0.20fF $ **FLOATING
C674 VDD.n248 GND 0.02fF $ **FLOATING
C675 VDD.n249 GND 0.02fF $ **FLOATING
C676 VDD.n250 GND 0.02fF $ **FLOATING
C677 VDD.n251 GND 0.06fF $ **FLOATING
C678 VDD.n252 GND 0.11fF $ **FLOATING
C679 VDD.n253 GND 0.06fF $ **FLOATING
C680 VDD.n254 GND 0.20fF $ **FLOATING
C681 VDD.n255 GND 0.02fF $ **FLOATING
C682 VDD.n256 GND 0.02fF $ **FLOATING
C683 VDD.n257 GND 0.01fF $ **FLOATING
C684 VDD.n258 GND 0.38fF $ **FLOATING
C685 VDD.t22 GND 0.09fF
C686 VDD.n259 GND 0.13fF $ **FLOATING
C687 VDD.n260 GND 0.02fF $ **FLOATING
C688 VDD.n261 GND 0.02fF $ **FLOATING
C689 VDD.n262 GND 0.02fF $ **FLOATING
C690 VDD.n263 GND 0.14fF $ **FLOATING
C691 VDD.n264 GND 0.02fF $ **FLOATING
C692 VDD.n265 GND 0.02fF $ **FLOATING
C693 VDD.n266 GND 0.02fF $ **FLOATING
C694 VDD.n267 GND 0.02fF $ **FLOATING
C695 VDD.n268 GND 0.02fF $ **FLOATING
C696 VDD.t0 GND 0.09fF
C697 VDD.n269 GND 0.13fF $ **FLOATING
C698 VDD.n270 GND 0.02fF $ **FLOATING
C699 VDD.n271 GND 0.02fF $ **FLOATING
C700 VDD.n272 GND 0.01fF $ **FLOATING
C701 VDD.n273 GND 0.14fF $ **FLOATING
C702 VDD.n274 GND 0.02fF $ **FLOATING
C703 VDD.n275 GND 0.02fF $ **FLOATING
C704 VDD.n276 GND 0.02fF $ **FLOATING
C705 VDD.t4 GND 0.09fF
C706 VDD.n277 GND 0.12fF $ **FLOATING
C707 VDD.n278 GND 0.02fF $ **FLOATING
C708 VDD.n279 GND 0.02fF $ **FLOATING
C709 VDD.n280 GND 0.02fF $ **FLOATING
C710 VDD.n281 GND 0.15fF $ **FLOATING
C711 VDD.n282 GND 0.02fF $ **FLOATING
C712 VDD.n283 GND 0.02fF $ **FLOATING
C713 VDD.n284 GND 0.02fF $ **FLOATING
C714 VDD.t2 GND 0.09fF
C715 VDD.n285 GND 0.13fF $ **FLOATING
C716 VDD.n286 GND 0.02fF $ **FLOATING
C717 VDD.n287 GND 0.02fF $ **FLOATING
C718 VDD.n288 GND 0.02fF $ **FLOATING
C719 VDD.n289 GND 0.38fF $ **FLOATING
C720 VDD.n290 GND 0.21fF $ **FLOATING
C721 VDD.n291 GND 0.02fF $ **FLOATING
C722 VDD.n292 GND 0.02fF $ **FLOATING
C723 VDD.n293 GND 0.01fF $ **FLOATING
C724 VDD.n294 GND 0.06fF $ **FLOATING
C725 VDD.n295 GND 0.18fF $ **FLOATING
C726 VDD.n296 GND 0.06fF $ **FLOATING
C727 VDD.n297 GND 0.38fF $ **FLOATING
C728 VDD.n298 GND 0.19fF $ **FLOATING
C729 VDD.n299 GND 0.02fF $ **FLOATING
C730 VDD.n300 GND 0.02fF $ **FLOATING
C731 VDD.n301 GND 0.01fF $ **FLOATING
C732 VDD.t26 GND 0.10fF
C733 VDD.n302 GND 0.12fF $ **FLOATING
C734 VDD.n303 GND 0.02fF $ **FLOATING
C735 VDD.n304 GND 0.02fF $ **FLOATING
C736 VDD.n305 GND 0.02fF $ **FLOATING
C737 VDD.n306 GND 0.15fF $ **FLOATING
C738 VDD.n307 GND 0.02fF $ **FLOATING
C739 VDD.n308 GND 0.02fF $ **FLOATING
C740 VDD.n309 GND 0.02fF $ **FLOATING
C741 VDD.t29 GND 0.09fF
C742 VDD.n310 GND 0.11fF $ **FLOATING
C743 VDD.n311 GND 0.02fF $ **FLOATING
C744 VDD.n312 GND 0.02fF $ **FLOATING
C745 VDD.n313 GND 0.02fF $ **FLOATING
C746 CMOS_AND_0/VDD GND 0.01fF $ **FLOATING
.ends

