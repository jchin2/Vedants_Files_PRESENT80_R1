magic
tech sky130A
timestamp 1672436480
<< end >>
