magic
tech sky130A
magscale 1 2
timestamp 1677186444
<< nwell >>
rect -389 1139 909 1369
rect 1169 1139 2121 1369
rect 2381 1139 3333 1369
rect -333 449 888 1139
rect 1225 449 2075 1139
rect 2402 449 3292 1139
rect -368 -1729 672 -1039
rect 1190 -1729 2080 -1039
rect 2402 -1729 3442 -1039
rect -389 -1959 693 -1729
rect 1169 -1959 2121 -1729
rect 2381 -1959 3463 -1729
<< pwell >>
rect -299 -219 874 215
rect 1259 -219 2031 215
rect 2416 -219 3278 215
rect -379 -371 910 -219
rect 1179 -371 2111 -219
rect 2391 -371 3464 -219
rect -354 -805 658 -371
rect 1204 -805 2066 -371
rect 2416 -805 3428 -371
<< nmos >>
rect -153 -111 -123 189
rect -3 -111 27 189
rect 147 -111 177 189
rect 297 -111 327 189
rect 698 -111 728 189
rect 1405 -111 1435 189
rect 1555 -111 1585 189
rect 1705 -111 1735 189
rect 1855 -111 1885 189
rect 2562 -111 2592 189
rect 2712 -111 2742 189
rect 3102 -111 3132 189
rect -208 -779 -178 -479
rect -58 -779 -28 -479
rect 92 -779 122 -479
rect 482 -779 512 -479
rect 1350 -779 1380 -479
rect 1500 -779 1530 -479
rect 1890 -779 1920 -479
rect 2562 -779 2592 -479
rect 2712 -779 2742 -479
rect 2862 -779 2892 -479
rect 3252 -779 3282 -479
<< pmos >>
rect -153 499 -123 1099
rect -3 499 27 1099
rect 147 499 177 1099
rect 297 499 327 1099
rect 698 499 728 1099
rect 1405 499 1435 1099
rect 1555 499 1585 1099
rect 1705 499 1735 1099
rect 1855 499 1885 1099
rect 2562 499 2592 1099
rect 2712 499 2742 1099
rect 3102 499 3132 1099
rect -208 -1689 -178 -1089
rect -58 -1689 -28 -1089
rect 92 -1689 122 -1089
rect 482 -1689 512 -1089
rect 1350 -1689 1380 -1089
rect 1500 -1689 1530 -1089
rect 1890 -1689 1920 -1089
rect 2562 -1689 2592 -1089
rect 2712 -1689 2742 -1089
rect 2862 -1689 2892 -1089
rect 3252 -1689 3282 -1089
<< ndiff >>
rect -273 158 -153 189
rect -273 124 -230 158
rect -196 124 -153 158
rect -273 90 -153 124
rect -273 56 -230 90
rect -196 56 -153 90
rect -273 22 -153 56
rect -273 -12 -230 22
rect -196 -12 -153 22
rect -273 -46 -153 -12
rect -273 -80 -230 -46
rect -196 -80 -153 -46
rect -273 -111 -153 -80
rect -123 -111 -3 189
rect 27 158 147 189
rect 27 124 70 158
rect 104 124 147 158
rect 27 90 147 124
rect 27 56 70 90
rect 104 56 147 90
rect 27 22 147 56
rect 27 -12 70 22
rect 104 -12 147 22
rect 27 -46 147 -12
rect 27 -80 70 -46
rect 104 -80 147 -46
rect 27 -111 147 -80
rect 177 -111 297 189
rect 327 158 447 189
rect 327 124 370 158
rect 404 124 447 158
rect 327 90 447 124
rect 327 56 370 90
rect 404 56 447 90
rect 327 22 447 56
rect 327 -12 370 22
rect 404 -12 447 22
rect 327 -46 447 -12
rect 327 -80 370 -46
rect 404 -80 447 -46
rect 327 -111 447 -80
rect 578 158 698 189
rect 578 124 621 158
rect 655 124 698 158
rect 578 90 698 124
rect 578 56 621 90
rect 655 56 698 90
rect 578 22 698 56
rect 578 -12 621 22
rect 655 -12 698 22
rect 578 -46 698 -12
rect 578 -80 621 -46
rect 655 -80 698 -46
rect 578 -111 698 -80
rect 728 158 848 189
rect 728 124 771 158
rect 805 124 848 158
rect 728 90 848 124
rect 728 56 771 90
rect 805 56 848 90
rect 728 22 848 56
rect 728 -12 771 22
rect 805 -12 848 22
rect 728 -46 848 -12
rect 728 -80 771 -46
rect 805 -80 848 -46
rect 728 -111 848 -80
rect 1285 158 1405 189
rect 1285 124 1328 158
rect 1362 124 1405 158
rect 1285 90 1405 124
rect 1285 56 1328 90
rect 1362 56 1405 90
rect 1285 22 1405 56
rect 1285 -12 1328 22
rect 1362 -12 1405 22
rect 1285 -46 1405 -12
rect 1285 -80 1328 -46
rect 1362 -80 1405 -46
rect 1285 -111 1405 -80
rect 1435 -111 1555 189
rect 1585 158 1705 189
rect 1585 124 1628 158
rect 1662 124 1705 158
rect 1585 90 1705 124
rect 1585 56 1628 90
rect 1662 56 1705 90
rect 1585 22 1705 56
rect 1585 -12 1628 22
rect 1662 -12 1705 22
rect 1585 -46 1705 -12
rect 1585 -80 1628 -46
rect 1662 -80 1705 -46
rect 1585 -111 1705 -80
rect 1735 -111 1855 189
rect 1885 158 2005 189
rect 1885 124 1928 158
rect 1962 124 2005 158
rect 1885 90 2005 124
rect 1885 56 1928 90
rect 1962 56 2005 90
rect 1885 22 2005 56
rect 1885 -12 1928 22
rect 1962 -12 2005 22
rect 1885 -46 2005 -12
rect 1885 -80 1928 -46
rect 1962 -80 2005 -46
rect 1885 -111 2005 -80
rect 2442 158 2562 189
rect 2442 124 2485 158
rect 2519 124 2562 158
rect 2442 90 2562 124
rect 2442 56 2485 90
rect 2519 56 2562 90
rect 2442 22 2562 56
rect 2442 -12 2485 22
rect 2519 -12 2562 22
rect 2442 -46 2562 -12
rect 2442 -80 2485 -46
rect 2519 -80 2562 -46
rect 2442 -111 2562 -80
rect 2592 -111 2712 189
rect 2742 158 2862 189
rect 2742 124 2785 158
rect 2819 124 2862 158
rect 2742 90 2862 124
rect 2742 56 2785 90
rect 2819 56 2862 90
rect 2742 22 2862 56
rect 2742 -12 2785 22
rect 2819 -12 2862 22
rect 2742 -46 2862 -12
rect 2742 -80 2785 -46
rect 2819 -80 2862 -46
rect 2742 -111 2862 -80
rect 2982 158 3102 189
rect 2982 124 3025 158
rect 3059 124 3102 158
rect 2982 90 3102 124
rect 2982 56 3025 90
rect 3059 56 3102 90
rect 2982 22 3102 56
rect 2982 -12 3025 22
rect 3059 -12 3102 22
rect 2982 -46 3102 -12
rect 2982 -80 3025 -46
rect 3059 -80 3102 -46
rect 2982 -111 3102 -80
rect 3132 158 3252 189
rect 3132 124 3175 158
rect 3209 124 3252 158
rect 3132 90 3252 124
rect 3132 56 3175 90
rect 3209 56 3252 90
rect 3132 22 3252 56
rect 3132 -12 3175 22
rect 3209 -12 3252 22
rect 3132 -46 3252 -12
rect 3132 -80 3175 -46
rect 3209 -80 3252 -46
rect 3132 -111 3252 -80
rect -328 -510 -208 -479
rect -328 -544 -285 -510
rect -251 -544 -208 -510
rect -328 -578 -208 -544
rect -328 -612 -285 -578
rect -251 -612 -208 -578
rect -328 -646 -208 -612
rect -328 -680 -285 -646
rect -251 -680 -208 -646
rect -328 -714 -208 -680
rect -328 -748 -285 -714
rect -251 -748 -208 -714
rect -328 -779 -208 -748
rect -178 -779 -58 -479
rect -28 -779 92 -479
rect 122 -510 242 -479
rect 122 -544 165 -510
rect 199 -544 242 -510
rect 122 -578 242 -544
rect 122 -612 165 -578
rect 199 -612 242 -578
rect 122 -646 242 -612
rect 122 -680 165 -646
rect 199 -680 242 -646
rect 122 -714 242 -680
rect 122 -748 165 -714
rect 199 -748 242 -714
rect 122 -779 242 -748
rect 362 -510 482 -479
rect 362 -544 405 -510
rect 439 -544 482 -510
rect 362 -578 482 -544
rect 362 -612 405 -578
rect 439 -612 482 -578
rect 362 -646 482 -612
rect 362 -680 405 -646
rect 439 -680 482 -646
rect 362 -714 482 -680
rect 362 -748 405 -714
rect 439 -748 482 -714
rect 362 -779 482 -748
rect 512 -510 632 -479
rect 512 -544 555 -510
rect 589 -544 632 -510
rect 512 -578 632 -544
rect 512 -612 555 -578
rect 589 -612 632 -578
rect 512 -646 632 -612
rect 512 -680 555 -646
rect 589 -680 632 -646
rect 512 -714 632 -680
rect 512 -748 555 -714
rect 589 -748 632 -714
rect 512 -779 632 -748
rect 1230 -510 1350 -479
rect 1230 -544 1273 -510
rect 1307 -544 1350 -510
rect 1230 -578 1350 -544
rect 1230 -612 1273 -578
rect 1307 -612 1350 -578
rect 1230 -646 1350 -612
rect 1230 -680 1273 -646
rect 1307 -680 1350 -646
rect 1230 -714 1350 -680
rect 1230 -748 1273 -714
rect 1307 -748 1350 -714
rect 1230 -779 1350 -748
rect 1380 -779 1500 -479
rect 1530 -510 1650 -479
rect 1530 -544 1573 -510
rect 1607 -544 1650 -510
rect 1530 -578 1650 -544
rect 1530 -612 1573 -578
rect 1607 -612 1650 -578
rect 1530 -646 1650 -612
rect 1530 -680 1573 -646
rect 1607 -680 1650 -646
rect 1530 -714 1650 -680
rect 1530 -748 1573 -714
rect 1607 -748 1650 -714
rect 1530 -779 1650 -748
rect 1770 -510 1890 -479
rect 1770 -544 1813 -510
rect 1847 -544 1890 -510
rect 1770 -578 1890 -544
rect 1770 -612 1813 -578
rect 1847 -612 1890 -578
rect 1770 -646 1890 -612
rect 1770 -680 1813 -646
rect 1847 -680 1890 -646
rect 1770 -714 1890 -680
rect 1770 -748 1813 -714
rect 1847 -748 1890 -714
rect 1770 -779 1890 -748
rect 1920 -510 2040 -479
rect 1920 -544 1963 -510
rect 1997 -544 2040 -510
rect 1920 -578 2040 -544
rect 1920 -612 1963 -578
rect 1997 -612 2040 -578
rect 1920 -646 2040 -612
rect 1920 -680 1963 -646
rect 1997 -680 2040 -646
rect 1920 -714 2040 -680
rect 1920 -748 1963 -714
rect 1997 -748 2040 -714
rect 1920 -779 2040 -748
rect 2442 -510 2562 -479
rect 2442 -544 2485 -510
rect 2519 -544 2562 -510
rect 2442 -578 2562 -544
rect 2442 -612 2485 -578
rect 2519 -612 2562 -578
rect 2442 -646 2562 -612
rect 2442 -680 2485 -646
rect 2519 -680 2562 -646
rect 2442 -714 2562 -680
rect 2442 -748 2485 -714
rect 2519 -748 2562 -714
rect 2442 -779 2562 -748
rect 2592 -510 2712 -479
rect 2592 -544 2635 -510
rect 2669 -544 2712 -510
rect 2592 -578 2712 -544
rect 2592 -612 2635 -578
rect 2669 -612 2712 -578
rect 2592 -646 2712 -612
rect 2592 -680 2635 -646
rect 2669 -680 2712 -646
rect 2592 -714 2712 -680
rect 2592 -748 2635 -714
rect 2669 -748 2712 -714
rect 2592 -779 2712 -748
rect 2742 -510 2862 -479
rect 2742 -544 2785 -510
rect 2819 -544 2862 -510
rect 2742 -578 2862 -544
rect 2742 -612 2785 -578
rect 2819 -612 2862 -578
rect 2742 -646 2862 -612
rect 2742 -680 2785 -646
rect 2819 -680 2862 -646
rect 2742 -714 2862 -680
rect 2742 -748 2785 -714
rect 2819 -748 2862 -714
rect 2742 -779 2862 -748
rect 2892 -510 3012 -479
rect 2892 -544 2935 -510
rect 2969 -544 3012 -510
rect 2892 -578 3012 -544
rect 2892 -612 2935 -578
rect 2969 -612 3012 -578
rect 2892 -646 3012 -612
rect 2892 -680 2935 -646
rect 2969 -680 3012 -646
rect 2892 -714 3012 -680
rect 2892 -748 2935 -714
rect 2969 -748 3012 -714
rect 2892 -779 3012 -748
rect 3132 -510 3252 -479
rect 3132 -544 3175 -510
rect 3209 -544 3252 -510
rect 3132 -578 3252 -544
rect 3132 -612 3175 -578
rect 3209 -612 3252 -578
rect 3132 -646 3252 -612
rect 3132 -680 3175 -646
rect 3209 -680 3252 -646
rect 3132 -714 3252 -680
rect 3132 -748 3175 -714
rect 3209 -748 3252 -714
rect 3132 -779 3252 -748
rect 3282 -510 3402 -479
rect 3282 -544 3325 -510
rect 3359 -544 3402 -510
rect 3282 -578 3402 -544
rect 3282 -612 3325 -578
rect 3359 -612 3402 -578
rect 3282 -646 3402 -612
rect 3282 -680 3325 -646
rect 3359 -680 3402 -646
rect 3282 -714 3402 -680
rect 3282 -748 3325 -714
rect 3359 -748 3402 -714
rect 3282 -779 3402 -748
<< pdiff >>
rect -273 1054 -153 1099
rect -273 1020 -230 1054
rect -196 1020 -153 1054
rect -273 986 -153 1020
rect -273 952 -230 986
rect -196 952 -153 986
rect -273 918 -153 952
rect -273 884 -230 918
rect -196 884 -153 918
rect -273 850 -153 884
rect -273 816 -230 850
rect -196 816 -153 850
rect -273 782 -153 816
rect -273 748 -230 782
rect -196 748 -153 782
rect -273 714 -153 748
rect -273 680 -230 714
rect -196 680 -153 714
rect -273 646 -153 680
rect -273 612 -230 646
rect -196 612 -153 646
rect -273 578 -153 612
rect -273 544 -230 578
rect -196 544 -153 578
rect -273 499 -153 544
rect -123 499 -3 1099
rect 27 1054 147 1099
rect 27 1020 70 1054
rect 104 1020 147 1054
rect 27 986 147 1020
rect 27 952 70 986
rect 104 952 147 986
rect 27 918 147 952
rect 27 884 70 918
rect 104 884 147 918
rect 27 850 147 884
rect 27 816 70 850
rect 104 816 147 850
rect 27 782 147 816
rect 27 748 70 782
rect 104 748 147 782
rect 27 714 147 748
rect 27 680 70 714
rect 104 680 147 714
rect 27 646 147 680
rect 27 612 70 646
rect 104 612 147 646
rect 27 578 147 612
rect 27 544 70 578
rect 104 544 147 578
rect 27 499 147 544
rect 177 499 297 1099
rect 327 1054 447 1099
rect 327 1020 370 1054
rect 404 1020 447 1054
rect 327 986 447 1020
rect 327 952 370 986
rect 404 952 447 986
rect 327 918 447 952
rect 327 884 370 918
rect 404 884 447 918
rect 327 850 447 884
rect 327 816 370 850
rect 404 816 447 850
rect 327 782 447 816
rect 327 748 370 782
rect 404 748 447 782
rect 327 714 447 748
rect 327 680 370 714
rect 404 680 447 714
rect 327 646 447 680
rect 327 612 370 646
rect 404 612 447 646
rect 327 578 447 612
rect 327 544 370 578
rect 404 544 447 578
rect 327 499 447 544
rect 578 1054 698 1099
rect 578 1020 621 1054
rect 655 1020 698 1054
rect 578 986 698 1020
rect 578 952 621 986
rect 655 952 698 986
rect 578 918 698 952
rect 578 884 621 918
rect 655 884 698 918
rect 578 850 698 884
rect 578 816 621 850
rect 655 816 698 850
rect 578 782 698 816
rect 578 748 621 782
rect 655 748 698 782
rect 578 714 698 748
rect 578 680 621 714
rect 655 680 698 714
rect 578 646 698 680
rect 578 612 621 646
rect 655 612 698 646
rect 578 578 698 612
rect 578 544 621 578
rect 655 544 698 578
rect 578 499 698 544
rect 728 1054 848 1099
rect 728 1020 771 1054
rect 805 1020 848 1054
rect 728 986 848 1020
rect 728 952 771 986
rect 805 952 848 986
rect 728 918 848 952
rect 728 884 771 918
rect 805 884 848 918
rect 728 850 848 884
rect 728 816 771 850
rect 805 816 848 850
rect 728 782 848 816
rect 728 748 771 782
rect 805 748 848 782
rect 728 714 848 748
rect 728 680 771 714
rect 805 680 848 714
rect 728 646 848 680
rect 728 612 771 646
rect 805 612 848 646
rect 728 578 848 612
rect 728 544 771 578
rect 805 544 848 578
rect 728 499 848 544
rect 1285 1054 1405 1099
rect 1285 1020 1328 1054
rect 1362 1020 1405 1054
rect 1285 986 1405 1020
rect 1285 952 1328 986
rect 1362 952 1405 986
rect 1285 918 1405 952
rect 1285 884 1328 918
rect 1362 884 1405 918
rect 1285 850 1405 884
rect 1285 816 1328 850
rect 1362 816 1405 850
rect 1285 782 1405 816
rect 1285 748 1328 782
rect 1362 748 1405 782
rect 1285 714 1405 748
rect 1285 680 1328 714
rect 1362 680 1405 714
rect 1285 646 1405 680
rect 1285 612 1328 646
rect 1362 612 1405 646
rect 1285 578 1405 612
rect 1285 544 1328 578
rect 1362 544 1405 578
rect 1285 499 1405 544
rect 1435 499 1555 1099
rect 1585 1054 1705 1099
rect 1585 1020 1628 1054
rect 1662 1020 1705 1054
rect 1585 986 1705 1020
rect 1585 952 1628 986
rect 1662 952 1705 986
rect 1585 918 1705 952
rect 1585 884 1628 918
rect 1662 884 1705 918
rect 1585 850 1705 884
rect 1585 816 1628 850
rect 1662 816 1705 850
rect 1585 782 1705 816
rect 1585 748 1628 782
rect 1662 748 1705 782
rect 1585 714 1705 748
rect 1585 680 1628 714
rect 1662 680 1705 714
rect 1585 646 1705 680
rect 1585 612 1628 646
rect 1662 612 1705 646
rect 1585 578 1705 612
rect 1585 544 1628 578
rect 1662 544 1705 578
rect 1585 499 1705 544
rect 1735 499 1855 1099
rect 1885 1054 2005 1099
rect 1885 1020 1928 1054
rect 1962 1020 2005 1054
rect 1885 986 2005 1020
rect 1885 952 1928 986
rect 1962 952 2005 986
rect 1885 918 2005 952
rect 1885 884 1928 918
rect 1962 884 2005 918
rect 1885 850 2005 884
rect 1885 816 1928 850
rect 1962 816 2005 850
rect 1885 782 2005 816
rect 1885 748 1928 782
rect 1962 748 2005 782
rect 1885 714 2005 748
rect 1885 680 1928 714
rect 1962 680 2005 714
rect 1885 646 2005 680
rect 1885 612 1928 646
rect 1962 612 2005 646
rect 1885 578 2005 612
rect 1885 544 1928 578
rect 1962 544 2005 578
rect 1885 499 2005 544
rect 2442 1054 2562 1099
rect 2442 1020 2485 1054
rect 2519 1020 2562 1054
rect 2442 986 2562 1020
rect 2442 952 2485 986
rect 2519 952 2562 986
rect 2442 918 2562 952
rect 2442 884 2485 918
rect 2519 884 2562 918
rect 2442 850 2562 884
rect 2442 816 2485 850
rect 2519 816 2562 850
rect 2442 782 2562 816
rect 2442 748 2485 782
rect 2519 748 2562 782
rect 2442 714 2562 748
rect 2442 680 2485 714
rect 2519 680 2562 714
rect 2442 646 2562 680
rect 2442 612 2485 646
rect 2519 612 2562 646
rect 2442 578 2562 612
rect 2442 544 2485 578
rect 2519 544 2562 578
rect 2442 499 2562 544
rect 2592 1054 2712 1099
rect 2592 1020 2635 1054
rect 2669 1020 2712 1054
rect 2592 986 2712 1020
rect 2592 952 2635 986
rect 2669 952 2712 986
rect 2592 918 2712 952
rect 2592 884 2635 918
rect 2669 884 2712 918
rect 2592 850 2712 884
rect 2592 816 2635 850
rect 2669 816 2712 850
rect 2592 782 2712 816
rect 2592 748 2635 782
rect 2669 748 2712 782
rect 2592 714 2712 748
rect 2592 680 2635 714
rect 2669 680 2712 714
rect 2592 646 2712 680
rect 2592 612 2635 646
rect 2669 612 2712 646
rect 2592 578 2712 612
rect 2592 544 2635 578
rect 2669 544 2712 578
rect 2592 499 2712 544
rect 2742 1054 2862 1099
rect 2742 1020 2785 1054
rect 2819 1020 2862 1054
rect 2742 986 2862 1020
rect 2742 952 2785 986
rect 2819 952 2862 986
rect 2742 918 2862 952
rect 2742 884 2785 918
rect 2819 884 2862 918
rect 2742 850 2862 884
rect 2742 816 2785 850
rect 2819 816 2862 850
rect 2742 782 2862 816
rect 2742 748 2785 782
rect 2819 748 2862 782
rect 2742 714 2862 748
rect 2742 680 2785 714
rect 2819 680 2862 714
rect 2742 646 2862 680
rect 2742 612 2785 646
rect 2819 612 2862 646
rect 2742 578 2862 612
rect 2742 544 2785 578
rect 2819 544 2862 578
rect 2742 499 2862 544
rect 2982 1054 3102 1099
rect 2982 1020 3025 1054
rect 3059 1020 3102 1054
rect 2982 986 3102 1020
rect 2982 952 3025 986
rect 3059 952 3102 986
rect 2982 918 3102 952
rect 2982 884 3025 918
rect 3059 884 3102 918
rect 2982 850 3102 884
rect 2982 816 3025 850
rect 3059 816 3102 850
rect 2982 782 3102 816
rect 2982 748 3025 782
rect 3059 748 3102 782
rect 2982 714 3102 748
rect 2982 680 3025 714
rect 3059 680 3102 714
rect 2982 646 3102 680
rect 2982 612 3025 646
rect 3059 612 3102 646
rect 2982 578 3102 612
rect 2982 544 3025 578
rect 3059 544 3102 578
rect 2982 499 3102 544
rect 3132 1054 3252 1099
rect 3132 1020 3175 1054
rect 3209 1020 3252 1054
rect 3132 986 3252 1020
rect 3132 952 3175 986
rect 3209 952 3252 986
rect 3132 918 3252 952
rect 3132 884 3175 918
rect 3209 884 3252 918
rect 3132 850 3252 884
rect 3132 816 3175 850
rect 3209 816 3252 850
rect 3132 782 3252 816
rect 3132 748 3175 782
rect 3209 748 3252 782
rect 3132 714 3252 748
rect 3132 680 3175 714
rect 3209 680 3252 714
rect 3132 646 3252 680
rect 3132 612 3175 646
rect 3209 612 3252 646
rect 3132 578 3252 612
rect 3132 544 3175 578
rect 3209 544 3252 578
rect 3132 499 3252 544
rect -328 -1134 -208 -1089
rect -328 -1168 -285 -1134
rect -251 -1168 -208 -1134
rect -328 -1202 -208 -1168
rect -328 -1236 -285 -1202
rect -251 -1236 -208 -1202
rect -328 -1270 -208 -1236
rect -328 -1304 -285 -1270
rect -251 -1304 -208 -1270
rect -328 -1338 -208 -1304
rect -328 -1372 -285 -1338
rect -251 -1372 -208 -1338
rect -328 -1406 -208 -1372
rect -328 -1440 -285 -1406
rect -251 -1440 -208 -1406
rect -328 -1474 -208 -1440
rect -328 -1508 -285 -1474
rect -251 -1508 -208 -1474
rect -328 -1542 -208 -1508
rect -328 -1576 -285 -1542
rect -251 -1576 -208 -1542
rect -328 -1610 -208 -1576
rect -328 -1644 -285 -1610
rect -251 -1644 -208 -1610
rect -328 -1689 -208 -1644
rect -178 -1134 -58 -1089
rect -178 -1168 -135 -1134
rect -101 -1168 -58 -1134
rect -178 -1202 -58 -1168
rect -178 -1236 -135 -1202
rect -101 -1236 -58 -1202
rect -178 -1270 -58 -1236
rect -178 -1304 -135 -1270
rect -101 -1304 -58 -1270
rect -178 -1338 -58 -1304
rect -178 -1372 -135 -1338
rect -101 -1372 -58 -1338
rect -178 -1406 -58 -1372
rect -178 -1440 -135 -1406
rect -101 -1440 -58 -1406
rect -178 -1474 -58 -1440
rect -178 -1508 -135 -1474
rect -101 -1508 -58 -1474
rect -178 -1542 -58 -1508
rect -178 -1576 -135 -1542
rect -101 -1576 -58 -1542
rect -178 -1610 -58 -1576
rect -178 -1644 -135 -1610
rect -101 -1644 -58 -1610
rect -178 -1689 -58 -1644
rect -28 -1134 92 -1089
rect -28 -1168 15 -1134
rect 49 -1168 92 -1134
rect -28 -1202 92 -1168
rect -28 -1236 15 -1202
rect 49 -1236 92 -1202
rect -28 -1270 92 -1236
rect -28 -1304 15 -1270
rect 49 -1304 92 -1270
rect -28 -1338 92 -1304
rect -28 -1372 15 -1338
rect 49 -1372 92 -1338
rect -28 -1406 92 -1372
rect -28 -1440 15 -1406
rect 49 -1440 92 -1406
rect -28 -1474 92 -1440
rect -28 -1508 15 -1474
rect 49 -1508 92 -1474
rect -28 -1542 92 -1508
rect -28 -1576 15 -1542
rect 49 -1576 92 -1542
rect -28 -1610 92 -1576
rect -28 -1644 15 -1610
rect 49 -1644 92 -1610
rect -28 -1689 92 -1644
rect 122 -1134 242 -1089
rect 122 -1168 165 -1134
rect 199 -1168 242 -1134
rect 122 -1202 242 -1168
rect 122 -1236 165 -1202
rect 199 -1236 242 -1202
rect 122 -1270 242 -1236
rect 122 -1304 165 -1270
rect 199 -1304 242 -1270
rect 122 -1338 242 -1304
rect 122 -1372 165 -1338
rect 199 -1372 242 -1338
rect 122 -1406 242 -1372
rect 122 -1440 165 -1406
rect 199 -1440 242 -1406
rect 122 -1474 242 -1440
rect 122 -1508 165 -1474
rect 199 -1508 242 -1474
rect 122 -1542 242 -1508
rect 122 -1576 165 -1542
rect 199 -1576 242 -1542
rect 122 -1610 242 -1576
rect 122 -1644 165 -1610
rect 199 -1644 242 -1610
rect 122 -1689 242 -1644
rect 362 -1134 482 -1089
rect 362 -1168 405 -1134
rect 439 -1168 482 -1134
rect 362 -1202 482 -1168
rect 362 -1236 405 -1202
rect 439 -1236 482 -1202
rect 362 -1270 482 -1236
rect 362 -1304 405 -1270
rect 439 -1304 482 -1270
rect 362 -1338 482 -1304
rect 362 -1372 405 -1338
rect 439 -1372 482 -1338
rect 362 -1406 482 -1372
rect 362 -1440 405 -1406
rect 439 -1440 482 -1406
rect 362 -1474 482 -1440
rect 362 -1508 405 -1474
rect 439 -1508 482 -1474
rect 362 -1542 482 -1508
rect 362 -1576 405 -1542
rect 439 -1576 482 -1542
rect 362 -1610 482 -1576
rect 362 -1644 405 -1610
rect 439 -1644 482 -1610
rect 362 -1689 482 -1644
rect 512 -1134 632 -1089
rect 512 -1168 555 -1134
rect 589 -1168 632 -1134
rect 512 -1202 632 -1168
rect 512 -1236 555 -1202
rect 589 -1236 632 -1202
rect 512 -1270 632 -1236
rect 512 -1304 555 -1270
rect 589 -1304 632 -1270
rect 512 -1338 632 -1304
rect 512 -1372 555 -1338
rect 589 -1372 632 -1338
rect 512 -1406 632 -1372
rect 512 -1440 555 -1406
rect 589 -1440 632 -1406
rect 512 -1474 632 -1440
rect 512 -1508 555 -1474
rect 589 -1508 632 -1474
rect 512 -1542 632 -1508
rect 512 -1576 555 -1542
rect 589 -1576 632 -1542
rect 512 -1610 632 -1576
rect 512 -1644 555 -1610
rect 589 -1644 632 -1610
rect 512 -1689 632 -1644
rect 1230 -1134 1350 -1089
rect 1230 -1168 1273 -1134
rect 1307 -1168 1350 -1134
rect 1230 -1202 1350 -1168
rect 1230 -1236 1273 -1202
rect 1307 -1236 1350 -1202
rect 1230 -1270 1350 -1236
rect 1230 -1304 1273 -1270
rect 1307 -1304 1350 -1270
rect 1230 -1338 1350 -1304
rect 1230 -1372 1273 -1338
rect 1307 -1372 1350 -1338
rect 1230 -1406 1350 -1372
rect 1230 -1440 1273 -1406
rect 1307 -1440 1350 -1406
rect 1230 -1474 1350 -1440
rect 1230 -1508 1273 -1474
rect 1307 -1508 1350 -1474
rect 1230 -1542 1350 -1508
rect 1230 -1576 1273 -1542
rect 1307 -1576 1350 -1542
rect 1230 -1610 1350 -1576
rect 1230 -1644 1273 -1610
rect 1307 -1644 1350 -1610
rect 1230 -1689 1350 -1644
rect 1380 -1134 1500 -1089
rect 1380 -1168 1423 -1134
rect 1457 -1168 1500 -1134
rect 1380 -1202 1500 -1168
rect 1380 -1236 1423 -1202
rect 1457 -1236 1500 -1202
rect 1380 -1270 1500 -1236
rect 1380 -1304 1423 -1270
rect 1457 -1304 1500 -1270
rect 1380 -1338 1500 -1304
rect 1380 -1372 1423 -1338
rect 1457 -1372 1500 -1338
rect 1380 -1406 1500 -1372
rect 1380 -1440 1423 -1406
rect 1457 -1440 1500 -1406
rect 1380 -1474 1500 -1440
rect 1380 -1508 1423 -1474
rect 1457 -1508 1500 -1474
rect 1380 -1542 1500 -1508
rect 1380 -1576 1423 -1542
rect 1457 -1576 1500 -1542
rect 1380 -1610 1500 -1576
rect 1380 -1644 1423 -1610
rect 1457 -1644 1500 -1610
rect 1380 -1689 1500 -1644
rect 1530 -1134 1650 -1089
rect 1530 -1168 1573 -1134
rect 1607 -1168 1650 -1134
rect 1530 -1202 1650 -1168
rect 1530 -1236 1573 -1202
rect 1607 -1236 1650 -1202
rect 1530 -1270 1650 -1236
rect 1530 -1304 1573 -1270
rect 1607 -1304 1650 -1270
rect 1530 -1338 1650 -1304
rect 1530 -1372 1573 -1338
rect 1607 -1372 1650 -1338
rect 1530 -1406 1650 -1372
rect 1530 -1440 1573 -1406
rect 1607 -1440 1650 -1406
rect 1530 -1474 1650 -1440
rect 1530 -1508 1573 -1474
rect 1607 -1508 1650 -1474
rect 1530 -1542 1650 -1508
rect 1530 -1576 1573 -1542
rect 1607 -1576 1650 -1542
rect 1530 -1610 1650 -1576
rect 1530 -1644 1573 -1610
rect 1607 -1644 1650 -1610
rect 1530 -1689 1650 -1644
rect 1770 -1134 1890 -1089
rect 1770 -1168 1813 -1134
rect 1847 -1168 1890 -1134
rect 1770 -1202 1890 -1168
rect 1770 -1236 1813 -1202
rect 1847 -1236 1890 -1202
rect 1770 -1270 1890 -1236
rect 1770 -1304 1813 -1270
rect 1847 -1304 1890 -1270
rect 1770 -1338 1890 -1304
rect 1770 -1372 1813 -1338
rect 1847 -1372 1890 -1338
rect 1770 -1406 1890 -1372
rect 1770 -1440 1813 -1406
rect 1847 -1440 1890 -1406
rect 1770 -1474 1890 -1440
rect 1770 -1508 1813 -1474
rect 1847 -1508 1890 -1474
rect 1770 -1542 1890 -1508
rect 1770 -1576 1813 -1542
rect 1847 -1576 1890 -1542
rect 1770 -1610 1890 -1576
rect 1770 -1644 1813 -1610
rect 1847 -1644 1890 -1610
rect 1770 -1689 1890 -1644
rect 1920 -1134 2040 -1089
rect 1920 -1168 1963 -1134
rect 1997 -1168 2040 -1134
rect 1920 -1202 2040 -1168
rect 1920 -1236 1963 -1202
rect 1997 -1236 2040 -1202
rect 1920 -1270 2040 -1236
rect 1920 -1304 1963 -1270
rect 1997 -1304 2040 -1270
rect 1920 -1338 2040 -1304
rect 1920 -1372 1963 -1338
rect 1997 -1372 2040 -1338
rect 1920 -1406 2040 -1372
rect 1920 -1440 1963 -1406
rect 1997 -1440 2040 -1406
rect 1920 -1474 2040 -1440
rect 1920 -1508 1963 -1474
rect 1997 -1508 2040 -1474
rect 1920 -1542 2040 -1508
rect 1920 -1576 1963 -1542
rect 1997 -1576 2040 -1542
rect 1920 -1610 2040 -1576
rect 1920 -1644 1963 -1610
rect 1997 -1644 2040 -1610
rect 1920 -1689 2040 -1644
rect 2442 -1134 2562 -1089
rect 2442 -1168 2485 -1134
rect 2519 -1168 2562 -1134
rect 2442 -1202 2562 -1168
rect 2442 -1236 2485 -1202
rect 2519 -1236 2562 -1202
rect 2442 -1270 2562 -1236
rect 2442 -1304 2485 -1270
rect 2519 -1304 2562 -1270
rect 2442 -1338 2562 -1304
rect 2442 -1372 2485 -1338
rect 2519 -1372 2562 -1338
rect 2442 -1406 2562 -1372
rect 2442 -1440 2485 -1406
rect 2519 -1440 2562 -1406
rect 2442 -1474 2562 -1440
rect 2442 -1508 2485 -1474
rect 2519 -1508 2562 -1474
rect 2442 -1542 2562 -1508
rect 2442 -1576 2485 -1542
rect 2519 -1576 2562 -1542
rect 2442 -1610 2562 -1576
rect 2442 -1644 2485 -1610
rect 2519 -1644 2562 -1610
rect 2442 -1689 2562 -1644
rect 2592 -1689 2712 -1089
rect 2742 -1689 2862 -1089
rect 2892 -1134 3012 -1089
rect 2892 -1168 2935 -1134
rect 2969 -1168 3012 -1134
rect 2892 -1202 3012 -1168
rect 2892 -1236 2935 -1202
rect 2969 -1236 3012 -1202
rect 2892 -1270 3012 -1236
rect 2892 -1304 2935 -1270
rect 2969 -1304 3012 -1270
rect 2892 -1338 3012 -1304
rect 2892 -1372 2935 -1338
rect 2969 -1372 3012 -1338
rect 2892 -1406 3012 -1372
rect 2892 -1440 2935 -1406
rect 2969 -1440 3012 -1406
rect 2892 -1474 3012 -1440
rect 2892 -1508 2935 -1474
rect 2969 -1508 3012 -1474
rect 2892 -1542 3012 -1508
rect 2892 -1576 2935 -1542
rect 2969 -1576 3012 -1542
rect 2892 -1610 3012 -1576
rect 2892 -1644 2935 -1610
rect 2969 -1644 3012 -1610
rect 2892 -1689 3012 -1644
rect 3132 -1134 3252 -1089
rect 3132 -1168 3175 -1134
rect 3209 -1168 3252 -1134
rect 3132 -1202 3252 -1168
rect 3132 -1236 3175 -1202
rect 3209 -1236 3252 -1202
rect 3132 -1270 3252 -1236
rect 3132 -1304 3175 -1270
rect 3209 -1304 3252 -1270
rect 3132 -1338 3252 -1304
rect 3132 -1372 3175 -1338
rect 3209 -1372 3252 -1338
rect 3132 -1406 3252 -1372
rect 3132 -1440 3175 -1406
rect 3209 -1440 3252 -1406
rect 3132 -1474 3252 -1440
rect 3132 -1508 3175 -1474
rect 3209 -1508 3252 -1474
rect 3132 -1542 3252 -1508
rect 3132 -1576 3175 -1542
rect 3209 -1576 3252 -1542
rect 3132 -1610 3252 -1576
rect 3132 -1644 3175 -1610
rect 3209 -1644 3252 -1610
rect 3132 -1689 3252 -1644
rect 3282 -1134 3402 -1089
rect 3282 -1168 3325 -1134
rect 3359 -1168 3402 -1134
rect 3282 -1202 3402 -1168
rect 3282 -1236 3325 -1202
rect 3359 -1236 3402 -1202
rect 3282 -1270 3402 -1236
rect 3282 -1304 3325 -1270
rect 3359 -1304 3402 -1270
rect 3282 -1338 3402 -1304
rect 3282 -1372 3325 -1338
rect 3359 -1372 3402 -1338
rect 3282 -1406 3402 -1372
rect 3282 -1440 3325 -1406
rect 3359 -1440 3402 -1406
rect 3282 -1474 3402 -1440
rect 3282 -1508 3325 -1474
rect 3359 -1508 3402 -1474
rect 3282 -1542 3402 -1508
rect 3282 -1576 3325 -1542
rect 3359 -1576 3402 -1542
rect 3282 -1610 3402 -1576
rect 3282 -1644 3325 -1610
rect 3359 -1644 3402 -1610
rect 3282 -1689 3402 -1644
<< ndiffc >>
rect -230 124 -196 158
rect -230 56 -196 90
rect -230 -12 -196 22
rect -230 -80 -196 -46
rect 70 124 104 158
rect 70 56 104 90
rect 70 -12 104 22
rect 70 -80 104 -46
rect 370 124 404 158
rect 370 56 404 90
rect 370 -12 404 22
rect 370 -80 404 -46
rect 621 124 655 158
rect 621 56 655 90
rect 621 -12 655 22
rect 621 -80 655 -46
rect 771 124 805 158
rect 771 56 805 90
rect 771 -12 805 22
rect 771 -80 805 -46
rect 1328 124 1362 158
rect 1328 56 1362 90
rect 1328 -12 1362 22
rect 1328 -80 1362 -46
rect 1628 124 1662 158
rect 1628 56 1662 90
rect 1628 -12 1662 22
rect 1628 -80 1662 -46
rect 1928 124 1962 158
rect 1928 56 1962 90
rect 1928 -12 1962 22
rect 1928 -80 1962 -46
rect 2485 124 2519 158
rect 2485 56 2519 90
rect 2485 -12 2519 22
rect 2485 -80 2519 -46
rect 2785 124 2819 158
rect 2785 56 2819 90
rect 2785 -12 2819 22
rect 2785 -80 2819 -46
rect 3025 124 3059 158
rect 3025 56 3059 90
rect 3025 -12 3059 22
rect 3025 -80 3059 -46
rect 3175 124 3209 158
rect 3175 56 3209 90
rect 3175 -12 3209 22
rect 3175 -80 3209 -46
rect -285 -544 -251 -510
rect -285 -612 -251 -578
rect -285 -680 -251 -646
rect -285 -748 -251 -714
rect 165 -544 199 -510
rect 165 -612 199 -578
rect 165 -680 199 -646
rect 165 -748 199 -714
rect 405 -544 439 -510
rect 405 -612 439 -578
rect 405 -680 439 -646
rect 405 -748 439 -714
rect 555 -544 589 -510
rect 555 -612 589 -578
rect 555 -680 589 -646
rect 555 -748 589 -714
rect 1273 -544 1307 -510
rect 1273 -612 1307 -578
rect 1273 -680 1307 -646
rect 1273 -748 1307 -714
rect 1573 -544 1607 -510
rect 1573 -612 1607 -578
rect 1573 -680 1607 -646
rect 1573 -748 1607 -714
rect 1813 -544 1847 -510
rect 1813 -612 1847 -578
rect 1813 -680 1847 -646
rect 1813 -748 1847 -714
rect 1963 -544 1997 -510
rect 1963 -612 1997 -578
rect 1963 -680 1997 -646
rect 1963 -748 1997 -714
rect 2485 -544 2519 -510
rect 2485 -612 2519 -578
rect 2485 -680 2519 -646
rect 2485 -748 2519 -714
rect 2635 -544 2669 -510
rect 2635 -612 2669 -578
rect 2635 -680 2669 -646
rect 2635 -748 2669 -714
rect 2785 -544 2819 -510
rect 2785 -612 2819 -578
rect 2785 -680 2819 -646
rect 2785 -748 2819 -714
rect 2935 -544 2969 -510
rect 2935 -612 2969 -578
rect 2935 -680 2969 -646
rect 2935 -748 2969 -714
rect 3175 -544 3209 -510
rect 3175 -612 3209 -578
rect 3175 -680 3209 -646
rect 3175 -748 3209 -714
rect 3325 -544 3359 -510
rect 3325 -612 3359 -578
rect 3325 -680 3359 -646
rect 3325 -748 3359 -714
<< pdiffc >>
rect -230 1020 -196 1054
rect -230 952 -196 986
rect -230 884 -196 918
rect -230 816 -196 850
rect -230 748 -196 782
rect -230 680 -196 714
rect -230 612 -196 646
rect -230 544 -196 578
rect 70 1020 104 1054
rect 70 952 104 986
rect 70 884 104 918
rect 70 816 104 850
rect 70 748 104 782
rect 70 680 104 714
rect 70 612 104 646
rect 70 544 104 578
rect 370 1020 404 1054
rect 370 952 404 986
rect 370 884 404 918
rect 370 816 404 850
rect 370 748 404 782
rect 370 680 404 714
rect 370 612 404 646
rect 370 544 404 578
rect 621 1020 655 1054
rect 621 952 655 986
rect 621 884 655 918
rect 621 816 655 850
rect 621 748 655 782
rect 621 680 655 714
rect 621 612 655 646
rect 621 544 655 578
rect 771 1020 805 1054
rect 771 952 805 986
rect 771 884 805 918
rect 771 816 805 850
rect 771 748 805 782
rect 771 680 805 714
rect 771 612 805 646
rect 771 544 805 578
rect 1328 1020 1362 1054
rect 1328 952 1362 986
rect 1328 884 1362 918
rect 1328 816 1362 850
rect 1328 748 1362 782
rect 1328 680 1362 714
rect 1328 612 1362 646
rect 1328 544 1362 578
rect 1628 1020 1662 1054
rect 1628 952 1662 986
rect 1628 884 1662 918
rect 1628 816 1662 850
rect 1628 748 1662 782
rect 1628 680 1662 714
rect 1628 612 1662 646
rect 1628 544 1662 578
rect 1928 1020 1962 1054
rect 1928 952 1962 986
rect 1928 884 1962 918
rect 1928 816 1962 850
rect 1928 748 1962 782
rect 1928 680 1962 714
rect 1928 612 1962 646
rect 1928 544 1962 578
rect 2485 1020 2519 1054
rect 2485 952 2519 986
rect 2485 884 2519 918
rect 2485 816 2519 850
rect 2485 748 2519 782
rect 2485 680 2519 714
rect 2485 612 2519 646
rect 2485 544 2519 578
rect 2635 1020 2669 1054
rect 2635 952 2669 986
rect 2635 884 2669 918
rect 2635 816 2669 850
rect 2635 748 2669 782
rect 2635 680 2669 714
rect 2635 612 2669 646
rect 2635 544 2669 578
rect 2785 1020 2819 1054
rect 2785 952 2819 986
rect 2785 884 2819 918
rect 2785 816 2819 850
rect 2785 748 2819 782
rect 2785 680 2819 714
rect 2785 612 2819 646
rect 2785 544 2819 578
rect 3025 1020 3059 1054
rect 3025 952 3059 986
rect 3025 884 3059 918
rect 3025 816 3059 850
rect 3025 748 3059 782
rect 3025 680 3059 714
rect 3025 612 3059 646
rect 3025 544 3059 578
rect 3175 1020 3209 1054
rect 3175 952 3209 986
rect 3175 884 3209 918
rect 3175 816 3209 850
rect 3175 748 3209 782
rect 3175 680 3209 714
rect 3175 612 3209 646
rect 3175 544 3209 578
rect -285 -1168 -251 -1134
rect -285 -1236 -251 -1202
rect -285 -1304 -251 -1270
rect -285 -1372 -251 -1338
rect -285 -1440 -251 -1406
rect -285 -1508 -251 -1474
rect -285 -1576 -251 -1542
rect -285 -1644 -251 -1610
rect -135 -1168 -101 -1134
rect -135 -1236 -101 -1202
rect -135 -1304 -101 -1270
rect -135 -1372 -101 -1338
rect -135 -1440 -101 -1406
rect -135 -1508 -101 -1474
rect -135 -1576 -101 -1542
rect -135 -1644 -101 -1610
rect 15 -1168 49 -1134
rect 15 -1236 49 -1202
rect 15 -1304 49 -1270
rect 15 -1372 49 -1338
rect 15 -1440 49 -1406
rect 15 -1508 49 -1474
rect 15 -1576 49 -1542
rect 15 -1644 49 -1610
rect 165 -1168 199 -1134
rect 165 -1236 199 -1202
rect 165 -1304 199 -1270
rect 165 -1372 199 -1338
rect 165 -1440 199 -1406
rect 165 -1508 199 -1474
rect 165 -1576 199 -1542
rect 165 -1644 199 -1610
rect 405 -1168 439 -1134
rect 405 -1236 439 -1202
rect 405 -1304 439 -1270
rect 405 -1372 439 -1338
rect 405 -1440 439 -1406
rect 405 -1508 439 -1474
rect 405 -1576 439 -1542
rect 405 -1644 439 -1610
rect 555 -1168 589 -1134
rect 555 -1236 589 -1202
rect 555 -1304 589 -1270
rect 555 -1372 589 -1338
rect 555 -1440 589 -1406
rect 555 -1508 589 -1474
rect 555 -1576 589 -1542
rect 555 -1644 589 -1610
rect 1273 -1168 1307 -1134
rect 1273 -1236 1307 -1202
rect 1273 -1304 1307 -1270
rect 1273 -1372 1307 -1338
rect 1273 -1440 1307 -1406
rect 1273 -1508 1307 -1474
rect 1273 -1576 1307 -1542
rect 1273 -1644 1307 -1610
rect 1423 -1168 1457 -1134
rect 1423 -1236 1457 -1202
rect 1423 -1304 1457 -1270
rect 1423 -1372 1457 -1338
rect 1423 -1440 1457 -1406
rect 1423 -1508 1457 -1474
rect 1423 -1576 1457 -1542
rect 1423 -1644 1457 -1610
rect 1573 -1168 1607 -1134
rect 1573 -1236 1607 -1202
rect 1573 -1304 1607 -1270
rect 1573 -1372 1607 -1338
rect 1573 -1440 1607 -1406
rect 1573 -1508 1607 -1474
rect 1573 -1576 1607 -1542
rect 1573 -1644 1607 -1610
rect 1813 -1168 1847 -1134
rect 1813 -1236 1847 -1202
rect 1813 -1304 1847 -1270
rect 1813 -1372 1847 -1338
rect 1813 -1440 1847 -1406
rect 1813 -1508 1847 -1474
rect 1813 -1576 1847 -1542
rect 1813 -1644 1847 -1610
rect 1963 -1168 1997 -1134
rect 1963 -1236 1997 -1202
rect 1963 -1304 1997 -1270
rect 1963 -1372 1997 -1338
rect 1963 -1440 1997 -1406
rect 1963 -1508 1997 -1474
rect 1963 -1576 1997 -1542
rect 1963 -1644 1997 -1610
rect 2485 -1168 2519 -1134
rect 2485 -1236 2519 -1202
rect 2485 -1304 2519 -1270
rect 2485 -1372 2519 -1338
rect 2485 -1440 2519 -1406
rect 2485 -1508 2519 -1474
rect 2485 -1576 2519 -1542
rect 2485 -1644 2519 -1610
rect 2935 -1168 2969 -1134
rect 2935 -1236 2969 -1202
rect 2935 -1304 2969 -1270
rect 2935 -1372 2969 -1338
rect 2935 -1440 2969 -1406
rect 2935 -1508 2969 -1474
rect 2935 -1576 2969 -1542
rect 2935 -1644 2969 -1610
rect 3175 -1168 3209 -1134
rect 3175 -1236 3209 -1202
rect 3175 -1304 3209 -1270
rect 3175 -1372 3209 -1338
rect 3175 -1440 3209 -1406
rect 3175 -1508 3209 -1474
rect 3175 -1576 3209 -1542
rect 3175 -1644 3209 -1610
rect 3325 -1168 3359 -1134
rect 3325 -1236 3359 -1202
rect 3325 -1304 3359 -1270
rect 3325 -1372 3359 -1338
rect 3325 -1440 3359 -1406
rect 3325 -1508 3359 -1474
rect 3325 -1576 3359 -1542
rect 3325 -1644 3359 -1610
<< psubdiff >>
rect -353 -278 884 -245
rect -353 -312 -330 -278
rect -296 -312 -258 -278
rect -224 -312 -186 -278
rect -152 -312 -114 -278
rect -80 -312 -42 -278
rect -8 -312 30 -278
rect 64 -312 102 -278
rect 136 -312 174 -278
rect 208 -312 246 -278
rect 280 -312 318 -278
rect 352 -312 390 -278
rect 424 -312 462 -278
rect 496 -312 534 -278
rect 568 -312 606 -278
rect 640 -312 678 -278
rect 712 -312 750 -278
rect 784 -312 822 -278
rect 856 -312 884 -278
rect -353 -345 884 -312
rect 1205 -278 2085 -245
rect 1205 -312 1228 -278
rect 1262 -312 1300 -278
rect 1334 -312 1372 -278
rect 1406 -312 1444 -278
rect 1478 -312 1516 -278
rect 1550 -312 1588 -278
rect 1622 -312 1660 -278
rect 1694 -312 1732 -278
rect 1766 -312 1804 -278
rect 1838 -312 1876 -278
rect 1910 -312 1948 -278
rect 1982 -312 2020 -278
rect 2054 -312 2085 -278
rect 1205 -345 2085 -312
rect 2417 -278 3438 -245
rect 2417 -312 2440 -278
rect 2474 -312 2512 -278
rect 2546 -312 2584 -278
rect 2618 -312 2656 -278
rect 2690 -312 2728 -278
rect 2762 -312 2800 -278
rect 2834 -312 2872 -278
rect 2906 -312 2944 -278
rect 2978 -312 3016 -278
rect 3050 -312 3088 -278
rect 3122 -312 3160 -278
rect 3194 -312 3232 -278
rect 3266 -312 3304 -278
rect 3338 -312 3376 -278
rect 3410 -312 3438 -278
rect 2417 -345 3438 -312
<< nsubdiff >>
rect -353 1300 873 1333
rect -353 1266 -330 1300
rect -296 1266 -258 1300
rect -224 1266 -186 1300
rect -152 1266 -114 1300
rect -80 1266 -42 1300
rect -8 1266 30 1300
rect 64 1266 102 1300
rect 136 1266 174 1300
rect 208 1266 246 1300
rect 280 1266 318 1300
rect 352 1266 390 1300
rect 424 1266 462 1300
rect 496 1266 534 1300
rect 568 1266 606 1300
rect 640 1266 678 1300
rect 712 1266 750 1300
rect 784 1266 822 1300
rect 856 1266 873 1300
rect -353 1233 873 1266
rect 1205 1300 2085 1333
rect 1205 1266 1228 1300
rect 1262 1266 1300 1300
rect 1334 1266 1372 1300
rect 1406 1266 1444 1300
rect 1478 1266 1516 1300
rect 1550 1266 1588 1300
rect 1622 1266 1660 1300
rect 1694 1266 1732 1300
rect 1766 1266 1804 1300
rect 1838 1266 1876 1300
rect 1910 1266 1948 1300
rect 1982 1266 2020 1300
rect 2054 1266 2085 1300
rect 1205 1233 2085 1266
rect 2417 1300 3297 1333
rect 2417 1266 2440 1300
rect 2474 1266 2512 1300
rect 2546 1266 2584 1300
rect 2618 1266 2656 1300
rect 2690 1266 2728 1300
rect 2762 1266 2800 1300
rect 2834 1266 2872 1300
rect 2906 1266 2944 1300
rect 2978 1266 3016 1300
rect 3050 1266 3088 1300
rect 3122 1266 3160 1300
rect 3194 1266 3232 1300
rect 3266 1266 3297 1300
rect 2417 1233 3297 1266
rect -353 -1856 657 -1823
rect -353 -1890 -330 -1856
rect -296 -1890 -258 -1856
rect -224 -1890 -186 -1856
rect -152 -1890 -114 -1856
rect -80 -1890 -42 -1856
rect -8 -1890 30 -1856
rect 64 -1890 102 -1856
rect 136 -1890 174 -1856
rect 208 -1890 246 -1856
rect 280 -1890 318 -1856
rect 352 -1890 390 -1856
rect 424 -1890 462 -1856
rect 496 -1890 534 -1856
rect 568 -1890 606 -1856
rect 640 -1890 657 -1856
rect -353 -1923 657 -1890
rect 1205 -1856 2085 -1823
rect 1205 -1890 1228 -1856
rect 1262 -1890 1300 -1856
rect 1334 -1890 1372 -1856
rect 1406 -1890 1444 -1856
rect 1478 -1890 1516 -1856
rect 1550 -1890 1588 -1856
rect 1622 -1890 1660 -1856
rect 1694 -1890 1732 -1856
rect 1766 -1890 1804 -1856
rect 1838 -1890 1876 -1856
rect 1910 -1890 1948 -1856
rect 1982 -1890 2020 -1856
rect 2054 -1890 2085 -1856
rect 1205 -1923 2085 -1890
rect 2417 -1856 3427 -1823
rect 2417 -1890 2440 -1856
rect 2474 -1890 2512 -1856
rect 2546 -1890 2584 -1856
rect 2618 -1890 2656 -1856
rect 2690 -1890 2728 -1856
rect 2762 -1890 2800 -1856
rect 2834 -1890 2872 -1856
rect 2906 -1890 2944 -1856
rect 2978 -1890 3016 -1856
rect 3050 -1890 3088 -1856
rect 3122 -1890 3160 -1856
rect 3194 -1890 3232 -1856
rect 3266 -1890 3304 -1856
rect 3338 -1890 3376 -1856
rect 3410 -1890 3427 -1856
rect 2417 -1923 3427 -1890
<< psubdiffcont >>
rect -330 -312 -296 -278
rect -258 -312 -224 -278
rect -186 -312 -152 -278
rect -114 -312 -80 -278
rect -42 -312 -8 -278
rect 30 -312 64 -278
rect 102 -312 136 -278
rect 174 -312 208 -278
rect 246 -312 280 -278
rect 318 -312 352 -278
rect 390 -312 424 -278
rect 462 -312 496 -278
rect 534 -312 568 -278
rect 606 -312 640 -278
rect 678 -312 712 -278
rect 750 -312 784 -278
rect 822 -312 856 -278
rect 1228 -312 1262 -278
rect 1300 -312 1334 -278
rect 1372 -312 1406 -278
rect 1444 -312 1478 -278
rect 1516 -312 1550 -278
rect 1588 -312 1622 -278
rect 1660 -312 1694 -278
rect 1732 -312 1766 -278
rect 1804 -312 1838 -278
rect 1876 -312 1910 -278
rect 1948 -312 1982 -278
rect 2020 -312 2054 -278
rect 2440 -312 2474 -278
rect 2512 -312 2546 -278
rect 2584 -312 2618 -278
rect 2656 -312 2690 -278
rect 2728 -312 2762 -278
rect 2800 -312 2834 -278
rect 2872 -312 2906 -278
rect 2944 -312 2978 -278
rect 3016 -312 3050 -278
rect 3088 -312 3122 -278
rect 3160 -312 3194 -278
rect 3232 -312 3266 -278
rect 3304 -312 3338 -278
rect 3376 -312 3410 -278
<< nsubdiffcont >>
rect -330 1266 -296 1300
rect -258 1266 -224 1300
rect -186 1266 -152 1300
rect -114 1266 -80 1300
rect -42 1266 -8 1300
rect 30 1266 64 1300
rect 102 1266 136 1300
rect 174 1266 208 1300
rect 246 1266 280 1300
rect 318 1266 352 1300
rect 390 1266 424 1300
rect 462 1266 496 1300
rect 534 1266 568 1300
rect 606 1266 640 1300
rect 678 1266 712 1300
rect 750 1266 784 1300
rect 822 1266 856 1300
rect 1228 1266 1262 1300
rect 1300 1266 1334 1300
rect 1372 1266 1406 1300
rect 1444 1266 1478 1300
rect 1516 1266 1550 1300
rect 1588 1266 1622 1300
rect 1660 1266 1694 1300
rect 1732 1266 1766 1300
rect 1804 1266 1838 1300
rect 1876 1266 1910 1300
rect 1948 1266 1982 1300
rect 2020 1266 2054 1300
rect 2440 1266 2474 1300
rect 2512 1266 2546 1300
rect 2584 1266 2618 1300
rect 2656 1266 2690 1300
rect 2728 1266 2762 1300
rect 2800 1266 2834 1300
rect 2872 1266 2906 1300
rect 2944 1266 2978 1300
rect 3016 1266 3050 1300
rect 3088 1266 3122 1300
rect 3160 1266 3194 1300
rect 3232 1266 3266 1300
rect -330 -1890 -296 -1856
rect -258 -1890 -224 -1856
rect -186 -1890 -152 -1856
rect -114 -1890 -80 -1856
rect -42 -1890 -8 -1856
rect 30 -1890 64 -1856
rect 102 -1890 136 -1856
rect 174 -1890 208 -1856
rect 246 -1890 280 -1856
rect 318 -1890 352 -1856
rect 390 -1890 424 -1856
rect 462 -1890 496 -1856
rect 534 -1890 568 -1856
rect 606 -1890 640 -1856
rect 1228 -1890 1262 -1856
rect 1300 -1890 1334 -1856
rect 1372 -1890 1406 -1856
rect 1444 -1890 1478 -1856
rect 1516 -1890 1550 -1856
rect 1588 -1890 1622 -1856
rect 1660 -1890 1694 -1856
rect 1732 -1890 1766 -1856
rect 1804 -1890 1838 -1856
rect 1876 -1890 1910 -1856
rect 1948 -1890 1982 -1856
rect 2020 -1890 2054 -1856
rect 2440 -1890 2474 -1856
rect 2512 -1890 2546 -1856
rect 2584 -1890 2618 -1856
rect 2656 -1890 2690 -1856
rect 2728 -1890 2762 -1856
rect 2800 -1890 2834 -1856
rect 2872 -1890 2906 -1856
rect 2944 -1890 2978 -1856
rect 3016 -1890 3050 -1856
rect 3088 -1890 3122 -1856
rect 3160 -1890 3194 -1856
rect 3232 -1890 3266 -1856
rect 3304 -1890 3338 -1856
rect 3376 -1890 3410 -1856
<< poly >>
rect 247 1186 327 1209
rect 247 1152 270 1186
rect 304 1152 327 1186
rect 247 1129 327 1152
rect 1805 1186 1885 1209
rect 1805 1152 1828 1186
rect 1862 1152 1885 1186
rect 1805 1129 1885 1152
rect -153 1099 -123 1129
rect -3 1099 27 1129
rect 147 1099 177 1129
rect 297 1099 327 1129
rect 698 1099 728 1129
rect 1405 1099 1435 1129
rect 1555 1099 1585 1129
rect 1705 1099 1735 1129
rect 1855 1099 1885 1129
rect 2562 1099 2592 1129
rect 2712 1099 2742 1129
rect 3102 1099 3132 1129
rect -153 475 -123 499
rect -233 452 -123 475
rect -233 418 -210 452
rect -176 418 -123 452
rect -233 398 -123 418
rect -233 395 -153 398
rect -3 356 27 499
rect -125 326 27 356
rect 147 356 177 499
rect 297 475 327 499
rect 297 452 407 475
rect 698 469 728 499
rect 1405 475 1435 499
rect 297 418 350 452
rect 384 418 407 452
rect 297 398 407 418
rect 327 395 407 398
rect 618 446 728 469
rect 618 412 641 446
rect 675 412 728 446
rect 618 389 728 412
rect 1325 452 1435 475
rect 1325 418 1348 452
rect 1382 418 1435 452
rect 1325 398 1435 418
rect 1325 395 1405 398
rect 147 326 299 356
rect -125 284 -95 326
rect -203 261 -95 284
rect -203 227 -180 261
rect -146 227 -95 261
rect -203 219 -95 227
rect -53 261 27 284
rect -53 227 -30 261
rect 4 227 27 261
rect -203 204 -123 219
rect -53 204 27 227
rect -153 189 -123 204
rect -3 189 27 204
rect 147 261 227 284
rect 147 227 170 261
rect 204 227 227 261
rect 147 204 227 227
rect 269 241 299 326
rect 269 211 327 241
rect 147 189 177 204
rect 297 189 327 211
rect 698 189 728 389
rect 1555 356 1585 499
rect 1433 326 1585 356
rect 1705 356 1735 499
rect 1855 475 1885 499
rect 1855 452 1965 475
rect 2562 469 2592 499
rect 1855 418 1908 452
rect 1942 418 1965 452
rect 1855 398 1965 418
rect 1885 395 1965 398
rect 2482 446 2592 469
rect 2482 412 2505 446
rect 2539 412 2592 446
rect 2482 389 2592 412
rect 1705 326 1857 356
rect 1433 284 1463 326
rect 1355 261 1463 284
rect 1355 227 1378 261
rect 1412 227 1463 261
rect 1355 219 1463 227
rect 1505 261 1585 284
rect 1505 227 1528 261
rect 1562 227 1585 261
rect 1355 204 1435 219
rect 1505 204 1585 227
rect 1405 189 1435 204
rect 1555 189 1585 204
rect 1705 261 1785 284
rect 1705 227 1728 261
rect 1762 227 1785 261
rect 1705 204 1785 227
rect 1827 241 1857 326
rect 1827 211 1885 241
rect 1705 189 1735 204
rect 1855 189 1885 211
rect 2562 189 2592 389
rect 2712 189 2742 499
rect 3102 469 3132 499
rect 3022 446 3132 469
rect 3022 412 3045 446
rect 3079 412 3132 446
rect 3022 389 3132 412
rect 3102 189 3132 389
rect -153 -141 -123 -111
rect -3 -141 27 -111
rect 147 -141 177 -111
rect 297 -141 327 -111
rect 698 -141 728 -111
rect 1405 -141 1435 -111
rect 1555 -141 1585 -111
rect 1705 -141 1735 -111
rect 1855 -141 1885 -111
rect 2562 -141 2592 -111
rect 2712 -141 2742 -111
rect 3102 -141 3132 -111
rect 247 -164 327 -141
rect 247 -198 270 -164
rect 304 -198 327 -164
rect 247 -221 327 -198
rect 1805 -164 1885 -141
rect 1805 -198 1828 -164
rect 1862 -198 1885 -164
rect 1805 -221 1885 -198
rect 2662 -164 2742 -141
rect 2662 -198 2685 -164
rect 2719 -198 2742 -164
rect 2662 -221 2742 -198
rect -108 -392 -28 -369
rect -108 -426 -85 -392
rect -51 -426 -28 -392
rect -108 -449 -28 -426
rect 1450 -392 1530 -369
rect 1450 -426 1473 -392
rect 1507 -426 1530 -392
rect 1450 -449 1530 -426
rect 2662 -392 2742 -369
rect 2662 -426 2685 -392
rect 2719 -426 2742 -392
rect 2662 -449 2742 -426
rect -208 -479 -178 -449
rect -58 -479 -28 -449
rect 92 -479 122 -449
rect 482 -479 512 -449
rect 1350 -479 1380 -449
rect 1500 -479 1530 -449
rect 1890 -479 1920 -449
rect 2562 -479 2592 -449
rect 2712 -479 2742 -449
rect 2862 -479 2892 -449
rect 3252 -479 3282 -449
rect -208 -969 -178 -779
rect -258 -992 -178 -969
rect -258 -1026 -235 -992
rect -201 -1026 -178 -992
rect -258 -1049 -178 -1026
rect -208 -1089 -178 -1049
rect -58 -1089 -28 -779
rect 92 -1089 122 -779
rect 482 -979 512 -779
rect 1350 -979 1380 -779
rect 402 -1002 512 -979
rect 402 -1036 425 -1002
rect 459 -1036 512 -1002
rect 402 -1059 512 -1036
rect 1270 -1002 1380 -979
rect 1270 -1036 1293 -1002
rect 1327 -1036 1380 -1002
rect 1270 -1059 1380 -1036
rect 482 -1089 512 -1059
rect 1350 -1089 1380 -1059
rect 1500 -1089 1530 -779
rect 1890 -979 1920 -779
rect 2562 -969 2592 -779
rect 1810 -1002 1920 -979
rect 1810 -1036 1833 -1002
rect 1867 -1036 1920 -1002
rect 1810 -1059 1920 -1036
rect 2512 -992 2592 -969
rect 2512 -1026 2535 -992
rect 2569 -1026 2592 -992
rect 2512 -1049 2592 -1026
rect 1890 -1089 1920 -1059
rect 2562 -1089 2592 -1049
rect 2712 -1089 2742 -779
rect 2862 -1089 2892 -779
rect 3252 -979 3282 -779
rect 3172 -1002 3282 -979
rect 3172 -1036 3195 -1002
rect 3229 -1036 3282 -1002
rect 3172 -1059 3282 -1036
rect 3252 -1089 3282 -1059
rect -208 -1719 -178 -1689
rect -58 -1719 -28 -1689
rect 92 -1719 122 -1689
rect 482 -1719 512 -1689
rect 1350 -1719 1380 -1689
rect 1500 -1719 1530 -1689
rect 1890 -1719 1920 -1689
rect 2562 -1719 2592 -1689
rect 2712 -1719 2742 -1689
rect 2862 -1719 2892 -1689
rect 3252 -1719 3282 -1689
rect 92 -1742 172 -1719
rect 92 -1776 115 -1742
rect 149 -1776 172 -1742
rect 92 -1799 172 -1776
rect 2832 -1742 2912 -1719
rect 2832 -1776 2855 -1742
rect 2889 -1776 2912 -1742
rect 2832 -1799 2912 -1776
<< polycont >>
rect 270 1152 304 1186
rect 1828 1152 1862 1186
rect -210 418 -176 452
rect 350 418 384 452
rect 641 412 675 446
rect 1348 418 1382 452
rect -180 227 -146 261
rect -30 227 4 261
rect 170 227 204 261
rect 1908 418 1942 452
rect 2505 412 2539 446
rect 1378 227 1412 261
rect 1528 227 1562 261
rect 1728 227 1762 261
rect 3045 412 3079 446
rect 270 -198 304 -164
rect 1828 -198 1862 -164
rect 2685 -198 2719 -164
rect -85 -426 -51 -392
rect 1473 -426 1507 -392
rect 2685 -426 2719 -392
rect -235 -1026 -201 -992
rect 425 -1036 459 -1002
rect 1293 -1036 1327 -1002
rect 1833 -1036 1867 -1002
rect 2535 -1026 2569 -992
rect 3195 -1036 3229 -1002
rect 115 -1776 149 -1742
rect 2855 -1776 2889 -1742
<< locali >>
rect -353 1300 873 1323
rect -1031 1258 -951 1281
rect -1031 1224 -1008 1258
rect -974 1224 -951 1258
rect -353 1266 -330 1300
rect -296 1266 -258 1300
rect -224 1266 -186 1300
rect -152 1266 -114 1300
rect -80 1266 -42 1300
rect -8 1266 30 1300
rect 64 1266 102 1300
rect 136 1266 174 1300
rect 208 1266 246 1300
rect 280 1266 318 1300
rect 352 1266 390 1300
rect 424 1266 462 1300
rect 496 1266 534 1300
rect 568 1266 606 1300
rect 640 1266 678 1300
rect 712 1266 750 1300
rect 784 1266 822 1300
rect 856 1266 873 1300
rect -353 1243 873 1266
rect 1205 1300 2085 1323
rect 1205 1266 1228 1300
rect 1262 1266 1300 1300
rect 1334 1266 1372 1300
rect 1406 1266 1444 1300
rect 1478 1266 1516 1300
rect 1550 1266 1588 1300
rect 1622 1266 1660 1300
rect 1694 1266 1732 1300
rect 1766 1266 1804 1300
rect 1838 1266 1876 1300
rect 1910 1266 1948 1300
rect 1982 1266 2020 1300
rect 2054 1266 2085 1300
rect 1205 1243 2085 1266
rect 2417 1300 3297 1323
rect 2417 1266 2440 1300
rect 2474 1266 2512 1300
rect 2546 1266 2584 1300
rect 2618 1266 2656 1300
rect 2690 1266 2728 1300
rect 2762 1266 2800 1300
rect 2834 1266 2872 1300
rect 2906 1266 2944 1300
rect 2978 1266 3016 1300
rect 3050 1266 3088 1300
rect 3122 1266 3160 1300
rect 3194 1266 3232 1300
rect 3266 1266 3297 1300
rect 2417 1243 3297 1266
rect -1031 1189 -951 1224
rect 247 1189 327 1209
rect -1031 1186 327 1189
rect -1031 1152 -1008 1186
rect -974 1152 270 1186
rect 304 1152 327 1186
rect -1031 1149 327 1152
rect -1031 1114 -951 1149
rect 247 1129 327 1149
rect 1660 1189 1740 1205
rect 1805 1189 1885 1209
rect 1660 1186 1885 1189
rect 1660 1182 1828 1186
rect 1660 1148 1683 1182
rect 1717 1152 1828 1182
rect 1862 1152 1885 1186
rect 1717 1149 1885 1152
rect 1717 1148 1740 1149
rect 1660 1125 1740 1148
rect 1805 1129 1885 1149
rect -1031 1080 -1008 1114
rect -974 1080 -951 1114
rect -1031 1057 -951 1080
rect -253 1068 -173 1079
rect -253 1020 -230 1068
rect -196 1020 -173 1068
rect -253 996 -173 1020
rect -253 952 -230 996
rect -196 952 -173 996
rect -253 924 -173 952
rect -253 884 -230 924
rect -196 884 -173 924
rect -253 852 -173 884
rect -253 816 -230 852
rect -196 816 -173 852
rect -253 782 -173 816
rect -253 746 -230 782
rect -196 746 -173 782
rect -253 714 -173 746
rect -253 674 -230 714
rect -196 674 -173 714
rect -253 646 -173 674
rect -253 602 -230 646
rect -196 602 -173 646
rect -253 578 -173 602
rect -917 524 -837 547
rect -917 490 -894 524
rect -860 490 -837 524
rect -253 530 -230 578
rect -196 530 -173 578
rect -253 519 -173 530
rect 47 1068 127 1079
rect 47 1020 70 1068
rect 104 1020 127 1068
rect 47 996 127 1020
rect 47 952 70 996
rect 104 952 127 996
rect 47 924 127 952
rect 47 884 70 924
rect 104 884 127 924
rect 47 852 127 884
rect 47 816 70 852
rect 104 816 127 852
rect 47 782 127 816
rect 47 746 70 782
rect 104 746 127 782
rect 47 714 127 746
rect 47 674 70 714
rect 104 674 127 714
rect 47 646 127 674
rect 47 602 70 646
rect 104 602 127 646
rect 47 578 127 602
rect 47 530 70 578
rect 104 530 127 578
rect 47 519 127 530
rect 347 1068 427 1079
rect 347 1020 370 1068
rect 404 1020 427 1068
rect 347 996 427 1020
rect 347 952 370 996
rect 404 952 427 996
rect 347 924 427 952
rect 347 884 370 924
rect 404 884 427 924
rect 347 852 427 884
rect 347 816 370 852
rect 404 816 427 852
rect 347 782 427 816
rect 347 746 370 782
rect 404 746 427 782
rect 347 714 427 746
rect 347 674 370 714
rect 404 674 427 714
rect 347 646 427 674
rect 347 602 370 646
rect 404 602 427 646
rect 347 578 427 602
rect 347 530 370 578
rect 404 530 427 578
rect 347 519 427 530
rect 598 1068 678 1079
rect 598 1020 621 1068
rect 655 1020 678 1068
rect 598 996 678 1020
rect 598 952 621 996
rect 655 952 678 996
rect 598 924 678 952
rect 598 884 621 924
rect 655 884 678 924
rect 598 852 678 884
rect 598 816 621 852
rect 655 816 678 852
rect 598 782 678 816
rect 598 746 621 782
rect 655 746 678 782
rect 598 714 678 746
rect 598 674 621 714
rect 655 674 678 714
rect 598 646 678 674
rect 598 602 621 646
rect 655 602 678 646
rect 598 578 678 602
rect 598 530 621 578
rect 655 530 678 578
rect 598 519 678 530
rect 748 1054 828 1079
rect 748 1020 771 1054
rect 805 1020 828 1054
rect 748 986 828 1020
rect 748 952 771 986
rect 805 952 828 986
rect 748 918 828 952
rect 748 884 771 918
rect 805 884 828 918
rect 748 850 828 884
rect 748 816 771 850
rect 805 816 828 850
rect 748 782 828 816
rect 748 748 771 782
rect 805 748 828 782
rect 748 714 828 748
rect 748 680 771 714
rect 805 680 828 714
rect 748 646 828 680
rect 748 612 771 646
rect 805 612 828 646
rect 748 578 828 612
rect 748 544 771 578
rect 805 544 828 578
rect 748 519 828 544
rect 1305 1068 1385 1079
rect 1305 1020 1328 1068
rect 1362 1020 1385 1068
rect 1305 996 1385 1020
rect 1305 952 1328 996
rect 1362 952 1385 996
rect 1305 924 1385 952
rect 1305 884 1328 924
rect 1362 884 1385 924
rect 1305 852 1385 884
rect 1305 816 1328 852
rect 1362 816 1385 852
rect 1305 782 1385 816
rect 1305 746 1328 782
rect 1362 746 1385 782
rect 1305 714 1385 746
rect 1305 674 1328 714
rect 1362 674 1385 714
rect 1305 646 1385 674
rect 1305 602 1328 646
rect 1362 602 1385 646
rect 1305 578 1385 602
rect 1305 530 1328 578
rect 1362 530 1385 578
rect 1305 519 1385 530
rect 1605 1068 1685 1079
rect 1605 1020 1628 1068
rect 1662 1020 1685 1068
rect 1605 996 1685 1020
rect 1605 952 1628 996
rect 1662 952 1685 996
rect 1605 924 1685 952
rect 1605 884 1628 924
rect 1662 884 1685 924
rect 1605 852 1685 884
rect 1605 816 1628 852
rect 1662 816 1685 852
rect 1605 782 1685 816
rect 1605 746 1628 782
rect 1662 746 1685 782
rect 1605 714 1685 746
rect 1605 674 1628 714
rect 1662 674 1685 714
rect 1605 646 1685 674
rect 1605 602 1628 646
rect 1662 602 1685 646
rect 1605 578 1685 602
rect 1605 530 1628 578
rect 1662 530 1685 578
rect 1605 519 1685 530
rect 1905 1068 1985 1079
rect 1905 1020 1928 1068
rect 1962 1020 1985 1068
rect 1905 996 1985 1020
rect 1905 952 1928 996
rect 1962 952 1985 996
rect 1905 924 1985 952
rect 1905 884 1928 924
rect 1962 884 1985 924
rect 1905 852 1985 884
rect 1905 816 1928 852
rect 1962 816 1985 852
rect 1905 782 1985 816
rect 1905 746 1928 782
rect 1962 746 1985 782
rect 1905 714 1985 746
rect 1905 674 1928 714
rect 1962 674 1985 714
rect 1905 646 1985 674
rect 1905 602 1928 646
rect 1962 602 1985 646
rect 1905 578 1985 602
rect 1905 530 1928 578
rect 1962 530 1985 578
rect 1905 519 1985 530
rect 2462 1068 2542 1079
rect 2462 1020 2485 1068
rect 2519 1020 2542 1068
rect 2462 996 2542 1020
rect 2462 952 2485 996
rect 2519 952 2542 996
rect 2462 924 2542 952
rect 2462 884 2485 924
rect 2519 884 2542 924
rect 2462 852 2542 884
rect 2462 816 2485 852
rect 2519 816 2542 852
rect 2462 782 2542 816
rect 2462 746 2485 782
rect 2519 746 2542 782
rect 2462 714 2542 746
rect 2462 674 2485 714
rect 2519 674 2542 714
rect 2462 646 2542 674
rect 2462 602 2485 646
rect 2519 602 2542 646
rect 2462 578 2542 602
rect 2462 530 2485 578
rect 2519 530 2542 578
rect 2462 519 2542 530
rect 2612 1054 2692 1079
rect 2612 1020 2635 1054
rect 2669 1020 2692 1054
rect 2612 986 2692 1020
rect 2612 952 2635 986
rect 2669 952 2692 986
rect 2612 918 2692 952
rect 2612 884 2635 918
rect 2669 884 2692 918
rect 2612 850 2692 884
rect 2612 816 2635 850
rect 2669 816 2692 850
rect 2612 782 2692 816
rect 2612 748 2635 782
rect 2669 748 2692 782
rect 2612 714 2692 748
rect 2612 680 2635 714
rect 2669 680 2692 714
rect 2612 646 2692 680
rect 2612 612 2635 646
rect 2669 612 2692 646
rect 2612 578 2692 612
rect 2612 544 2635 578
rect 2669 544 2692 578
rect 2612 519 2692 544
rect 2762 1068 2842 1079
rect 2762 1020 2785 1068
rect 2819 1020 2842 1068
rect 2762 996 2842 1020
rect 2762 952 2785 996
rect 2819 952 2842 996
rect 2762 924 2842 952
rect 2762 884 2785 924
rect 2819 884 2842 924
rect 2762 852 2842 884
rect 2762 816 2785 852
rect 2819 816 2842 852
rect 2762 782 2842 816
rect 2762 746 2785 782
rect 2819 746 2842 782
rect 2762 714 2842 746
rect 2762 674 2785 714
rect 2819 674 2842 714
rect 2762 646 2842 674
rect 2762 602 2785 646
rect 2819 602 2842 646
rect 2762 578 2842 602
rect 2762 530 2785 578
rect 2819 530 2842 578
rect 2762 519 2842 530
rect 3002 1068 3082 1079
rect 3002 1020 3025 1068
rect 3059 1020 3082 1068
rect 3002 996 3082 1020
rect 3002 952 3025 996
rect 3059 952 3082 996
rect 3002 924 3082 952
rect 3002 884 3025 924
rect 3059 884 3082 924
rect 3002 852 3082 884
rect 3002 816 3025 852
rect 3059 816 3082 852
rect 3002 782 3082 816
rect 3002 746 3025 782
rect 3059 746 3082 782
rect 3002 714 3082 746
rect 3002 674 3025 714
rect 3059 674 3082 714
rect 3002 646 3082 674
rect 3002 602 3025 646
rect 3059 602 3082 646
rect 3002 578 3082 602
rect 3002 530 3025 578
rect 3059 530 3082 578
rect 3002 519 3082 530
rect 3152 1054 3232 1079
rect 3152 1020 3175 1054
rect 3209 1020 3232 1054
rect 3152 986 3232 1020
rect 3152 952 3175 986
rect 3209 952 3232 986
rect 3152 918 3232 952
rect 3152 884 3175 918
rect 3209 884 3232 918
rect 3152 850 3232 884
rect 3152 816 3175 850
rect 3209 816 3232 850
rect 3152 782 3232 816
rect 3152 748 3175 782
rect 3209 748 3232 782
rect 3152 714 3232 748
rect 3152 680 3175 714
rect 3209 680 3232 714
rect 3152 646 3232 680
rect 3152 612 3175 646
rect 3209 612 3232 646
rect 3152 578 3232 612
rect 3152 544 3175 578
rect 3209 544 3232 578
rect 3152 519 3232 544
rect -917 455 -837 490
rect -233 455 -153 475
rect -917 452 207 455
rect -917 418 -894 452
rect -860 418 -210 452
rect -176 418 207 452
rect -917 415 207 418
rect -917 380 -837 415
rect -233 395 -153 415
rect -1487 333 -1407 356
rect -1487 299 -1464 333
rect -1430 299 -1407 333
rect -917 346 -894 380
rect -860 346 -837 380
rect -917 323 -837 346
rect -1487 264 -1407 299
rect 167 284 207 415
rect 327 452 407 475
rect 327 418 350 452
rect 384 418 407 452
rect 618 449 698 469
rect 327 395 407 418
rect 496 446 698 449
rect 496 412 641 446
rect 675 412 698 446
rect 496 409 698 412
rect 496 363 536 409
rect 618 389 698 409
rect 476 340 556 363
rect 476 306 499 340
rect 533 306 556 340
rect -203 264 -123 284
rect -1487 261 -123 264
rect -1487 227 -1464 261
rect -1430 227 -180 261
rect -146 227 -123 261
rect -1487 224 -123 227
rect -1487 189 -1407 224
rect -203 204 -123 224
rect -53 261 27 284
rect -53 227 -30 261
rect 4 227 27 261
rect -53 204 27 227
rect 147 261 227 284
rect 476 283 556 306
rect 147 227 170 261
rect 204 227 227 261
rect 147 204 227 227
rect -1487 155 -1464 189
rect -1430 155 -1407 189
rect 768 169 808 519
rect 1325 455 1405 475
rect 1325 452 1765 455
rect 1325 418 1348 452
rect 1382 418 1765 452
rect 1325 415 1765 418
rect 1325 395 1405 415
rect 1725 284 1765 415
rect 1885 452 1965 475
rect 1885 418 1908 452
rect 1942 418 1965 452
rect 1885 395 1965 418
rect 2482 446 2562 469
rect 2482 412 2505 446
rect 2539 412 2562 446
rect 2482 389 2562 412
rect 2632 449 2672 519
rect 3022 449 3102 469
rect 2632 446 3102 449
rect 2632 412 3045 446
rect 3079 412 3102 446
rect 2632 409 3102 412
rect 2056 360 2136 383
rect 2056 326 2079 360
rect 2113 326 2136 360
rect 2056 303 2136 326
rect 1355 261 1435 284
rect 1355 227 1378 261
rect 1412 227 1435 261
rect 1355 204 1435 227
rect 1505 261 1585 284
rect 1505 227 1528 261
rect 1562 227 1585 261
rect 1505 204 1585 227
rect 1705 261 1785 284
rect 1705 227 1728 261
rect 1762 227 1785 261
rect 1705 204 1785 227
rect -1487 132 -1407 155
rect -253 158 -173 169
rect -253 94 -230 158
rect -196 94 -173 158
rect -253 90 -173 94
rect -253 -12 -230 90
rect -196 -12 -173 90
rect -253 -16 -173 -12
rect -1373 -92 -1293 -69
rect -253 -80 -230 -16
rect -196 -80 -173 -16
rect -253 -91 -173 -80
rect 47 158 127 169
rect 47 94 70 158
rect 104 94 127 158
rect 47 90 127 94
rect 47 -12 70 90
rect 104 -12 127 90
rect 47 -16 127 -12
rect 47 -80 70 -16
rect 104 -80 127 -16
rect 47 -91 127 -80
rect 347 158 427 169
rect 347 94 370 158
rect 404 94 427 158
rect 347 90 427 94
rect 347 -12 370 90
rect 404 -12 427 90
rect 347 -16 427 -12
rect 347 -80 370 -16
rect 404 -80 427 -16
rect 347 -91 427 -80
rect 598 158 678 169
rect 598 94 621 158
rect 655 94 678 158
rect 598 90 678 94
rect 598 -12 621 90
rect 655 -12 678 90
rect 598 -16 678 -12
rect 598 -80 621 -16
rect 655 -80 678 -16
rect 598 -91 678 -80
rect 748 158 828 169
rect 748 124 771 158
rect 805 124 828 158
rect 748 90 828 124
rect 748 56 771 90
rect 805 56 828 90
rect 748 22 828 56
rect 748 -12 771 22
rect 805 -12 828 22
rect 748 -46 828 -12
rect 748 -80 771 -46
rect 805 -51 828 -46
rect 1305 158 1385 169
rect 1305 94 1328 158
rect 1362 94 1385 158
rect 1305 90 1385 94
rect 1305 -12 1328 90
rect 1362 -12 1385 90
rect 1305 -16 1385 -12
rect 805 -80 958 -51
rect 748 -91 958 -80
rect 1305 -80 1328 -16
rect 1362 -80 1385 -16
rect 1305 -91 1385 -80
rect 1605 158 1685 169
rect 1605 94 1628 158
rect 1662 94 1685 158
rect 1605 90 1685 94
rect 1605 -12 1628 90
rect 1662 -12 1685 90
rect 1605 -16 1685 -12
rect 1605 -80 1628 -16
rect 1662 -80 1685 -16
rect 1605 -91 1685 -80
rect 1905 158 1985 169
rect 1905 94 1928 158
rect 1962 94 1985 158
rect 1905 90 1985 94
rect 1905 -12 1928 90
rect 1962 -12 1985 90
rect 1905 -16 1985 -12
rect 1905 -80 1928 -16
rect 1962 -80 1985 -16
rect 1905 -91 1985 -80
rect -1373 -126 -1350 -92
rect -1316 -126 -1293 -92
rect -1373 -161 -1293 -126
rect -649 -149 -421 -109
rect -649 -161 -609 -149
rect -1373 -164 -609 -161
rect -1373 -198 -1350 -164
rect -1316 -198 -609 -164
rect -461 -161 -421 -149
rect 247 -161 327 -141
rect -461 -164 327 -161
rect -1373 -201 -609 -198
rect -1373 -236 -1293 -201
rect -1373 -270 -1350 -236
rect -1316 -270 -1293 -236
rect -1373 -293 -1293 -270
rect -575 -206 -495 -183
rect -461 -198 270 -164
rect 304 -198 327 -164
rect -461 -201 327 -198
rect -575 -240 -552 -206
rect -518 -240 -495 -206
rect 247 -221 327 -201
rect -575 -255 -495 -240
rect -575 -278 884 -255
rect -575 -312 -552 -278
rect -518 -312 -330 -278
rect -296 -312 -258 -278
rect -224 -312 -186 -278
rect -152 -312 -114 -278
rect -80 -312 -42 -278
rect -8 -312 30 -278
rect 64 -312 102 -278
rect 136 -312 174 -278
rect 208 -312 246 -278
rect 280 -312 318 -278
rect 352 -312 390 -278
rect 424 -312 462 -278
rect 496 -312 534 -278
rect 568 -312 606 -278
rect 640 -312 678 -278
rect 712 -312 750 -278
rect 784 -312 822 -278
rect 856 -312 884 -278
rect -575 -335 884 -312
rect -1259 -372 -1179 -349
rect -1259 -406 -1236 -372
rect -1202 -406 -1179 -372
rect -1259 -441 -1179 -406
rect -575 -350 -495 -335
rect -575 -384 -552 -350
rect -518 -384 -495 -350
rect -575 -407 -495 -384
rect -108 -391 -28 -369
rect -461 -392 -28 -391
rect -461 -426 -85 -392
rect -51 -393 -28 -392
rect 556 -393 636 -373
rect -51 -396 636 -393
rect -51 -426 579 -396
rect -461 -430 579 -426
rect 613 -430 636 -396
rect 918 -389 958 -91
rect 1660 -160 1740 -137
rect 1660 -194 1683 -160
rect 1717 -161 1740 -160
rect 1805 -161 1885 -141
rect 1717 -164 1885 -161
rect 1717 -194 1828 -164
rect 1660 -198 1828 -194
rect 1862 -198 1885 -164
rect 1660 -201 1885 -198
rect 2077 -161 2117 303
rect 2782 169 2822 409
rect 3022 389 3102 409
rect 3172 431 3212 519
rect 3172 408 3319 431
rect 3172 374 3262 408
rect 3296 374 3319 408
rect 3172 336 3319 374
rect 3172 302 3262 336
rect 3296 302 3319 336
rect 3172 279 3319 302
rect 3172 169 3212 279
rect 2462 158 2542 169
rect 2462 94 2485 158
rect 2519 94 2542 158
rect 2462 90 2542 94
rect 2462 -12 2485 90
rect 2519 -12 2542 90
rect 2462 -16 2542 -12
rect 2462 -80 2485 -16
rect 2519 -80 2542 -16
rect 2462 -91 2542 -80
rect 2762 158 2842 169
rect 2762 124 2785 158
rect 2819 124 2842 158
rect 2762 90 2842 124
rect 2762 56 2785 90
rect 2819 56 2842 90
rect 2762 22 2842 56
rect 2762 -12 2785 22
rect 2819 -12 2842 22
rect 2762 -46 2842 -12
rect 2762 -80 2785 -46
rect 2819 -80 2842 -46
rect 2762 -91 2842 -80
rect 3002 158 3082 169
rect 3002 94 3025 158
rect 3059 94 3082 158
rect 3002 90 3082 94
rect 3002 -12 3025 90
rect 3059 -12 3082 90
rect 3002 -16 3082 -12
rect 3002 -80 3025 -16
rect 3059 -80 3082 -16
rect 3002 -91 3082 -80
rect 3152 158 3232 169
rect 3152 124 3175 158
rect 3209 124 3232 158
rect 3152 90 3232 124
rect 3152 56 3175 90
rect 3209 56 3232 90
rect 3152 22 3232 56
rect 3152 -12 3175 22
rect 3209 -12 3232 22
rect 3152 -46 3232 -12
rect 3152 -80 3175 -46
rect 3209 -80 3232 -46
rect 3152 -91 3232 -80
rect 2662 -161 2742 -141
rect 2077 -164 2742 -161
rect 2077 -198 2685 -164
rect 2719 -198 2742 -164
rect 2077 -201 2742 -198
rect 1660 -217 1740 -201
rect 1805 -221 1885 -201
rect 2662 -221 2742 -201
rect 1205 -278 2085 -255
rect 1205 -312 1228 -278
rect 1262 -312 1300 -278
rect 1334 -312 1372 -278
rect 1406 -312 1444 -278
rect 1478 -312 1516 -278
rect 1550 -312 1588 -278
rect 1622 -312 1660 -278
rect 1694 -312 1732 -278
rect 1766 -312 1804 -278
rect 1838 -312 1876 -278
rect 1910 -312 1948 -278
rect 1982 -312 2020 -278
rect 2054 -312 2085 -278
rect 1205 -335 2085 -312
rect 2417 -278 3438 -255
rect 2417 -312 2440 -278
rect 2474 -312 2512 -278
rect 2546 -312 2584 -278
rect 2618 -312 2656 -278
rect 2690 -312 2728 -278
rect 2762 -312 2800 -278
rect 2834 -312 2872 -278
rect 2906 -312 2944 -278
rect 2978 -312 3016 -278
rect 3050 -312 3088 -278
rect 3122 -312 3160 -278
rect 3194 -312 3232 -278
rect 3266 -312 3304 -278
rect 3338 -312 3376 -278
rect 3410 -312 3438 -278
rect 2417 -335 3438 -312
rect 1450 -389 1530 -369
rect 918 -392 1530 -389
rect 918 -426 1473 -392
rect 1507 -426 1530 -392
rect 918 -429 1530 -426
rect -461 -431 636 -430
rect -461 -441 -421 -431
rect -1259 -444 -421 -441
rect -1259 -478 -1236 -444
rect -1202 -478 -421 -444
rect -108 -433 636 -431
rect -108 -449 -28 -433
rect 556 -453 636 -433
rect 1450 -449 1530 -429
rect 2662 -392 2742 -369
rect 2662 -426 2685 -392
rect 2719 -393 2742 -392
rect 3239 -393 3319 -373
rect 2719 -396 3319 -393
rect 2719 -426 3262 -396
rect 2662 -430 3262 -426
rect 3296 -430 3319 -396
rect 2662 -433 3319 -430
rect 2662 -449 2742 -433
rect 3239 -453 3319 -433
rect -1259 -481 -421 -478
rect -1259 -516 -1179 -481
rect -1259 -550 -1236 -516
rect -1202 -550 -1179 -516
rect -1259 -573 -1179 -550
rect -308 -510 -228 -499
rect -308 -574 -285 -510
rect -251 -574 -228 -510
rect -308 -578 -228 -574
rect -308 -680 -285 -578
rect -251 -680 -228 -578
rect -308 -684 -228 -680
rect -308 -748 -285 -684
rect -251 -748 -228 -684
rect -308 -759 -228 -748
rect 142 -510 222 -499
rect 142 -544 165 -510
rect 199 -544 222 -510
rect 142 -578 222 -544
rect 142 -612 165 -578
rect 199 -612 222 -578
rect 142 -646 222 -612
rect 142 -680 165 -646
rect 199 -680 222 -646
rect 142 -714 222 -680
rect 142 -748 165 -714
rect 199 -748 222 -714
rect 142 -759 222 -748
rect 382 -510 462 -499
rect 382 -574 405 -510
rect 439 -574 462 -510
rect 382 -578 462 -574
rect 382 -680 405 -578
rect 439 -680 462 -578
rect 382 -684 462 -680
rect 382 -748 405 -684
rect 439 -748 462 -684
rect 382 -759 462 -748
rect 532 -510 612 -499
rect 532 -544 555 -510
rect 589 -544 612 -510
rect 532 -578 612 -544
rect 532 -612 555 -578
rect 589 -612 612 -578
rect 532 -646 612 -612
rect 532 -680 555 -646
rect 589 -680 612 -646
rect 532 -714 612 -680
rect 532 -748 555 -714
rect 589 -748 612 -714
rect 532 -759 612 -748
rect 1250 -510 1330 -499
rect 1250 -574 1273 -510
rect 1307 -574 1330 -510
rect 1250 -578 1330 -574
rect 1250 -680 1273 -578
rect 1307 -680 1330 -578
rect 1250 -684 1330 -680
rect 1250 -748 1273 -684
rect 1307 -748 1330 -684
rect 1250 -759 1330 -748
rect 1550 -510 1630 -499
rect 1550 -544 1573 -510
rect 1607 -544 1630 -510
rect 1550 -578 1630 -544
rect 1550 -612 1573 -578
rect 1607 -612 1630 -578
rect 1550 -646 1630 -612
rect 1550 -680 1573 -646
rect 1607 -680 1630 -646
rect 1550 -714 1630 -680
rect 1550 -748 1573 -714
rect 1607 -748 1630 -714
rect 1550 -759 1630 -748
rect 1790 -510 1870 -499
rect 1790 -574 1813 -510
rect 1847 -574 1870 -510
rect 1790 -578 1870 -574
rect 1790 -680 1813 -578
rect 1847 -680 1870 -578
rect 1790 -684 1870 -680
rect 1790 -748 1813 -684
rect 1847 -748 1870 -684
rect 1790 -759 1870 -748
rect 1940 -510 2020 -499
rect 1940 -544 1963 -510
rect 1997 -544 2020 -510
rect 1940 -578 2020 -544
rect 1940 -612 1963 -578
rect 1997 -612 2020 -578
rect 1940 -646 2020 -612
rect 1940 -680 1963 -646
rect 1997 -680 2020 -646
rect 1940 -714 2020 -680
rect 1940 -748 1963 -714
rect 1997 -748 2020 -714
rect 1940 -759 2020 -748
rect 2462 -510 2542 -499
rect 2462 -544 2485 -510
rect 2519 -544 2542 -510
rect 2462 -578 2542 -544
rect 2462 -612 2485 -578
rect 2519 -612 2542 -578
rect 2462 -646 2542 -612
rect 2462 -680 2485 -646
rect 2519 -680 2542 -646
rect 2462 -714 2542 -680
rect 2462 -748 2485 -714
rect 2519 -748 2542 -714
rect 2462 -759 2542 -748
rect 2612 -510 2692 -499
rect 2612 -574 2635 -510
rect 2669 -574 2692 -510
rect 2612 -578 2692 -574
rect 2612 -680 2635 -578
rect 2669 -680 2692 -578
rect 2612 -684 2692 -680
rect 2612 -748 2635 -684
rect 2669 -748 2692 -684
rect 2612 -759 2692 -748
rect 2762 -510 2842 -499
rect 2762 -544 2785 -510
rect 2819 -544 2842 -510
rect 2762 -578 2842 -544
rect 2762 -612 2785 -578
rect 2819 -612 2842 -578
rect 2762 -646 2842 -612
rect 2762 -680 2785 -646
rect 2819 -680 2842 -646
rect 2762 -714 2842 -680
rect 2762 -748 2785 -714
rect 2819 -748 2842 -714
rect 2762 -759 2842 -748
rect 2912 -510 2992 -499
rect 2912 -574 2935 -510
rect 2969 -574 2992 -510
rect 2912 -578 2992 -574
rect 2912 -680 2935 -578
rect 2969 -680 2992 -578
rect 2912 -684 2992 -680
rect 2912 -748 2935 -684
rect 2969 -748 2992 -684
rect 2912 -759 2992 -748
rect 3152 -510 3232 -499
rect 3152 -574 3175 -510
rect 3209 -574 3232 -510
rect 3152 -578 3232 -574
rect 3152 -680 3175 -578
rect 3209 -680 3232 -578
rect 3152 -684 3232 -680
rect 3152 -748 3175 -684
rect 3209 -748 3232 -684
rect 3152 -759 3232 -748
rect 3302 -510 3382 -499
rect 3302 -544 3325 -510
rect 3359 -544 3382 -510
rect 3302 -578 3382 -544
rect 3302 -612 3325 -578
rect 3359 -612 3382 -578
rect 3302 -646 3382 -612
rect 3302 -680 3325 -646
rect 3359 -680 3382 -646
rect 3302 -714 3382 -680
rect 3302 -748 3325 -714
rect 3359 -748 3382 -714
rect 3302 -759 3382 -748
rect -1373 -920 -1293 -897
rect -1373 -954 -1350 -920
rect -1316 -954 -1293 -920
rect -1373 -989 -1293 -954
rect -258 -989 -178 -969
rect -1373 -992 -178 -989
rect -1373 -1026 -1350 -992
rect -1316 -1026 -235 -992
rect -201 -1026 -178 -992
rect 162 -999 202 -759
rect 402 -999 482 -979
rect -1373 -1029 -178 -1026
rect -1373 -1064 -1293 -1029
rect -258 -1049 -178 -1029
rect 12 -1002 482 -999
rect 12 -1036 425 -1002
rect 459 -1036 482 -1002
rect 12 -1039 482 -1036
rect -1373 -1098 -1350 -1064
rect -1316 -1098 -1293 -1064
rect -1373 -1121 -1293 -1098
rect 12 -1109 52 -1039
rect 402 -1059 482 -1039
rect 552 -1109 592 -759
rect 1270 -1002 1350 -979
rect 1570 -999 1610 -759
rect 1810 -999 1890 -979
rect 1270 -1036 1293 -1002
rect 1327 -1036 1350 -1002
rect 1270 -1059 1350 -1036
rect 1420 -1002 1890 -999
rect 1420 -1036 1833 -1002
rect 1867 -1036 1890 -1002
rect 1420 -1039 1890 -1036
rect 1420 -1109 1460 -1039
rect 1810 -1059 1890 -1039
rect 1960 -989 2000 -759
rect 2482 -793 2522 -759
rect 2782 -793 2822 -759
rect 2482 -833 2822 -793
rect 2512 -989 2592 -969
rect 1960 -992 2592 -989
rect 1960 -1026 2535 -992
rect 2569 -1026 2592 -992
rect 1960 -1029 2592 -1026
rect 1960 -1109 2000 -1029
rect 2512 -1049 2592 -1029
rect 2782 -999 2822 -833
rect 3322 -860 3362 -759
rect 3303 -883 3383 -860
rect 3303 -917 3326 -883
rect 3360 -917 3383 -883
rect 3303 -955 3383 -917
rect 3172 -999 3252 -979
rect 2782 -1002 3252 -999
rect 2782 -1036 3195 -1002
rect 3229 -1036 3252 -1002
rect 3303 -989 3326 -955
rect 3360 -989 3383 -955
rect 3303 -1012 3383 -989
rect 2782 -1039 3252 -1036
rect 2932 -1109 2972 -1039
rect 3172 -1059 3252 -1039
rect 3322 -1109 3362 -1012
rect -308 -1134 -228 -1109
rect -308 -1168 -285 -1134
rect -251 -1168 -228 -1134
rect -308 -1202 -228 -1168
rect -308 -1236 -285 -1202
rect -251 -1236 -228 -1202
rect -308 -1270 -228 -1236
rect -308 -1304 -285 -1270
rect -251 -1304 -228 -1270
rect -308 -1338 -228 -1304
rect -308 -1372 -285 -1338
rect -251 -1372 -228 -1338
rect -308 -1406 -228 -1372
rect -308 -1440 -285 -1406
rect -251 -1440 -228 -1406
rect -308 -1474 -228 -1440
rect -308 -1508 -285 -1474
rect -251 -1508 -228 -1474
rect -308 -1542 -228 -1508
rect -308 -1576 -285 -1542
rect -251 -1576 -228 -1542
rect -308 -1610 -228 -1576
rect -308 -1644 -285 -1610
rect -251 -1644 -228 -1610
rect -308 -1669 -228 -1644
rect -158 -1120 -78 -1109
rect -158 -1168 -135 -1120
rect -101 -1168 -78 -1120
rect -158 -1192 -78 -1168
rect -158 -1236 -135 -1192
rect -101 -1236 -78 -1192
rect -158 -1264 -78 -1236
rect -158 -1304 -135 -1264
rect -101 -1304 -78 -1264
rect -158 -1336 -78 -1304
rect -158 -1372 -135 -1336
rect -101 -1372 -78 -1336
rect -158 -1406 -78 -1372
rect -158 -1442 -135 -1406
rect -101 -1442 -78 -1406
rect -158 -1474 -78 -1442
rect -158 -1514 -135 -1474
rect -101 -1514 -78 -1474
rect -158 -1542 -78 -1514
rect -158 -1586 -135 -1542
rect -101 -1586 -78 -1542
rect -158 -1610 -78 -1586
rect -158 -1658 -135 -1610
rect -101 -1658 -78 -1610
rect -158 -1669 -78 -1658
rect -8 -1134 72 -1109
rect -8 -1168 15 -1134
rect 49 -1168 72 -1134
rect -8 -1202 72 -1168
rect -8 -1236 15 -1202
rect 49 -1236 72 -1202
rect -8 -1270 72 -1236
rect -8 -1304 15 -1270
rect 49 -1304 72 -1270
rect -8 -1338 72 -1304
rect -8 -1372 15 -1338
rect 49 -1372 72 -1338
rect -8 -1406 72 -1372
rect -8 -1440 15 -1406
rect 49 -1440 72 -1406
rect -8 -1474 72 -1440
rect -8 -1508 15 -1474
rect 49 -1508 72 -1474
rect -8 -1542 72 -1508
rect -8 -1576 15 -1542
rect 49 -1576 72 -1542
rect -8 -1610 72 -1576
rect -8 -1644 15 -1610
rect 49 -1644 72 -1610
rect -8 -1669 72 -1644
rect 142 -1120 222 -1109
rect 142 -1168 165 -1120
rect 199 -1168 222 -1120
rect 142 -1192 222 -1168
rect 142 -1236 165 -1192
rect 199 -1236 222 -1192
rect 142 -1264 222 -1236
rect 142 -1304 165 -1264
rect 199 -1304 222 -1264
rect 142 -1336 222 -1304
rect 142 -1372 165 -1336
rect 199 -1372 222 -1336
rect 142 -1406 222 -1372
rect 142 -1442 165 -1406
rect 199 -1442 222 -1406
rect 142 -1474 222 -1442
rect 142 -1514 165 -1474
rect 199 -1514 222 -1474
rect 142 -1542 222 -1514
rect 142 -1586 165 -1542
rect 199 -1586 222 -1542
rect 142 -1610 222 -1586
rect 142 -1658 165 -1610
rect 199 -1658 222 -1610
rect 142 -1669 222 -1658
rect 382 -1120 462 -1109
rect 382 -1168 405 -1120
rect 439 -1168 462 -1120
rect 382 -1192 462 -1168
rect 382 -1236 405 -1192
rect 439 -1236 462 -1192
rect 382 -1264 462 -1236
rect 382 -1304 405 -1264
rect 439 -1304 462 -1264
rect 382 -1336 462 -1304
rect 382 -1372 405 -1336
rect 439 -1372 462 -1336
rect 382 -1406 462 -1372
rect 382 -1442 405 -1406
rect 439 -1442 462 -1406
rect 382 -1474 462 -1442
rect 382 -1514 405 -1474
rect 439 -1514 462 -1474
rect 382 -1542 462 -1514
rect 382 -1586 405 -1542
rect 439 -1586 462 -1542
rect 382 -1610 462 -1586
rect 382 -1658 405 -1610
rect 439 -1658 462 -1610
rect 382 -1669 462 -1658
rect 532 -1134 612 -1109
rect 532 -1168 555 -1134
rect 589 -1168 612 -1134
rect 532 -1202 612 -1168
rect 532 -1236 555 -1202
rect 589 -1236 612 -1202
rect 532 -1270 612 -1236
rect 532 -1304 555 -1270
rect 589 -1304 612 -1270
rect 532 -1338 612 -1304
rect 532 -1372 555 -1338
rect 589 -1372 612 -1338
rect 532 -1406 612 -1372
rect 532 -1440 555 -1406
rect 589 -1440 612 -1406
rect 532 -1474 612 -1440
rect 532 -1508 555 -1474
rect 589 -1508 612 -1474
rect 532 -1542 612 -1508
rect 532 -1576 555 -1542
rect 589 -1576 612 -1542
rect 532 -1610 612 -1576
rect 532 -1644 555 -1610
rect 589 -1644 612 -1610
rect 532 -1669 612 -1644
rect 1250 -1120 1330 -1109
rect 1250 -1168 1273 -1120
rect 1307 -1168 1330 -1120
rect 1250 -1192 1330 -1168
rect 1250 -1236 1273 -1192
rect 1307 -1236 1330 -1192
rect 1250 -1264 1330 -1236
rect 1250 -1304 1273 -1264
rect 1307 -1304 1330 -1264
rect 1250 -1336 1330 -1304
rect 1250 -1372 1273 -1336
rect 1307 -1372 1330 -1336
rect 1250 -1406 1330 -1372
rect 1250 -1442 1273 -1406
rect 1307 -1442 1330 -1406
rect 1250 -1474 1330 -1442
rect 1250 -1514 1273 -1474
rect 1307 -1514 1330 -1474
rect 1250 -1542 1330 -1514
rect 1250 -1586 1273 -1542
rect 1307 -1586 1330 -1542
rect 1250 -1610 1330 -1586
rect 1250 -1658 1273 -1610
rect 1307 -1658 1330 -1610
rect 1250 -1669 1330 -1658
rect 1400 -1134 1480 -1109
rect 1400 -1168 1423 -1134
rect 1457 -1168 1480 -1134
rect 1400 -1202 1480 -1168
rect 1400 -1236 1423 -1202
rect 1457 -1236 1480 -1202
rect 1400 -1270 1480 -1236
rect 1400 -1304 1423 -1270
rect 1457 -1304 1480 -1270
rect 1400 -1338 1480 -1304
rect 1400 -1372 1423 -1338
rect 1457 -1372 1480 -1338
rect 1400 -1406 1480 -1372
rect 1400 -1440 1423 -1406
rect 1457 -1440 1480 -1406
rect 1400 -1474 1480 -1440
rect 1400 -1508 1423 -1474
rect 1457 -1508 1480 -1474
rect 1400 -1542 1480 -1508
rect 1400 -1576 1423 -1542
rect 1457 -1576 1480 -1542
rect 1400 -1610 1480 -1576
rect 1400 -1644 1423 -1610
rect 1457 -1644 1480 -1610
rect 1400 -1669 1480 -1644
rect 1550 -1120 1630 -1109
rect 1550 -1168 1573 -1120
rect 1607 -1168 1630 -1120
rect 1550 -1192 1630 -1168
rect 1550 -1236 1573 -1192
rect 1607 -1236 1630 -1192
rect 1550 -1264 1630 -1236
rect 1550 -1304 1573 -1264
rect 1607 -1304 1630 -1264
rect 1550 -1336 1630 -1304
rect 1550 -1372 1573 -1336
rect 1607 -1372 1630 -1336
rect 1550 -1406 1630 -1372
rect 1550 -1442 1573 -1406
rect 1607 -1442 1630 -1406
rect 1550 -1474 1630 -1442
rect 1550 -1514 1573 -1474
rect 1607 -1514 1630 -1474
rect 1550 -1542 1630 -1514
rect 1550 -1586 1573 -1542
rect 1607 -1586 1630 -1542
rect 1550 -1610 1630 -1586
rect 1550 -1658 1573 -1610
rect 1607 -1658 1630 -1610
rect 1550 -1669 1630 -1658
rect 1790 -1120 1870 -1109
rect 1790 -1168 1813 -1120
rect 1847 -1168 1870 -1120
rect 1790 -1192 1870 -1168
rect 1790 -1236 1813 -1192
rect 1847 -1236 1870 -1192
rect 1790 -1264 1870 -1236
rect 1790 -1304 1813 -1264
rect 1847 -1304 1870 -1264
rect 1790 -1336 1870 -1304
rect 1790 -1372 1813 -1336
rect 1847 -1372 1870 -1336
rect 1790 -1406 1870 -1372
rect 1790 -1442 1813 -1406
rect 1847 -1442 1870 -1406
rect 1790 -1474 1870 -1442
rect 1790 -1514 1813 -1474
rect 1847 -1514 1870 -1474
rect 1790 -1542 1870 -1514
rect 1790 -1586 1813 -1542
rect 1847 -1586 1870 -1542
rect 1790 -1610 1870 -1586
rect 1790 -1658 1813 -1610
rect 1847 -1658 1870 -1610
rect 1790 -1669 1870 -1658
rect 1940 -1134 2020 -1109
rect 1940 -1168 1963 -1134
rect 1997 -1168 2020 -1134
rect 1940 -1202 2020 -1168
rect 1940 -1236 1963 -1202
rect 1997 -1236 2020 -1202
rect 1940 -1270 2020 -1236
rect 1940 -1304 1963 -1270
rect 1997 -1304 2020 -1270
rect 1940 -1338 2020 -1304
rect 1940 -1372 1963 -1338
rect 1997 -1372 2020 -1338
rect 1940 -1406 2020 -1372
rect 1940 -1440 1963 -1406
rect 1997 -1440 2020 -1406
rect 1940 -1474 2020 -1440
rect 1940 -1508 1963 -1474
rect 1997 -1508 2020 -1474
rect 1940 -1542 2020 -1508
rect 1940 -1576 1963 -1542
rect 1997 -1576 2020 -1542
rect 1940 -1610 2020 -1576
rect 1940 -1644 1963 -1610
rect 1997 -1644 2020 -1610
rect 1940 -1669 2020 -1644
rect 2462 -1120 2542 -1109
rect 2462 -1168 2485 -1120
rect 2519 -1168 2542 -1120
rect 2462 -1192 2542 -1168
rect 2462 -1236 2485 -1192
rect 2519 -1236 2542 -1192
rect 2462 -1264 2542 -1236
rect 2462 -1304 2485 -1264
rect 2519 -1304 2542 -1264
rect 2462 -1336 2542 -1304
rect 2462 -1372 2485 -1336
rect 2519 -1372 2542 -1336
rect 2462 -1406 2542 -1372
rect 2462 -1442 2485 -1406
rect 2519 -1442 2542 -1406
rect 2462 -1474 2542 -1442
rect 2462 -1514 2485 -1474
rect 2519 -1514 2542 -1474
rect 2462 -1542 2542 -1514
rect 2462 -1586 2485 -1542
rect 2519 -1586 2542 -1542
rect 2462 -1610 2542 -1586
rect 2462 -1658 2485 -1610
rect 2519 -1658 2542 -1610
rect 2462 -1669 2542 -1658
rect 2912 -1134 2992 -1109
rect 2912 -1168 2935 -1134
rect 2969 -1168 2992 -1134
rect 2912 -1202 2992 -1168
rect 2912 -1236 2935 -1202
rect 2969 -1236 2992 -1202
rect 2912 -1270 2992 -1236
rect 2912 -1304 2935 -1270
rect 2969 -1304 2992 -1270
rect 2912 -1338 2992 -1304
rect 2912 -1372 2935 -1338
rect 2969 -1372 2992 -1338
rect 2912 -1406 2992 -1372
rect 2912 -1440 2935 -1406
rect 2969 -1440 2992 -1406
rect 2912 -1474 2992 -1440
rect 2912 -1508 2935 -1474
rect 2969 -1508 2992 -1474
rect 2912 -1542 2992 -1508
rect 2912 -1576 2935 -1542
rect 2969 -1576 2992 -1542
rect 2912 -1610 2992 -1576
rect 2912 -1644 2935 -1610
rect 2969 -1644 2992 -1610
rect 2912 -1669 2992 -1644
rect 3152 -1120 3232 -1109
rect 3152 -1168 3175 -1120
rect 3209 -1168 3232 -1120
rect 3152 -1192 3232 -1168
rect 3152 -1236 3175 -1192
rect 3209 -1236 3232 -1192
rect 3152 -1264 3232 -1236
rect 3152 -1304 3175 -1264
rect 3209 -1304 3232 -1264
rect 3152 -1336 3232 -1304
rect 3152 -1372 3175 -1336
rect 3209 -1372 3232 -1336
rect 3152 -1406 3232 -1372
rect 3152 -1442 3175 -1406
rect 3209 -1442 3232 -1406
rect 3152 -1474 3232 -1442
rect 3152 -1514 3175 -1474
rect 3209 -1514 3232 -1474
rect 3152 -1542 3232 -1514
rect 3152 -1586 3175 -1542
rect 3209 -1586 3232 -1542
rect 3152 -1610 3232 -1586
rect 3152 -1658 3175 -1610
rect 3209 -1658 3232 -1610
rect 3152 -1669 3232 -1658
rect 3302 -1134 3382 -1109
rect 3302 -1168 3325 -1134
rect 3359 -1168 3382 -1134
rect 3302 -1202 3382 -1168
rect 3302 -1236 3325 -1202
rect 3359 -1236 3382 -1202
rect 3302 -1270 3382 -1236
rect 3302 -1304 3325 -1270
rect 3359 -1304 3382 -1270
rect 3302 -1338 3382 -1304
rect 3302 -1372 3325 -1338
rect 3359 -1372 3382 -1338
rect 3302 -1406 3382 -1372
rect 3302 -1440 3325 -1406
rect 3359 -1440 3382 -1406
rect 3302 -1474 3382 -1440
rect 3302 -1508 3325 -1474
rect 3359 -1508 3382 -1474
rect 3302 -1542 3382 -1508
rect 3302 -1576 3325 -1542
rect 3359 -1576 3382 -1542
rect 3302 -1610 3382 -1576
rect 3302 -1644 3325 -1610
rect 3359 -1644 3382 -1610
rect 3302 -1669 3382 -1644
rect -288 -1709 -248 -1669
rect 12 -1709 52 -1669
rect -288 -1749 52 -1709
rect 92 -1739 172 -1719
rect 230 -1738 310 -1715
rect 230 -1739 253 -1738
rect 92 -1742 253 -1739
rect 92 -1776 115 -1742
rect 149 -1772 253 -1742
rect 287 -1772 310 -1738
rect 149 -1776 310 -1772
rect 92 -1779 310 -1776
rect 552 -1739 592 -1669
rect 2832 -1739 2912 -1719
rect 552 -1742 2912 -1739
rect 552 -1776 2855 -1742
rect 2889 -1776 2912 -1742
rect 552 -1779 2912 -1776
rect 92 -1799 172 -1779
rect 230 -1795 310 -1779
rect 2832 -1799 2912 -1779
rect -353 -1856 657 -1833
rect -353 -1890 -330 -1856
rect -296 -1890 -258 -1856
rect -224 -1890 -186 -1856
rect -152 -1890 -114 -1856
rect -80 -1890 -42 -1856
rect -8 -1890 30 -1856
rect 64 -1890 102 -1856
rect 136 -1890 174 -1856
rect 208 -1890 246 -1856
rect 280 -1890 318 -1856
rect 352 -1890 390 -1856
rect 424 -1890 462 -1856
rect 496 -1890 534 -1856
rect 568 -1890 606 -1856
rect 640 -1890 657 -1856
rect -353 -1913 657 -1890
rect 1205 -1856 2085 -1833
rect 1205 -1890 1228 -1856
rect 1262 -1890 1300 -1856
rect 1334 -1890 1372 -1856
rect 1406 -1890 1444 -1856
rect 1478 -1890 1516 -1856
rect 1550 -1890 1588 -1856
rect 1622 -1890 1660 -1856
rect 1694 -1890 1732 -1856
rect 1766 -1890 1804 -1856
rect 1838 -1890 1876 -1856
rect 1910 -1890 1948 -1856
rect 1982 -1890 2020 -1856
rect 2054 -1890 2085 -1856
rect 1205 -1913 2085 -1890
rect 2417 -1856 3427 -1833
rect 2417 -1890 2440 -1856
rect 2474 -1890 2512 -1856
rect 2546 -1890 2584 -1856
rect 2618 -1890 2656 -1856
rect 2690 -1890 2728 -1856
rect 2762 -1890 2800 -1856
rect 2834 -1890 2872 -1856
rect 2906 -1890 2944 -1856
rect 2978 -1890 3016 -1856
rect 3050 -1890 3088 -1856
rect 3122 -1890 3160 -1856
rect 3194 -1890 3232 -1856
rect 3266 -1890 3304 -1856
rect 3338 -1890 3376 -1856
rect 3410 -1890 3427 -1856
rect 2417 -1913 3427 -1890
<< viali >>
rect -1008 1224 -974 1258
rect -330 1266 -296 1300
rect -258 1266 -224 1300
rect -186 1266 -152 1300
rect -114 1266 -80 1300
rect -42 1266 -8 1300
rect 30 1266 64 1300
rect 102 1266 136 1300
rect 174 1266 208 1300
rect 246 1266 280 1300
rect 318 1266 352 1300
rect 390 1266 424 1300
rect 462 1266 496 1300
rect 534 1266 568 1300
rect 606 1266 640 1300
rect 678 1266 712 1300
rect 750 1266 784 1300
rect 822 1266 856 1300
rect 1228 1266 1262 1300
rect 1300 1266 1334 1300
rect 1372 1266 1406 1300
rect 1444 1266 1478 1300
rect 1516 1266 1550 1300
rect 1588 1266 1622 1300
rect 1660 1266 1694 1300
rect 1732 1266 1766 1300
rect 1804 1266 1838 1300
rect 1876 1266 1910 1300
rect 1948 1266 1982 1300
rect 2020 1266 2054 1300
rect 2440 1266 2474 1300
rect 2512 1266 2546 1300
rect 2584 1266 2618 1300
rect 2656 1266 2690 1300
rect 2728 1266 2762 1300
rect 2800 1266 2834 1300
rect 2872 1266 2906 1300
rect 2944 1266 2978 1300
rect 3016 1266 3050 1300
rect 3088 1266 3122 1300
rect 3160 1266 3194 1300
rect 3232 1266 3266 1300
rect -1008 1152 -974 1186
rect 1683 1148 1717 1182
rect -1008 1080 -974 1114
rect -230 1054 -196 1068
rect -230 1034 -196 1054
rect -230 986 -196 996
rect -230 962 -196 986
rect -230 918 -196 924
rect -230 890 -196 918
rect -230 850 -196 852
rect -230 818 -196 850
rect -230 748 -196 780
rect -230 746 -196 748
rect -230 680 -196 708
rect -230 674 -196 680
rect -230 612 -196 636
rect -230 602 -196 612
rect -894 490 -860 524
rect -230 544 -196 564
rect -230 530 -196 544
rect 70 1054 104 1068
rect 70 1034 104 1054
rect 70 986 104 996
rect 70 962 104 986
rect 70 918 104 924
rect 70 890 104 918
rect 70 850 104 852
rect 70 818 104 850
rect 70 748 104 780
rect 70 746 104 748
rect 70 680 104 708
rect 70 674 104 680
rect 70 612 104 636
rect 70 602 104 612
rect 70 544 104 564
rect 70 530 104 544
rect 370 1054 404 1068
rect 370 1034 404 1054
rect 370 986 404 996
rect 370 962 404 986
rect 370 918 404 924
rect 370 890 404 918
rect 370 850 404 852
rect 370 818 404 850
rect 370 748 404 780
rect 370 746 404 748
rect 370 680 404 708
rect 370 674 404 680
rect 370 612 404 636
rect 370 602 404 612
rect 370 544 404 564
rect 370 530 404 544
rect 621 1054 655 1068
rect 621 1034 655 1054
rect 621 986 655 996
rect 621 962 655 986
rect 621 918 655 924
rect 621 890 655 918
rect 621 850 655 852
rect 621 818 655 850
rect 621 748 655 780
rect 621 746 655 748
rect 621 680 655 708
rect 621 674 655 680
rect 621 612 655 636
rect 621 602 655 612
rect 621 544 655 564
rect 621 530 655 544
rect 1328 1054 1362 1068
rect 1328 1034 1362 1054
rect 1328 986 1362 996
rect 1328 962 1362 986
rect 1328 918 1362 924
rect 1328 890 1362 918
rect 1328 850 1362 852
rect 1328 818 1362 850
rect 1328 748 1362 780
rect 1328 746 1362 748
rect 1328 680 1362 708
rect 1328 674 1362 680
rect 1328 612 1362 636
rect 1328 602 1362 612
rect 1328 544 1362 564
rect 1328 530 1362 544
rect 1628 1054 1662 1068
rect 1628 1034 1662 1054
rect 1628 986 1662 996
rect 1628 962 1662 986
rect 1628 918 1662 924
rect 1628 890 1662 918
rect 1628 850 1662 852
rect 1628 818 1662 850
rect 1628 748 1662 780
rect 1628 746 1662 748
rect 1628 680 1662 708
rect 1628 674 1662 680
rect 1628 612 1662 636
rect 1628 602 1662 612
rect 1628 544 1662 564
rect 1628 530 1662 544
rect 1928 1054 1962 1068
rect 1928 1034 1962 1054
rect 1928 986 1962 996
rect 1928 962 1962 986
rect 1928 918 1962 924
rect 1928 890 1962 918
rect 1928 850 1962 852
rect 1928 818 1962 850
rect 1928 748 1962 780
rect 1928 746 1962 748
rect 1928 680 1962 708
rect 1928 674 1962 680
rect 1928 612 1962 636
rect 1928 602 1962 612
rect 1928 544 1962 564
rect 1928 530 1962 544
rect 2485 1054 2519 1068
rect 2485 1034 2519 1054
rect 2485 986 2519 996
rect 2485 962 2519 986
rect 2485 918 2519 924
rect 2485 890 2519 918
rect 2485 850 2519 852
rect 2485 818 2519 850
rect 2485 748 2519 780
rect 2485 746 2519 748
rect 2485 680 2519 708
rect 2485 674 2519 680
rect 2485 612 2519 636
rect 2485 602 2519 612
rect 2485 544 2519 564
rect 2485 530 2519 544
rect 2785 1054 2819 1068
rect 2785 1034 2819 1054
rect 2785 986 2819 996
rect 2785 962 2819 986
rect 2785 918 2819 924
rect 2785 890 2819 918
rect 2785 850 2819 852
rect 2785 818 2819 850
rect 2785 748 2819 780
rect 2785 746 2819 748
rect 2785 680 2819 708
rect 2785 674 2819 680
rect 2785 612 2819 636
rect 2785 602 2819 612
rect 2785 544 2819 564
rect 2785 530 2819 544
rect 3025 1054 3059 1068
rect 3025 1034 3059 1054
rect 3025 986 3059 996
rect 3025 962 3059 986
rect 3025 918 3059 924
rect 3025 890 3059 918
rect 3025 850 3059 852
rect 3025 818 3059 850
rect 3025 748 3059 780
rect 3025 746 3059 748
rect 3025 680 3059 708
rect 3025 674 3059 680
rect 3025 612 3059 636
rect 3025 602 3059 612
rect 3025 544 3059 564
rect 3025 530 3059 544
rect -894 418 -860 452
rect -1464 299 -1430 333
rect -894 346 -860 380
rect 350 418 384 452
rect 499 306 533 340
rect -1464 227 -1430 261
rect -30 227 4 261
rect -1464 155 -1430 189
rect 1348 418 1382 452
rect 1908 418 1942 452
rect 2505 412 2539 446
rect 2079 326 2113 360
rect 1378 227 1412 261
rect 1528 227 1562 261
rect -230 124 -196 128
rect -230 94 -196 124
rect -230 22 -196 56
rect -230 -46 -196 -16
rect -230 -50 -196 -46
rect 70 124 104 128
rect 70 94 104 124
rect 70 22 104 56
rect 70 -46 104 -16
rect 70 -50 104 -46
rect 370 124 404 128
rect 370 94 404 124
rect 370 22 404 56
rect 370 -46 404 -16
rect 370 -50 404 -46
rect 621 124 655 128
rect 621 94 655 124
rect 621 22 655 56
rect 621 -46 655 -16
rect 621 -50 655 -46
rect 1328 124 1362 128
rect 1328 94 1362 124
rect 1328 22 1362 56
rect 1328 -46 1362 -16
rect 1328 -50 1362 -46
rect 1628 124 1662 128
rect 1628 94 1662 124
rect 1628 22 1662 56
rect 1628 -46 1662 -16
rect 1628 -50 1662 -46
rect 1928 124 1962 128
rect 1928 94 1962 124
rect 1928 22 1962 56
rect 1928 -46 1962 -16
rect 1928 -50 1962 -46
rect -1350 -126 -1316 -92
rect -1350 -198 -1316 -164
rect -1350 -270 -1316 -236
rect -552 -240 -518 -206
rect -552 -312 -518 -278
rect -330 -312 -296 -278
rect -258 -312 -224 -278
rect -186 -312 -152 -278
rect -114 -312 -80 -278
rect -42 -312 -8 -278
rect 30 -312 64 -278
rect 102 -312 136 -278
rect 174 -312 208 -278
rect 246 -312 280 -278
rect 318 -312 352 -278
rect 390 -312 424 -278
rect 462 -312 496 -278
rect 534 -312 568 -278
rect 606 -312 640 -278
rect 678 -312 712 -278
rect 750 -312 784 -278
rect 822 -312 856 -278
rect -1236 -406 -1202 -372
rect -552 -384 -518 -350
rect 579 -430 613 -396
rect 1683 -194 1717 -160
rect 3262 374 3296 408
rect 3262 302 3296 336
rect 2485 124 2519 128
rect 2485 94 2519 124
rect 2485 22 2519 56
rect 2485 -46 2519 -16
rect 2485 -50 2519 -46
rect 3025 124 3059 128
rect 3025 94 3059 124
rect 3025 22 3059 56
rect 3025 -46 3059 -16
rect 3025 -50 3059 -46
rect 1228 -312 1262 -278
rect 1300 -312 1334 -278
rect 1372 -312 1406 -278
rect 1444 -312 1478 -278
rect 1516 -312 1550 -278
rect 1588 -312 1622 -278
rect 1660 -312 1694 -278
rect 1732 -312 1766 -278
rect 1804 -312 1838 -278
rect 1876 -312 1910 -278
rect 1948 -312 1982 -278
rect 2020 -312 2054 -278
rect 2440 -312 2474 -278
rect 2512 -312 2546 -278
rect 2584 -312 2618 -278
rect 2656 -312 2690 -278
rect 2728 -312 2762 -278
rect 2800 -312 2834 -278
rect 2872 -312 2906 -278
rect 2944 -312 2978 -278
rect 3016 -312 3050 -278
rect 3088 -312 3122 -278
rect 3160 -312 3194 -278
rect 3232 -312 3266 -278
rect 3304 -312 3338 -278
rect 3376 -312 3410 -278
rect -1236 -478 -1202 -444
rect 3262 -430 3296 -396
rect -1236 -550 -1202 -516
rect -285 -544 -251 -540
rect -285 -574 -251 -544
rect -285 -646 -251 -612
rect -285 -714 -251 -684
rect -285 -718 -251 -714
rect 405 -544 439 -540
rect 405 -574 439 -544
rect 405 -646 439 -612
rect 405 -714 439 -684
rect 405 -718 439 -714
rect 1273 -544 1307 -540
rect 1273 -574 1307 -544
rect 1273 -646 1307 -612
rect 1273 -714 1307 -684
rect 1273 -718 1307 -714
rect 1813 -544 1847 -540
rect 1813 -574 1847 -544
rect 1813 -646 1847 -612
rect 1813 -714 1847 -684
rect 1813 -718 1847 -714
rect 2635 -544 2669 -540
rect 2635 -574 2669 -544
rect 2635 -646 2669 -612
rect 2635 -714 2669 -684
rect 2635 -718 2669 -714
rect 2935 -544 2969 -540
rect 2935 -574 2969 -544
rect 2935 -646 2969 -612
rect 2935 -714 2969 -684
rect 2935 -718 2969 -714
rect 3175 -544 3209 -540
rect 3175 -574 3209 -544
rect 3175 -646 3209 -612
rect 3175 -714 3209 -684
rect 3175 -718 3209 -714
rect -1350 -954 -1316 -920
rect -1350 -1026 -1316 -992
rect -1350 -1098 -1316 -1064
rect 1293 -1036 1327 -1002
rect 3326 -917 3360 -883
rect 3326 -989 3360 -955
rect -135 -1134 -101 -1120
rect -135 -1154 -101 -1134
rect -135 -1202 -101 -1192
rect -135 -1226 -101 -1202
rect -135 -1270 -101 -1264
rect -135 -1298 -101 -1270
rect -135 -1338 -101 -1336
rect -135 -1370 -101 -1338
rect -135 -1440 -101 -1408
rect -135 -1442 -101 -1440
rect -135 -1508 -101 -1480
rect -135 -1514 -101 -1508
rect -135 -1576 -101 -1552
rect -135 -1586 -101 -1576
rect -135 -1644 -101 -1624
rect -135 -1658 -101 -1644
rect 165 -1134 199 -1120
rect 165 -1154 199 -1134
rect 165 -1202 199 -1192
rect 165 -1226 199 -1202
rect 165 -1270 199 -1264
rect 165 -1298 199 -1270
rect 165 -1338 199 -1336
rect 165 -1370 199 -1338
rect 165 -1440 199 -1408
rect 165 -1442 199 -1440
rect 165 -1508 199 -1480
rect 165 -1514 199 -1508
rect 165 -1576 199 -1552
rect 165 -1586 199 -1576
rect 165 -1644 199 -1624
rect 165 -1658 199 -1644
rect 405 -1134 439 -1120
rect 405 -1154 439 -1134
rect 405 -1202 439 -1192
rect 405 -1226 439 -1202
rect 405 -1270 439 -1264
rect 405 -1298 439 -1270
rect 405 -1338 439 -1336
rect 405 -1370 439 -1338
rect 405 -1440 439 -1408
rect 405 -1442 439 -1440
rect 405 -1508 439 -1480
rect 405 -1514 439 -1508
rect 405 -1576 439 -1552
rect 405 -1586 439 -1576
rect 405 -1644 439 -1624
rect 405 -1658 439 -1644
rect 1273 -1134 1307 -1120
rect 1273 -1154 1307 -1134
rect 1273 -1202 1307 -1192
rect 1273 -1226 1307 -1202
rect 1273 -1270 1307 -1264
rect 1273 -1298 1307 -1270
rect 1273 -1338 1307 -1336
rect 1273 -1370 1307 -1338
rect 1273 -1440 1307 -1408
rect 1273 -1442 1307 -1440
rect 1273 -1508 1307 -1480
rect 1273 -1514 1307 -1508
rect 1273 -1576 1307 -1552
rect 1273 -1586 1307 -1576
rect 1273 -1644 1307 -1624
rect 1273 -1658 1307 -1644
rect 1573 -1134 1607 -1120
rect 1573 -1154 1607 -1134
rect 1573 -1202 1607 -1192
rect 1573 -1226 1607 -1202
rect 1573 -1270 1607 -1264
rect 1573 -1298 1607 -1270
rect 1573 -1338 1607 -1336
rect 1573 -1370 1607 -1338
rect 1573 -1440 1607 -1408
rect 1573 -1442 1607 -1440
rect 1573 -1508 1607 -1480
rect 1573 -1514 1607 -1508
rect 1573 -1576 1607 -1552
rect 1573 -1586 1607 -1576
rect 1573 -1644 1607 -1624
rect 1573 -1658 1607 -1644
rect 1813 -1134 1847 -1120
rect 1813 -1154 1847 -1134
rect 1813 -1202 1847 -1192
rect 1813 -1226 1847 -1202
rect 1813 -1270 1847 -1264
rect 1813 -1298 1847 -1270
rect 1813 -1338 1847 -1336
rect 1813 -1370 1847 -1338
rect 1813 -1440 1847 -1408
rect 1813 -1442 1847 -1440
rect 1813 -1508 1847 -1480
rect 1813 -1514 1847 -1508
rect 1813 -1576 1847 -1552
rect 1813 -1586 1847 -1576
rect 1813 -1644 1847 -1624
rect 1813 -1658 1847 -1644
rect 2485 -1134 2519 -1120
rect 2485 -1154 2519 -1134
rect 2485 -1202 2519 -1192
rect 2485 -1226 2519 -1202
rect 2485 -1270 2519 -1264
rect 2485 -1298 2519 -1270
rect 2485 -1338 2519 -1336
rect 2485 -1370 2519 -1338
rect 2485 -1440 2519 -1408
rect 2485 -1442 2519 -1440
rect 2485 -1508 2519 -1480
rect 2485 -1514 2519 -1508
rect 2485 -1576 2519 -1552
rect 2485 -1586 2519 -1576
rect 2485 -1644 2519 -1624
rect 2485 -1658 2519 -1644
rect 3175 -1134 3209 -1120
rect 3175 -1154 3209 -1134
rect 3175 -1202 3209 -1192
rect 3175 -1226 3209 -1202
rect 3175 -1270 3209 -1264
rect 3175 -1298 3209 -1270
rect 3175 -1338 3209 -1336
rect 3175 -1370 3209 -1338
rect 3175 -1440 3209 -1408
rect 3175 -1442 3209 -1440
rect 3175 -1508 3209 -1480
rect 3175 -1514 3209 -1508
rect 3175 -1576 3209 -1552
rect 3175 -1586 3209 -1576
rect 3175 -1644 3209 -1624
rect 3175 -1658 3209 -1644
rect 253 -1772 287 -1738
rect -330 -1890 -296 -1856
rect -258 -1890 -224 -1856
rect -186 -1890 -152 -1856
rect -114 -1890 -80 -1856
rect -42 -1890 -8 -1856
rect 30 -1890 64 -1856
rect 102 -1890 136 -1856
rect 174 -1890 208 -1856
rect 246 -1890 280 -1856
rect 318 -1890 352 -1856
rect 390 -1890 424 -1856
rect 462 -1890 496 -1856
rect 534 -1890 568 -1856
rect 606 -1890 640 -1856
rect 1228 -1890 1262 -1856
rect 1300 -1890 1334 -1856
rect 1372 -1890 1406 -1856
rect 1444 -1890 1478 -1856
rect 1516 -1890 1550 -1856
rect 1588 -1890 1622 -1856
rect 1660 -1890 1694 -1856
rect 1732 -1890 1766 -1856
rect 1804 -1890 1838 -1856
rect 1876 -1890 1910 -1856
rect 1948 -1890 1982 -1856
rect 2020 -1890 2054 -1856
rect 2440 -1890 2474 -1856
rect 2512 -1890 2546 -1856
rect 2584 -1890 2618 -1856
rect 2656 -1890 2690 -1856
rect 2728 -1890 2762 -1856
rect 2800 -1890 2834 -1856
rect 2872 -1890 2906 -1856
rect 2944 -1890 2978 -1856
rect 3016 -1890 3050 -1856
rect 3088 -1890 3122 -1856
rect 3160 -1890 3194 -1856
rect 3232 -1890 3266 -1856
rect 3304 -1890 3338 -1856
rect 3376 -1890 3410 -1856
<< metal1 >>
rect -1487 333 -1407 1333
rect -1487 299 -1464 333
rect -1430 299 -1407 333
rect -1487 261 -1407 299
rect -1487 227 -1464 261
rect -1430 227 -1407 261
rect -1487 189 -1407 227
rect -1487 155 -1464 189
rect -1430 155 -1407 189
rect -1487 -1924 -1407 155
rect -1373 -92 -1293 1333
rect -1373 -126 -1350 -92
rect -1316 -126 -1293 -92
rect -1373 -164 -1293 -126
rect -1373 -198 -1350 -164
rect -1316 -198 -1293 -164
rect -1373 -236 -1293 -198
rect -1373 -270 -1350 -236
rect -1316 -270 -1293 -236
rect -1373 -920 -1293 -270
rect -1373 -954 -1350 -920
rect -1316 -954 -1293 -920
rect -1373 -992 -1293 -954
rect -1373 -1026 -1350 -992
rect -1316 -1026 -1293 -992
rect -1373 -1064 -1293 -1026
rect -1373 -1098 -1350 -1064
rect -1316 -1098 -1293 -1064
rect -1373 -1924 -1293 -1098
rect -1259 -372 -1179 1333
rect -1259 -406 -1236 -372
rect -1202 -406 -1179 -372
rect -1259 -444 -1179 -406
rect -1259 -478 -1236 -444
rect -1202 -478 -1179 -444
rect -1259 -516 -1179 -478
rect -1259 -550 -1236 -516
rect -1202 -550 -1179 -516
rect -1259 -1924 -1179 -550
rect -1145 -407 -1065 1333
rect -1145 -459 -1131 -407
rect -1079 -459 -1065 -407
rect -1145 -475 -1065 -459
rect -1145 -527 -1131 -475
rect -1079 -527 -1065 -475
rect -1145 -543 -1065 -527
rect -1145 -595 -1131 -543
rect -1079 -595 -1065 -543
rect -1145 -1924 -1065 -595
rect -1031 1258 -951 1333
rect -1031 1224 -1008 1258
rect -974 1224 -951 1258
rect -1031 1186 -951 1224
rect -1031 1152 -1008 1186
rect -974 1152 -951 1186
rect -1031 1114 -951 1152
rect -1031 1080 -1008 1114
rect -974 1080 -951 1114
rect -1031 -1923 -951 1080
rect -917 524 -837 1333
rect -917 490 -894 524
rect -860 490 -837 524
rect -917 452 -837 490
rect -917 418 -894 452
rect -860 418 -837 452
rect -917 380 -837 418
rect -917 346 -894 380
rect -860 346 -837 380
rect -917 -563 -837 346
rect -917 -615 -903 -563
rect -851 -615 -837 -563
rect -917 -631 -837 -615
rect -917 -683 -903 -631
rect -851 -683 -837 -631
rect -917 -699 -837 -683
rect -917 -751 -903 -699
rect -851 -751 -837 -699
rect -917 -1924 -837 -751
rect -803 1259 -723 1333
rect -803 1207 -789 1259
rect -737 1207 -723 1259
rect -803 1191 -723 1207
rect -803 1139 -789 1191
rect -737 1139 -723 1191
rect -803 1123 -723 1139
rect -803 1071 -789 1123
rect -737 1071 -723 1123
rect -803 -926 -723 1071
rect -803 -978 -789 -926
rect -737 -978 -723 -926
rect -803 -994 -723 -978
rect -803 -1046 -789 -994
rect -737 -1046 -723 -994
rect -803 -1062 -723 -1046
rect -803 -1114 -789 -1062
rect -737 -1114 -723 -1062
rect -803 -1923 -723 -1114
rect -689 -87 -609 1333
rect -689 -139 -675 -87
rect -623 -139 -609 -87
rect -689 -155 -609 -139
rect -689 -207 -675 -155
rect -623 -207 -609 -155
rect -689 -223 -609 -207
rect -689 -275 -675 -223
rect -623 -275 -609 -223
rect -689 -1665 -609 -275
rect -689 -1717 -675 -1665
rect -623 -1717 -609 -1665
rect -689 -1733 -609 -1717
rect -689 -1785 -675 -1733
rect -623 -1785 -609 -1733
rect -689 -1801 -609 -1785
rect -689 -1853 -675 -1801
rect -623 -1853 -609 -1801
rect -689 -1923 -609 -1853
rect -575 -206 -495 1333
rect -575 -240 -552 -206
rect -518 -240 -495 -206
rect -575 -278 -495 -240
rect -575 -312 -552 -278
rect -518 -312 -495 -278
rect -575 -350 -495 -312
rect -575 -384 -552 -350
rect -518 -384 -495 -350
rect -575 -1923 -495 -384
rect -461 1300 3297 1333
rect -461 1266 -330 1300
rect -296 1266 -258 1300
rect -224 1266 -186 1300
rect -152 1266 -114 1300
rect -80 1266 -42 1300
rect -8 1266 30 1300
rect 64 1266 102 1300
rect 136 1266 174 1300
rect 208 1266 246 1300
rect 280 1266 318 1300
rect 352 1266 390 1300
rect 424 1266 462 1300
rect 496 1266 534 1300
rect 568 1266 606 1300
rect 640 1266 678 1300
rect 712 1266 750 1300
rect 784 1266 822 1300
rect 856 1266 1228 1300
rect 1262 1266 1300 1300
rect 1334 1266 1372 1300
rect 1406 1266 1444 1300
rect 1478 1266 1516 1300
rect 1550 1266 1588 1300
rect 1622 1266 1660 1300
rect 1694 1266 1732 1300
rect 1766 1266 1804 1300
rect 1838 1266 1876 1300
rect 1910 1266 1948 1300
rect 1982 1266 2020 1300
rect 2054 1266 2440 1300
rect 2474 1266 2512 1300
rect 2546 1266 2584 1300
rect 2618 1266 2656 1300
rect 2690 1266 2728 1300
rect 2762 1266 2800 1300
rect 2834 1266 2872 1300
rect 2906 1266 2944 1300
rect 2978 1266 3016 1300
rect 3050 1266 3088 1300
rect 3122 1266 3160 1300
rect 3194 1266 3232 1300
rect 3266 1266 3297 1300
rect -461 1233 3297 1266
rect -461 -1823 -381 1233
rect -233 1079 -193 1233
rect 367 1079 407 1233
rect 618 1079 658 1233
rect 1325 1079 1365 1233
rect 1660 1191 1740 1205
rect 1660 1139 1674 1191
rect 1726 1139 1740 1191
rect 1660 1125 1740 1139
rect 1925 1079 1965 1233
rect 2482 1079 2522 1233
rect 2783 1079 2823 1233
rect 3022 1079 3062 1233
rect -253 1068 -173 1079
rect -253 1034 -230 1068
rect -196 1034 -173 1068
rect -253 996 -173 1034
rect -253 962 -230 996
rect -196 962 -173 996
rect -253 924 -173 962
rect -253 890 -230 924
rect -196 890 -173 924
rect -253 852 -173 890
rect -253 818 -230 852
rect -196 818 -173 852
rect -253 780 -173 818
rect -253 746 -230 780
rect -196 746 -173 780
rect -253 708 -173 746
rect -253 674 -230 708
rect -196 674 -173 708
rect -253 636 -173 674
rect -253 602 -230 636
rect -196 602 -173 636
rect -253 564 -173 602
rect -253 530 -230 564
rect -196 530 -173 564
rect -253 519 -173 530
rect 47 1077 127 1079
rect 47 1025 61 1077
rect 113 1025 127 1077
rect 47 1005 127 1025
rect 47 953 61 1005
rect 113 953 127 1005
rect 47 933 127 953
rect 47 881 61 933
rect 113 881 127 933
rect 47 861 127 881
rect 47 809 61 861
rect 113 809 127 861
rect 47 789 127 809
rect 47 737 61 789
rect 113 737 127 789
rect 47 717 127 737
rect 47 665 61 717
rect 113 665 127 717
rect 47 645 127 665
rect 47 593 61 645
rect 113 593 127 645
rect 47 573 127 593
rect 47 521 61 573
rect 113 521 127 573
rect 47 519 127 521
rect 347 1068 427 1079
rect 347 1034 370 1068
rect 404 1034 427 1068
rect 347 996 427 1034
rect 347 962 370 996
rect 404 962 427 996
rect 347 924 427 962
rect 347 890 370 924
rect 404 890 427 924
rect 347 852 427 890
rect 347 818 370 852
rect 404 818 427 852
rect 347 780 427 818
rect 347 746 370 780
rect 404 746 427 780
rect 347 708 427 746
rect 347 674 370 708
rect 404 674 427 708
rect 347 636 427 674
rect 347 602 370 636
rect 404 602 427 636
rect 347 564 427 602
rect 347 530 370 564
rect 404 530 427 564
rect 347 519 427 530
rect 598 1068 678 1079
rect 598 1034 621 1068
rect 655 1034 678 1068
rect 598 996 678 1034
rect 598 962 621 996
rect 655 962 678 996
rect 598 924 678 962
rect 598 890 621 924
rect 655 890 678 924
rect 598 852 678 890
rect 598 818 621 852
rect 655 818 678 852
rect 598 780 678 818
rect 598 746 621 780
rect 655 746 678 780
rect 598 708 678 746
rect 598 674 621 708
rect 655 674 678 708
rect 598 636 678 674
rect 598 602 621 636
rect 655 602 678 636
rect 598 564 678 602
rect 598 530 621 564
rect 655 530 678 564
rect 598 519 678 530
rect 1305 1068 1385 1079
rect 1305 1034 1328 1068
rect 1362 1034 1385 1068
rect 1305 996 1385 1034
rect 1305 962 1328 996
rect 1362 962 1385 996
rect 1305 924 1385 962
rect 1305 890 1328 924
rect 1362 890 1385 924
rect 1305 852 1385 890
rect 1305 818 1328 852
rect 1362 818 1385 852
rect 1305 780 1385 818
rect 1305 746 1328 780
rect 1362 746 1385 780
rect 1305 708 1385 746
rect 1305 674 1328 708
rect 1362 674 1385 708
rect 1305 636 1385 674
rect 1305 602 1328 636
rect 1362 602 1385 636
rect 1305 564 1385 602
rect 1305 530 1328 564
rect 1362 530 1385 564
rect 1305 519 1385 530
rect 1605 1077 1685 1079
rect 1605 1025 1619 1077
rect 1671 1025 1685 1077
rect 1605 1005 1685 1025
rect 1605 953 1619 1005
rect 1671 953 1685 1005
rect 1605 933 1685 953
rect 1605 881 1619 933
rect 1671 881 1685 933
rect 1605 861 1685 881
rect 1605 809 1619 861
rect 1671 809 1685 861
rect 1605 789 1685 809
rect 1605 737 1619 789
rect 1671 737 1685 789
rect 1605 717 1685 737
rect 1605 665 1619 717
rect 1671 665 1685 717
rect 1605 645 1685 665
rect 1605 593 1619 645
rect 1671 593 1685 645
rect 1605 573 1685 593
rect 1605 521 1619 573
rect 1671 521 1685 573
rect 1605 519 1685 521
rect 1905 1068 1985 1079
rect 1905 1034 1928 1068
rect 1962 1034 1985 1068
rect 1905 996 1985 1034
rect 1905 962 1928 996
rect 1962 962 1985 996
rect 1905 924 1985 962
rect 1905 890 1928 924
rect 1962 890 1985 924
rect 1905 852 1985 890
rect 1905 818 1928 852
rect 1962 818 1985 852
rect 1905 780 1985 818
rect 1905 746 1928 780
rect 1962 746 1985 780
rect 1905 708 1985 746
rect 1905 674 1928 708
rect 1962 674 1985 708
rect 1905 636 1985 674
rect 1905 602 1928 636
rect 1962 602 1985 636
rect 1905 564 1985 602
rect 1905 530 1928 564
rect 1962 530 1985 564
rect 1905 519 1985 530
rect 2462 1068 2542 1079
rect 2462 1034 2485 1068
rect 2519 1034 2542 1068
rect 2462 996 2542 1034
rect 2462 962 2485 996
rect 2519 962 2542 996
rect 2462 924 2542 962
rect 2462 890 2485 924
rect 2519 890 2542 924
rect 2462 852 2542 890
rect 2462 818 2485 852
rect 2519 818 2542 852
rect 2462 780 2542 818
rect 2462 746 2485 780
rect 2519 746 2542 780
rect 2462 708 2542 746
rect 2462 674 2485 708
rect 2519 674 2542 708
rect 2462 636 2542 674
rect 2462 602 2485 636
rect 2519 602 2542 636
rect 2462 564 2542 602
rect 2462 530 2485 564
rect 2519 530 2542 564
rect 2462 519 2542 530
rect 2762 1068 2842 1079
rect 2762 1034 2785 1068
rect 2819 1034 2842 1068
rect 2762 996 2842 1034
rect 2762 962 2785 996
rect 2819 962 2842 996
rect 2762 924 2842 962
rect 2762 890 2785 924
rect 2819 890 2842 924
rect 2762 852 2842 890
rect 2762 818 2785 852
rect 2819 818 2842 852
rect 2762 780 2842 818
rect 2762 746 2785 780
rect 2819 746 2842 780
rect 2762 708 2842 746
rect 2762 674 2785 708
rect 2819 674 2842 708
rect 2762 636 2842 674
rect 2762 602 2785 636
rect 2819 602 2842 636
rect 2762 564 2842 602
rect 2762 530 2785 564
rect 2819 530 2842 564
rect 2762 519 2842 530
rect 3002 1068 3082 1079
rect 3002 1034 3025 1068
rect 3059 1034 3082 1068
rect 3002 996 3082 1034
rect 3002 962 3025 996
rect 3059 962 3082 996
rect 3002 924 3082 962
rect 3002 890 3025 924
rect 3059 890 3082 924
rect 3002 852 3082 890
rect 3002 818 3025 852
rect 3059 818 3082 852
rect 3002 780 3082 818
rect 3002 746 3025 780
rect 3059 746 3082 780
rect 3002 708 3082 746
rect 3002 674 3025 708
rect 3059 674 3082 708
rect 3002 636 3082 674
rect 3002 602 3025 636
rect 3059 602 3082 636
rect 3002 564 3082 602
rect 3002 530 3025 564
rect 3059 530 3082 564
rect 3002 519 3082 530
rect 327 452 407 475
rect 327 418 350 452
rect 384 418 407 452
rect 327 395 407 418
rect 1325 461 1405 475
rect 1325 409 1339 461
rect 1391 409 1405 461
rect 1325 395 1405 409
rect 1885 452 1965 475
rect 1885 418 1908 452
rect 1942 418 1965 452
rect 1885 395 1965 418
rect 2482 455 2562 469
rect 2482 403 2496 455
rect 2548 403 2562 455
rect -53 264 27 284
rect 347 264 386 395
rect 476 349 556 363
rect 476 297 490 349
rect 542 297 556 349
rect 476 283 556 297
rect -53 261 386 264
rect -53 227 -30 261
rect 4 227 386 261
rect -53 224 386 227
rect 1355 270 1435 284
rect -53 204 27 224
rect 1355 218 1369 270
rect 1421 218 1435 270
rect 1355 204 1435 218
rect 1505 264 1585 284
rect 1905 264 1944 395
rect 2482 389 2562 403
rect 3239 417 3319 431
rect 2056 369 2136 383
rect 2056 317 2070 369
rect 2122 317 2136 369
rect 2056 303 2136 317
rect 3239 365 3253 417
rect 3305 365 3319 417
rect 3239 345 3319 365
rect 3239 293 3253 345
rect 3305 293 3319 345
rect 3239 279 3319 293
rect 1505 261 1944 264
rect 1505 227 1528 261
rect 1562 227 1944 261
rect 1505 224 1944 227
rect 1505 204 1585 224
rect -253 128 -173 169
rect -253 94 -230 128
rect -196 94 -173 128
rect -253 56 -173 94
rect -253 22 -230 56
rect -196 22 -173 56
rect -253 -16 -173 22
rect -253 -50 -230 -16
rect -196 -50 -173 -16
rect -253 -91 -173 -50
rect 47 137 127 169
rect 47 85 61 137
rect 113 85 127 137
rect 47 65 127 85
rect 47 13 61 65
rect 113 13 127 65
rect 47 -7 127 13
rect 47 -59 61 -7
rect 113 -59 127 -7
rect 47 -91 127 -59
rect 347 128 427 169
rect 347 94 370 128
rect 404 94 427 128
rect 347 56 427 94
rect 347 22 370 56
rect 404 22 427 56
rect 347 -16 427 22
rect 347 -50 370 -16
rect 404 -50 427 -16
rect 347 -91 427 -50
rect 598 128 678 169
rect 598 94 621 128
rect 655 94 678 128
rect 598 56 678 94
rect 598 22 621 56
rect 655 22 678 56
rect 598 -16 678 22
rect 598 -50 621 -16
rect 655 -50 678 -16
rect 598 -91 678 -50
rect 1305 128 1385 169
rect 1305 94 1328 128
rect 1362 94 1385 128
rect 1305 56 1385 94
rect 1305 22 1328 56
rect 1362 22 1385 56
rect 1305 -16 1385 22
rect 1305 -50 1328 -16
rect 1362 -50 1385 -16
rect 1305 -91 1385 -50
rect 1605 137 1685 169
rect 1605 85 1619 137
rect 1671 85 1685 137
rect 1605 65 1685 85
rect 1605 13 1619 65
rect 1671 13 1685 65
rect 1605 -7 1685 13
rect 1605 -59 1619 -7
rect 1671 -59 1685 -7
rect 1605 -91 1685 -59
rect 1905 128 1985 169
rect 1905 94 1928 128
rect 1962 94 1985 128
rect 1905 56 1985 94
rect 1905 22 1928 56
rect 1962 22 1985 56
rect 1905 -16 1985 22
rect 1905 -50 1928 -16
rect 1962 -50 1985 -16
rect 1905 -91 1985 -50
rect 2462 128 2542 169
rect 2462 94 2485 128
rect 2519 94 2542 128
rect 2462 56 2542 94
rect 2462 22 2485 56
rect 2519 22 2542 56
rect 2462 -16 2542 22
rect 2462 -50 2485 -16
rect 2519 -50 2542 -16
rect 2462 -91 2542 -50
rect 3002 128 3082 169
rect 3002 94 3025 128
rect 3059 94 3082 128
rect 3002 56 3082 94
rect 3002 22 3025 56
rect 3059 22 3082 56
rect 3002 -16 3082 22
rect 3002 -50 3025 -16
rect 3059 -50 3082 -16
rect 3002 -91 3082 -50
rect -233 -245 -193 -91
rect 367 -245 407 -91
rect 618 -245 658 -91
rect 1325 -245 1365 -91
rect 1660 -151 1740 -137
rect 1660 -203 1674 -151
rect 1726 -203 1740 -151
rect 1660 -217 1740 -203
rect 1925 -245 1965 -91
rect 2482 -245 2522 -91
rect 3022 -245 3062 -91
rect -353 -278 3438 -245
rect -353 -312 -330 -278
rect -296 -312 -258 -278
rect -224 -312 -186 -278
rect -152 -312 -114 -278
rect -80 -312 -42 -278
rect -8 -312 30 -278
rect 64 -312 102 -278
rect 136 -312 174 -278
rect 208 -312 246 -278
rect 280 -312 318 -278
rect 352 -312 390 -278
rect 424 -312 462 -278
rect 496 -312 534 -278
rect 568 -312 606 -278
rect 640 -312 678 -278
rect 712 -312 750 -278
rect 784 -312 822 -278
rect 856 -312 1228 -278
rect 1262 -312 1300 -278
rect 1334 -312 1372 -278
rect 1406 -312 1444 -278
rect 1478 -312 1516 -278
rect 1550 -312 1588 -278
rect 1622 -312 1660 -278
rect 1694 -312 1732 -278
rect 1766 -312 1804 -278
rect 1838 -312 1876 -278
rect 1910 -312 1948 -278
rect 1982 -312 2020 -278
rect 2054 -312 2440 -278
rect 2474 -312 2512 -278
rect 2546 -312 2584 -278
rect 2618 -312 2656 -278
rect 2690 -312 2728 -278
rect 2762 -312 2800 -278
rect 2834 -312 2872 -278
rect 2906 -312 2944 -278
rect 2978 -312 3016 -278
rect 3050 -312 3088 -278
rect 3122 -312 3160 -278
rect 3194 -312 3232 -278
rect 3266 -312 3304 -278
rect 3338 -312 3376 -278
rect 3410 -312 3438 -278
rect -353 -345 3438 -312
rect -288 -499 -248 -345
rect 402 -499 442 -345
rect 556 -387 636 -373
rect 556 -439 570 -387
rect 622 -439 636 -387
rect 556 -453 636 -439
rect 1270 -499 1310 -345
rect 1810 -499 1850 -345
rect 2632 -499 2672 -345
rect 2932 -499 2972 -345
rect 3171 -499 3211 -345
rect 3239 -387 3319 -373
rect 3239 -439 3253 -387
rect 3305 -439 3319 -387
rect 3239 -453 3319 -439
rect -308 -540 -228 -499
rect -308 -574 -285 -540
rect -251 -574 -228 -540
rect -308 -612 -228 -574
rect -308 -646 -285 -612
rect -251 -646 -228 -612
rect -308 -684 -228 -646
rect -308 -718 -285 -684
rect -251 -718 -228 -684
rect -308 -759 -228 -718
rect 382 -540 462 -499
rect 382 -574 405 -540
rect 439 -574 462 -540
rect 382 -612 462 -574
rect 382 -646 405 -612
rect 439 -646 462 -612
rect 382 -684 462 -646
rect 382 -718 405 -684
rect 439 -718 462 -684
rect 382 -759 462 -718
rect 1250 -540 1330 -499
rect 1250 -574 1273 -540
rect 1307 -574 1330 -540
rect 1250 -612 1330 -574
rect 1250 -646 1273 -612
rect 1307 -646 1330 -612
rect 1250 -684 1330 -646
rect 1250 -718 1273 -684
rect 1307 -718 1330 -684
rect 1250 -759 1330 -718
rect 1790 -540 1870 -499
rect 1790 -574 1813 -540
rect 1847 -574 1870 -540
rect 1790 -612 1870 -574
rect 1790 -646 1813 -612
rect 1847 -646 1870 -612
rect 1790 -684 1870 -646
rect 1790 -718 1813 -684
rect 1847 -718 1870 -684
rect 1790 -759 1870 -718
rect 2612 -540 2692 -499
rect 2612 -574 2635 -540
rect 2669 -574 2692 -540
rect 2612 -612 2692 -574
rect 2612 -646 2635 -612
rect 2669 -646 2692 -612
rect 2612 -684 2692 -646
rect 2612 -718 2635 -684
rect 2669 -718 2692 -684
rect 2612 -759 2692 -718
rect 2912 -540 2992 -499
rect 2912 -574 2935 -540
rect 2969 -574 2992 -540
rect 2912 -612 2992 -574
rect 2912 -646 2935 -612
rect 2969 -646 2992 -612
rect 2912 -684 2992 -646
rect 2912 -718 2935 -684
rect 2969 -718 2992 -684
rect 2912 -759 2992 -718
rect 3152 -540 3232 -499
rect 3152 -574 3175 -540
rect 3209 -574 3232 -540
rect 3152 -612 3232 -574
rect 3152 -646 3175 -612
rect 3209 -646 3232 -612
rect 3152 -684 3232 -646
rect 3152 -718 3175 -684
rect 3209 -718 3232 -684
rect 3152 -759 3232 -718
rect 3303 -874 3383 -860
rect 3303 -926 3317 -874
rect 3369 -926 3383 -874
rect 3303 -946 3383 -926
rect 1270 -993 1350 -979
rect 1270 -1045 1284 -993
rect 1336 -1045 1350 -993
rect 3303 -998 3317 -946
rect 3369 -998 3383 -946
rect 3303 -1012 3383 -998
rect 1270 -1059 1350 -1045
rect -158 -1120 -78 -1109
rect -158 -1154 -135 -1120
rect -101 -1154 -78 -1120
rect -158 -1192 -78 -1154
rect -158 -1226 -135 -1192
rect -101 -1226 -78 -1192
rect -158 -1264 -78 -1226
rect -158 -1298 -135 -1264
rect -101 -1298 -78 -1264
rect -158 -1336 -78 -1298
rect -158 -1370 -135 -1336
rect -101 -1370 -78 -1336
rect -158 -1408 -78 -1370
rect -158 -1442 -135 -1408
rect -101 -1442 -78 -1408
rect -158 -1480 -78 -1442
rect -158 -1514 -135 -1480
rect -101 -1514 -78 -1480
rect -158 -1552 -78 -1514
rect -158 -1586 -135 -1552
rect -101 -1586 -78 -1552
rect -158 -1624 -78 -1586
rect -158 -1658 -135 -1624
rect -101 -1658 -78 -1624
rect -158 -1669 -78 -1658
rect 142 -1120 222 -1109
rect 142 -1154 165 -1120
rect 199 -1154 222 -1120
rect 142 -1192 222 -1154
rect 142 -1226 165 -1192
rect 199 -1226 222 -1192
rect 142 -1264 222 -1226
rect 142 -1298 165 -1264
rect 199 -1298 222 -1264
rect 142 -1336 222 -1298
rect 142 -1370 165 -1336
rect 199 -1370 222 -1336
rect 142 -1408 222 -1370
rect 142 -1442 165 -1408
rect 199 -1442 222 -1408
rect 142 -1480 222 -1442
rect 142 -1514 165 -1480
rect 199 -1514 222 -1480
rect 142 -1552 222 -1514
rect 142 -1586 165 -1552
rect 199 -1586 222 -1552
rect 142 -1624 222 -1586
rect 142 -1658 165 -1624
rect 199 -1658 222 -1624
rect 142 -1669 222 -1658
rect 382 -1120 462 -1109
rect 382 -1154 405 -1120
rect 439 -1154 462 -1120
rect 382 -1192 462 -1154
rect 382 -1226 405 -1192
rect 439 -1226 462 -1192
rect 382 -1264 462 -1226
rect 382 -1298 405 -1264
rect 439 -1298 462 -1264
rect 382 -1336 462 -1298
rect 382 -1370 405 -1336
rect 439 -1370 462 -1336
rect 382 -1408 462 -1370
rect 382 -1442 405 -1408
rect 439 -1442 462 -1408
rect 382 -1480 462 -1442
rect 382 -1514 405 -1480
rect 439 -1514 462 -1480
rect 382 -1552 462 -1514
rect 382 -1586 405 -1552
rect 439 -1586 462 -1552
rect 382 -1624 462 -1586
rect 382 -1658 405 -1624
rect 439 -1658 462 -1624
rect 382 -1669 462 -1658
rect 1250 -1120 1330 -1109
rect 1250 -1154 1273 -1120
rect 1307 -1154 1330 -1120
rect 1250 -1192 1330 -1154
rect 1250 -1226 1273 -1192
rect 1307 -1226 1330 -1192
rect 1250 -1264 1330 -1226
rect 1250 -1298 1273 -1264
rect 1307 -1298 1330 -1264
rect 1250 -1336 1330 -1298
rect 1250 -1370 1273 -1336
rect 1307 -1370 1330 -1336
rect 1250 -1408 1330 -1370
rect 1250 -1442 1273 -1408
rect 1307 -1442 1330 -1408
rect 1250 -1480 1330 -1442
rect 1250 -1514 1273 -1480
rect 1307 -1514 1330 -1480
rect 1250 -1552 1330 -1514
rect 1250 -1586 1273 -1552
rect 1307 -1586 1330 -1552
rect 1250 -1624 1330 -1586
rect 1250 -1658 1273 -1624
rect 1307 -1658 1330 -1624
rect 1250 -1669 1330 -1658
rect 1550 -1120 1630 -1109
rect 1550 -1154 1573 -1120
rect 1607 -1154 1630 -1120
rect 1550 -1192 1630 -1154
rect 1550 -1226 1573 -1192
rect 1607 -1226 1630 -1192
rect 1550 -1264 1630 -1226
rect 1550 -1298 1573 -1264
rect 1607 -1298 1630 -1264
rect 1550 -1336 1630 -1298
rect 1550 -1370 1573 -1336
rect 1607 -1370 1630 -1336
rect 1550 -1408 1630 -1370
rect 1550 -1442 1573 -1408
rect 1607 -1442 1630 -1408
rect 1550 -1480 1630 -1442
rect 1550 -1514 1573 -1480
rect 1607 -1514 1630 -1480
rect 1550 -1552 1630 -1514
rect 1550 -1586 1573 -1552
rect 1607 -1586 1630 -1552
rect 1550 -1624 1630 -1586
rect 1550 -1658 1573 -1624
rect 1607 -1658 1630 -1624
rect 1550 -1669 1630 -1658
rect 1790 -1120 1870 -1109
rect 1790 -1154 1813 -1120
rect 1847 -1154 1870 -1120
rect 1790 -1192 1870 -1154
rect 1790 -1226 1813 -1192
rect 1847 -1226 1870 -1192
rect 1790 -1264 1870 -1226
rect 1790 -1298 1813 -1264
rect 1847 -1298 1870 -1264
rect 1790 -1336 1870 -1298
rect 1790 -1370 1813 -1336
rect 1847 -1370 1870 -1336
rect 1790 -1408 1870 -1370
rect 1790 -1442 1813 -1408
rect 1847 -1442 1870 -1408
rect 1790 -1480 1870 -1442
rect 1790 -1514 1813 -1480
rect 1847 -1514 1870 -1480
rect 1790 -1552 1870 -1514
rect 1790 -1586 1813 -1552
rect 1847 -1586 1870 -1552
rect 1790 -1624 1870 -1586
rect 1790 -1658 1813 -1624
rect 1847 -1658 1870 -1624
rect 1790 -1669 1870 -1658
rect 2462 -1120 2542 -1109
rect 2462 -1154 2485 -1120
rect 2519 -1154 2542 -1120
rect 2462 -1192 2542 -1154
rect 2462 -1226 2485 -1192
rect 2519 -1226 2542 -1192
rect 2462 -1264 2542 -1226
rect 2462 -1298 2485 -1264
rect 2519 -1298 2542 -1264
rect 2462 -1336 2542 -1298
rect 2462 -1370 2485 -1336
rect 2519 -1370 2542 -1336
rect 2462 -1408 2542 -1370
rect 2462 -1442 2485 -1408
rect 2519 -1442 2542 -1408
rect 2462 -1480 2542 -1442
rect 2462 -1514 2485 -1480
rect 2519 -1514 2542 -1480
rect 2462 -1552 2542 -1514
rect 2462 -1586 2485 -1552
rect 2519 -1586 2542 -1552
rect 2462 -1624 2542 -1586
rect 2462 -1658 2485 -1624
rect 2519 -1658 2542 -1624
rect 2462 -1669 2542 -1658
rect 3152 -1120 3232 -1109
rect 3152 -1154 3175 -1120
rect 3209 -1154 3232 -1120
rect 3152 -1192 3232 -1154
rect 3152 -1226 3175 -1192
rect 3209 -1226 3232 -1192
rect 3152 -1264 3232 -1226
rect 3152 -1298 3175 -1264
rect 3209 -1298 3232 -1264
rect 3152 -1336 3232 -1298
rect 3152 -1370 3175 -1336
rect 3209 -1370 3232 -1336
rect 3152 -1408 3232 -1370
rect 3152 -1442 3175 -1408
rect 3209 -1442 3232 -1408
rect 3152 -1480 3232 -1442
rect 3152 -1514 3175 -1480
rect 3209 -1514 3232 -1480
rect 3152 -1552 3232 -1514
rect 3152 -1586 3175 -1552
rect 3209 -1586 3232 -1552
rect 3152 -1624 3232 -1586
rect 3152 -1658 3175 -1624
rect 3209 -1658 3232 -1624
rect 3152 -1669 3232 -1658
rect -138 -1823 -98 -1669
rect 162 -1823 202 -1669
rect 230 -1729 310 -1715
rect 230 -1781 244 -1729
rect 296 -1781 310 -1729
rect 230 -1795 310 -1781
rect 402 -1823 442 -1669
rect 1270 -1823 1310 -1669
rect 1571 -1823 1611 -1669
rect 1810 -1823 1850 -1669
rect 2482 -1823 2522 -1669
rect 3173 -1823 3213 -1669
rect -461 -1856 3427 -1823
rect -461 -1890 -330 -1856
rect -296 -1890 -258 -1856
rect -224 -1890 -186 -1856
rect -152 -1890 -114 -1856
rect -80 -1890 -42 -1856
rect -8 -1890 30 -1856
rect 64 -1890 102 -1856
rect 136 -1890 174 -1856
rect 208 -1890 246 -1856
rect 280 -1890 318 -1856
rect 352 -1890 390 -1856
rect 424 -1890 462 -1856
rect 496 -1890 534 -1856
rect 568 -1890 606 -1856
rect 640 -1890 1228 -1856
rect 1262 -1890 1300 -1856
rect 1334 -1890 1372 -1856
rect 1406 -1890 1444 -1856
rect 1478 -1890 1516 -1856
rect 1550 -1890 1588 -1856
rect 1622 -1890 1660 -1856
rect 1694 -1890 1732 -1856
rect 1766 -1890 1804 -1856
rect 1838 -1890 1876 -1856
rect 1910 -1890 1948 -1856
rect 1982 -1890 2020 -1856
rect 2054 -1890 2440 -1856
rect 2474 -1890 2512 -1856
rect 2546 -1890 2584 -1856
rect 2618 -1890 2656 -1856
rect 2690 -1890 2728 -1856
rect 2762 -1890 2800 -1856
rect 2834 -1890 2872 -1856
rect 2906 -1890 2944 -1856
rect 2978 -1890 3016 -1856
rect 3050 -1890 3088 -1856
rect 3122 -1890 3160 -1856
rect 3194 -1890 3232 -1856
rect 3266 -1890 3304 -1856
rect 3338 -1890 3376 -1856
rect 3410 -1890 3427 -1856
rect -461 -1923 3427 -1890
<< via1 >>
rect -1131 -459 -1079 -407
rect -1131 -527 -1079 -475
rect -1131 -595 -1079 -543
rect -903 -615 -851 -563
rect -903 -683 -851 -631
rect -903 -751 -851 -699
rect -789 1207 -737 1259
rect -789 1139 -737 1191
rect -789 1071 -737 1123
rect -789 -978 -737 -926
rect -789 -1046 -737 -994
rect -789 -1114 -737 -1062
rect -675 -139 -623 -87
rect -675 -207 -623 -155
rect -675 -275 -623 -223
rect -675 -1717 -623 -1665
rect -675 -1785 -623 -1733
rect -675 -1853 -623 -1801
rect 1674 1182 1726 1191
rect 1674 1148 1683 1182
rect 1683 1148 1717 1182
rect 1717 1148 1726 1182
rect 1674 1139 1726 1148
rect 61 1068 113 1077
rect 61 1034 70 1068
rect 70 1034 104 1068
rect 104 1034 113 1068
rect 61 1025 113 1034
rect 61 996 113 1005
rect 61 962 70 996
rect 70 962 104 996
rect 104 962 113 996
rect 61 953 113 962
rect 61 924 113 933
rect 61 890 70 924
rect 70 890 104 924
rect 104 890 113 924
rect 61 881 113 890
rect 61 852 113 861
rect 61 818 70 852
rect 70 818 104 852
rect 104 818 113 852
rect 61 809 113 818
rect 61 780 113 789
rect 61 746 70 780
rect 70 746 104 780
rect 104 746 113 780
rect 61 737 113 746
rect 61 708 113 717
rect 61 674 70 708
rect 70 674 104 708
rect 104 674 113 708
rect 61 665 113 674
rect 61 636 113 645
rect 61 602 70 636
rect 70 602 104 636
rect 104 602 113 636
rect 61 593 113 602
rect 61 564 113 573
rect 61 530 70 564
rect 70 530 104 564
rect 104 530 113 564
rect 61 521 113 530
rect 1619 1068 1671 1077
rect 1619 1034 1628 1068
rect 1628 1034 1662 1068
rect 1662 1034 1671 1068
rect 1619 1025 1671 1034
rect 1619 996 1671 1005
rect 1619 962 1628 996
rect 1628 962 1662 996
rect 1662 962 1671 996
rect 1619 953 1671 962
rect 1619 924 1671 933
rect 1619 890 1628 924
rect 1628 890 1662 924
rect 1662 890 1671 924
rect 1619 881 1671 890
rect 1619 852 1671 861
rect 1619 818 1628 852
rect 1628 818 1662 852
rect 1662 818 1671 852
rect 1619 809 1671 818
rect 1619 780 1671 789
rect 1619 746 1628 780
rect 1628 746 1662 780
rect 1662 746 1671 780
rect 1619 737 1671 746
rect 1619 708 1671 717
rect 1619 674 1628 708
rect 1628 674 1662 708
rect 1662 674 1671 708
rect 1619 665 1671 674
rect 1619 636 1671 645
rect 1619 602 1628 636
rect 1628 602 1662 636
rect 1662 602 1671 636
rect 1619 593 1671 602
rect 1619 564 1671 573
rect 1619 530 1628 564
rect 1628 530 1662 564
rect 1662 530 1671 564
rect 1619 521 1671 530
rect 1339 452 1391 461
rect 1339 418 1348 452
rect 1348 418 1382 452
rect 1382 418 1391 452
rect 1339 409 1391 418
rect 2496 446 2548 455
rect 2496 412 2505 446
rect 2505 412 2539 446
rect 2539 412 2548 446
rect 2496 403 2548 412
rect 490 340 542 349
rect 490 306 499 340
rect 499 306 533 340
rect 533 306 542 340
rect 490 297 542 306
rect 1369 261 1421 270
rect 1369 227 1378 261
rect 1378 227 1412 261
rect 1412 227 1421 261
rect 1369 218 1421 227
rect 2070 360 2122 369
rect 2070 326 2079 360
rect 2079 326 2113 360
rect 2113 326 2122 360
rect 2070 317 2122 326
rect 3253 408 3305 417
rect 3253 374 3262 408
rect 3262 374 3296 408
rect 3296 374 3305 408
rect 3253 365 3305 374
rect 3253 336 3305 345
rect 3253 302 3262 336
rect 3262 302 3296 336
rect 3296 302 3305 336
rect 3253 293 3305 302
rect 61 128 113 137
rect 61 94 70 128
rect 70 94 104 128
rect 104 94 113 128
rect 61 85 113 94
rect 61 56 113 65
rect 61 22 70 56
rect 70 22 104 56
rect 104 22 113 56
rect 61 13 113 22
rect 61 -16 113 -7
rect 61 -50 70 -16
rect 70 -50 104 -16
rect 104 -50 113 -16
rect 61 -59 113 -50
rect 1619 128 1671 137
rect 1619 94 1628 128
rect 1628 94 1662 128
rect 1662 94 1671 128
rect 1619 85 1671 94
rect 1619 56 1671 65
rect 1619 22 1628 56
rect 1628 22 1662 56
rect 1662 22 1671 56
rect 1619 13 1671 22
rect 1619 -16 1671 -7
rect 1619 -50 1628 -16
rect 1628 -50 1662 -16
rect 1662 -50 1671 -16
rect 1619 -59 1671 -50
rect 1674 -160 1726 -151
rect 1674 -194 1683 -160
rect 1683 -194 1717 -160
rect 1717 -194 1726 -160
rect 1674 -203 1726 -194
rect 570 -396 622 -387
rect 570 -430 579 -396
rect 579 -430 613 -396
rect 613 -430 622 -396
rect 570 -439 622 -430
rect 3253 -396 3305 -387
rect 3253 -430 3262 -396
rect 3262 -430 3296 -396
rect 3296 -430 3305 -396
rect 3253 -439 3305 -430
rect 3317 -883 3369 -874
rect 3317 -917 3326 -883
rect 3326 -917 3360 -883
rect 3360 -917 3369 -883
rect 3317 -926 3369 -917
rect 1284 -1002 1336 -993
rect 1284 -1036 1293 -1002
rect 1293 -1036 1327 -1002
rect 1327 -1036 1336 -1002
rect 1284 -1045 1336 -1036
rect 3317 -955 3369 -946
rect 3317 -989 3326 -955
rect 3326 -989 3360 -955
rect 3360 -989 3369 -955
rect 3317 -998 3369 -989
rect 244 -1738 296 -1729
rect 244 -1772 253 -1738
rect 253 -1772 287 -1738
rect 287 -1772 296 -1738
rect 244 -1781 296 -1772
<< metal2 >>
rect -803 1259 -723 1273
rect -803 1207 -789 1259
rect -737 1207 -723 1259
rect -803 1191 -723 1207
rect -803 1139 -789 1191
rect -737 1185 -723 1191
rect 1660 1191 1740 1205
rect 1660 1185 1674 1191
rect -737 1145 1674 1185
rect -737 1139 -723 1145
rect -803 1123 -723 1139
rect 1660 1139 1674 1145
rect 1726 1139 1740 1191
rect 1660 1125 1740 1139
rect -803 1071 -789 1123
rect -737 1071 -723 1123
rect -803 1057 -723 1071
rect 47 1077 127 1079
rect 47 1025 61 1077
rect 113 1025 127 1077
rect 47 1005 127 1025
rect 47 953 61 1005
rect 113 953 127 1005
rect 47 933 127 953
rect 47 881 61 933
rect 113 881 127 933
rect 47 861 127 881
rect 47 809 61 861
rect 113 809 127 861
rect 47 789 127 809
rect 47 737 61 789
rect 113 737 127 789
rect 47 717 127 737
rect 47 665 61 717
rect 113 665 127 717
rect 47 645 127 665
rect 47 593 61 645
rect 113 593 127 645
rect 47 573 127 593
rect 47 521 61 573
rect 113 521 127 573
rect 47 519 127 521
rect 1605 1077 1685 1079
rect 1605 1025 1619 1077
rect 1671 1025 1685 1077
rect 1605 1005 1685 1025
rect 1605 953 1619 1005
rect 1671 953 1685 1005
rect 1605 933 1685 953
rect 1605 881 1619 933
rect 1671 881 1685 933
rect 1605 861 1685 881
rect 1605 809 1619 861
rect 1671 809 1685 861
rect 1605 789 1685 809
rect 1605 737 1619 789
rect 1671 737 1685 789
rect 1605 717 1685 737
rect 1605 665 1619 717
rect 1671 665 1685 717
rect 1605 645 1685 665
rect 1605 593 1619 645
rect 1671 593 1685 645
rect 1605 573 1685 593
rect 1605 521 1619 573
rect 1671 521 1685 573
rect 1605 519 1685 521
rect 67 363 107 519
rect 1325 461 1405 475
rect 1325 455 1339 461
rect 980 415 1339 455
rect 67 349 556 363
rect 67 323 490 349
rect 67 169 107 323
rect 476 297 490 323
rect 542 297 556 349
rect 476 283 556 297
rect 47 137 127 169
rect 47 85 61 137
rect 113 85 127 137
rect 47 65 127 85
rect 47 13 61 65
rect 113 13 127 65
rect 47 -7 127 13
rect 47 -59 61 -7
rect 113 -59 127 -7
rect -689 -87 -609 -73
rect -689 -139 -675 -87
rect -623 -139 -609 -87
rect 47 -91 127 -59
rect -689 -155 -609 -139
rect -689 -207 -675 -155
rect -623 -161 -609 -155
rect 980 -161 1020 415
rect 1325 409 1339 415
rect 1391 409 1405 461
rect 1325 395 1405 409
rect 1625 363 1665 519
rect 2482 455 2562 469
rect 2482 449 2496 455
rect 2164 409 2496 449
rect 2056 369 2136 383
rect 2056 363 2070 369
rect 1625 323 2070 363
rect 1355 270 1435 284
rect 1355 218 1369 270
rect 1421 218 1435 270
rect 1355 204 1435 218
rect -623 -201 1020 -161
rect -623 -207 -609 -201
rect -689 -223 -609 -207
rect -689 -275 -675 -223
rect -623 -275 -609 -223
rect -689 -289 -609 -275
rect 556 -387 636 -373
rect -1145 -407 -1065 -393
rect -1145 -459 -1131 -407
rect -1079 -459 -1065 -407
rect 556 -439 570 -387
rect 622 -393 636 -387
rect 1375 -393 1415 204
rect 1625 169 1665 323
rect 2056 317 2070 323
rect 2122 317 2136 369
rect 2056 303 2136 317
rect 1605 137 1685 169
rect 1605 85 1619 137
rect 1671 85 1685 137
rect 1605 65 1685 85
rect 1605 13 1619 65
rect 1671 13 1685 65
rect 1605 -7 1685 13
rect 1605 -59 1619 -7
rect 1671 -59 1685 -7
rect 1605 -91 1685 -59
rect 1660 -151 1740 -137
rect 1660 -203 1674 -151
rect 1726 -203 1740 -151
rect 1660 -217 1740 -203
rect 622 -433 1415 -393
rect 622 -439 636 -433
rect 556 -453 636 -439
rect -1145 -475 -1065 -459
rect -1145 -527 -1131 -475
rect -1079 -481 -1065 -475
rect 1680 -481 1720 -217
rect -1079 -521 1720 -481
rect -1079 -527 -1065 -521
rect -1145 -543 -1065 -527
rect -1145 -595 -1131 -543
rect -1079 -595 -1065 -543
rect 2164 -549 2204 409
rect 2482 403 2496 409
rect 2548 403 2562 455
rect 2482 389 2562 403
rect 3239 417 3319 431
rect 3239 365 3253 417
rect 3305 365 3319 417
rect 3239 345 3319 365
rect 3239 293 3253 345
rect 3305 293 3319 345
rect 3239 279 3319 293
rect 3259 -373 3299 279
rect 3239 -387 3319 -373
rect 3239 -439 3253 -387
rect 3305 -439 3319 -387
rect 3239 -453 3319 -439
rect -1145 -609 -1065 -595
rect -917 -563 2204 -549
rect -917 -615 -903 -563
rect -851 -589 2204 -563
rect -851 -615 -837 -589
rect -917 -631 -837 -615
rect -917 -683 -903 -631
rect -851 -683 -837 -631
rect -917 -699 -837 -683
rect -917 -751 -903 -699
rect -851 -751 -837 -699
rect -917 -765 -837 -751
rect 3303 -874 3383 -860
rect -803 -926 -723 -912
rect -803 -978 -789 -926
rect -737 -978 -723 -926
rect -803 -994 -723 -978
rect 3303 -926 3317 -874
rect 3369 -916 3383 -874
rect 3369 -926 3428 -916
rect 3303 -946 3428 -926
rect -803 -1046 -789 -994
rect -737 -1000 -723 -994
rect 1270 -993 1350 -979
rect 1270 -1000 1284 -993
rect -737 -1040 1284 -1000
rect -737 -1046 -723 -1040
rect -803 -1062 -723 -1046
rect 1270 -1045 1284 -1040
rect 1336 -1045 1350 -993
rect 3303 -998 3317 -946
rect 3369 -956 3428 -946
rect 3369 -998 3383 -956
rect 3303 -1012 3383 -998
rect 1270 -1059 1350 -1045
rect -803 -1114 -789 -1062
rect -737 -1114 -723 -1062
rect -803 -1128 -723 -1114
rect -689 -1665 -609 -1651
rect -689 -1717 -675 -1665
rect -623 -1717 -609 -1665
rect -689 -1733 -609 -1717
rect -689 -1785 -675 -1733
rect -623 -1739 -609 -1733
rect 230 -1729 310 -1715
rect 230 -1739 244 -1729
rect -623 -1779 244 -1739
rect -623 -1785 -609 -1779
rect -689 -1801 -609 -1785
rect 230 -1781 244 -1779
rect 296 -1781 310 -1729
rect 230 -1795 310 -1781
rect -689 -1853 -675 -1801
rect -623 -1853 -609 -1801
rect -689 -1867 -609 -1853
<< labels >>
flabel metal1 s -552 -312 -518 -278 2 FreeSans 2500 0 0 0 GND
port 1 nsew
flabel metal1 s -1477 1267 -1416 1327 2 FreeSans 3126 0 0 0 x0
port 2 nsew
flabel metal1 s -1364 1206 -1303 1266 2 FreeSans 3126 0 0 0 x0_bar
port 3 nsew
flabel metal1 s -1249 1267 -1188 1327 2 FreeSans 3126 0 0 0 x1
port 4 nsew
flabel metal1 s -1135 1206 -1074 1266 2 FreeSans 3126 0 0 0 x1_bar
port 5 nsew
flabel metal1 s -1021 1268 -960 1328 2 FreeSans 3126 0 0 0 x2
port 6 nsew
flabel metal1 s -908 1207 -847 1267 2 FreeSans 3126 0 0 0 x2_bar
port 7 nsew
flabel metal1 s -793 1268 -732 1328 2 FreeSans 3126 0 0 0 x3
port 8 nsew
flabel metal1 s -443 1267 -409 1301 2 FreeSans 2500 0 0 0 VDD
port 9 nsew
flabel metal1 s -678 1208 -617 1268 2 FreeSans 3126 0 0 0 x3_bar
port 10 nsew
flabel metal2 s 3326 -917 3360 -883 2 FreeSans 2500 0 0 0 s1
port 11 nsew
flabel locali 1963 -1036 1997 -1002 4 FreeSans 2000 0 0 0 CMOS_AND_1/AND
flabel locali 1473 -426 1507 -392 4 FreeSans 2000 0 0 0 CMOS_AND_1/A
flabel locali 1293 -1036 1327 -1002 4 FreeSans 2000 0 0 0 CMOS_AND_1/B
rlabel metal1 1585 -315 1625 -275 2 CMOS_AND_1/GND!
rlabel metal1 1585 -1893 1625 -1853 2 CMOS_AND_1/VDD
flabel locali 3175 412 3209 446 2 FreeSans 2000 0 0 0 CMOS_AND_0/AND
flabel locali 2685 -198 2719 -164 2 FreeSans 2000 0 0 0 CMOS_AND_0/A
flabel locali 2505 412 2539 446 2 FreeSans 2000 0 0 0 CMOS_AND_0/B
rlabel metal1 2797 -315 2837 -275 4 CMOS_AND_0/GND!
rlabel metal1 2797 1263 2837 1303 4 CMOS_AND_0/VDD
flabel locali 2535 -1026 2569 -992 4 FreeSans 2000 0 0 0 CMOS_3in_OR_0/A
flabel locali 2685 -426 2719 -392 4 FreeSans 2000 0 0 0 CMOS_3in_OR_0/B
flabel locali 2855 -1776 2889 -1742 4 FreeSans 2000 0 0 0 CMOS_3in_OR_0/C
flabel locali 3325 -923 3359 -889 4 FreeSans 2000 0 0 0 CMOS_3in_OR_0/OR
rlabel metal1 2797 -315 2837 -275 2 CMOS_3in_OR_0/GND!
rlabel metal1 2797 -1893 2837 -1853 2 CMOS_3in_OR_0/VDD
flabel locali 115 -1776 149 -1742 4 FreeSans 2000 0 0 0 CMOS_3in_AND_0/A
flabel locali -85 -426 -51 -392 4 FreeSans 2000 0 0 0 CMOS_3in_AND_0/B
flabel locali -235 -1026 -201 -992 4 FreeSans 2000 0 0 0 CMOS_3in_AND_0/C
flabel locali 555 -941 589 -907 4 FreeSans 2000 0 0 0 CMOS_3in_AND_0/OUT
rlabel metal1 27 -1893 67 -1853 2 CMOS_3in_AND_0/VDD
rlabel metal1 27 -315 67 -275 2 CMOS_3in_AND_0/GND!
flabel locali 1828 1152 1862 1186 2 FreeSans 2500 0 0 0 CMOS_XOR_0/B
flabel locali 1828 -198 1862 -164 2 FreeSans 2500 0 0 0 CMOS_XOR_0/A_bar
flabel locali 1378 227 1412 261 2 FreeSans 2500 0 0 0 CMOS_XOR_0/A
rlabel locali 1342 410 1391 457 4 CMOS_XOR_0/B_bar
rlabel metal1 1585 -315 1625 -275 4 CMOS_XOR_0/GND!
rlabel metal1 1585 1263 1625 1303 4 CMOS_XOR_0/VDD
flabel metal2 1985 325 2021 361 2 FreeSans 2500 0 0 0 CMOS_XOR_0/XOR
flabel locali 771 317 805 351 2 FreeSans 2500 0 0 0 CMOS_XNOR_0/XNOR
flabel locali 270 1152 304 1186 2 FreeSans 3126 0 0 0 CMOS_XNOR_0/B
flabel locali 270 -198 304 -164 2 FreeSans 3126 0 0 0 CMOS_XNOR_0/A_bar
flabel locali -180 227 -146 261 2 FreeSans 3126 0 0 0 CMOS_XNOR_0/A
rlabel locali -216 410 -167 457 4 CMOS_XNOR_0/B_bar
rlabel metal1 27 -315 67 -275 4 CMOS_XNOR_0/GND!
rlabel metal1 27 1263 67 1303 4 CMOS_XNOR_0/VDD
<< end >>
