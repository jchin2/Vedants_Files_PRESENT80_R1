magic
tech sky130A
magscale 1 2
timestamp 1676578411
<< nwell >>
rect -1231 2000 -279 2230
rect -1210 1310 -320 2000
<< pwell >>
rect -1196 718 -334 1152
rect -1221 566 -289 718
<< nmos >>
rect -1050 826 -1020 1126
rect -900 826 -870 1126
rect -510 826 -480 1126
<< pmos >>
rect -1050 1360 -1020 1960
rect -900 1360 -870 1960
rect -510 1360 -480 1960
<< ndiff >>
rect -1170 1095 -1050 1126
rect -1170 1061 -1127 1095
rect -1093 1061 -1050 1095
rect -1170 1027 -1050 1061
rect -1170 993 -1127 1027
rect -1093 993 -1050 1027
rect -1170 959 -1050 993
rect -1170 925 -1127 959
rect -1093 925 -1050 959
rect -1170 891 -1050 925
rect -1170 857 -1127 891
rect -1093 857 -1050 891
rect -1170 826 -1050 857
rect -1020 1095 -900 1126
rect -1020 1061 -977 1095
rect -943 1061 -900 1095
rect -1020 1027 -900 1061
rect -1020 993 -977 1027
rect -943 993 -900 1027
rect -1020 959 -900 993
rect -1020 925 -977 959
rect -943 925 -900 959
rect -1020 891 -900 925
rect -1020 857 -977 891
rect -943 857 -900 891
rect -1020 826 -900 857
rect -870 1095 -750 1126
rect -870 1061 -827 1095
rect -793 1061 -750 1095
rect -870 1027 -750 1061
rect -870 993 -827 1027
rect -793 993 -750 1027
rect -870 959 -750 993
rect -870 925 -827 959
rect -793 925 -750 959
rect -870 891 -750 925
rect -870 857 -827 891
rect -793 857 -750 891
rect -870 826 -750 857
rect -630 1095 -510 1126
rect -630 1061 -587 1095
rect -553 1061 -510 1095
rect -630 1027 -510 1061
rect -630 993 -587 1027
rect -553 993 -510 1027
rect -630 959 -510 993
rect -630 925 -587 959
rect -553 925 -510 959
rect -630 891 -510 925
rect -630 857 -587 891
rect -553 857 -510 891
rect -630 826 -510 857
rect -480 1095 -360 1126
rect -480 1061 -437 1095
rect -403 1061 -360 1095
rect -480 1027 -360 1061
rect -480 993 -437 1027
rect -403 993 -360 1027
rect -480 959 -360 993
rect -480 925 -437 959
rect -403 925 -360 959
rect -480 891 -360 925
rect -480 857 -437 891
rect -403 857 -360 891
rect -480 826 -360 857
<< pdiff >>
rect -1170 1915 -1050 1960
rect -1170 1881 -1127 1915
rect -1093 1881 -1050 1915
rect -1170 1847 -1050 1881
rect -1170 1813 -1127 1847
rect -1093 1813 -1050 1847
rect -1170 1779 -1050 1813
rect -1170 1745 -1127 1779
rect -1093 1745 -1050 1779
rect -1170 1711 -1050 1745
rect -1170 1677 -1127 1711
rect -1093 1677 -1050 1711
rect -1170 1643 -1050 1677
rect -1170 1609 -1127 1643
rect -1093 1609 -1050 1643
rect -1170 1575 -1050 1609
rect -1170 1541 -1127 1575
rect -1093 1541 -1050 1575
rect -1170 1507 -1050 1541
rect -1170 1473 -1127 1507
rect -1093 1473 -1050 1507
rect -1170 1439 -1050 1473
rect -1170 1405 -1127 1439
rect -1093 1405 -1050 1439
rect -1170 1360 -1050 1405
rect -1020 1360 -900 1960
rect -870 1915 -750 1960
rect -870 1881 -827 1915
rect -793 1881 -750 1915
rect -870 1847 -750 1881
rect -870 1813 -827 1847
rect -793 1813 -750 1847
rect -870 1779 -750 1813
rect -870 1745 -827 1779
rect -793 1745 -750 1779
rect -870 1711 -750 1745
rect -870 1677 -827 1711
rect -793 1677 -750 1711
rect -870 1643 -750 1677
rect -870 1609 -827 1643
rect -793 1609 -750 1643
rect -870 1575 -750 1609
rect -870 1541 -827 1575
rect -793 1541 -750 1575
rect -870 1507 -750 1541
rect -870 1473 -827 1507
rect -793 1473 -750 1507
rect -870 1439 -750 1473
rect -870 1405 -827 1439
rect -793 1405 -750 1439
rect -870 1360 -750 1405
rect -630 1915 -510 1960
rect -630 1881 -587 1915
rect -553 1881 -510 1915
rect -630 1847 -510 1881
rect -630 1813 -587 1847
rect -553 1813 -510 1847
rect -630 1779 -510 1813
rect -630 1745 -587 1779
rect -553 1745 -510 1779
rect -630 1711 -510 1745
rect -630 1677 -587 1711
rect -553 1677 -510 1711
rect -630 1643 -510 1677
rect -630 1609 -587 1643
rect -553 1609 -510 1643
rect -630 1575 -510 1609
rect -630 1541 -587 1575
rect -553 1541 -510 1575
rect -630 1507 -510 1541
rect -630 1473 -587 1507
rect -553 1473 -510 1507
rect -630 1439 -510 1473
rect -630 1405 -587 1439
rect -553 1405 -510 1439
rect -630 1360 -510 1405
rect -480 1915 -360 1960
rect -480 1881 -437 1915
rect -403 1881 -360 1915
rect -480 1847 -360 1881
rect -480 1813 -437 1847
rect -403 1813 -360 1847
rect -480 1779 -360 1813
rect -480 1745 -437 1779
rect -403 1745 -360 1779
rect -480 1711 -360 1745
rect -480 1677 -437 1711
rect -403 1677 -360 1711
rect -480 1643 -360 1677
rect -480 1609 -437 1643
rect -403 1609 -360 1643
rect -480 1575 -360 1609
rect -480 1541 -437 1575
rect -403 1541 -360 1575
rect -480 1507 -360 1541
rect -480 1473 -437 1507
rect -403 1473 -360 1507
rect -480 1439 -360 1473
rect -480 1405 -437 1439
rect -403 1405 -360 1439
rect -480 1360 -360 1405
<< ndiffc >>
rect -1127 1061 -1093 1095
rect -1127 993 -1093 1027
rect -1127 925 -1093 959
rect -1127 857 -1093 891
rect -977 1061 -943 1095
rect -977 993 -943 1027
rect -977 925 -943 959
rect -977 857 -943 891
rect -827 1061 -793 1095
rect -827 993 -793 1027
rect -827 925 -793 959
rect -827 857 -793 891
rect -587 1061 -553 1095
rect -587 993 -553 1027
rect -587 925 -553 959
rect -587 857 -553 891
rect -437 1061 -403 1095
rect -437 993 -403 1027
rect -437 925 -403 959
rect -437 857 -403 891
<< pdiffc >>
rect -1127 1881 -1093 1915
rect -1127 1813 -1093 1847
rect -1127 1745 -1093 1779
rect -1127 1677 -1093 1711
rect -1127 1609 -1093 1643
rect -1127 1541 -1093 1575
rect -1127 1473 -1093 1507
rect -1127 1405 -1093 1439
rect -827 1881 -793 1915
rect -827 1813 -793 1847
rect -827 1745 -793 1779
rect -827 1677 -793 1711
rect -827 1609 -793 1643
rect -827 1541 -793 1575
rect -827 1473 -793 1507
rect -827 1405 -793 1439
rect -587 1881 -553 1915
rect -587 1813 -553 1847
rect -587 1745 -553 1779
rect -587 1677 -553 1711
rect -587 1609 -553 1643
rect -587 1541 -553 1575
rect -587 1473 -553 1507
rect -587 1405 -553 1439
rect -437 1881 -403 1915
rect -437 1813 -403 1847
rect -437 1745 -403 1779
rect -437 1677 -403 1711
rect -437 1609 -403 1643
rect -437 1541 -403 1575
rect -437 1473 -403 1507
rect -437 1405 -403 1439
<< psubdiff >>
rect -1195 659 -315 692
rect -1195 625 -1172 659
rect -1138 625 -1100 659
rect -1066 625 -1028 659
rect -994 625 -956 659
rect -922 625 -884 659
rect -850 625 -812 659
rect -778 625 -740 659
rect -706 625 -668 659
rect -634 625 -596 659
rect -562 625 -524 659
rect -490 625 -452 659
rect -418 625 -380 659
rect -346 625 -315 659
rect -1195 592 -315 625
<< nsubdiff >>
rect -1195 2161 -315 2194
rect -1195 2127 -1172 2161
rect -1138 2127 -1100 2161
rect -1066 2127 -1028 2161
rect -994 2127 -956 2161
rect -922 2127 -884 2161
rect -850 2127 -812 2161
rect -778 2127 -740 2161
rect -706 2127 -668 2161
rect -634 2127 -596 2161
rect -562 2127 -524 2161
rect -490 2127 -452 2161
rect -418 2127 -380 2161
rect -346 2127 -315 2161
rect -1195 2094 -315 2127
<< psubdiffcont >>
rect -1172 625 -1138 659
rect -1100 625 -1066 659
rect -1028 625 -994 659
rect -956 625 -922 659
rect -884 625 -850 659
rect -812 625 -778 659
rect -740 625 -706 659
rect -668 625 -634 659
rect -596 625 -562 659
rect -524 625 -490 659
rect -452 625 -418 659
rect -380 625 -346 659
<< nsubdiffcont >>
rect -1172 2127 -1138 2161
rect -1100 2127 -1066 2161
rect -1028 2127 -994 2161
rect -956 2127 -922 2161
rect -884 2127 -850 2161
rect -812 2127 -778 2161
rect -740 2127 -706 2161
rect -668 2127 -634 2161
rect -596 2127 -562 2161
rect -524 2127 -490 2161
rect -452 2127 -418 2161
rect -380 2127 -346 2161
<< poly >>
rect -1050 1960 -1020 1990
rect -900 1960 -870 1990
rect -510 1960 -480 1990
rect -1050 1330 -1020 1360
rect -1130 1307 -1020 1330
rect -1130 1273 -1107 1307
rect -1073 1273 -1020 1307
rect -1130 1250 -1020 1273
rect -1050 1126 -1020 1250
rect -900 1126 -870 1360
rect -510 1330 -480 1360
rect -590 1307 -480 1330
rect -590 1273 -567 1307
rect -533 1273 -480 1307
rect -590 1250 -480 1273
rect -510 1126 -480 1250
rect -1050 796 -1020 826
rect -900 796 -870 826
rect -510 796 -480 826
rect -950 773 -870 796
rect -950 739 -927 773
rect -893 739 -870 773
rect -950 716 -870 739
<< polycont >>
rect -1107 1273 -1073 1307
rect -567 1273 -533 1307
rect -927 739 -893 773
<< locali >>
rect -1195 2161 -315 2184
rect -1195 2127 -1172 2161
rect -1138 2127 -1100 2161
rect -1066 2127 -1028 2161
rect -994 2127 -956 2161
rect -922 2127 -884 2161
rect -850 2127 -812 2161
rect -778 2127 -740 2161
rect -706 2127 -668 2161
rect -634 2127 -596 2161
rect -562 2127 -524 2161
rect -490 2127 -452 2161
rect -418 2127 -380 2161
rect -346 2127 -315 2161
rect -1195 2104 -315 2127
rect -1150 1929 -1070 1940
rect -1150 1881 -1127 1929
rect -1093 1881 -1070 1929
rect -1150 1857 -1070 1881
rect -1150 1813 -1127 1857
rect -1093 1813 -1070 1857
rect -1150 1785 -1070 1813
rect -1150 1745 -1127 1785
rect -1093 1745 -1070 1785
rect -1150 1713 -1070 1745
rect -1150 1677 -1127 1713
rect -1093 1677 -1070 1713
rect -1150 1643 -1070 1677
rect -1150 1607 -1127 1643
rect -1093 1607 -1070 1643
rect -1150 1575 -1070 1607
rect -1150 1535 -1127 1575
rect -1093 1535 -1070 1575
rect -1150 1507 -1070 1535
rect -1150 1463 -1127 1507
rect -1093 1463 -1070 1507
rect -1150 1439 -1070 1463
rect -1150 1391 -1127 1439
rect -1093 1391 -1070 1439
rect -1150 1380 -1070 1391
rect -850 1915 -770 1940
rect -850 1881 -827 1915
rect -793 1881 -770 1915
rect -850 1847 -770 1881
rect -850 1813 -827 1847
rect -793 1813 -770 1847
rect -850 1779 -770 1813
rect -850 1745 -827 1779
rect -793 1745 -770 1779
rect -850 1711 -770 1745
rect -850 1677 -827 1711
rect -793 1677 -770 1711
rect -850 1643 -770 1677
rect -850 1609 -827 1643
rect -793 1609 -770 1643
rect -850 1575 -770 1609
rect -850 1541 -827 1575
rect -793 1541 -770 1575
rect -850 1507 -770 1541
rect -850 1473 -827 1507
rect -793 1473 -770 1507
rect -850 1439 -770 1473
rect -850 1405 -827 1439
rect -793 1405 -770 1439
rect -850 1380 -770 1405
rect -610 1929 -530 1940
rect -610 1881 -587 1929
rect -553 1881 -530 1929
rect -610 1857 -530 1881
rect -610 1813 -587 1857
rect -553 1813 -530 1857
rect -610 1785 -530 1813
rect -610 1745 -587 1785
rect -553 1745 -530 1785
rect -610 1713 -530 1745
rect -610 1677 -587 1713
rect -553 1677 -530 1713
rect -610 1643 -530 1677
rect -610 1607 -587 1643
rect -553 1607 -530 1643
rect -610 1575 -530 1607
rect -610 1535 -587 1575
rect -553 1535 -530 1575
rect -610 1507 -530 1535
rect -610 1463 -587 1507
rect -553 1463 -530 1507
rect -610 1439 -530 1463
rect -610 1391 -587 1439
rect -553 1391 -530 1439
rect -610 1380 -530 1391
rect -460 1915 -380 1940
rect -460 1881 -437 1915
rect -403 1881 -380 1915
rect -460 1847 -380 1881
rect -460 1813 -437 1847
rect -403 1813 -380 1847
rect -460 1779 -380 1813
rect -460 1745 -437 1779
rect -403 1745 -380 1779
rect -460 1711 -380 1745
rect -460 1677 -437 1711
rect -403 1677 -380 1711
rect -460 1643 -380 1677
rect -460 1609 -437 1643
rect -403 1609 -380 1643
rect -460 1575 -380 1609
rect -460 1541 -437 1575
rect -403 1541 -380 1575
rect -460 1507 -380 1541
rect -460 1473 -437 1507
rect -403 1473 -380 1507
rect -460 1439 -380 1473
rect -460 1405 -437 1439
rect -403 1405 -380 1439
rect -460 1380 -380 1405
rect -1130 1307 -1050 1330
rect -830 1310 -790 1380
rect -590 1310 -510 1330
rect -1130 1273 -1107 1307
rect -1073 1273 -1050 1307
rect -1130 1250 -1050 1273
rect -980 1307 -510 1310
rect -980 1273 -567 1307
rect -533 1273 -510 1307
rect -980 1270 -510 1273
rect -980 1106 -940 1270
rect -590 1250 -510 1270
rect -440 1106 -400 1380
rect -1150 1095 -1070 1106
rect -1150 1031 -1127 1095
rect -1093 1031 -1070 1095
rect -1150 1027 -1070 1031
rect -1150 925 -1127 1027
rect -1093 925 -1070 1027
rect -1150 921 -1070 925
rect -1150 857 -1127 921
rect -1093 857 -1070 921
rect -1150 846 -1070 857
rect -1000 1095 -920 1106
rect -1000 1061 -977 1095
rect -943 1061 -920 1095
rect -1000 1027 -920 1061
rect -1000 993 -977 1027
rect -943 993 -920 1027
rect -1000 959 -920 993
rect -1000 925 -977 959
rect -943 925 -920 959
rect -1000 891 -920 925
rect -1000 857 -977 891
rect -943 857 -920 891
rect -1000 846 -920 857
rect -850 1095 -770 1106
rect -850 1031 -827 1095
rect -793 1031 -770 1095
rect -850 1027 -770 1031
rect -850 925 -827 1027
rect -793 925 -770 1027
rect -850 921 -770 925
rect -850 857 -827 921
rect -793 857 -770 921
rect -850 846 -770 857
rect -610 1095 -530 1106
rect -610 1031 -587 1095
rect -553 1031 -530 1095
rect -610 1027 -530 1031
rect -610 925 -587 1027
rect -553 925 -530 1027
rect -610 921 -530 925
rect -610 857 -587 921
rect -553 857 -530 921
rect -610 846 -530 857
rect -460 1095 -380 1106
rect -460 1061 -437 1095
rect -403 1061 -380 1095
rect -460 1027 -380 1061
rect -460 993 -437 1027
rect -403 993 -380 1027
rect -460 959 -380 993
rect -460 925 -437 959
rect -403 925 -380 959
rect -460 891 -380 925
rect -460 857 -437 891
rect -403 857 -380 891
rect -460 846 -380 857
rect -950 773 -870 796
rect -950 739 -927 773
rect -893 739 -870 773
rect -950 716 -870 739
rect -1195 659 -315 682
rect -1195 625 -1172 659
rect -1138 625 -1100 659
rect -1066 625 -1028 659
rect -994 625 -956 659
rect -922 625 -884 659
rect -850 625 -812 659
rect -778 625 -740 659
rect -706 625 -668 659
rect -634 625 -596 659
rect -562 625 -524 659
rect -490 625 -452 659
rect -418 625 -380 659
rect -346 625 -315 659
rect -1195 602 -315 625
<< viali >>
rect -1172 2127 -1138 2161
rect -1100 2127 -1066 2161
rect -1028 2127 -994 2161
rect -956 2127 -922 2161
rect -884 2127 -850 2161
rect -812 2127 -778 2161
rect -740 2127 -706 2161
rect -668 2127 -634 2161
rect -596 2127 -562 2161
rect -524 2127 -490 2161
rect -452 2127 -418 2161
rect -380 2127 -346 2161
rect -1127 1915 -1093 1929
rect -1127 1895 -1093 1915
rect -1127 1847 -1093 1857
rect -1127 1823 -1093 1847
rect -1127 1779 -1093 1785
rect -1127 1751 -1093 1779
rect -1127 1711 -1093 1713
rect -1127 1679 -1093 1711
rect -1127 1609 -1093 1641
rect -1127 1607 -1093 1609
rect -1127 1541 -1093 1569
rect -1127 1535 -1093 1541
rect -1127 1473 -1093 1497
rect -1127 1463 -1093 1473
rect -1127 1405 -1093 1425
rect -1127 1391 -1093 1405
rect -587 1915 -553 1929
rect -587 1895 -553 1915
rect -587 1847 -553 1857
rect -587 1823 -553 1847
rect -587 1779 -553 1785
rect -587 1751 -553 1779
rect -587 1711 -553 1713
rect -587 1679 -553 1711
rect -587 1609 -553 1641
rect -587 1607 -553 1609
rect -587 1541 -553 1569
rect -587 1535 -553 1541
rect -587 1473 -553 1497
rect -587 1463 -553 1473
rect -587 1405 -553 1425
rect -587 1391 -553 1405
rect -1127 1061 -1093 1065
rect -1127 1031 -1093 1061
rect -1127 959 -1093 993
rect -1127 891 -1093 921
rect -1127 887 -1093 891
rect -827 1061 -793 1065
rect -827 1031 -793 1061
rect -827 959 -793 993
rect -827 891 -793 921
rect -827 887 -793 891
rect -587 1061 -553 1065
rect -587 1031 -553 1061
rect -587 959 -553 993
rect -587 891 -553 921
rect -587 887 -553 891
rect -1172 625 -1138 659
rect -1100 625 -1066 659
rect -1028 625 -994 659
rect -956 625 -922 659
rect -884 625 -850 659
rect -812 625 -778 659
rect -740 625 -706 659
rect -668 625 -634 659
rect -596 625 -562 659
rect -524 625 -490 659
rect -452 625 -418 659
rect -380 625 -346 659
<< metal1 >>
rect -1195 2161 -315 2194
rect -1195 2127 -1172 2161
rect -1138 2127 -1100 2161
rect -1066 2127 -1028 2161
rect -994 2127 -956 2161
rect -922 2127 -884 2161
rect -850 2127 -812 2161
rect -778 2127 -740 2161
rect -706 2127 -668 2161
rect -634 2127 -596 2161
rect -562 2127 -524 2161
rect -490 2127 -452 2161
rect -418 2127 -380 2161
rect -346 2127 -315 2161
rect -1195 2094 -315 2127
rect -1130 1940 -1090 2094
rect -590 1940 -550 2094
rect -1150 1929 -1070 1940
rect -1150 1895 -1127 1929
rect -1093 1895 -1070 1929
rect -1150 1857 -1070 1895
rect -1150 1823 -1127 1857
rect -1093 1823 -1070 1857
rect -1150 1785 -1070 1823
rect -1150 1751 -1127 1785
rect -1093 1751 -1070 1785
rect -1150 1713 -1070 1751
rect -1150 1679 -1127 1713
rect -1093 1679 -1070 1713
rect -1150 1641 -1070 1679
rect -1150 1607 -1127 1641
rect -1093 1607 -1070 1641
rect -1150 1569 -1070 1607
rect -1150 1535 -1127 1569
rect -1093 1535 -1070 1569
rect -1150 1497 -1070 1535
rect -1150 1463 -1127 1497
rect -1093 1463 -1070 1497
rect -1150 1425 -1070 1463
rect -1150 1391 -1127 1425
rect -1093 1391 -1070 1425
rect -1150 1380 -1070 1391
rect -610 1929 -530 1940
rect -610 1895 -587 1929
rect -553 1895 -530 1929
rect -610 1857 -530 1895
rect -610 1823 -587 1857
rect -553 1823 -530 1857
rect -610 1785 -530 1823
rect -610 1751 -587 1785
rect -553 1751 -530 1785
rect -610 1713 -530 1751
rect -610 1679 -587 1713
rect -553 1679 -530 1713
rect -610 1641 -530 1679
rect -610 1607 -587 1641
rect -553 1607 -530 1641
rect -610 1569 -530 1607
rect -610 1535 -587 1569
rect -553 1535 -530 1569
rect -610 1497 -530 1535
rect -610 1463 -587 1497
rect -553 1463 -530 1497
rect -610 1425 -530 1463
rect -610 1391 -587 1425
rect -553 1391 -530 1425
rect -610 1380 -530 1391
rect -1150 1065 -1070 1106
rect -1150 1031 -1127 1065
rect -1093 1031 -1070 1065
rect -1150 993 -1070 1031
rect -1150 959 -1127 993
rect -1093 959 -1070 993
rect -1150 921 -1070 959
rect -1150 887 -1127 921
rect -1093 887 -1070 921
rect -1150 846 -1070 887
rect -850 1065 -770 1106
rect -850 1031 -827 1065
rect -793 1031 -770 1065
rect -850 993 -770 1031
rect -850 959 -827 993
rect -793 959 -770 993
rect -850 921 -770 959
rect -850 887 -827 921
rect -793 887 -770 921
rect -850 846 -770 887
rect -610 1065 -530 1106
rect -610 1031 -587 1065
rect -553 1031 -530 1065
rect -610 993 -530 1031
rect -610 959 -587 993
rect -553 959 -530 993
rect -610 921 -530 959
rect -610 887 -587 921
rect -553 887 -530 921
rect -610 846 -530 887
rect -1130 692 -1090 846
rect -830 692 -790 846
rect -590 692 -550 846
rect -1195 659 -315 692
rect -1195 625 -1172 659
rect -1138 625 -1100 659
rect -1066 625 -1028 659
rect -994 625 -956 659
rect -922 625 -884 659
rect -850 625 -812 659
rect -778 625 -740 659
rect -706 625 -668 659
rect -634 625 -596 659
rect -562 625 -524 659
rect -490 625 -452 659
rect -418 625 -380 659
rect -346 625 -315 659
rect -1195 592 -315 625
<< labels >>
rlabel metal1 s -815 622 -775 662 4 GND!
port 1 nsew
rlabel metal1 s -815 2124 -775 2164 4 VDD
port 2 nsew
flabel locali s -437 1273 -403 1307 2 FreeSans 2000 0 0 0 OR
port 3 nsew
flabel locali s -1107 1273 -1073 1307 2 FreeSans 2000 0 0 0 A
port 4 nsew
flabel locali s -927 739 -893 773 2 FreeSans 2000 0 0 0 B
port 5 nsew
<< properties >>
string path -2.850 9.700 -2.850 10.470 
<< end >>
