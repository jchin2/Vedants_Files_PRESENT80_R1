magic
tech sky130A
timestamp 1676418097
<< error_p >>
rect -745 410 -150 755
rect -725 205 -665 355
rect -650 205 -590 355
rect -575 205 -515 355
rect -500 205 -440 355
rect -425 205 -365 355
rect -305 205 -245 355
rect -230 205 -170 355
<< nwell >>
rect -745 410 -150 755
<< nmos >>
rect -665 205 -650 355
rect -590 205 -575 355
rect -515 205 -500 355
rect -440 205 -425 355
rect -245 205 -230 355
<< pmos >>
rect -665 435 -650 735
rect -590 435 -575 735
rect -515 435 -500 735
rect -440 435 -425 735
rect -245 435 -230 735
<< ndiff >>
rect -725 340 -665 355
rect -725 220 -705 340
rect -685 220 -665 340
rect -725 205 -665 220
rect -650 205 -590 355
rect -575 205 -515 355
rect -500 205 -440 355
rect -425 340 -365 355
rect -425 220 -405 340
rect -385 220 -365 340
rect -425 205 -365 220
rect -305 340 -245 355
rect -305 220 -285 340
rect -265 220 -245 340
rect -305 205 -245 220
rect -230 340 -170 355
rect -230 220 -210 340
rect -190 220 -170 340
rect -230 205 -170 220
<< pdiff >>
rect -725 720 -665 735
rect -725 450 -705 720
rect -685 450 -665 720
rect -725 435 -665 450
rect -650 720 -590 735
rect -650 450 -630 720
rect -610 450 -590 720
rect -650 435 -590 450
rect -575 720 -515 735
rect -575 450 -555 720
rect -535 450 -515 720
rect -575 435 -515 450
rect -500 720 -440 735
rect -500 450 -480 720
rect -460 450 -440 720
rect -500 435 -440 450
rect -425 720 -365 735
rect -425 450 -405 720
rect -385 450 -365 720
rect -425 435 -365 450
rect -305 720 -245 735
rect -305 450 -285 720
rect -265 450 -245 720
rect -305 435 -245 450
rect -230 715 -170 735
rect -230 455 -210 715
rect -190 455 -170 715
rect -230 435 -170 455
<< ndiffc >>
rect -705 220 -685 340
rect -405 220 -385 340
rect -285 220 -265 340
rect -210 220 -190 340
<< pdiffc >>
rect -705 450 -685 720
rect -630 450 -610 720
rect -555 450 -535 720
rect -480 450 -460 720
rect -405 450 -385 720
rect -285 450 -265 720
rect -210 455 -190 715
<< poly >>
rect -690 780 -650 790
rect -690 760 -680 780
rect -660 760 -650 780
rect -690 750 -650 760
rect -665 735 -650 750
rect -590 735 -575 750
rect -515 735 -500 750
rect -440 735 -425 750
rect -245 735 -230 750
rect -665 355 -650 435
rect -590 415 -575 435
rect -615 405 -575 415
rect -615 385 -605 405
rect -585 385 -575 405
rect -615 375 -575 385
rect -590 355 -575 375
rect -515 355 -500 435
rect -440 355 -425 435
rect -245 420 -230 435
rect -285 410 -230 420
rect -285 390 -275 410
rect -255 390 -230 410
rect -285 380 -230 390
rect -245 355 -230 380
rect -665 190 -650 205
rect -590 190 -575 205
rect -515 190 -500 205
rect -540 180 -500 190
rect -540 160 -530 180
rect -510 160 -500 180
rect -540 150 -500 160
rect -440 140 -425 205
rect -245 190 -230 205
rect -455 130 -415 140
rect -455 110 -445 130
rect -425 110 -415 130
rect -455 100 -415 110
<< polycont >>
rect -680 760 -660 780
rect -605 385 -585 405
rect -275 390 -255 410
rect -530 160 -510 180
rect -445 110 -425 130
<< locali >>
rect -690 780 -650 790
rect -690 760 -680 780
rect -660 760 -650 780
rect -690 750 -650 760
rect -630 745 -460 765
rect -630 725 -610 745
rect -480 725 -460 745
rect -715 720 -675 725
rect -715 450 -705 720
rect -685 450 -675 720
rect -715 445 -675 450
rect -640 720 -600 725
rect -640 450 -630 720
rect -610 450 -600 720
rect -640 445 -600 450
rect -565 720 -525 725
rect -565 450 -555 720
rect -535 450 -525 720
rect -565 445 -525 450
rect -490 720 -450 725
rect -490 450 -480 720
rect -460 450 -450 720
rect -490 445 -450 450
rect -415 720 -375 725
rect -415 450 -405 720
rect -385 450 -375 720
rect -415 445 -375 450
rect -295 720 -255 725
rect -295 450 -285 720
rect -265 450 -255 720
rect -295 445 -255 450
rect -220 715 -180 725
rect -220 455 -210 715
rect -190 455 -180 715
rect -220 445 -180 455
rect -615 405 -575 415
rect -615 385 -605 405
rect -585 385 -575 405
rect -480 410 -460 445
rect -285 410 -245 420
rect -480 390 -275 410
rect -255 390 -245 410
rect -615 375 -575 385
rect -405 345 -385 390
rect -285 380 -245 390
rect -210 345 -190 445
rect -715 340 -675 345
rect -715 220 -705 340
rect -685 220 -675 340
rect -715 215 -675 220
rect -415 340 -375 345
rect -415 220 -405 340
rect -385 220 -375 340
rect -415 215 -375 220
rect -295 340 -255 345
rect -295 220 -285 340
rect -265 220 -255 340
rect -295 215 -255 220
rect -220 340 -180 345
rect -220 220 -210 340
rect -190 220 -180 340
rect -220 215 -180 220
rect -540 180 -500 190
rect -540 160 -530 180
rect -510 160 -500 180
rect -540 150 -500 160
rect -455 130 -415 140
rect -455 110 -445 130
rect -425 110 -415 130
rect -455 100 -415 110
<< viali >>
rect -705 450 -685 720
rect -555 450 -535 720
rect -405 450 -385 720
rect -285 450 -265 720
rect -705 220 -685 340
rect -285 220 -265 340
<< metal1 >>
rect -715 720 -675 725
rect -715 450 -705 720
rect -685 450 -675 720
rect -715 445 -675 450
rect -565 720 -525 725
rect -565 450 -555 720
rect -535 450 -525 720
rect -565 445 -525 450
rect -415 720 -375 725
rect -415 450 -405 720
rect -385 450 -375 720
rect -415 445 -375 450
rect -295 720 -255 725
rect -295 450 -285 720
rect -265 450 -255 720
rect -295 445 -255 450
rect -715 340 -675 345
rect -715 220 -705 340
rect -685 220 -675 340
rect -715 215 -675 220
rect -295 340 -255 345
rect -295 220 -285 340
rect -265 220 -255 340
rect -295 215 -255 220
<< end >>
