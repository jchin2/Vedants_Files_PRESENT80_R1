* NGSPICE file created from CMOS_s3.ext - technology: sky130A

.subckt CMOS_AND GND AND A B VDD
X0 a_n265_0# B VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=5.4e+12p ps=2.16e+07u w=3e+06u l=150000u
X1 VDD A a_n265_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2 a_n265_0# A a_n265_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X3 AND a_n265_0# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X4 a_n265_n610# B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X5 AND a_n265_0# GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt CMOS_3in_OR GND A B C OR VDD
X0 a_n480_n610# B GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+12p pd=8.4e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X1 OR a_n480_n610# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X2 a_n480_n610# C a_n180_0# VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X3 GND A a_n480_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 OR a_n480_n610# GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n330_0# A VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X6 a_n180_0# B a_n330_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X7 GND C a_n480_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt CMOS_XNOR GND XNOR B A_bar A B_bar VDD
X0 XNOR a_n233_n610# GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=2.7e+12p ps=1.26e+07u w=1.5e+06u l=150000u
X1 a_n383_n610# A GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n233_n610# B a_n383_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n383_0# B_bar VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=5.4e+12p ps=2.16e+07u w=3e+06u l=150000u
X4 a_n233_n610# A a_n383_0# VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X5 a_n83_0# A_bar a_n233_n610# VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X6 a_n83_n610# B_bar a_n233_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X7 GND A_bar a_n83_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 XNOR a_n233_n610# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=0p ps=0u w=3e+06u l=150000u
X9 VDD B a_n83_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
.ends

.subckt CMOS_3in_AND GND A B C OUT VDD
X0 a_n180_n610# B a_n330_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X1 OUT a_n480_0# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=5.4e+12p ps=2.16e+07u w=3e+06u l=150000u
X2 VDD A a_n480_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.6e+12p ps=1.44e+07u w=3e+06u l=150000u
X3 a_n330_n610# C GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X4 OUT a_n480_0# GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 VDD C a_n480_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X6 a_n480_0# B VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X7 a_n480_0# A a_n180_n610# GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt CMOS_XOR GND XOR B A_bar A B_bar VDD
X0 a_90_0# A_bar XOR VDD sky130_fd_pr__pfet_01v8 ad=1.8e+12p pd=7.2e+06u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X1 VDD B a_90_0# VDD sky130_fd_pr__pfet_01v8 ad=3.6e+12p pd=1.44e+07u as=0p ps=0u w=3e+06u l=150000u
X2 a_n210_n610# A GND GND sky130_fd_pr__nfet_01v8 ad=9e+11p pd=4.2e+06u as=1.8e+12p ps=8.4e+06u w=1.5e+06u l=150000u
X3 GND A_bar a_90_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X4 XOR A a_n210_0# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.8e+12p ps=7.2e+06u w=3e+06u l=150000u
X5 a_n210_0# B_bar VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X6 a_90_n610# B_bar XOR GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9e+11p ps=4.2e+06u w=1.5e+06u l=150000u
X7 XOR B a_n210_n610# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt CMOS_s3 GND x0 x0_bar x1 x1_bar x2 x2_bar x3 VDD x3_bar s3
XCMOS_AND_0 GND CMOS_AND_0/AND CMOS_AND_0/A x1 VDD CMOS_AND
XCMOS_AND_1 GND CMOS_AND_1/AND CMOS_AND_1/A x3_bar VDD CMOS_AND
XCMOS_3in_OR_0 GND CMOS_AND_1/AND CMOS_AND_0/AND CMOS_3in_OR_0/C s3 VDD CMOS_3in_OR
XCMOS_XNOR_0 GND CMOS_AND_1/A x0 x1_bar x1 x0_bar VDD CMOS_XNOR
XCMOS_3in_AND_0 GND x2_bar x0 x3 CMOS_3in_OR_0/C VDD CMOS_3in_AND
XCMOS_XOR_0 GND CMOS_AND_0/A x3 x2_bar x2 x3_bar VDD CMOS_XOR
.ends

