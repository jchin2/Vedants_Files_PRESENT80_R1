magic
tech sky130A
magscale 1 2
timestamp 1676578218
<< nwell >>
rect -2556 1280 -1604 1510
rect -2500 590 -1650 1280
<< pwell >>
rect -2466 -78 -1694 356
rect -2546 -230 -1614 -78
<< nmos >>
rect -2320 30 -2290 330
rect -2170 30 -2140 330
rect -2020 30 -1990 330
rect -1870 30 -1840 330
<< pmos >>
rect -2320 640 -2290 1240
rect -2170 640 -2140 1240
rect -2020 640 -1990 1240
rect -1870 640 -1840 1240
<< ndiff >>
rect -2440 299 -2320 330
rect -2440 265 -2397 299
rect -2363 265 -2320 299
rect -2440 231 -2320 265
rect -2440 197 -2397 231
rect -2363 197 -2320 231
rect -2440 163 -2320 197
rect -2440 129 -2397 163
rect -2363 129 -2320 163
rect -2440 95 -2320 129
rect -2440 61 -2397 95
rect -2363 61 -2320 95
rect -2440 30 -2320 61
rect -2290 30 -2170 330
rect -2140 299 -2020 330
rect -2140 265 -2097 299
rect -2063 265 -2020 299
rect -2140 231 -2020 265
rect -2140 197 -2097 231
rect -2063 197 -2020 231
rect -2140 163 -2020 197
rect -2140 129 -2097 163
rect -2063 129 -2020 163
rect -2140 95 -2020 129
rect -2140 61 -2097 95
rect -2063 61 -2020 95
rect -2140 30 -2020 61
rect -1990 30 -1870 330
rect -1840 299 -1720 330
rect -1840 265 -1797 299
rect -1763 265 -1720 299
rect -1840 231 -1720 265
rect -1840 197 -1797 231
rect -1763 197 -1720 231
rect -1840 163 -1720 197
rect -1840 129 -1797 163
rect -1763 129 -1720 163
rect -1840 95 -1720 129
rect -1840 61 -1797 95
rect -1763 61 -1720 95
rect -1840 30 -1720 61
<< pdiff >>
rect -2440 1195 -2320 1240
rect -2440 1161 -2397 1195
rect -2363 1161 -2320 1195
rect -2440 1127 -2320 1161
rect -2440 1093 -2397 1127
rect -2363 1093 -2320 1127
rect -2440 1059 -2320 1093
rect -2440 1025 -2397 1059
rect -2363 1025 -2320 1059
rect -2440 991 -2320 1025
rect -2440 957 -2397 991
rect -2363 957 -2320 991
rect -2440 923 -2320 957
rect -2440 889 -2397 923
rect -2363 889 -2320 923
rect -2440 855 -2320 889
rect -2440 821 -2397 855
rect -2363 821 -2320 855
rect -2440 787 -2320 821
rect -2440 753 -2397 787
rect -2363 753 -2320 787
rect -2440 719 -2320 753
rect -2440 685 -2397 719
rect -2363 685 -2320 719
rect -2440 640 -2320 685
rect -2290 640 -2170 1240
rect -2140 1195 -2020 1240
rect -2140 1161 -2097 1195
rect -2063 1161 -2020 1195
rect -2140 1127 -2020 1161
rect -2140 1093 -2097 1127
rect -2063 1093 -2020 1127
rect -2140 1059 -2020 1093
rect -2140 1025 -2097 1059
rect -2063 1025 -2020 1059
rect -2140 991 -2020 1025
rect -2140 957 -2097 991
rect -2063 957 -2020 991
rect -2140 923 -2020 957
rect -2140 889 -2097 923
rect -2063 889 -2020 923
rect -2140 855 -2020 889
rect -2140 821 -2097 855
rect -2063 821 -2020 855
rect -2140 787 -2020 821
rect -2140 753 -2097 787
rect -2063 753 -2020 787
rect -2140 719 -2020 753
rect -2140 685 -2097 719
rect -2063 685 -2020 719
rect -2140 640 -2020 685
rect -1990 640 -1870 1240
rect -1840 1195 -1720 1240
rect -1840 1161 -1797 1195
rect -1763 1161 -1720 1195
rect -1840 1127 -1720 1161
rect -1840 1093 -1797 1127
rect -1763 1093 -1720 1127
rect -1840 1059 -1720 1093
rect -1840 1025 -1797 1059
rect -1763 1025 -1720 1059
rect -1840 991 -1720 1025
rect -1840 957 -1797 991
rect -1763 957 -1720 991
rect -1840 923 -1720 957
rect -1840 889 -1797 923
rect -1763 889 -1720 923
rect -1840 855 -1720 889
rect -1840 821 -1797 855
rect -1763 821 -1720 855
rect -1840 787 -1720 821
rect -1840 753 -1797 787
rect -1763 753 -1720 787
rect -1840 719 -1720 753
rect -1840 685 -1797 719
rect -1763 685 -1720 719
rect -1840 640 -1720 685
<< ndiffc >>
rect -2397 265 -2363 299
rect -2397 197 -2363 231
rect -2397 129 -2363 163
rect -2397 61 -2363 95
rect -2097 265 -2063 299
rect -2097 197 -2063 231
rect -2097 129 -2063 163
rect -2097 61 -2063 95
rect -1797 265 -1763 299
rect -1797 197 -1763 231
rect -1797 129 -1763 163
rect -1797 61 -1763 95
<< pdiffc >>
rect -2397 1161 -2363 1195
rect -2397 1093 -2363 1127
rect -2397 1025 -2363 1059
rect -2397 957 -2363 991
rect -2397 889 -2363 923
rect -2397 821 -2363 855
rect -2397 753 -2363 787
rect -2397 685 -2363 719
rect -2097 1161 -2063 1195
rect -2097 1093 -2063 1127
rect -2097 1025 -2063 1059
rect -2097 957 -2063 991
rect -2097 889 -2063 923
rect -2097 821 -2063 855
rect -2097 753 -2063 787
rect -2097 685 -2063 719
rect -1797 1161 -1763 1195
rect -1797 1093 -1763 1127
rect -1797 1025 -1763 1059
rect -1797 957 -1763 991
rect -1797 889 -1763 923
rect -1797 821 -1763 855
rect -1797 753 -1763 787
rect -1797 685 -1763 719
<< psubdiff >>
rect -2520 -137 -1640 -104
rect -2520 -171 -2497 -137
rect -2463 -171 -2425 -137
rect -2391 -171 -2353 -137
rect -2319 -171 -2281 -137
rect -2247 -171 -2209 -137
rect -2175 -171 -2137 -137
rect -2103 -171 -2065 -137
rect -2031 -171 -1993 -137
rect -1959 -171 -1921 -137
rect -1887 -171 -1849 -137
rect -1815 -171 -1777 -137
rect -1743 -171 -1705 -137
rect -1671 -171 -1640 -137
rect -2520 -204 -1640 -171
<< nsubdiff >>
rect -2520 1441 -1640 1474
rect -2520 1407 -2497 1441
rect -2463 1407 -2425 1441
rect -2391 1407 -2353 1441
rect -2319 1407 -2281 1441
rect -2247 1407 -2209 1441
rect -2175 1407 -2137 1441
rect -2103 1407 -2065 1441
rect -2031 1407 -1993 1441
rect -1959 1407 -1921 1441
rect -1887 1407 -1849 1441
rect -1815 1407 -1777 1441
rect -1743 1407 -1705 1441
rect -1671 1407 -1640 1441
rect -2520 1374 -1640 1407
<< psubdiffcont >>
rect -2497 -171 -2463 -137
rect -2425 -171 -2391 -137
rect -2353 -171 -2319 -137
rect -2281 -171 -2247 -137
rect -2209 -171 -2175 -137
rect -2137 -171 -2103 -137
rect -2065 -171 -2031 -137
rect -1993 -171 -1959 -137
rect -1921 -171 -1887 -137
rect -1849 -171 -1815 -137
rect -1777 -171 -1743 -137
rect -1705 -171 -1671 -137
<< nsubdiffcont >>
rect -2497 1407 -2463 1441
rect -2425 1407 -2391 1441
rect -2353 1407 -2319 1441
rect -2281 1407 -2247 1441
rect -2209 1407 -2175 1441
rect -2137 1407 -2103 1441
rect -2065 1407 -2031 1441
rect -1993 1407 -1959 1441
rect -1921 1407 -1887 1441
rect -1849 1407 -1815 1441
rect -1777 1407 -1743 1441
rect -1705 1407 -1671 1441
<< poly >>
rect -1920 1327 -1840 1350
rect -1920 1293 -1897 1327
rect -1863 1293 -1840 1327
rect -1920 1270 -1840 1293
rect -2320 1240 -2290 1270
rect -2170 1240 -2140 1270
rect -2020 1240 -1990 1270
rect -1870 1240 -1840 1270
rect -2320 616 -2290 640
rect -2400 593 -2290 616
rect -2400 559 -2377 593
rect -2343 559 -2290 593
rect -2400 539 -2290 559
rect -2400 536 -2320 539
rect -2170 497 -2140 640
rect -2292 467 -2140 497
rect -2020 497 -1990 640
rect -1870 616 -1840 640
rect -1870 593 -1760 616
rect -1870 559 -1817 593
rect -1783 559 -1760 593
rect -1870 539 -1760 559
rect -1840 536 -1760 539
rect -2020 467 -1868 497
rect -2292 425 -2262 467
rect -2370 402 -2262 425
rect -2370 368 -2347 402
rect -2313 368 -2262 402
rect -2370 360 -2262 368
rect -2220 402 -2140 425
rect -2220 368 -2197 402
rect -2163 368 -2140 402
rect -2370 345 -2290 360
rect -2220 345 -2140 368
rect -2320 330 -2290 345
rect -2170 330 -2140 345
rect -2020 402 -1940 425
rect -2020 368 -1997 402
rect -1963 368 -1940 402
rect -2020 345 -1940 368
rect -1898 382 -1868 467
rect -1898 352 -1840 382
rect -2020 330 -1990 345
rect -1870 330 -1840 352
rect -2320 0 -2290 30
rect -2170 0 -2140 30
rect -2020 0 -1990 30
rect -1870 0 -1840 30
rect -1920 -23 -1840 0
rect -1920 -57 -1897 -23
rect -1863 -57 -1840 -23
rect -1920 -80 -1840 -57
<< polycont >>
rect -1897 1293 -1863 1327
rect -2377 559 -2343 593
rect -1817 559 -1783 593
rect -2347 368 -2313 402
rect -2197 368 -2163 402
rect -1997 368 -1963 402
rect -1897 -57 -1863 -23
<< locali >>
rect -2520 1441 -1640 1464
rect -2520 1407 -2497 1441
rect -2463 1407 -2425 1441
rect -2391 1407 -2353 1441
rect -2319 1407 -2281 1441
rect -2247 1407 -2209 1441
rect -2175 1407 -2137 1441
rect -2103 1407 -2065 1441
rect -2031 1407 -1993 1441
rect -1959 1407 -1921 1441
rect -1887 1407 -1849 1441
rect -1815 1407 -1777 1441
rect -1743 1407 -1705 1441
rect -1671 1407 -1640 1441
rect -2520 1384 -1640 1407
rect -1920 1327 -1840 1350
rect -1920 1293 -1897 1327
rect -1863 1293 -1840 1327
rect -1920 1270 -1840 1293
rect -2420 1209 -2340 1220
rect -2420 1161 -2397 1209
rect -2363 1161 -2340 1209
rect -2420 1137 -2340 1161
rect -2420 1093 -2397 1137
rect -2363 1093 -2340 1137
rect -2420 1065 -2340 1093
rect -2420 1025 -2397 1065
rect -2363 1025 -2340 1065
rect -2420 993 -2340 1025
rect -2420 957 -2397 993
rect -2363 957 -2340 993
rect -2420 923 -2340 957
rect -2420 887 -2397 923
rect -2363 887 -2340 923
rect -2420 855 -2340 887
rect -2420 815 -2397 855
rect -2363 815 -2340 855
rect -2420 787 -2340 815
rect -2420 743 -2397 787
rect -2363 743 -2340 787
rect -2420 719 -2340 743
rect -2420 671 -2397 719
rect -2363 671 -2340 719
rect -2420 660 -2340 671
rect -2120 1209 -2040 1220
rect -2120 1161 -2097 1209
rect -2063 1161 -2040 1209
rect -2120 1137 -2040 1161
rect -2120 1093 -2097 1137
rect -2063 1093 -2040 1137
rect -2120 1065 -2040 1093
rect -2120 1025 -2097 1065
rect -2063 1025 -2040 1065
rect -2120 993 -2040 1025
rect -2120 957 -2097 993
rect -2063 957 -2040 993
rect -2120 923 -2040 957
rect -2120 887 -2097 923
rect -2063 887 -2040 923
rect -2120 855 -2040 887
rect -2120 815 -2097 855
rect -2063 815 -2040 855
rect -2120 787 -2040 815
rect -2120 743 -2097 787
rect -2063 743 -2040 787
rect -2120 719 -2040 743
rect -2120 671 -2097 719
rect -2063 671 -2040 719
rect -2120 660 -2040 671
rect -1820 1209 -1740 1220
rect -1820 1161 -1797 1209
rect -1763 1161 -1740 1209
rect -1820 1137 -1740 1161
rect -1820 1093 -1797 1137
rect -1763 1093 -1740 1137
rect -1820 1065 -1740 1093
rect -1820 1025 -1797 1065
rect -1763 1025 -1740 1065
rect -1820 993 -1740 1025
rect -1820 957 -1797 993
rect -1763 957 -1740 993
rect -1820 923 -1740 957
rect -1820 887 -1797 923
rect -1763 887 -1740 923
rect -1820 855 -1740 887
rect -1820 815 -1797 855
rect -1763 815 -1740 855
rect -1820 787 -1740 815
rect -1820 743 -1797 787
rect -1763 743 -1740 787
rect -1820 719 -1740 743
rect -1820 671 -1797 719
rect -1763 671 -1740 719
rect -1820 660 -1740 671
rect -2400 596 -2320 616
rect -2400 593 -1960 596
rect -2400 559 -2377 593
rect -2343 559 -1960 593
rect -2400 556 -1960 559
rect -2400 536 -2320 556
rect -2000 425 -1960 556
rect -1840 593 -1760 616
rect -1840 559 -1817 593
rect -1783 559 -1760 593
rect -1840 536 -1760 559
rect -2370 402 -2290 425
rect -2370 368 -2347 402
rect -2313 368 -2290 402
rect -2370 345 -2290 368
rect -2220 402 -2140 425
rect -2220 368 -2197 402
rect -2163 368 -2140 402
rect -2220 345 -2140 368
rect -2020 402 -1940 425
rect -2020 368 -1997 402
rect -1963 368 -1940 402
rect -2020 345 -1940 368
rect -2420 299 -2340 310
rect -2420 235 -2397 299
rect -2363 235 -2340 299
rect -2420 231 -2340 235
rect -2420 129 -2397 231
rect -2363 129 -2340 231
rect -2420 125 -2340 129
rect -2420 61 -2397 125
rect -2363 61 -2340 125
rect -2420 50 -2340 61
rect -2120 299 -2040 310
rect -2120 235 -2097 299
rect -2063 235 -2040 299
rect -2120 231 -2040 235
rect -2120 129 -2097 231
rect -2063 129 -2040 231
rect -2120 125 -2040 129
rect -2120 61 -2097 125
rect -2063 61 -2040 125
rect -2120 50 -2040 61
rect -1820 299 -1740 310
rect -1820 235 -1797 299
rect -1763 235 -1740 299
rect -1820 231 -1740 235
rect -1820 129 -1797 231
rect -1763 129 -1740 231
rect -1820 125 -1740 129
rect -1820 61 -1797 125
rect -1763 61 -1740 125
rect -1820 50 -1740 61
rect -1920 -23 -1840 0
rect -1920 -57 -1897 -23
rect -1863 -57 -1840 -23
rect -1920 -80 -1840 -57
rect -2520 -137 -1640 -114
rect -2520 -171 -2497 -137
rect -2463 -171 -2425 -137
rect -2391 -171 -2353 -137
rect -2319 -171 -2281 -137
rect -2247 -171 -2209 -137
rect -2175 -171 -2137 -137
rect -2103 -171 -2065 -137
rect -2031 -171 -1993 -137
rect -1959 -171 -1921 -137
rect -1887 -171 -1849 -137
rect -1815 -171 -1777 -137
rect -1743 -171 -1705 -137
rect -1671 -171 -1640 -137
rect -2520 -194 -1640 -171
<< viali >>
rect -2497 1407 -2463 1441
rect -2425 1407 -2391 1441
rect -2353 1407 -2319 1441
rect -2281 1407 -2247 1441
rect -2209 1407 -2175 1441
rect -2137 1407 -2103 1441
rect -2065 1407 -2031 1441
rect -1993 1407 -1959 1441
rect -1921 1407 -1887 1441
rect -1849 1407 -1815 1441
rect -1777 1407 -1743 1441
rect -1705 1407 -1671 1441
rect -2397 1195 -2363 1209
rect -2397 1175 -2363 1195
rect -2397 1127 -2363 1137
rect -2397 1103 -2363 1127
rect -2397 1059 -2363 1065
rect -2397 1031 -2363 1059
rect -2397 991 -2363 993
rect -2397 959 -2363 991
rect -2397 889 -2363 921
rect -2397 887 -2363 889
rect -2397 821 -2363 849
rect -2397 815 -2363 821
rect -2397 753 -2363 777
rect -2397 743 -2363 753
rect -2397 685 -2363 705
rect -2397 671 -2363 685
rect -2097 1195 -2063 1209
rect -2097 1175 -2063 1195
rect -2097 1127 -2063 1137
rect -2097 1103 -2063 1127
rect -2097 1059 -2063 1065
rect -2097 1031 -2063 1059
rect -2097 991 -2063 993
rect -2097 959 -2063 991
rect -2097 889 -2063 921
rect -2097 887 -2063 889
rect -2097 821 -2063 849
rect -2097 815 -2063 821
rect -2097 753 -2063 777
rect -2097 743 -2063 753
rect -2097 685 -2063 705
rect -2097 671 -2063 685
rect -1797 1195 -1763 1209
rect -1797 1175 -1763 1195
rect -1797 1127 -1763 1137
rect -1797 1103 -1763 1127
rect -1797 1059 -1763 1065
rect -1797 1031 -1763 1059
rect -1797 991 -1763 993
rect -1797 959 -1763 991
rect -1797 889 -1763 921
rect -1797 887 -1763 889
rect -1797 821 -1763 849
rect -1797 815 -1763 821
rect -1797 753 -1763 777
rect -1797 743 -1763 753
rect -1797 685 -1763 705
rect -1797 671 -1763 685
rect -1817 559 -1783 593
rect -2197 368 -2163 402
rect -2397 265 -2363 269
rect -2397 235 -2363 265
rect -2397 163 -2363 197
rect -2397 95 -2363 125
rect -2397 91 -2363 95
rect -2097 265 -2063 269
rect -2097 235 -2063 265
rect -2097 163 -2063 197
rect -2097 95 -2063 125
rect -2097 91 -2063 95
rect -1797 265 -1763 269
rect -1797 235 -1763 265
rect -1797 163 -1763 197
rect -1797 95 -1763 125
rect -1797 91 -1763 95
rect -2497 -171 -2463 -137
rect -2425 -171 -2391 -137
rect -2353 -171 -2319 -137
rect -2281 -171 -2247 -137
rect -2209 -171 -2175 -137
rect -2137 -171 -2103 -137
rect -2065 -171 -2031 -137
rect -1993 -171 -1959 -137
rect -1921 -171 -1887 -137
rect -1849 -171 -1815 -137
rect -1777 -171 -1743 -137
rect -1705 -171 -1671 -137
<< metal1 >>
rect -2520 1441 -1640 1474
rect -2520 1407 -2497 1441
rect -2463 1407 -2425 1441
rect -2391 1407 -2353 1441
rect -2319 1407 -2281 1441
rect -2247 1407 -2209 1441
rect -2175 1407 -2137 1441
rect -2103 1407 -2065 1441
rect -2031 1407 -1993 1441
rect -1959 1407 -1921 1441
rect -1887 1407 -1849 1441
rect -1815 1407 -1777 1441
rect -1743 1407 -1705 1441
rect -1671 1407 -1640 1441
rect -2520 1374 -1640 1407
rect -2400 1220 -2360 1374
rect -1800 1220 -1760 1374
rect -2420 1209 -2340 1220
rect -2420 1175 -2397 1209
rect -2363 1175 -2340 1209
rect -2420 1137 -2340 1175
rect -2420 1103 -2397 1137
rect -2363 1103 -2340 1137
rect -2420 1065 -2340 1103
rect -2420 1031 -2397 1065
rect -2363 1031 -2340 1065
rect -2420 993 -2340 1031
rect -2420 959 -2397 993
rect -2363 959 -2340 993
rect -2420 921 -2340 959
rect -2420 887 -2397 921
rect -2363 887 -2340 921
rect -2420 849 -2340 887
rect -2420 815 -2397 849
rect -2363 815 -2340 849
rect -2420 777 -2340 815
rect -2420 743 -2397 777
rect -2363 743 -2340 777
rect -2420 705 -2340 743
rect -2420 671 -2397 705
rect -2363 671 -2340 705
rect -2420 660 -2340 671
rect -2120 1218 -2040 1220
rect -2120 1166 -2106 1218
rect -2054 1166 -2040 1218
rect -2120 1146 -2040 1166
rect -2120 1094 -2106 1146
rect -2054 1094 -2040 1146
rect -2120 1074 -2040 1094
rect -2120 1022 -2106 1074
rect -2054 1022 -2040 1074
rect -2120 1002 -2040 1022
rect -2120 950 -2106 1002
rect -2054 950 -2040 1002
rect -2120 930 -2040 950
rect -2120 878 -2106 930
rect -2054 878 -2040 930
rect -2120 858 -2040 878
rect -2120 806 -2106 858
rect -2054 806 -2040 858
rect -2120 786 -2040 806
rect -2120 734 -2106 786
rect -2054 734 -2040 786
rect -2120 714 -2040 734
rect -2120 662 -2106 714
rect -2054 662 -2040 714
rect -2120 660 -2040 662
rect -1820 1209 -1740 1220
rect -1820 1175 -1797 1209
rect -1763 1175 -1740 1209
rect -1820 1137 -1740 1175
rect -1820 1103 -1797 1137
rect -1763 1103 -1740 1137
rect -1820 1065 -1740 1103
rect -1820 1031 -1797 1065
rect -1763 1031 -1740 1065
rect -1820 993 -1740 1031
rect -1820 959 -1797 993
rect -1763 959 -1740 993
rect -1820 921 -1740 959
rect -1820 887 -1797 921
rect -1763 887 -1740 921
rect -1820 849 -1740 887
rect -1820 815 -1797 849
rect -1763 815 -1740 849
rect -1820 777 -1740 815
rect -1820 743 -1797 777
rect -1763 743 -1740 777
rect -1820 705 -1740 743
rect -1820 671 -1797 705
rect -1763 671 -1740 705
rect -1820 660 -1740 671
rect -1840 593 -1760 616
rect -1840 559 -1817 593
rect -1783 559 -1760 593
rect -1840 536 -1760 559
rect -2220 405 -2140 425
rect -1820 405 -1781 536
rect -2220 402 -1781 405
rect -2220 368 -2197 402
rect -2163 368 -1781 402
rect -2220 365 -1781 368
rect -2220 345 -2140 365
rect -2420 269 -2340 310
rect -2420 235 -2397 269
rect -2363 235 -2340 269
rect -2420 197 -2340 235
rect -2420 163 -2397 197
rect -2363 163 -2340 197
rect -2420 125 -2340 163
rect -2420 91 -2397 125
rect -2363 91 -2340 125
rect -2420 50 -2340 91
rect -2120 278 -2040 310
rect -2120 226 -2106 278
rect -2054 226 -2040 278
rect -2120 206 -2040 226
rect -2120 154 -2106 206
rect -2054 154 -2040 206
rect -2120 134 -2040 154
rect -2120 82 -2106 134
rect -2054 82 -2040 134
rect -2120 50 -2040 82
rect -1820 269 -1740 310
rect -1820 235 -1797 269
rect -1763 235 -1740 269
rect -1820 197 -1740 235
rect -1820 163 -1797 197
rect -1763 163 -1740 197
rect -1820 125 -1740 163
rect -1820 91 -1797 125
rect -1763 91 -1740 125
rect -1820 50 -1740 91
rect -2400 -104 -2360 50
rect -1800 -104 -1760 50
rect -2520 -137 -1640 -104
rect -2520 -171 -2497 -137
rect -2463 -171 -2425 -137
rect -2391 -171 -2353 -137
rect -2319 -171 -2281 -137
rect -2247 -171 -2209 -137
rect -2175 -171 -2137 -137
rect -2103 -171 -2065 -137
rect -2031 -171 -1993 -137
rect -1959 -171 -1921 -137
rect -1887 -171 -1849 -137
rect -1815 -171 -1777 -137
rect -1743 -171 -1705 -137
rect -1671 -171 -1640 -137
rect -2520 -204 -1640 -171
<< via1 >>
rect -2106 1209 -2054 1218
rect -2106 1175 -2097 1209
rect -2097 1175 -2063 1209
rect -2063 1175 -2054 1209
rect -2106 1166 -2054 1175
rect -2106 1137 -2054 1146
rect -2106 1103 -2097 1137
rect -2097 1103 -2063 1137
rect -2063 1103 -2054 1137
rect -2106 1094 -2054 1103
rect -2106 1065 -2054 1074
rect -2106 1031 -2097 1065
rect -2097 1031 -2063 1065
rect -2063 1031 -2054 1065
rect -2106 1022 -2054 1031
rect -2106 993 -2054 1002
rect -2106 959 -2097 993
rect -2097 959 -2063 993
rect -2063 959 -2054 993
rect -2106 950 -2054 959
rect -2106 921 -2054 930
rect -2106 887 -2097 921
rect -2097 887 -2063 921
rect -2063 887 -2054 921
rect -2106 878 -2054 887
rect -2106 849 -2054 858
rect -2106 815 -2097 849
rect -2097 815 -2063 849
rect -2063 815 -2054 849
rect -2106 806 -2054 815
rect -2106 777 -2054 786
rect -2106 743 -2097 777
rect -2097 743 -2063 777
rect -2063 743 -2054 777
rect -2106 734 -2054 743
rect -2106 705 -2054 714
rect -2106 671 -2097 705
rect -2097 671 -2063 705
rect -2063 671 -2054 705
rect -2106 662 -2054 671
rect -2106 269 -2054 278
rect -2106 235 -2097 269
rect -2097 235 -2063 269
rect -2063 235 -2054 269
rect -2106 226 -2054 235
rect -2106 197 -2054 206
rect -2106 163 -2097 197
rect -2097 163 -2063 197
rect -2063 163 -2054 197
rect -2106 154 -2054 163
rect -2106 125 -2054 134
rect -2106 91 -2097 125
rect -2097 91 -2063 125
rect -2063 91 -2054 125
rect -2106 82 -2054 91
<< metal2 >>
rect -2120 1218 -2040 1220
rect -2120 1166 -2106 1218
rect -2054 1166 -2040 1218
rect -2120 1146 -2040 1166
rect -2120 1094 -2106 1146
rect -2054 1094 -2040 1146
rect -2120 1074 -2040 1094
rect -2120 1022 -2106 1074
rect -2054 1022 -2040 1074
rect -2120 1002 -2040 1022
rect -2120 950 -2106 1002
rect -2054 950 -2040 1002
rect -2120 930 -2040 950
rect -2120 878 -2106 930
rect -2054 878 -2040 930
rect -2120 858 -2040 878
rect -2120 806 -2106 858
rect -2054 806 -2040 858
rect -2120 786 -2040 806
rect -2120 734 -2106 786
rect -2054 734 -2040 786
rect -2120 714 -2040 734
rect -2120 662 -2106 714
rect -2054 662 -2040 714
rect -2120 660 -2040 662
rect -2100 504 -2060 660
rect -2100 464 -1650 504
rect -2100 310 -2060 464
rect -2120 278 -2040 310
rect -2120 226 -2106 278
rect -2054 226 -2040 278
rect -2120 206 -2040 226
rect -2120 154 -2106 206
rect -2054 154 -2040 206
rect -2120 134 -2040 154
rect -2120 82 -2106 134
rect -2054 82 -2040 134
rect -2120 50 -2040 82
<< labels >>
rlabel metal1 s -2140 -174 -2100 -134 4 GND!
port 1 nsew
rlabel metal1 s -2140 1404 -2100 1444 4 VDD
port 2 nsew
flabel locali s -1897 1293 -1863 1327 2 FreeSans 2500 0 0 0 B
port 3 nsew
flabel locali s -1897 -57 -1863 -23 2 FreeSans 2500 0 0 0 A_bar
port 4 nsew
flabel locali s -2347 368 -2313 402 2 FreeSans 2500 0 0 0 A
port 5 nsew
rlabel locali s -2383 551 -2334 598 4 B_bar
port 6 nsew
flabel metal2 s -1740 466 -1704 502 2 FreeSans 2500 0 0 0 XOR
port 7 nsew
<< end >>
